magic
tech sky130A
magscale 1 2
timestamp 1699069426
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1931 203
rect 29 -17 63 21
<< locali >>
rect 1833 59 1903 93
rect 1869 93 1903 127
rect 1869 127 1915 161
rect 1881 161 1915 315
rect 1869 315 1915 349
rect 1869 349 1903 451
rect 1833 451 1903 485
rect 1605 215 1761 249
rect 1605 249 1639 255
rect 1685 249 1719 255
rect 1605 255 1639 299
rect 1593 299 1639 333
rect 1593 333 1627 391
rect 29 215 117 249
rect 29 249 63 323
rect 307 199 341 215
rect 305 215 341 255
rect 307 255 341 265
<< obsli1 >>
rect 121 435 155 527
rect 63 527 121 561
rect 155 527 213 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 749 375 951 409
rect 749 409 783 493
rect 917 409 951 493
rect 189 67 267 101
rect 233 101 267 357
rect 205 357 267 391
rect 205 391 239 493
rect 1569 59 1719 93
rect 1685 93 1719 143
rect 1685 143 1831 177
rect 1797 177 1831 199
rect 1797 199 1841 265
rect 1797 265 1831 289
rect 1777 289 1831 323
rect 1797 323 1831 367
rect 1669 367 1831 401
rect 1669 401 1703 493
rect 405 51 439 127
rect 377 127 439 161
rect 377 161 411 375
rect 377 375 439 409
rect 405 409 439 493
rect 1105 51 1139 127
rect 1041 127 1139 161
rect 1041 161 1075 199
rect 779 199 813 215
rect 1041 199 1075 215
rect 779 215 815 265
rect 1041 215 1075 265
rect 781 265 815 299
rect 1041 265 1075 299
rect 781 299 1075 333
rect 1041 333 1075 357
rect 1041 357 1123 391
rect 1089 391 1123 451
rect 1089 451 1167 485
rect 1185 59 1415 93
rect 1381 93 1415 127
rect 1381 127 1547 161
rect 1513 161 1547 199
rect 1513 199 1565 265
rect 1513 265 1547 357
rect 1405 357 1547 391
rect 1405 391 1439 451
rect 1281 451 1439 485
rect 29 51 71 125
rect 37 125 71 143
rect 37 143 195 177
rect 161 177 195 199
rect 161 199 197 265
rect 161 265 195 289
rect 121 289 195 323
rect 121 323 155 367
rect 21 367 155 401
rect 21 401 87 485
rect 569 59 743 93
rect 709 93 743 127
rect 709 127 1003 161
rect 709 161 743 199
rect 969 161 1003 199
rect 709 199 743 249
rect 969 199 1005 249
rect 709 249 743 265
rect 971 249 1005 265
rect 709 265 743 299
rect 681 299 743 333
rect 681 333 715 443
rect 485 443 715 477
rect 1147 199 1181 215
rect 1339 199 1373 215
rect 1147 215 1191 265
rect 1329 215 1373 265
rect 1157 265 1191 357
rect 1329 265 1363 357
rect 1157 357 1363 391
rect 447 199 481 215
rect 639 199 673 215
rect 447 215 483 265
rect 613 215 673 265
rect 449 265 483 299
rect 613 265 647 299
rect 449 299 647 333
rect 581 333 615 391
rect 1435 199 1469 215
rect 1409 215 1469 265
rect 1409 265 1443 323
rect 1243 199 1277 215
rect 1225 215 1277 265
rect 1225 265 1259 323
rect 489 85 523 127
rect 489 127 575 161
rect 541 161 575 199
rect 541 199 577 249
rect 543 249 577 265
rect 875 199 909 221
rect 857 221 909 255
rect 875 255 909 265
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 527 29 561
rect 309 427 343 527
rect 339 527 397 561
rect 247 527 305 561
rect 1021 427 1055 527
rect 983 527 1041 561
rect 891 527 949 561
rect 1765 435 1799 527
rect 1719 527 1777 561
rect 1627 527 1685 561
rect 1481 435 1619 527
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1351 527 1409 561
rect 1259 527 1317 561
rect 1167 527 1225 561
rect 1075 527 1133 561
rect 817 451 883 527
rect 799 527 857 561
rect 707 527 765 561
rect 615 527 673 561
rect 523 527 581 561
rect 431 527 489 561
rect 1719 -17 1777 17
rect 1765 17 1799 109
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1465 17 1531 93
rect 1351 -17 1409 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 901 17 1071 93
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 309 17 343 109
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 121 17 155 109
rect 0 -17 29 17
<< obsli1c >>
rect 121 527 155 561
rect 765 527 799 561
rect 1685 527 1719 561
rect 489 527 523 561
rect 1317 527 1351 561
rect 1133 527 1167 561
rect 1593 527 1627 561
rect 397 527 431 561
rect 857 527 891 561
rect 305 527 339 561
rect 581 527 615 561
rect 1409 527 1443 561
rect 949 527 983 561
rect 1869 527 1903 561
rect 673 527 707 561
rect 29 527 63 561
rect 1041 527 1075 561
rect 1501 527 1535 561
rect 213 527 247 561
rect 1225 527 1259 561
rect 1777 527 1811 561
rect 213 -17 247 17
rect 1869 -17 1903 17
rect 1777 -17 1811 17
rect 765 -17 799 17
rect 1133 -17 1167 17
rect 1501 -17 1535 17
rect 1409 -17 1443 17
rect 581 -17 615 17
rect 1041 -17 1075 17
rect 1225 -17 1259 17
rect 673 -17 707 17
rect 1317 -17 1351 17
rect 29 -17 63 17
rect 1593 -17 1627 17
rect 949 -17 983 17
rect 121 -17 155 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 857 -17 891 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 496 1932 527
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 561 1932 592
rect 0 -48 1932 -17
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 17 1932 48
<< obsm1 >>
rect 201 351 259 360
rect 569 351 627 360
rect 1305 351 1363 360
rect 201 360 1363 388
rect 201 388 259 397
rect 569 388 627 397
rect 1305 388 1363 397
rect 1397 283 1455 292
rect 1765 283 1823 292
rect 1397 292 1823 320
rect 1397 320 1455 329
rect 1765 320 1823 329
rect 109 283 167 292
rect 1213 283 1271 292
rect 109 292 1271 320
rect 109 320 167 329
rect 1213 320 1271 329
rect 845 215 903 224
rect 1673 215 1731 224
rect 845 224 1731 252
rect 845 252 903 261
rect 1673 252 1731 261
rect 17 79 75 88
rect 477 79 535 88
rect 17 88 535 116
rect 17 116 75 125
rect 477 116 535 125
<< labels >>
rlabel locali s 29 215 117 249 6 CLK
port 1 nsew signal input
rlabel locali s 29 249 63 323 6 CLK
port 1 nsew signal input
rlabel locali s 307 199 341 215 6 D
port 2 nsew signal input
rlabel locali s 305 215 341 255 6 D
port 2 nsew signal input
rlabel locali s 307 255 341 265 6 D
port 2 nsew signal input
rlabel locali s 1605 215 1761 249 6 RESET_B
port 3 nsew signal input
rlabel locali s 1605 249 1639 255 6 RESET_B
port 3 nsew signal input
rlabel locali s 1685 249 1719 255 6 RESET_B
port 3 nsew signal input
rlabel locali s 1605 255 1639 299 6 RESET_B
port 3 nsew signal input
rlabel locali s 1593 299 1639 333 6 RESET_B
port 3 nsew signal input
rlabel locali s 1593 333 1627 391 6 RESET_B
port 3 nsew signal input
rlabel locali s 1833 59 1903 93 6 Q
port 8 nsew signal output
rlabel locali s 1869 93 1903 127 6 Q
port 8 nsew signal output
rlabel locali s 1869 127 1915 161 6 Q
port 8 nsew signal output
rlabel locali s 1881 161 1915 315 6 Q
port 8 nsew signal output
rlabel locali s 1869 315 1915 349 6 Q
port 8 nsew signal output
rlabel locali s 1869 349 1903 451 6 Q
port 8 nsew signal output
rlabel locali s 1833 451 1903 485 6 Q
port 8 nsew signal output
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1931 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1970 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 -48 1932 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 6 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ht_sc_tt05.gds
string GDS_START 23860
string GDS_END 37716
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
