magic
tech sky130A
magscale 1 2
timestamp 1698685089
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 827 203
rect 29 -17 63 21
<< scnmos >>
rect 81 47 111 177
rect 173 47 203 177
rect 257 47 287 177
rect 341 47 371 177
rect 425 47 455 177
rect 509 47 539 177
rect 601 47 631 177
rect 717 47 747 177
<< scpmoshvt >>
rect 81 297 111 497
rect 173 297 203 497
rect 257 297 287 497
rect 341 297 371 497
rect 425 297 455 497
rect 509 297 539 497
rect 601 297 631 497
rect 717 297 747 497
<< ndiff >>
rect 747 47 799 59
rect 747 59 757 93
rect 791 59 799 93
rect 747 93 799 127
rect 747 127 757 161
rect 791 127 799 161
rect 747 161 799 177
rect 631 47 717 59
rect 631 59 673 93
rect 707 59 717 93
rect 631 93 717 127
rect 631 127 673 161
rect 707 127 717 161
rect 631 161 717 177
rect 539 47 601 59
rect 539 59 557 93
rect 591 59 601 93
rect 539 93 601 177
rect 455 47 509 177
rect 371 47 425 59
rect 371 59 381 93
rect 415 59 425 93
rect 371 93 425 177
rect 287 47 341 177
rect 203 47 257 59
rect 203 59 213 93
rect 247 59 257 93
rect 203 93 257 177
rect 111 47 173 177
rect 29 47 81 59
rect 29 59 37 93
rect 71 59 81 93
rect 29 93 81 177
<< pdiff >>
rect 631 297 717 315
rect 631 315 673 349
rect 707 315 717 349
rect 631 349 717 383
rect 631 383 673 417
rect 707 383 717 417
rect 631 417 717 451
rect 631 451 673 485
rect 707 451 717 485
rect 631 485 717 497
rect 539 297 601 383
rect 539 383 557 417
rect 591 383 601 417
rect 539 417 601 451
rect 539 451 557 485
rect 591 451 601 485
rect 539 485 601 497
rect 455 297 509 497
rect 371 297 425 383
rect 371 383 381 417
rect 415 383 425 417
rect 371 417 425 451
rect 371 451 381 485
rect 415 451 425 485
rect 371 485 425 497
rect 287 297 341 497
rect 203 297 257 451
rect 203 451 213 485
rect 247 451 257 485
rect 203 485 257 497
rect 111 297 173 497
rect 29 297 81 383
rect 29 383 37 417
rect 71 383 81 417
rect 29 417 81 451
rect 29 451 37 485
rect 71 451 81 485
rect 29 485 81 497
rect 747 297 799 315
rect 747 315 757 349
rect 791 315 799 349
rect 747 349 799 383
rect 747 383 757 417
rect 791 383 799 417
rect 747 417 799 451
rect 747 451 757 485
rect 791 451 799 485
rect 747 485 799 497
<< ndiffc >>
rect 757 127 791 161
rect 673 127 707 161
rect 37 59 71 93
rect 673 59 707 93
rect 381 59 415 93
rect 757 59 791 93
rect 213 59 247 93
rect 557 59 591 93
<< pdiffc >>
rect 757 451 791 485
rect 381 451 415 485
rect 673 451 707 485
rect 213 451 247 485
rect 557 451 591 485
rect 37 451 71 485
rect 757 383 791 417
rect 381 383 415 417
rect 557 383 591 417
rect 37 383 71 417
rect 673 383 707 417
rect 757 315 791 349
rect 673 315 707 349
<< poly >>
rect 509 497 539 523
rect 425 497 455 523
rect 341 497 371 523
rect 81 497 111 523
rect 257 497 287 523
rect 173 497 203 523
rect 717 497 747 523
rect 601 497 631 523
rect 173 177 203 199
rect 257 177 287 199
rect 173 199 287 215
rect 173 215 211 249
rect 245 215 287 249
rect 173 249 287 265
rect 173 265 203 297
rect 257 265 287 297
rect 601 177 631 199
rect 717 177 747 199
rect 601 199 747 215
rect 601 215 611 249
rect 645 215 747 249
rect 601 249 747 265
rect 601 265 631 297
rect 717 265 747 297
rect 509 177 539 199
rect 497 199 551 215
rect 497 215 507 249
rect 541 215 551 249
rect 497 249 551 265
rect 509 265 539 297
rect 341 177 371 199
rect 425 177 455 199
rect 341 199 455 215
rect 341 215 379 249
rect 413 215 455 249
rect 341 249 455 265
rect 341 265 371 297
rect 425 265 455 297
rect 81 177 111 199
rect 77 199 131 215
rect 77 215 87 249
rect 121 215 131 249
rect 77 249 131 265
rect 81 265 111 297
rect 173 21 203 47
rect 81 21 111 47
rect 257 21 287 47
rect 341 21 371 47
rect 425 21 455 47
rect 509 21 539 47
rect 601 21 631 47
rect 717 21 747 47
<< polycont >>
rect 507 215 541 249
rect 87 215 121 249
rect 211 215 245 249
rect 379 215 413 249
rect 611 215 645 249
<< locali >>
rect 197 451 213 485
rect 247 451 263 485
rect 197 485 263 527
rect 155 527 213 561
rect 247 527 305 561
rect 799 527 828 561
rect 17 59 37 93
rect 71 59 87 93
rect 365 59 381 93
rect 415 59 431 93
rect 17 93 87 127
rect 365 93 431 127
rect 17 127 623 161
rect 17 161 51 199
rect 589 161 623 199
rect 17 199 51 215
rect 589 199 645 215
rect 17 215 51 249
rect 589 215 611 249
rect 17 249 51 265
rect 611 249 645 265
rect 17 265 51 383
rect 17 383 37 417
rect 71 383 381 417
rect 415 383 431 417
rect 17 417 87 451
rect 365 417 431 451
rect 17 451 37 485
rect 71 451 87 485
rect 365 451 381 485
rect 415 451 431 485
rect 657 59 673 93
rect 707 59 723 93
rect 657 93 723 127
rect 657 127 673 161
rect 707 127 723 161
rect 689 161 723 315
rect 657 315 673 349
rect 707 315 723 349
rect 657 349 723 383
rect 657 383 673 417
rect 707 383 723 417
rect 657 417 723 451
rect 657 451 673 485
rect 707 451 723 485
rect 757 417 791 451
rect 757 349 791 383
rect 87 199 149 215
rect 121 215 149 221
rect 121 221 155 249
rect 489 221 507 249
rect 87 249 155 265
rect 489 249 541 265
rect 121 265 155 315
rect 489 265 523 315
rect 121 315 523 349
rect 757 299 791 315
rect 413 221 431 249
rect 379 249 431 255
rect 379 255 413 265
rect 245 221 339 249
rect 211 249 339 255
rect 211 255 245 265
rect 379 199 413 215
rect 507 199 541 215
rect 211 199 245 215
rect 757 161 791 177
rect 757 93 791 127
rect 799 -17 828 17
rect 63 527 121 561
rect 0 527 29 561
rect 757 485 791 527
rect 707 527 765 561
rect 615 527 673 561
rect 541 383 557 417
rect 591 383 607 417
rect 541 417 607 451
rect 541 451 557 485
rect 591 451 607 485
rect 541 485 607 527
rect 523 527 581 561
rect 431 527 489 561
rect 339 527 397 561
rect 707 -17 765 17
rect 757 17 791 59
rect 523 -17 581 17
rect 615 -17 673 17
rect 541 17 607 59
rect 541 59 557 93
rect 591 59 607 93
rect 431 -17 489 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 197 17 263 59
rect 197 59 213 93
rect 247 59 263 93
rect 0 -17 29 17
rect 63 -17 121 17
<< viali >>
rect 305 527 339 561
rect 765 527 799 561
rect 213 527 247 561
rect 673 527 707 561
rect 121 527 155 561
rect 581 527 615 561
rect 29 527 63 561
rect 489 527 523 561
rect 397 527 431 561
rect 121 -17 155 17
rect 765 -17 799 17
rect 397 -17 431 17
rect 29 -17 63 17
rect 673 -17 707 17
rect 305 -17 339 17
rect 581 -17 615 17
rect 213 -17 247 17
rect 489 -17 523 17
<< metal1 >>
rect 0 496 828 527
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 561 828 592
rect 0 -48 828 -17
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 17 828 48
<< labels >>
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 A
port 5 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 B
port 6 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel locali s 489 289 523 323 0 FreeSans 200 0 0 0 C
port 7 nsew signal input
flabel locali s 673 85 707 119 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 -48 828 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 4 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 maj3_2
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ht_sc_tt05.gds
string GDS_START 7312
string GDS_END 13152
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
