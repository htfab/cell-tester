magic
tech sky130A
magscale 1 2
timestamp 1698890999
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 1 21 1379 203
rect 29 -17 63 21
<< locali >>
rect 1273 59 1363 119
rect 1329 119 1363 357
rect 1273 357 1363 485
rect 31 199 65 221
rect 29 221 65 265
rect 29 265 63 323
rect 303 215 369 255
rect 1133 85 1167 215
rect 1133 215 1201 249
rect 1133 249 1167 255
<< obsli1 >>
rect 105 451 171 527
rect 63 527 121 561
rect 155 527 213 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 309 51 343 143
rect 309 143 439 177
rect 405 177 439 199
rect 405 199 481 265
rect 405 265 439 289
rect 309 289 439 323
rect 309 323 343 493
rect 21 127 155 161
rect 121 161 155 199
rect 121 199 197 265
rect 121 265 159 323
rect 121 323 155 375
rect 21 375 155 409
rect 37 409 71 493
rect 205 351 251 493
rect 605 127 671 143
rect 605 143 891 177
rect 857 177 891 289
rect 857 289 895 323
rect 857 323 891 357
rect 841 357 891 391
rect 841 391 875 451
rect 713 451 875 485
rect 1093 451 1159 485
rect 497 451 671 485
rect 977 59 1063 93
rect 977 93 1011 143
rect 941 143 1011 177
rect 941 177 975 199
rect 939 199 975 215
rect 1259 199 1293 215
rect 939 215 975 265
rect 1257 215 1293 265
rect 941 265 975 289
rect 1257 265 1291 289
rect 941 289 975 323
rect 1133 289 1291 323
rect 941 323 975 357
rect 1133 323 1167 357
rect 941 357 1167 391
rect 489 85 551 119
rect 517 119 551 215
rect 517 215 605 249
rect 755 215 821 249
rect 517 249 551 357
rect 773 249 807 357
rect 489 357 807 391
rect 647 215 713 255
rect 673 255 711 323
rect 1027 215 1093 249
rect 1041 249 1075 289
rect 1041 289 1079 323
rect 205 51 251 125
rect 1351 -17 1380 17
rect 713 59 875 93
rect 0 527 29 561
rect 909 435 1047 527
rect 891 527 949 561
rect 983 527 1041 561
rect 799 527 857 561
rect 707 527 765 561
rect 615 527 673 561
rect 523 527 581 561
rect 1205 435 1239 527
rect 1167 527 1225 561
rect 1075 527 1133 561
rect 405 367 439 527
rect 431 527 489 561
rect 339 527 397 561
rect 247 527 305 561
rect 1259 -17 1317 17
rect 1167 -17 1225 17
rect 1205 17 1239 109
rect 1075 -17 1133 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 909 17 943 109
rect 799 -17 857 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 389 17 455 93
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 105 17 171 93
rect 0 -17 29 17
<< obsli1c >>
rect 305 527 339 561
rect 29 527 63 561
rect 213 527 247 561
rect 121 527 155 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 857 -17 891 17
rect 1133 -17 1167 17
rect 673 -17 707 17
rect 949 -17 983 17
rect 581 -17 615 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 121 -17 155 17
rect 29 -17 63 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 1041 -17 1075 17
rect 765 -17 799 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 496 1380 527
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 561 1380 592
rect 0 -48 1380 -17
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 17 1380 48
<< obsm1 >>
rect 201 351 259 360
rect 477 351 535 360
rect 201 360 535 388
rect 201 388 259 397
rect 477 388 535 397
rect 845 283 903 292
rect 1029 283 1087 292
rect 845 292 1087 320
rect 845 320 903 329
rect 1029 320 1087 329
rect 109 283 167 292
rect 661 283 719 292
rect 109 292 719 320
rect 109 320 167 329
rect 661 320 719 329
rect 201 79 259 88
rect 477 79 535 88
rect 201 88 535 116
rect 201 116 259 125
rect 477 116 535 125
<< labels >>
rlabel locali s 31 199 65 221 6 GATE
port 5 nsew signal input
rlabel locali s 29 221 65 265 6 GATE
port 5 nsew signal input
rlabel locali s 29 265 63 323 6 GATE
port 5 nsew signal input
rlabel locali s 303 215 369 255 6 D
port 6 nsew signal input
rlabel locali s 1133 85 1167 215 6 RESET_B
port 7 nsew signal input
rlabel locali s 1133 215 1201 249 6 RESET_B
port 7 nsew signal input
rlabel locali s 1133 249 1167 255 6 RESET_B
port 7 nsew signal input
rlabel locali s 1273 59 1363 119 6 Q
port 8 nsew signal output
rlabel locali s 1329 119 1363 357 6 Q
port 8 nsew signal output
rlabel locali s 1273 357 1363 485 6 Q
port 8 nsew signal output
rlabel pwell s 30 -17 64 21 6 VNB
port 1 nsew ground bidirectional
rlabel pwell s 1 21 1379 203 6 VNB
port 1 nsew ground bidirectional
rlabel nwell s -38 261 1418 582 6 VPB
port 2 nsew power bidirectional
rlabel metal1 s 0 -48 1380 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1380 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1380 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ht_sc_tt05.gds
string GDS_START 13210
string GDS_END 24074
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
