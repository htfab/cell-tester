magic
tech sky130A
magscale 1 2
timestamp 1698676621
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 1 21 1379 203
rect 29 -17 63 21
<< scnmos >>
rect 1055 47 1085 177
rect 1151 47 1181 177
rect 1247 47 1277 177
rect 79 47 109 177
rect 163 47 193 177
rect 351 47 381 177
rect 447 47 477 177
rect 555 47 585 177
rect 663 47 693 177
rect 771 47 801 177
rect 867 47 897 177
<< scpmoshvt >>
rect 1055 297 1085 497
rect 1151 297 1181 497
rect 1247 297 1277 497
rect 79 297 109 497
rect 163 297 193 497
rect 351 297 381 497
rect 447 297 477 497
rect 555 297 585 497
rect 663 297 693 497
rect 771 297 801 497
rect 867 297 897 497
<< ndiff >>
rect 801 47 867 59
rect 801 59 823 93
rect 857 59 867 93
rect 801 93 867 177
rect 897 47 949 59
rect 897 59 907 93
rect 941 59 949 93
rect 897 93 949 177
rect 693 47 771 59
rect 693 59 727 93
rect 761 59 771 93
rect 693 93 771 177
rect 585 47 663 127
rect 585 127 619 161
rect 653 127 663 161
rect 585 161 663 177
rect 477 47 555 177
rect 381 47 447 59
rect 381 59 403 93
rect 437 59 447 93
rect 381 93 447 177
rect 193 47 245 67
rect 193 67 203 101
rect 237 67 245 101
rect 193 101 245 177
rect 109 47 163 59
rect 109 59 119 93
rect 153 59 163 93
rect 109 93 163 177
rect 1277 47 1329 59
rect 1277 59 1287 93
rect 1321 59 1329 93
rect 1277 93 1329 177
rect 1181 47 1247 59
rect 1181 59 1203 93
rect 1237 59 1247 93
rect 1181 93 1247 177
rect 1085 47 1151 177
rect 1003 47 1055 59
rect 1003 59 1011 93
rect 1045 59 1055 93
rect 1003 93 1055 177
rect 27 47 79 127
rect 27 127 35 161
rect 69 127 79 161
rect 27 161 79 177
rect 299 47 351 67
rect 299 67 307 101
rect 341 67 351 101
rect 299 101 351 177
<< pdiff >>
rect 801 297 867 497
rect 897 297 949 451
rect 897 451 907 485
rect 941 451 949 485
rect 897 485 949 497
rect 299 297 351 375
rect 299 375 307 409
rect 341 375 351 409
rect 299 409 351 443
rect 299 443 307 477
rect 341 443 351 477
rect 299 477 351 497
rect 27 297 79 375
rect 27 375 35 409
rect 69 375 79 409
rect 27 409 79 443
rect 27 443 35 477
rect 69 443 79 477
rect 27 477 79 497
rect 1003 297 1055 451
rect 1003 451 1011 485
rect 1045 451 1055 485
rect 1003 485 1055 497
rect 1085 297 1151 357
rect 1085 357 1107 391
rect 1141 357 1151 391
rect 1085 391 1151 451
rect 1085 451 1107 485
rect 1141 451 1151 485
rect 1085 485 1151 497
rect 1181 297 1247 451
rect 1181 451 1203 485
rect 1237 451 1247 485
rect 1181 485 1247 497
rect 1277 297 1329 383
rect 1277 383 1287 417
rect 1321 383 1329 417
rect 1277 417 1329 451
rect 1277 451 1287 485
rect 1321 451 1329 485
rect 1277 485 1329 497
rect 109 297 163 451
rect 109 451 119 485
rect 153 451 163 485
rect 109 485 163 497
rect 193 297 245 375
rect 193 375 203 409
rect 237 375 245 409
rect 193 409 245 443
rect 193 443 203 477
rect 237 443 245 477
rect 193 477 245 497
rect 381 297 447 383
rect 381 383 403 417
rect 437 383 447 417
rect 381 417 447 451
rect 381 451 403 485
rect 437 451 447 485
rect 381 485 447 497
rect 477 297 555 451
rect 477 451 511 485
rect 545 451 555 485
rect 477 485 555 497
rect 585 297 663 451
rect 585 451 619 485
rect 653 451 663 485
rect 585 485 663 497
rect 693 297 771 451
rect 693 451 727 485
rect 761 451 771 485
rect 693 485 771 497
<< ndiffc >>
rect 619 127 653 161
rect 35 127 69 161
rect 307 67 341 101
rect 203 67 237 101
rect 727 59 761 93
rect 1011 59 1045 93
rect 1287 59 1321 93
rect 907 59 941 93
rect 1203 59 1237 93
rect 119 59 153 93
rect 823 59 857 93
rect 403 59 437 93
<< pdiffc >>
rect 1011 451 1045 485
rect 511 451 545 485
rect 1203 451 1237 485
rect 403 451 437 485
rect 619 451 653 485
rect 119 451 153 485
rect 907 451 941 485
rect 1107 451 1141 485
rect 727 451 761 485
rect 1287 451 1321 485
rect 35 443 69 477
rect 203 443 237 477
rect 307 443 341 477
rect 1287 383 1321 417
rect 403 383 437 417
rect 35 375 69 409
rect 307 375 341 409
rect 203 375 237 409
rect 1107 357 1141 391
<< poly >>
rect 163 497 193 523
rect 1247 497 1277 523
rect 1151 497 1181 523
rect 1055 497 1085 523
rect 867 497 897 523
rect 771 497 801 523
rect 663 497 693 523
rect 555 497 585 523
rect 447 497 477 523
rect 351 497 381 523
rect 79 497 109 523
rect 1055 177 1085 199
rect 1031 199 1085 215
rect 1031 215 1041 249
rect 1075 215 1085 249
rect 1031 249 1085 265
rect 1055 265 1085 297
rect 79 177 109 199
rect 19 199 109 215
rect 19 215 29 249
rect 63 215 109 249
rect 19 249 109 265
rect 79 265 109 297
rect 867 177 897 199
rect 867 199 973 215
rect 867 215 929 249
rect 963 215 973 249
rect 867 249 973 265
rect 867 265 897 297
rect 771 177 801 199
rect 759 199 813 215
rect 759 215 769 249
rect 803 215 813 249
rect 759 249 813 265
rect 771 265 801 297
rect 663 177 693 199
rect 651 199 705 215
rect 651 215 661 249
rect 695 215 705 249
rect 651 249 705 265
rect 663 265 693 297
rect 555 177 585 199
rect 543 199 597 215
rect 543 215 553 249
rect 587 215 597 249
rect 543 249 597 265
rect 555 265 585 297
rect 351 177 381 199
rect 307 199 381 215
rect 307 215 317 249
rect 351 215 381 249
rect 307 249 381 265
rect 351 265 381 297
rect 163 177 193 199
rect 151 199 205 215
rect 151 215 161 249
rect 195 215 205 249
rect 151 249 205 265
rect 163 265 193 297
rect 1151 177 1181 199
rect 1139 199 1193 215
rect 1139 215 1149 249
rect 1183 215 1193 249
rect 1139 249 1193 265
rect 1151 265 1181 297
rect 447 177 477 199
rect 435 199 489 215
rect 435 215 445 249
rect 479 215 489 249
rect 435 249 489 265
rect 447 265 477 297
rect 1247 177 1277 199
rect 1247 199 1301 215
rect 1247 215 1257 249
rect 1291 215 1301 249
rect 1247 249 1301 265
rect 1247 265 1277 297
rect 79 21 109 47
rect 867 21 897 47
rect 771 21 801 47
rect 663 21 693 47
rect 555 21 585 47
rect 447 21 477 47
rect 351 21 381 47
rect 1247 21 1277 47
rect 1151 21 1181 47
rect 1055 21 1085 47
rect 163 21 193 47
<< polycont >>
rect 553 215 587 249
rect 661 215 695 249
rect 769 215 803 249
rect 317 215 351 249
rect 1257 215 1291 249
rect 929 215 963 249
rect 1149 215 1183 249
rect 445 215 479 249
rect 29 215 63 249
rect 161 215 195 249
rect 1041 215 1075 249
<< locali >>
rect 103 451 119 485
rect 153 451 169 485
rect 103 485 169 527
rect 63 527 121 561
rect 155 527 213 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 35 477 69 493
rect 307 477 341 493
rect 203 351 249 357
rect 203 357 213 375
rect 247 357 249 375
rect 247 375 249 391
rect 237 391 249 409
rect 203 409 249 443
rect 237 443 249 477
rect 203 477 249 493
rect 545 451 619 485
rect 1271 59 1287 93
rect 1321 59 1361 93
rect 1271 93 1361 119
rect 1327 119 1361 357
rect 1271 357 1361 383
rect 1271 383 1287 417
rect 1321 383 1361 417
rect 1271 417 1361 451
rect 1271 451 1287 485
rect 1321 451 1361 485
rect 603 127 619 143
rect 653 127 669 143
rect 603 143 619 161
rect 653 143 889 161
rect 603 161 889 177
rect 855 177 889 289
rect 855 289 857 323
rect 855 323 889 357
rect 839 357 889 391
rect 839 391 873 451
rect 761 451 873 485
rect 1141 451 1157 485
rect 653 451 669 485
rect 495 451 511 485
rect 711 451 727 485
rect 1091 451 1107 485
rect 403 417 437 451
rect 1203 435 1237 451
rect 307 409 341 443
rect 69 127 153 161
rect 119 161 153 199
rect 119 199 195 215
rect 119 215 161 249
rect 119 249 195 265
rect 119 265 157 289
rect 119 289 121 323
rect 155 289 157 323
rect 119 323 153 375
rect 19 375 35 409
rect 69 375 153 409
rect 35 409 69 443
rect 523 85 549 119
rect 515 119 549 215
rect 515 215 553 249
rect 803 215 819 249
rect 515 249 549 357
rect 771 249 805 357
rect 523 357 805 391
rect 975 59 1011 93
rect 975 93 1009 143
rect 931 143 1009 177
rect 931 177 965 199
rect 929 199 965 215
rect 963 215 965 249
rect 929 249 965 265
rect 931 265 965 357
rect 931 357 1107 391
rect 1257 199 1291 215
rect 1255 215 1257 249
rect 1255 249 1291 265
rect 1255 265 1289 289
rect 1131 289 1289 323
rect 1131 323 1165 357
rect 1141 357 1165 391
rect 403 367 437 383
rect 307 101 341 143
rect 307 143 437 177
rect 403 177 437 199
rect 403 199 479 215
rect 403 215 445 249
rect 403 249 479 265
rect 403 265 437 289
rect 307 289 437 323
rect 307 323 341 375
rect 1025 215 1041 249
rect 1039 249 1073 289
rect 1039 289 1041 323
rect 645 215 661 249
rect 695 215 711 249
rect 645 249 711 255
rect 671 255 709 289
rect 671 289 673 323
rect 707 289 709 323
rect 27 221 29 249
rect 63 221 65 249
rect 27 249 65 323
rect 1075 289 1077 323
rect 301 215 317 249
rect 351 215 367 249
rect 301 249 367 255
rect 1131 85 1169 215
rect 1131 215 1149 249
rect 1131 249 1169 255
rect 1183 215 1199 249
rect 1075 215 1091 249
rect 587 215 603 249
rect 753 215 769 249
rect 29 199 63 215
rect 19 127 35 161
rect 203 51 249 67
rect 237 67 249 85
rect 247 85 249 101
rect 203 101 213 119
rect 247 101 249 119
rect 203 119 249 125
rect 1203 93 1237 109
rect 907 93 941 109
rect 1351 -17 1380 17
rect 761 59 823 93
rect 1045 59 1061 93
rect 857 59 873 93
rect 711 59 727 93
rect 307 51 341 67
rect 0 527 29 561
rect 403 485 437 527
rect 431 527 489 561
rect 339 527 397 561
rect 247 527 305 561
rect 907 435 1045 451
rect 941 451 1011 485
rect 907 485 1045 527
rect 891 527 949 561
rect 983 527 1041 561
rect 799 527 857 561
rect 707 527 765 561
rect 615 527 673 561
rect 523 527 581 561
rect 1203 485 1237 527
rect 1167 527 1225 561
rect 1075 527 1133 561
rect 487 357 489 391
rect 891 289 893 323
rect 487 85 489 119
rect 1259 -17 1317 17
rect 1167 -17 1225 17
rect 1203 17 1237 59
rect 1075 -17 1133 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 907 17 941 59
rect 799 -17 857 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 387 17 453 59
rect 387 59 403 93
rect 437 59 453 93
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 103 17 169 59
rect 103 59 119 93
rect 153 59 169 93
rect 0 -17 29 17
<< viali >>
rect 1317 527 1351 561
rect 1225 527 1259 561
rect 1133 527 1167 561
rect 1041 527 1075 561
rect 949 527 983 561
rect 857 527 891 561
rect 765 527 799 561
rect 673 527 707 561
rect 581 527 615 561
rect 489 527 523 561
rect 397 527 431 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 527 63 561
rect 213 357 247 391
rect 489 357 523 391
rect 673 289 707 323
rect 857 289 891 323
rect 1041 289 1075 323
rect 121 289 155 323
rect 489 85 523 119
rect 213 85 247 119
rect 857 -17 891 17
rect 1133 -17 1167 17
rect 673 -17 707 17
rect 949 -17 983 17
rect 581 -17 615 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 121 -17 155 17
rect 29 -17 63 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 1041 -17 1075 17
rect 765 -17 799 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 496 1380 527
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 561 1380 592
rect 201 351 259 357
rect 477 351 535 357
rect 201 357 213 360
rect 247 357 259 360
rect 477 357 489 360
rect 523 357 535 360
rect 201 360 213 388
rect 247 360 489 388
rect 523 360 535 388
rect 201 388 213 391
rect 247 388 259 391
rect 477 388 489 391
rect 523 388 535 391
rect 201 391 259 397
rect 477 391 535 397
rect 845 283 903 289
rect 1029 283 1087 289
rect 845 289 857 292
rect 891 289 903 292
rect 1029 289 1041 292
rect 1075 289 1087 292
rect 845 292 857 320
rect 891 292 1041 320
rect 1075 292 1087 320
rect 845 320 857 323
rect 891 320 903 323
rect 1029 320 1041 323
rect 1075 320 1087 323
rect 845 323 903 329
rect 1029 323 1087 329
rect 109 283 167 289
rect 661 283 719 289
rect 109 289 121 292
rect 155 289 167 292
rect 661 289 673 292
rect 707 289 719 292
rect 109 292 121 320
rect 155 292 673 320
rect 707 292 719 320
rect 109 320 121 323
rect 155 320 167 323
rect 661 320 673 323
rect 707 320 719 323
rect 109 323 167 329
rect 661 323 719 329
rect 201 79 259 85
rect 477 79 535 85
rect 201 85 213 88
rect 247 85 259 88
rect 477 85 489 88
rect 523 85 535 88
rect 201 88 213 116
rect 247 88 489 116
rect 523 88 535 116
rect 201 116 213 119
rect 247 116 259 119
rect 477 116 489 119
rect 523 116 535 119
rect 201 119 259 125
rect 477 119 535 125
rect 0 -48 1380 -17
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 17 1380 48
<< labels >>
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 GATE
port 5 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 GATE
port 5 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 D
port 6 nsew signal input
flabel locali s 1133 85 1167 119 0 FreeSans 200 0 0 0 RESET_B
port 7 nsew signal input
flabel locali s 1133 153 1167 187 0 FreeSans 200 0 0 0 RESET_B
port 7 nsew signal input
flabel locali s 1133 221 1167 255 0 FreeSans 200 0 0 0 RESET_B
port 7 nsew signal input
flabel locali s 1317 85 1351 119 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1317 357 1351 391 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1317 425 1351 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 -48 1380 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1380 592 1 VPWR
port 4 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 dlrtp_1
<< properties >>
string FIXED_BBOX 0 0 1380 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ht_sc_tt05.gds
string GDS_START 13210
string GDS_END 24074
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
