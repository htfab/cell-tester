magic
tech sky130A
magscale 1 2
timestamp 1699069426
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1931 203
rect 29 -17 63 21
<< scnmos >>
rect 1809 47 1839 177
rect 1065 47 1095 175
rect 1713 47 1743 131
rect 1629 47 1659 131
rect 793 47 823 131
rect 877 47 907 131
rect 353 47 383 131
rect 1425 47 1455 131
rect 81 47 111 131
rect 165 47 195 131
rect 1161 47 1191 119
rect 1245 47 1275 119
rect 545 47 575 119
rect 629 47 659 119
<< scpmoshvt >>
rect 81 369 111 497
rect 165 369 195 497
rect 353 413 383 497
rect 449 413 479 497
rect 545 413 575 497
rect 793 413 823 497
rect 877 413 907 497
rect 1629 413 1659 497
rect 1713 413 1743 497
rect 1809 297 1839 497
rect 1065 329 1095 497
rect 1245 413 1275 497
rect 1341 413 1371 497
rect 1425 413 1455 497
<< ndiff >>
rect 1743 47 1809 59
rect 1743 59 1765 93
rect 1799 59 1809 93
rect 1743 93 1809 131
rect 1758 131 1809 177
rect 1839 47 1891 59
rect 1839 59 1849 93
rect 1883 59 1891 93
rect 1839 93 1891 177
rect 1095 47 1161 67
rect 1095 67 1105 101
rect 1139 67 1161 101
rect 1095 101 1161 119
rect 1095 119 1146 175
rect 1013 47 1065 59
rect 1013 59 1021 93
rect 1055 59 1065 93
rect 1013 93 1065 175
rect 195 47 247 67
rect 195 67 205 101
rect 239 67 247 101
rect 195 101 247 131
rect 111 47 165 59
rect 111 59 121 93
rect 155 59 165 93
rect 111 93 165 131
rect 1455 47 1523 59
rect 1455 59 1481 93
rect 1515 59 1523 93
rect 1455 93 1523 131
rect 383 47 545 67
rect 383 67 405 101
rect 439 67 545 101
rect 383 101 545 119
rect 383 119 530 131
rect 907 47 959 59
rect 907 59 917 93
rect 951 59 959 93
rect 907 93 959 131
rect 823 47 877 131
rect 659 47 793 119
rect 674 119 793 131
rect 301 47 353 59
rect 301 59 309 93
rect 343 59 353 93
rect 301 93 353 131
rect 1275 47 1425 119
rect 1290 119 1425 131
rect 29 47 81 67
rect 29 67 37 101
rect 71 67 81 101
rect 29 101 81 131
rect 1577 47 1629 59
rect 1577 59 1585 93
rect 1619 59 1629 93
rect 1577 93 1629 131
rect 1659 47 1713 131
rect 1191 47 1245 59
rect 1191 59 1201 93
rect 1235 59 1245 93
rect 1191 93 1245 119
rect 575 47 629 59
rect 575 59 585 93
rect 619 59 629 93
rect 575 93 629 119
<< pdiff >>
rect 1371 413 1425 497
rect 1455 413 1523 451
rect 1455 451 1481 485
rect 1515 451 1523 485
rect 1455 485 1523 497
rect 1013 329 1065 443
rect 1013 443 1021 477
rect 1055 443 1065 477
rect 1013 477 1065 497
rect 1577 413 1629 451
rect 1577 451 1585 485
rect 1619 451 1629 485
rect 1577 485 1629 497
rect 301 413 353 443
rect 301 443 309 477
rect 343 443 353 477
rect 301 477 353 497
rect 29 369 81 383
rect 29 383 37 417
rect 71 383 81 417
rect 29 417 81 451
rect 29 451 37 485
rect 71 451 81 485
rect 29 485 81 497
rect 111 369 165 451
rect 111 451 121 485
rect 155 451 165 485
rect 111 485 165 497
rect 195 369 247 443
rect 195 443 205 477
rect 239 443 247 477
rect 195 477 247 497
rect 383 413 449 443
rect 383 443 405 477
rect 439 443 449 477
rect 383 477 449 497
rect 479 413 545 443
rect 479 443 501 477
rect 535 443 545 477
rect 479 477 545 497
rect 823 413 877 451
rect 823 451 833 485
rect 867 451 877 485
rect 823 485 877 497
rect 907 413 959 443
rect 907 443 917 477
rect 951 443 959 477
rect 907 477 959 497
rect 1659 413 1713 443
rect 1659 443 1669 477
rect 1703 443 1713 477
rect 1659 477 1713 497
rect 1758 297 1809 413
rect 1743 413 1809 451
rect 1743 451 1765 485
rect 1799 451 1809 485
rect 1743 485 1809 497
rect 1839 297 1891 451
rect 1839 451 1849 485
rect 1883 451 1891 485
rect 1839 485 1891 497
rect 1095 329 1230 413
rect 1095 413 1245 451
rect 1095 451 1117 485
rect 1151 451 1245 485
rect 1095 485 1245 497
rect 1275 413 1341 451
rect 1275 451 1297 485
rect 1331 451 1341 485
rect 1275 485 1341 497
rect 575 413 793 443
rect 575 443 749 477
rect 783 443 793 477
rect 575 477 793 497
<< ndiffc >>
rect 37 67 71 101
rect 205 67 239 101
rect 1105 67 1139 101
rect 405 67 439 101
rect 1481 59 1515 93
rect 121 59 155 93
rect 917 59 951 93
rect 1585 59 1619 93
rect 1021 59 1055 93
rect 309 59 343 93
rect 1765 59 1799 93
rect 1201 59 1235 93
rect 1849 59 1883 93
rect 585 59 619 93
<< pdiffc >>
rect 37 451 71 485
rect 121 451 155 485
rect 833 451 867 485
rect 1117 451 1151 485
rect 1297 451 1331 485
rect 1585 451 1619 485
rect 1765 451 1799 485
rect 1849 451 1883 485
rect 1481 451 1515 485
rect 309 443 343 477
rect 501 443 535 477
rect 1669 443 1703 477
rect 1021 443 1055 477
rect 405 443 439 477
rect 205 443 239 477
rect 749 443 783 477
rect 917 443 951 477
rect 37 383 71 417
<< poly >>
rect 1713 497 1743 523
rect 449 497 479 523
rect 1425 497 1455 523
rect 165 497 195 523
rect 793 497 823 523
rect 1245 497 1275 523
rect 1341 497 1371 523
rect 545 497 575 523
rect 877 497 907 523
rect 1629 497 1659 523
rect 81 497 111 523
rect 353 497 383 523
rect 1809 497 1839 523
rect 1065 497 1095 523
rect 1629 131 1659 199
rect 1521 199 1659 215
rect 1521 215 1531 249
rect 1565 215 1659 249
rect 1521 249 1659 265
rect 1629 265 1659 413
rect 1713 131 1743 199
rect 1701 199 1755 215
rect 1701 215 1711 249
rect 1745 215 1755 249
rect 1701 249 1755 265
rect 1713 265 1743 413
rect 1425 131 1455 199
rect 1425 199 1479 215
rect 1425 215 1435 249
rect 1469 215 1479 249
rect 1425 249 1479 265
rect 1425 265 1455 413
rect 1329 199 1383 215
rect 1329 215 1339 249
rect 1373 215 1383 249
rect 1329 249 1383 265
rect 1341 265 1371 413
rect 1245 119 1275 199
rect 1233 199 1287 215
rect 1233 215 1243 249
rect 1277 215 1287 249
rect 1233 249 1287 265
rect 1245 265 1275 413
rect 353 131 383 199
rect 297 199 383 215
rect 297 215 307 249
rect 341 215 383 249
rect 297 249 383 265
rect 353 265 383 413
rect 437 199 491 215
rect 437 215 447 249
rect 481 215 491 249
rect 437 249 491 265
rect 449 265 479 413
rect 545 119 575 199
rect 533 199 587 215
rect 533 215 543 249
rect 577 215 587 249
rect 533 249 587 265
rect 545 265 575 413
rect 793 131 823 199
rect 769 199 823 215
rect 769 215 779 249
rect 813 215 823 249
rect 769 249 823 265
rect 793 265 823 413
rect 877 131 907 199
rect 865 199 919 215
rect 865 215 875 249
rect 909 215 919 249
rect 865 249 919 265
rect 877 265 907 413
rect 81 131 111 199
rect 57 199 111 215
rect 57 215 67 249
rect 101 215 111 249
rect 57 249 111 265
rect 81 265 111 369
rect 165 131 195 199
rect 153 199 207 215
rect 153 215 163 249
rect 197 215 207 249
rect 153 249 207 265
rect 165 265 195 369
rect 1065 175 1095 199
rect 961 199 1095 215
rect 961 215 971 249
rect 1005 215 1095 249
rect 961 249 1095 265
rect 1065 265 1095 329
rect 1809 177 1839 199
rect 1797 199 1851 215
rect 1797 215 1807 249
rect 1841 215 1851 249
rect 1797 249 1851 265
rect 1809 265 1839 297
rect 1161 119 1191 199
rect 1137 199 1191 215
rect 1137 215 1147 249
rect 1181 215 1191 249
rect 1137 249 1191 265
rect 629 119 659 199
rect 629 199 683 215
rect 629 215 639 249
rect 673 215 683 249
rect 629 249 683 265
rect 81 21 111 47
rect 877 21 907 47
rect 793 21 823 47
rect 629 21 659 47
rect 545 21 575 47
rect 353 21 383 47
rect 1425 21 1455 47
rect 1245 21 1275 47
rect 1161 21 1191 47
rect 1065 21 1095 47
rect 1809 21 1839 47
rect 1713 21 1743 47
rect 1629 21 1659 47
rect 165 21 195 47
<< polycont >>
rect 1147 215 1181 249
rect 543 215 577 249
rect 163 215 197 249
rect 67 215 101 249
rect 639 215 673 249
rect 1711 215 1745 249
rect 307 215 341 249
rect 1435 215 1469 249
rect 1339 215 1373 249
rect 1531 215 1565 249
rect 1807 215 1841 249
rect 779 215 813 249
rect 1243 215 1277 249
rect 447 215 481 249
rect 875 215 909 249
rect 971 215 1005 249
<< locali >>
rect 121 485 155 527
rect 63 527 121 561
rect 155 527 213 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 749 477 783 493
rect 917 477 951 493
rect 205 477 239 493
rect 1669 477 1703 493
rect 405 477 439 493
rect 1105 101 1139 127
rect 1041 127 1139 161
rect 1041 161 1075 215
rect 813 215 815 249
rect 1041 215 1075 249
rect 779 249 815 265
rect 1041 249 1075 265
rect 781 265 815 299
rect 1041 265 1075 299
rect 781 299 1075 333
rect 1041 333 1075 357
rect 1041 357 1123 391
rect 1089 391 1123 451
rect 1089 451 1117 485
rect 1235 59 1415 93
rect 1381 93 1415 127
rect 1381 127 1547 161
rect 1513 161 1547 199
rect 1513 199 1565 215
rect 1513 215 1531 249
rect 1513 249 1565 265
rect 1513 265 1547 357
rect 1405 357 1547 391
rect 1405 391 1439 451
rect 1331 451 1439 485
rect 1883 59 1903 93
rect 1869 93 1903 127
rect 1869 127 1915 161
rect 1881 161 1915 315
rect 1869 315 1915 349
rect 1869 349 1903 451
rect 1883 451 1903 485
rect 1151 451 1167 485
rect 1833 451 1849 485
rect 1281 451 1297 485
rect 619 59 743 93
rect 709 93 743 127
rect 709 127 1003 161
rect 709 161 743 199
rect 969 161 1003 199
rect 709 199 743 215
rect 969 199 1005 215
rect 709 215 743 249
rect 969 215 971 249
rect 709 249 743 265
rect 971 249 1005 265
rect 709 265 743 299
rect 681 299 743 333
rect 681 333 715 443
rect 535 443 715 477
rect 485 443 501 477
rect 1765 435 1799 451
rect 121 435 155 451
rect 239 67 267 101
rect 233 101 267 357
rect 247 357 267 391
rect 309 427 343 443
rect 405 101 439 127
rect 377 127 439 161
rect 377 161 411 375
rect 377 375 439 409
rect 405 409 439 443
rect 1021 427 1055 443
rect 749 375 951 409
rect 749 409 783 443
rect 917 409 951 443
rect 1605 215 1711 221
rect 1605 221 1685 249
rect 1605 249 1639 299
rect 1593 299 1639 333
rect 1593 333 1627 391
rect 639 199 673 215
rect 481 215 483 249
rect 613 215 639 249
rect 447 249 483 265
rect 613 249 673 265
rect 449 265 483 299
rect 613 265 647 299
rect 449 299 647 333
rect 581 333 615 357
rect 1181 215 1191 249
rect 1147 249 1191 265
rect 1157 265 1191 357
rect 1157 357 1317 391
rect 29 215 67 249
rect 29 249 63 323
rect 1619 59 1719 93
rect 1685 93 1719 143
rect 1685 143 1831 177
rect 1797 177 1831 199
rect 1797 199 1841 215
rect 1797 215 1807 249
rect 1797 249 1841 265
rect 1797 265 1831 289
rect 1811 289 1831 323
rect 1797 323 1831 367
rect 1669 367 1831 401
rect 1669 401 1703 443
rect 63 101 71 119
rect 29 119 71 125
rect 37 125 71 143
rect 37 143 195 177
rect 161 177 195 199
rect 161 199 197 215
rect 161 215 163 249
rect 161 249 197 265
rect 161 265 195 289
rect 155 289 195 323
rect 121 323 155 367
rect 21 367 155 383
rect 21 383 37 401
rect 71 383 155 401
rect 21 401 37 417
rect 71 401 87 417
rect 21 417 87 451
rect 21 451 37 485
rect 71 451 87 485
rect 1435 199 1469 215
rect 1409 215 1435 249
rect 1409 249 1469 265
rect 1409 265 1443 289
rect 1243 199 1277 215
rect 1225 215 1243 249
rect 1225 249 1277 265
rect 1225 265 1259 289
rect 891 249 909 255
rect 875 255 909 265
rect 307 199 341 215
rect 305 215 307 249
rect 305 249 341 255
rect 307 255 341 265
rect 489 119 523 127
rect 489 127 575 161
rect 541 161 575 199
rect 541 199 577 215
rect 541 215 543 249
rect 543 249 577 265
rect 101 215 117 249
rect 1745 215 1761 249
rect 875 199 909 215
rect 779 199 813 215
rect 447 199 481 215
rect 1147 199 1181 215
rect 1765 93 1799 109
rect 309 93 343 109
rect 121 93 155 109
rect 189 67 205 101
rect 1185 59 1201 93
rect 1903 -17 1932 17
rect 1569 59 1585 93
rect 1833 59 1849 93
rect 569 59 585 93
rect 405 51 439 67
rect 1105 51 1139 67
rect 0 527 29 561
rect 1021 477 1055 527
rect 983 527 1041 561
rect 891 527 949 561
rect 1481 435 1619 451
rect 1515 451 1585 485
rect 1481 485 1619 527
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1351 527 1409 561
rect 1259 527 1317 561
rect 1167 527 1225 561
rect 1075 527 1133 561
rect 1765 485 1799 527
rect 1719 527 1777 561
rect 1627 527 1685 561
rect 309 477 343 527
rect 339 527 397 561
rect 247 527 305 561
rect 817 451 833 485
rect 867 451 883 485
rect 817 485 883 527
rect 799 527 857 561
rect 707 527 765 561
rect 615 527 673 561
rect 523 527 581 561
rect 431 527 489 561
rect 205 357 213 391
rect 205 391 239 443
rect 1339 199 1373 215
rect 1329 215 1339 249
rect 1329 249 1373 265
rect 1329 265 1363 357
rect 1351 357 1363 391
rect 29 51 71 67
rect 29 67 37 85
rect 1811 -17 1869 17
rect 1719 -17 1777 17
rect 1765 17 1799 59
rect 1627 -17 1685 17
rect 1535 -17 1593 17
rect 1443 -17 1501 17
rect 1465 17 1531 59
rect 1465 59 1481 93
rect 1515 59 1531 93
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 901 17 1071 59
rect 901 59 917 93
rect 951 59 1021 93
rect 1055 59 1071 93
rect 799 -17 857 17
rect 707 -17 765 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 309 17 343 59
rect 247 -17 305 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 121 17 155 59
rect 0 -17 29 17
<< viali >>
rect 1869 527 1903 561
rect 673 527 707 561
rect 29 527 63 561
rect 1041 527 1075 561
rect 1501 527 1535 561
rect 213 527 247 561
rect 1225 527 1259 561
rect 1777 527 1811 561
rect 1409 527 1443 561
rect 949 527 983 561
rect 581 527 615 561
rect 305 527 339 561
rect 857 527 891 561
rect 397 527 431 561
rect 1593 527 1627 561
rect 1133 527 1167 561
rect 1317 527 1351 561
rect 489 527 523 561
rect 1685 527 1719 561
rect 121 527 155 561
rect 765 527 799 561
rect 581 357 615 391
rect 1317 357 1351 391
rect 213 357 247 391
rect 1777 289 1811 323
rect 1409 289 1443 323
rect 1225 289 1259 323
rect 121 289 155 323
rect 857 221 891 255
rect 1685 221 1719 255
rect 489 85 523 119
rect 29 85 63 119
rect 1317 -17 1351 17
rect 1685 -17 1719 17
rect 857 -17 891 17
rect 489 -17 523 17
rect 397 -17 431 17
rect 305 -17 339 17
rect 121 -17 155 17
rect 949 -17 983 17
rect 1593 -17 1627 17
rect 29 -17 63 17
rect 213 -17 247 17
rect 673 -17 707 17
rect 1225 -17 1259 17
rect 1041 -17 1075 17
rect 581 -17 615 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1133 -17 1167 17
rect 765 -17 799 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 496 1932 527
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 561 1932 592
rect 201 351 259 357
rect 569 351 627 357
rect 1305 351 1363 357
rect 201 357 213 360
rect 247 357 259 360
rect 569 357 581 360
rect 615 357 627 360
rect 1305 357 1317 360
rect 1351 357 1363 360
rect 201 360 213 388
rect 247 360 581 388
rect 615 360 1317 388
rect 1351 360 1363 388
rect 201 388 213 391
rect 247 388 259 391
rect 569 388 581 391
rect 615 388 627 391
rect 1305 388 1317 391
rect 1351 388 1363 391
rect 201 391 259 397
rect 569 391 627 397
rect 1305 391 1363 397
rect 109 283 167 289
rect 1213 283 1271 289
rect 109 289 121 292
rect 155 289 167 292
rect 1213 289 1225 292
rect 1259 289 1271 292
rect 109 292 121 320
rect 155 292 1225 320
rect 1259 292 1271 320
rect 109 320 121 323
rect 155 320 167 323
rect 1213 320 1225 323
rect 1259 320 1271 323
rect 109 323 167 329
rect 1213 323 1271 329
rect 1397 283 1455 289
rect 1765 283 1823 289
rect 1397 289 1409 292
rect 1443 289 1455 292
rect 1765 289 1777 292
rect 1811 289 1823 292
rect 1397 292 1409 320
rect 1443 292 1777 320
rect 1811 292 1823 320
rect 1397 320 1409 323
rect 1443 320 1455 323
rect 1765 320 1777 323
rect 1811 320 1823 323
rect 1397 323 1455 329
rect 1765 323 1823 329
rect 845 215 903 221
rect 1673 215 1731 221
rect 845 221 857 224
rect 891 221 903 224
rect 1673 221 1685 224
rect 1719 221 1731 224
rect 845 224 857 252
rect 891 224 1685 252
rect 1719 224 1731 252
rect 845 252 857 255
rect 891 252 903 255
rect 1673 252 1685 255
rect 1719 252 1731 255
rect 845 255 903 261
rect 1673 255 1731 261
rect 17 79 75 85
rect 477 79 535 85
rect 17 85 29 88
rect 63 85 75 88
rect 477 85 489 88
rect 523 85 535 88
rect 17 88 29 116
rect 63 88 489 116
rect 523 88 535 116
rect 17 116 29 119
rect 63 116 75 119
rect 477 116 489 119
rect 523 116 535 119
rect 17 119 75 125
rect 477 119 535 125
rect 0 -48 1932 -17
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 17 1932 48
<< labels >>
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 CLK
port 1 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 1593 357 1627 391 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1869 85 1903 119 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1869 357 1903 391 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1869 425 1903 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 -48 1932 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 1 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 dfrtp_1
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ht_sc_tt05.gds
string GDS_START 23860
string GDS_END 37716
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
