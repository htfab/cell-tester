magic
tech sky130A
magscale 1 2
timestamp 1698685450
<< viali >>
rect 8033 21641 8067 21675
rect 13737 21641 13771 21675
rect 18889 21641 18923 21675
rect 23397 21641 23431 21675
rect 25697 21641 25731 21675
rect 27813 21641 27847 21675
rect 29653 21641 29687 21675
rect 22017 21573 22051 21607
rect 30389 21573 30423 21607
rect 1445 21487 1479 21521
rect 1685 21505 1719 21539
rect 3065 21505 3099 21539
rect 3712 21505 3746 21539
rect 6288 21505 6322 21539
rect 8728 21505 8762 21539
rect 8880 21487 8914 21521
rect 9137 21505 9171 21539
rect 11624 21505 11658 21539
rect 16313 21505 16347 21539
rect 17141 21505 17175 21539
rect 20821 21505 20855 21539
rect 22410 21505 22444 21539
rect 22569 21505 22603 21539
rect 23857 21505 23891 21539
rect 24501 21505 24535 21539
rect 24777 21505 24811 21539
rect 26433 21505 26467 21539
rect 949 21437 983 21471
rect 3249 21437 3283 21471
rect 3985 21437 4019 21471
rect 5641 21437 5675 21471
rect 5825 21437 5859 21471
rect 6561 21437 6595 21471
rect 8217 21437 8251 21471
rect 8401 21437 8435 21471
rect 10793 21437 10827 21471
rect 11161 21437 11195 21471
rect 11897 21437 11931 21471
rect 14289 21437 14323 21471
rect 14565 21437 14599 21471
rect 16129 21437 16163 21471
rect 16865 21437 16899 21471
rect 18797 21437 18831 21471
rect 19441 21437 19475 21471
rect 19717 21437 19751 21471
rect 21373 21437 21407 21471
rect 21557 21437 21591 21471
rect 22293 21437 22327 21471
rect 23581 21437 23615 21471
rect 24041 21437 24075 21471
rect 24894 21437 24928 21471
rect 25053 21437 25087 21471
rect 25789 21437 25823 21471
rect 26709 21437 26743 21471
rect 28273 21437 28307 21471
rect 29101 21437 29135 21471
rect 29285 21437 29319 21471
rect 29377 21437 29411 21471
rect 30573 21437 30607 21471
rect 5365 21369 5399 21403
rect 13645 21369 13679 21403
rect 15945 21369 15979 21403
rect 18521 21369 18555 21403
rect 26065 21369 26099 21403
rect 29929 21369 29963 21403
rect 1415 21301 1449 21335
rect 3715 21301 3749 21335
rect 5457 21301 5491 21335
rect 6291 21301 6325 21335
rect 7665 21301 7699 21335
rect 10241 21301 10275 21335
rect 10609 21301 10643 21335
rect 11627 21301 11661 21335
rect 13001 21301 13035 21335
rect 23213 21301 23247 21335
rect 28549 21301 28583 21335
rect 30021 21301 30055 21335
rect 1415 21097 1449 21131
rect 3623 21097 3657 21131
rect 6291 21097 6325 21131
rect 9965 21097 9999 21131
rect 14289 21097 14323 21131
rect 14749 21097 14783 21131
rect 15209 21097 15243 21131
rect 15669 21097 15703 21131
rect 17141 21097 17175 21131
rect 18613 21097 18647 21131
rect 20821 21097 20855 21131
rect 23121 21097 23155 21131
rect 25329 21097 25363 21131
rect 25697 21097 25731 21131
rect 5273 21029 5307 21063
rect 10425 21029 10459 21063
rect 26065 21029 26099 21063
rect 1685 20961 1719 20995
rect 5365 20961 5399 20995
rect 5825 20961 5859 20995
rect 11713 20961 11747 20995
rect 13277 20961 13311 20995
rect 16313 20961 16347 20995
rect 16681 20961 16715 20995
rect 17049 20961 17083 20995
rect 17509 20961 17543 20995
rect 21005 20961 21039 20995
rect 23305 20961 23339 20995
rect 25513 20961 25547 20995
rect 25881 20961 25915 20995
rect 26157 20961 26191 20995
rect 28692 20961 28726 20995
rect 949 20893 983 20927
rect 1455 20893 1489 20927
rect 3157 20893 3191 20927
rect 3620 20893 3654 20927
rect 3893 20893 3927 20927
rect 6288 20893 6322 20927
rect 6561 20893 6595 20927
rect 8125 20893 8159 20927
rect 8452 20893 8486 20927
rect 8631 20893 8665 20927
rect 8861 20893 8895 20927
rect 10977 20893 11011 20927
rect 11304 20893 11338 20927
rect 11440 20893 11474 20927
rect 17233 20893 17267 20927
rect 18981 20893 19015 20927
rect 19257 20893 19291 20927
rect 21281 20893 21315 20927
rect 21557 20893 21591 20927
rect 23489 20893 23523 20927
rect 23765 20893 23799 20927
rect 26433 20893 26467 20927
rect 26709 20893 26743 20927
rect 28365 20893 28399 20927
rect 28871 20893 28905 20927
rect 29101 20893 29135 20927
rect 2973 20757 3007 20791
rect 5549 20757 5583 20791
rect 7849 20757 7883 20791
rect 10517 20757 10551 20791
rect 12817 20757 12851 20791
rect 13369 20757 13403 20791
rect 27997 20757 28031 20791
rect 30205 20757 30239 20791
rect 2973 20553 3007 20587
rect 7941 20553 7975 20587
rect 16037 20553 16071 20587
rect 19073 20553 19107 20587
rect 30205 20553 30239 20587
rect 11069 20485 11103 20519
rect 1276 20417 1310 20451
rect 1445 20399 1479 20433
rect 1685 20417 1719 20451
rect 4399 20417 4433 20451
rect 6607 20417 6641 20451
rect 8999 20417 9033 20451
rect 11716 20417 11750 20451
rect 14105 20417 14139 20451
rect 16129 20417 16163 20451
rect 18705 20417 18739 20451
rect 19349 20417 19383 20451
rect 21833 20417 21867 20451
rect 24133 20417 24167 20451
rect 26709 20417 26743 20451
rect 27036 20417 27070 20451
rect 27215 20417 27249 20451
rect 949 20349 983 20383
rect 3341 20349 3375 20383
rect 3893 20349 3927 20383
rect 4629 20349 4663 20383
rect 6101 20349 6135 20383
rect 6428 20349 6462 20383
rect 6837 20349 6871 20383
rect 8493 20349 8527 20383
rect 9229 20349 9263 20383
rect 10793 20349 10827 20383
rect 11253 20349 11287 20383
rect 11989 20349 12023 20383
rect 14289 20349 14323 20383
rect 16405 20349 16439 20383
rect 17969 20349 18003 20383
rect 18889 20349 18923 20383
rect 21373 20349 21407 20383
rect 21557 20349 21591 20383
rect 23376 20349 23410 20383
rect 23581 20349 23615 20383
rect 23857 20349 23891 20383
rect 25881 20349 25915 20383
rect 27445 20349 27479 20383
rect 29469 20349 29503 20383
rect 29837 20349 29871 20383
rect 3709 20281 3743 20315
rect 10609 20281 10643 20315
rect 13829 20281 13863 20315
rect 14565 20281 14599 20315
rect 19625 20281 19659 20315
rect 26157 20281 26191 20315
rect 29101 20281 29135 20315
rect 30113 20281 30147 20315
rect 4359 20213 4393 20247
rect 5917 20213 5951 20247
rect 8959 20213 8993 20247
rect 11719 20213 11753 20247
rect 13093 20213 13127 20247
rect 17509 20213 17543 20247
rect 18061 20213 18095 20247
rect 21189 20213 21223 20247
rect 25697 20213 25731 20247
rect 26249 20213 26283 20247
rect 28549 20213 28583 20247
rect 29929 20213 29963 20247
rect 1415 20009 1449 20043
rect 2973 20009 3007 20043
rect 6291 20009 6325 20043
rect 21833 20009 21867 20043
rect 24041 20009 24075 20043
rect 27813 20009 27847 20043
rect 10609 19941 10643 19975
rect 19901 19941 19935 19975
rect 26065 19941 26099 19975
rect 3433 19873 3467 19907
rect 3852 19873 3886 19907
rect 5641 19873 5675 19907
rect 8125 19873 8159 19907
rect 10977 19873 11011 19907
rect 11529 19873 11563 19907
rect 11621 19873 11655 19907
rect 11713 19873 11747 19907
rect 14289 19873 14323 19907
rect 14565 19873 14599 19907
rect 16405 19873 16439 19907
rect 18153 19873 18187 19907
rect 21373 19873 21407 19907
rect 22017 19873 22051 19907
rect 22201 19873 22235 19907
rect 24225 19873 24259 19907
rect 24685 19873 24719 19907
rect 26422 19873 26456 19907
rect 26709 19873 26743 19907
rect 28365 19873 28399 19907
rect 949 19805 983 19839
rect 1445 19823 1479 19857
rect 1685 19805 1719 19839
rect 3525 19805 3559 19839
rect 4031 19805 4065 19839
rect 4261 19805 4295 19839
rect 5825 19805 5859 19839
rect 6288 19807 6322 19841
rect 6561 19805 6595 19839
rect 8493 19805 8527 19839
rect 8820 19805 8854 19839
rect 8956 19805 8990 19839
rect 9229 19805 9263 19839
rect 12081 19805 12115 19839
rect 12408 19805 12442 19839
rect 12587 19805 12621 19839
rect 12817 19805 12851 19839
rect 16129 19805 16163 19839
rect 17877 19805 17911 19839
rect 21005 19805 21039 19839
rect 22477 19805 22511 19839
rect 24409 19805 24443 19839
rect 28457 19805 28491 19839
rect 28784 19805 28818 19839
rect 28920 19805 28954 19839
rect 29193 19805 29227 19839
rect 7849 19737 7883 19771
rect 28181 19737 28215 19771
rect 3249 19669 3283 19703
rect 8309 19669 8343 19703
rect 11897 19669 11931 19703
rect 13921 19669 13955 19703
rect 15853 19669 15887 19703
rect 17693 19669 17727 19703
rect 19257 19669 19291 19703
rect 21465 19669 21499 19703
rect 30297 19669 30331 19703
rect 2789 19465 2823 19499
rect 4629 19465 4663 19499
rect 10241 19465 10275 19499
rect 14013 19465 14047 19499
rect 22017 19465 22051 19499
rect 22569 19397 22603 19431
rect 1455 19329 1489 19363
rect 3893 19329 3927 19363
rect 5828 19329 5862 19363
rect 8864 19329 8898 19363
rect 11256 19329 11290 19363
rect 14197 19329 14231 19363
rect 14473 19329 14507 19363
rect 16221 19329 16255 19363
rect 18153 19329 18187 19363
rect 18705 19329 18739 19363
rect 23581 19329 23615 19363
rect 26709 19329 26743 19363
rect 27215 19329 27249 19363
rect 29009 19329 29043 19363
rect 949 19261 983 19295
rect 1685 19261 1719 19295
rect 3617 19261 3651 19295
rect 3709 19261 3743 19295
rect 4353 19261 4387 19295
rect 5273 19261 5307 19295
rect 5365 19261 5399 19295
rect 6101 19261 6135 19295
rect 7757 19261 7791 19295
rect 8401 19261 8435 19295
rect 9137 19261 9171 19295
rect 10793 19261 10827 19295
rect 11529 19261 11563 19295
rect 13185 19261 13219 19295
rect 15945 19261 15979 19295
rect 17877 19261 17911 19295
rect 18061 19261 18095 19295
rect 18981 19261 19015 19295
rect 20453 19261 20487 19295
rect 20729 19261 20763 19295
rect 23305 19261 23339 19295
rect 23397 19261 23431 19295
rect 27036 19261 27070 19295
rect 27445 19261 27479 19295
rect 29285 19261 29319 19295
rect 4905 19193 4939 19227
rect 8033 19193 8067 19227
rect 13737 19193 13771 19227
rect 17601 19193 17635 19227
rect 22293 19193 22327 19227
rect 24133 19193 24167 19227
rect 30297 19193 30331 19227
rect 1415 19125 1449 19159
rect 3433 19125 3467 19159
rect 5831 19125 5865 19159
rect 7205 19125 7239 19159
rect 8867 19125 8901 19159
rect 11259 19125 11293 19159
rect 12633 19125 12667 19159
rect 13001 19125 13035 19159
rect 15761 19125 15795 19159
rect 18337 19125 18371 19159
rect 20085 19125 20119 19159
rect 22937 19125 22971 19159
rect 24409 19125 24443 19159
rect 24961 19125 24995 19159
rect 25421 19125 25455 19159
rect 25881 19125 25915 19159
rect 26341 19125 26375 19159
rect 28549 19125 28583 19159
rect 29929 19125 29963 19159
rect 30113 19125 30147 19159
rect 30389 19125 30423 19159
rect 3157 18921 3191 18955
rect 8493 18921 8527 18955
rect 12363 18921 12397 18955
rect 13921 18921 13955 18955
rect 17693 18921 17727 18955
rect 22661 18921 22695 18955
rect 23305 18921 23339 18955
rect 23765 18921 23799 18955
rect 28923 18921 28957 18955
rect 30297 18921 30331 18955
rect 4169 18853 4203 18887
rect 4721 18853 4755 18887
rect 5089 18853 5123 18887
rect 5273 18853 5307 18887
rect 8125 18853 8159 18887
rect 10793 18853 10827 18887
rect 1225 18785 1259 18819
rect 1317 18785 1351 18819
rect 3893 18785 3927 18819
rect 6009 18785 6043 18819
rect 6336 18785 6370 18819
rect 8401 18785 8435 18819
rect 9004 18785 9038 18819
rect 10977 18785 11011 18819
rect 11529 18785 11563 18819
rect 11897 18785 11931 18819
rect 12633 18785 12667 18819
rect 14565 18785 14599 18819
rect 16405 18785 16439 18819
rect 17877 18785 17911 18819
rect 18153 18785 18187 18819
rect 19901 18785 19935 18819
rect 20269 18785 20303 18819
rect 20545 18785 20579 18819
rect 23029 18785 23063 18819
rect 23673 18785 23707 18819
rect 24460 18785 24494 18819
rect 26617 18785 26651 18819
rect 28457 18785 28491 18819
rect 1644 18717 1678 18751
rect 1823 18719 1857 18753
rect 2053 18717 2087 18751
rect 6472 18717 6506 18751
rect 6745 18717 6779 18751
rect 8677 18717 8711 18751
rect 9183 18717 9217 18751
rect 9413 18717 9447 18751
rect 11161 18717 11195 18751
rect 12403 18719 12437 18753
rect 14289 18717 14323 18751
rect 16129 18717 16163 18751
rect 19993 18717 20027 18751
rect 21281 18717 21315 18751
rect 21557 18717 21591 18751
rect 24133 18717 24167 18751
rect 24639 18717 24673 18751
rect 24869 18717 24903 18751
rect 26893 18717 26927 18751
rect 28920 18717 28954 18751
rect 29193 18717 29227 18751
rect 11713 18649 11747 18683
rect 1041 18581 1075 18615
rect 3801 18581 3835 18615
rect 5549 18581 5583 18615
rect 15853 18581 15887 18615
rect 19257 18581 19291 18615
rect 20637 18581 20671 18615
rect 25973 18581 26007 18615
rect 28365 18581 28399 18615
rect 2973 18377 3007 18411
rect 5917 18377 5951 18411
rect 10609 18377 10643 18411
rect 13093 18377 13127 18411
rect 14105 18377 14139 18411
rect 20269 18377 20303 18411
rect 23581 18377 23615 18411
rect 23857 18377 23891 18411
rect 3525 18309 3559 18343
rect 16313 18309 16347 18343
rect 22845 18309 22879 18343
rect 24593 18309 24627 18343
rect 949 18241 983 18275
rect 1445 18223 1479 18257
rect 1685 18241 1719 18275
rect 4399 18241 4433 18275
rect 6564 18241 6598 18275
rect 9048 18241 9082 18275
rect 11759 18241 11793 18275
rect 14936 18239 14970 18273
rect 17141 18241 17175 18275
rect 18705 18241 18739 18275
rect 18981 18241 19015 18275
rect 21143 18241 21177 18275
rect 21373 18241 21407 18275
rect 25375 18241 25409 18275
rect 29009 18241 29043 18275
rect 3341 18173 3375 18207
rect 3893 18173 3927 18207
rect 4629 18173 4663 18207
rect 6101 18173 6135 18207
rect 6837 18173 6871 18207
rect 8585 18173 8619 18207
rect 9321 18173 9355 18207
rect 10977 18173 11011 18207
rect 11253 18173 11287 18207
rect 11989 18173 12023 18207
rect 14013 18173 14047 18207
rect 14473 18173 14507 18207
rect 15209 18173 15243 18207
rect 16865 18173 16899 18207
rect 20637 18173 20671 18207
rect 23029 18173 23063 18207
rect 23305 18173 23339 18207
rect 24041 18173 24075 18207
rect 24869 18173 24903 18207
rect 25605 18173 25639 18207
rect 27077 18173 27111 18207
rect 27353 18173 27387 18207
rect 29285 18173 29319 18207
rect 30573 18173 30607 18207
rect 8217 18105 8251 18139
rect 11161 18105 11195 18139
rect 13645 18105 13679 18139
rect 24409 18105 24443 18139
rect 1415 18037 1449 18071
rect 4359 18037 4393 18071
rect 6567 18037 6601 18071
rect 9051 18037 9085 18071
rect 11719 18037 11753 18071
rect 13737 18037 13771 18071
rect 14939 18037 14973 18071
rect 18429 18037 18463 18071
rect 21103 18037 21137 18071
rect 22477 18037 22511 18071
rect 25335 18037 25369 18071
rect 26709 18037 26743 18071
rect 28457 18037 28491 18071
rect 30113 18037 30147 18071
rect 30297 18037 30331 18071
rect 30389 18037 30423 18071
rect 1041 17833 1075 17867
rect 3157 17833 3191 17867
rect 3991 17833 4025 17867
rect 6935 17833 6969 17867
rect 14295 17833 14329 17867
rect 15669 17833 15703 17867
rect 17049 17833 17083 17867
rect 25973 17833 26007 17867
rect 27813 17833 27847 17867
rect 28831 17833 28865 17867
rect 30205 17833 30239 17867
rect 5641 17765 5675 17799
rect 10793 17765 10827 17799
rect 16221 17765 16255 17799
rect 1225 17697 1259 17731
rect 1317 17697 1351 17731
rect 1644 17697 1678 17731
rect 5917 17697 5951 17731
rect 8585 17697 8619 17731
rect 11161 17697 11195 17731
rect 11580 17697 11614 17731
rect 13461 17697 13495 17731
rect 16589 17697 16623 17731
rect 16957 17697 16991 17731
rect 19717 17697 19751 17731
rect 21097 17697 21131 17731
rect 23673 17697 23707 17731
rect 24041 17697 24075 17731
rect 26709 17697 26743 17731
rect 1813 17647 1847 17681
rect 2053 17629 2087 17663
rect 3525 17629 3559 17663
rect 4031 17629 4065 17663
rect 4261 17629 4295 17663
rect 6469 17629 6503 17663
rect 6932 17629 6966 17663
rect 7205 17629 7239 17663
rect 8677 17629 8711 17663
rect 9004 17629 9038 17663
rect 9140 17631 9174 17665
rect 9413 17629 9447 17663
rect 11253 17629 11287 17663
rect 11759 17631 11793 17665
rect 11989 17629 12023 17663
rect 13829 17629 13863 17663
rect 14335 17629 14369 17663
rect 14565 17629 14599 17663
rect 17141 17629 17175 17663
rect 17468 17629 17502 17663
rect 17647 17629 17681 17663
rect 17877 17629 17911 17663
rect 19441 17629 19475 17663
rect 21281 17629 21315 17663
rect 21608 17629 21642 17663
rect 21787 17629 21821 17663
rect 22017 17629 22051 17663
rect 24133 17629 24167 17663
rect 24460 17629 24494 17663
rect 24596 17631 24630 17665
rect 24869 17629 24903 17663
rect 26433 17629 26467 17663
rect 28365 17629 28399 17663
rect 28871 17629 28905 17663
rect 29101 17629 29135 17663
rect 23489 17561 23523 17595
rect 6193 17493 6227 17527
rect 10977 17493 11011 17527
rect 13093 17493 13127 17527
rect 13645 17493 13679 17527
rect 18981 17493 19015 17527
rect 23121 17493 23155 17527
rect 23857 17493 23891 17527
rect 2789 17289 2823 17323
rect 5917 17289 5951 17323
rect 8125 17289 8159 17323
rect 10517 17289 10551 17323
rect 13737 17289 13771 17323
rect 15577 17289 15611 17323
rect 18245 17289 18279 17323
rect 20269 17289 20303 17323
rect 14105 17221 14139 17255
rect 15945 17221 15979 17255
rect 23397 17221 23431 17255
rect 26709 17221 26743 17255
rect 949 17153 983 17187
rect 1455 17153 1489 17187
rect 3893 17153 3927 17187
rect 4399 17153 4433 17187
rect 6101 17153 6135 17187
rect 6564 17153 6598 17187
rect 6837 17153 6871 17187
rect 8677 17153 8711 17187
rect 9004 17153 9038 17187
rect 9183 17151 9217 17185
rect 9413 17153 9447 17187
rect 11759 17151 11793 17185
rect 16911 17153 16945 17187
rect 18981 17153 19015 17187
rect 21143 17153 21177 17187
rect 21373 17153 21407 17187
rect 24593 17153 24627 17187
rect 25196 17153 25230 17187
rect 25332 17153 25366 17187
rect 25605 17153 25639 17187
rect 27353 17153 27387 17187
rect 1685 17085 1719 17119
rect 3249 17085 3283 17119
rect 4629 17085 4663 17119
rect 8585 17085 8619 17119
rect 10977 17085 11011 17119
rect 11253 17085 11287 17119
rect 11989 17085 12023 17119
rect 13645 17085 13679 17119
rect 14289 17085 14323 17119
rect 14473 17085 14507 17119
rect 14749 17085 14783 17119
rect 15853 17085 15887 17119
rect 16129 17085 16163 17119
rect 16405 17085 16439 17119
rect 17141 17085 17175 17119
rect 18705 17085 18739 17119
rect 20637 17085 20671 17119
rect 23581 17085 23615 17119
rect 24041 17085 24075 17119
rect 24317 17085 24351 17119
rect 24869 17085 24903 17119
rect 27077 17085 27111 17119
rect 29561 17085 29595 17119
rect 29837 17085 29871 17119
rect 30113 17085 30147 17119
rect 3525 17017 3559 17051
rect 11161 17017 11195 17051
rect 22937 17017 22971 17051
rect 28733 17017 28767 17051
rect 29101 17017 29135 17051
rect 1415 16949 1449 16983
rect 4359 16949 4393 16983
rect 6567 16949 6601 16983
rect 8401 16949 8435 16983
rect 11719 16949 11753 16983
rect 13093 16949 13127 16983
rect 15393 16949 15427 16983
rect 15669 16949 15703 16983
rect 16871 16949 16905 16983
rect 21103 16949 21137 16983
rect 22477 16949 22511 16983
rect 23213 16949 23247 16983
rect 23857 16949 23891 16983
rect 29929 16949 29963 16983
rect 30389 16949 30423 16983
rect 949 16745 983 16779
rect 3065 16745 3099 16779
rect 7665 16745 7699 16779
rect 8033 16745 8067 16779
rect 11897 16745 11931 16779
rect 13461 16745 13495 16779
rect 15669 16745 15703 16779
rect 16313 16745 16347 16779
rect 16681 16745 16715 16779
rect 18981 16745 19015 16779
rect 23121 16745 23155 16779
rect 23955 16745 23989 16779
rect 28273 16745 28307 16779
rect 30389 16745 30423 16779
rect 5641 16677 5675 16711
rect 11161 16677 11195 16711
rect 21097 16677 21131 16711
rect 30297 16677 30331 16711
rect 1133 16609 1167 16643
rect 4261 16609 4295 16643
rect 6152 16609 6186 16643
rect 6561 16609 6595 16643
rect 8217 16609 8251 16643
rect 8493 16609 8527 16643
rect 8585 16609 8619 16643
rect 9321 16609 9355 16643
rect 12081 16609 12115 16643
rect 12357 16609 12391 16643
rect 13185 16609 13219 16643
rect 13645 16609 13679 16643
rect 14565 16609 14599 16643
rect 16221 16609 16255 16643
rect 16865 16609 16899 16643
rect 17141 16609 17175 16643
rect 19717 16609 19751 16643
rect 22017 16609 22051 16643
rect 24225 16609 24259 16643
rect 25789 16609 25823 16643
rect 26760 16609 26794 16643
rect 28917 16609 28951 16643
rect 30573 16609 30607 16643
rect 1225 16541 1259 16575
rect 1552 16541 1586 16575
rect 1721 16559 1755 16593
rect 1961 16541 1995 16575
rect 3525 16541 3559 16575
rect 3852 16541 3886 16575
rect 3988 16541 4022 16575
rect 5825 16541 5859 16575
rect 6331 16543 6365 16577
rect 8912 16541 8946 16575
rect 9091 16543 9125 16577
rect 11437 16541 11471 16575
rect 13837 16541 13871 16575
rect 14156 16541 14190 16575
rect 14335 16541 14369 16575
rect 17468 16541 17502 16575
rect 17637 16559 17671 16593
rect 17877 16541 17911 16575
rect 19441 16541 19475 16575
rect 21281 16541 21315 16575
rect 21608 16541 21642 16575
rect 21777 16559 21811 16593
rect 23489 16541 23523 16575
rect 23968 16543 24002 16577
rect 26433 16541 26467 16575
rect 26896 16543 26930 16577
rect 27169 16541 27203 16575
rect 28641 16541 28675 16575
rect 25973 16473 26007 16507
rect 8309 16405 8343 16439
rect 10425 16405 10459 16439
rect 13369 16405 13403 16439
rect 25329 16405 25363 16439
rect 2789 16201 2823 16235
rect 7941 16201 7975 16235
rect 13093 16201 13127 16235
rect 14105 16201 14139 16235
rect 14473 16201 14507 16235
rect 17509 16201 17543 16235
rect 17785 16201 17819 16235
rect 18429 16201 18463 16235
rect 5825 16133 5859 16167
rect 17233 16133 17267 16167
rect 25697 16133 25731 16167
rect 30389 16133 30423 16167
rect 1455 16065 1489 16099
rect 4307 16065 4341 16099
rect 6428 16065 6462 16099
rect 6607 16063 6641 16097
rect 9081 16047 9115 16081
rect 9321 16065 9355 16099
rect 11580 16065 11614 16099
rect 11759 16065 11793 16099
rect 14749 16065 14783 16099
rect 15255 16065 15289 16099
rect 19211 16065 19245 16099
rect 20821 16065 20855 16099
rect 22063 16065 22097 16099
rect 24184 16065 24218 16099
rect 24320 16063 24354 16097
rect 24593 16065 24627 16099
rect 26065 16065 26099 16099
rect 26528 16065 26562 16099
rect 26801 16065 26835 16099
rect 949 15997 983 16031
rect 1685 15997 1719 16031
rect 3341 15997 3375 16031
rect 3801 15997 3835 16031
rect 4537 15997 4571 16031
rect 6101 15997 6135 16031
rect 6837 15997 6871 16031
rect 8585 15997 8619 16031
rect 8912 15997 8946 16031
rect 11161 15997 11195 16031
rect 11253 15997 11287 16031
rect 11989 15997 12023 16031
rect 14289 15997 14323 16031
rect 14657 15997 14691 16031
rect 15485 15997 15519 16031
rect 16957 15997 16991 16031
rect 17417 15997 17451 16031
rect 17693 15997 17727 16031
rect 17969 15997 18003 16031
rect 18705 15997 18739 16031
rect 19441 15997 19475 16031
rect 20913 15997 20947 16031
rect 21557 15997 21591 16031
rect 22293 15997 22327 16031
rect 23857 15997 23891 16031
rect 28733 15997 28767 16031
rect 29101 15997 29135 16031
rect 29193 15997 29227 16031
rect 29377 15997 29411 16031
rect 29847 15997 29881 16031
rect 30573 15997 30607 16031
rect 13645 15929 13679 15963
rect 18153 15929 18187 15963
rect 21189 15929 21223 15963
rect 23673 15929 23707 15963
rect 28365 15929 28399 15963
rect 30113 15929 30147 15963
rect 1415 15861 1449 15895
rect 3617 15861 3651 15895
rect 4267 15861 4301 15895
rect 10425 15861 10459 15895
rect 10977 15861 11011 15895
rect 13737 15861 13771 15895
rect 15215 15861 15249 15895
rect 16589 15861 16623 15895
rect 17141 15861 17175 15895
rect 19171 15861 19205 15895
rect 22023 15861 22057 15895
rect 26531 15861 26565 15895
rect 27905 15861 27939 15895
rect 29653 15861 29687 15895
rect 3157 15657 3191 15691
rect 5549 15657 5583 15691
rect 12087 15657 12121 15691
rect 13461 15657 13495 15691
rect 17141 15657 17175 15691
rect 21005 15657 21039 15691
rect 23955 15657 23989 15691
rect 28273 15657 28307 15691
rect 30389 15657 30423 15691
rect 15945 15589 15979 15623
rect 26249 15589 26283 15623
rect 1225 15521 1259 15555
rect 4261 15521 4295 15555
rect 5917 15521 5951 15555
rect 6704 15521 6738 15555
rect 11069 15521 11103 15555
rect 14156 15521 14190 15555
rect 16129 15521 16163 15555
rect 16681 15521 16715 15555
rect 16957 15521 16991 15555
rect 17560 15521 17594 15555
rect 19717 15521 19751 15555
rect 25881 15521 25915 15555
rect 26433 15521 26467 15555
rect 26760 15521 26794 15555
rect 27169 15521 27203 15555
rect 28917 15521 28951 15555
rect 30573 15521 30607 15555
rect 1317 15453 1351 15487
rect 1644 15453 1678 15487
rect 1813 15471 1847 15505
rect 2053 15453 2087 15487
rect 3525 15453 3559 15487
rect 3852 15453 3886 15487
rect 3988 15455 4022 15489
rect 6377 15453 6411 15487
rect 6840 15471 6874 15505
rect 7113 15453 7147 15487
rect 8585 15453 8619 15487
rect 8912 15453 8946 15487
rect 9081 15471 9115 15505
rect 9321 15453 9355 15487
rect 11621 15453 11655 15487
rect 12127 15453 12161 15487
rect 12357 15453 12391 15487
rect 13829 15453 13863 15487
rect 14335 15453 14369 15487
rect 14565 15453 14599 15487
rect 16405 15453 16439 15487
rect 17233 15453 17267 15487
rect 17739 15453 17773 15487
rect 17969 15453 18003 15487
rect 19441 15453 19475 15487
rect 21281 15453 21315 15487
rect 21608 15453 21642 15487
rect 21787 15453 21821 15487
rect 21971 15453 22005 15487
rect 23489 15453 23523 15487
rect 23952 15455 23986 15489
rect 24225 15453 24259 15487
rect 26896 15453 26930 15487
rect 28641 15453 28675 15487
rect 11253 15385 11287 15419
rect 16865 15385 16899 15419
rect 1041 15317 1075 15351
rect 6193 15317 6227 15351
rect 8217 15317 8251 15351
rect 10425 15317 10459 15351
rect 16313 15317 16347 15351
rect 19073 15317 19107 15351
rect 23121 15317 23155 15351
rect 25329 15317 25363 15351
rect 30021 15317 30055 15351
rect 2789 15113 2823 15147
rect 5825 15113 5859 15147
rect 7941 15113 7975 15147
rect 16037 15113 16071 15147
rect 19257 15113 19291 15147
rect 19533 15113 19567 15147
rect 22201 15113 22235 15147
rect 23029 15113 23063 15147
rect 27905 15113 27939 15147
rect 10425 15045 10459 15079
rect 10977 15045 11011 15079
rect 18245 15045 18279 15079
rect 22477 15045 22511 15079
rect 29745 15045 29779 15079
rect 949 14977 983 15011
rect 1455 14977 1489 15011
rect 3801 14977 3835 15011
rect 4307 14977 4341 15011
rect 6607 14977 6641 15011
rect 8585 14977 8619 15011
rect 9081 14959 9115 14993
rect 11580 14977 11614 15011
rect 11759 14977 11793 15011
rect 11989 14977 12023 15011
rect 14703 14977 14737 15011
rect 16405 14977 16439 15011
rect 16911 14977 16945 15011
rect 19901 14977 19935 15011
rect 20407 14977 20441 15011
rect 20637 14977 20671 15011
rect 24184 14977 24218 15011
rect 24353 14977 24387 15011
rect 26528 14977 26562 15011
rect 29377 14977 29411 15011
rect 1685 14909 1719 14943
rect 3249 14909 3283 14943
rect 4128 14909 4162 14943
rect 4537 14909 4571 14943
rect 6101 14909 6135 14943
rect 6837 14909 6871 14943
rect 9321 14909 9355 14943
rect 11161 14909 11195 14943
rect 11253 14909 11287 14943
rect 13645 14909 13679 14943
rect 14197 14909 14231 14943
rect 14933 14909 14967 14943
rect 17141 14909 17175 14943
rect 18705 14909 18739 14943
rect 19441 14909 19475 14943
rect 19717 14909 19751 14943
rect 22385 14909 22419 14943
rect 22661 14909 22695 14943
rect 22937 14909 22971 14943
rect 23213 14909 23247 14943
rect 23673 14909 23707 14943
rect 23857 14909 23891 14943
rect 24593 14909 24627 14943
rect 26065 14909 26099 14943
rect 26801 14909 26835 14943
rect 28733 14909 28767 14943
rect 29561 14909 29595 14943
rect 3525 14841 3559 14875
rect 18981 14841 19015 14875
rect 28365 14841 28399 14875
rect 29101 14841 29135 14875
rect 30205 14841 30239 14875
rect 1415 14773 1449 14807
rect 6567 14773 6601 14807
rect 9051 14773 9085 14807
rect 13093 14773 13127 14807
rect 13921 14773 13955 14807
rect 14663 14773 14697 14807
rect 16871 14773 16905 14807
rect 20367 14773 20401 14807
rect 21741 14773 21775 14807
rect 22753 14773 22787 14807
rect 23489 14773 23523 14807
rect 25697 14773 25731 14807
rect 26531 14773 26565 14807
rect 30481 14773 30515 14807
rect 3985 14569 4019 14603
rect 4445 14569 4479 14603
rect 4721 14569 4755 14603
rect 4997 14569 5031 14603
rect 5457 14569 5491 14603
rect 6101 14569 6135 14603
rect 6377 14569 6411 14603
rect 9413 14569 9447 14603
rect 9689 14569 9723 14603
rect 9965 14569 9999 14603
rect 10333 14569 10367 14603
rect 13461 14569 13495 14603
rect 14295 14569 14329 14603
rect 16865 14569 16899 14603
rect 20085 14569 20119 14603
rect 20269 14569 20303 14603
rect 23765 14569 23799 14603
rect 24507 14569 24541 14603
rect 26065 14569 26099 14603
rect 28555 14569 28589 14603
rect 29929 14569 29963 14603
rect 11345 14501 11379 14535
rect 26893 14501 26927 14535
rect 27537 14501 27571 14535
rect 1133 14433 1167 14467
rect 1409 14433 1443 14467
rect 1501 14433 1535 14467
rect 3893 14433 3927 14467
rect 4169 14433 4203 14467
rect 4629 14433 4663 14467
rect 4905 14433 4939 14467
rect 5181 14433 5215 14467
rect 5641 14433 5675 14467
rect 6009 14433 6043 14467
rect 6285 14433 6319 14467
rect 6561 14433 6595 14467
rect 6653 14433 6687 14467
rect 8861 14433 8895 14467
rect 9137 14433 9171 14467
rect 9597 14433 9631 14467
rect 9873 14433 9907 14467
rect 10149 14433 10183 14467
rect 10517 14433 10551 14467
rect 10793 14433 10827 14467
rect 11069 14433 11103 14467
rect 11621 14433 11655 14467
rect 11948 14433 11982 14467
rect 15945 14433 15979 14467
rect 16221 14433 16255 14467
rect 16681 14433 16715 14467
rect 17468 14433 17502 14467
rect 19533 14433 19567 14467
rect 19809 14433 19843 14467
rect 20453 14433 20487 14467
rect 20737 14433 20771 14467
rect 21097 14433 21131 14467
rect 22017 14433 22051 14467
rect 23673 14433 23707 14467
rect 23949 14433 23983 14467
rect 24777 14433 24811 14467
rect 26617 14433 26651 14467
rect 27353 14433 27387 14467
rect 28089 14433 28123 14467
rect 30297 14433 30331 14467
rect 1828 14365 1862 14399
rect 2007 14367 2041 14401
rect 2237 14365 2271 14399
rect 3617 14365 3651 14399
rect 6980 14365 7014 14399
rect 7159 14365 7193 14399
rect 7389 14365 7423 14399
rect 12117 14367 12151 14401
rect 12311 14365 12345 14399
rect 13829 14365 13863 14399
rect 14335 14365 14369 14399
rect 14565 14365 14599 14399
rect 17141 14365 17175 14399
rect 17647 14365 17681 14399
rect 17877 14365 17911 14399
rect 21281 14365 21315 14399
rect 21608 14365 21642 14399
rect 21787 14365 21821 14399
rect 24041 14365 24075 14399
rect 24504 14365 24538 14399
rect 28595 14365 28629 14399
rect 28825 14365 28859 14399
rect 949 14297 983 14331
rect 18981 14297 19015 14331
rect 19349 14297 19383 14331
rect 20545 14297 20579 14331
rect 27813 14297 27847 14331
rect 1225 14229 1259 14263
rect 3709 14229 3743 14263
rect 5825 14229 5859 14263
rect 8677 14229 8711 14263
rect 10609 14229 10643 14263
rect 16497 14229 16531 14263
rect 19625 14229 19659 14263
rect 20913 14229 20947 14263
rect 23305 14229 23339 14263
rect 23489 14229 23523 14263
rect 27169 14229 27203 14263
rect 30481 14229 30515 14263
rect 7941 14025 7975 14059
rect 13093 14025 13127 14059
rect 13645 14025 13679 14059
rect 18245 14025 18279 14059
rect 23581 14025 23615 14059
rect 26065 14025 26099 14059
rect 28549 14025 28583 14059
rect 30113 14025 30147 14059
rect 10885 13957 10919 13991
rect 13921 13957 13955 13991
rect 16037 13957 16071 13991
rect 18705 13957 18739 13991
rect 18981 13957 19015 13991
rect 21649 13957 21683 13991
rect 26617 13957 26651 13991
rect 29285 13957 29319 13991
rect 30297 13957 30331 13991
rect 949 13889 983 13923
rect 1276 13889 1310 13923
rect 1445 13871 1479 13905
rect 4264 13889 4298 13923
rect 6607 13889 6641 13923
rect 8864 13889 8898 13923
rect 10517 13889 10551 13923
rect 11580 13889 11614 13923
rect 11759 13889 11793 13923
rect 14703 13889 14737 13923
rect 16405 13889 16439 13923
rect 16732 13889 16766 13923
rect 16911 13889 16945 13923
rect 17141 13889 17175 13923
rect 19441 13889 19475 13923
rect 20315 13889 20349 13923
rect 22293 13889 22327 13923
rect 24041 13889 24075 13923
rect 24368 13889 24402 13923
rect 24547 13887 24581 13921
rect 24777 13889 24811 13923
rect 26709 13889 26743 13923
rect 27215 13889 27249 13923
rect 27445 13889 27479 13923
rect 1685 13821 1719 13855
rect 3065 13821 3099 13855
rect 3433 13821 3467 13855
rect 3709 13821 3743 13855
rect 3801 13821 3835 13855
rect 4537 13821 4571 13855
rect 5917 13821 5951 13855
rect 6101 13821 6135 13855
rect 6837 13821 6871 13855
rect 8401 13821 8435 13855
rect 9137 13821 9171 13855
rect 11069 13821 11103 13855
rect 11253 13821 11287 13855
rect 11989 13821 12023 13855
rect 13829 13821 13863 13855
rect 14105 13821 14139 13855
rect 14197 13821 14231 13855
rect 14933 13821 14967 13855
rect 18889 13821 18923 13855
rect 19165 13821 19199 13855
rect 19809 13821 19843 13855
rect 20545 13821 20579 13855
rect 22017 13821 22051 13855
rect 26433 13821 26467 13855
rect 27036 13821 27070 13855
rect 29101 13821 29135 13855
rect 29837 13821 29871 13855
rect 30481 13821 30515 13855
rect 10609 13753 10643 13787
rect 29469 13753 29503 13787
rect 3249 13685 3283 13719
rect 3525 13685 3559 13719
rect 4267 13685 4301 13719
rect 6567 13685 6601 13719
rect 8867 13685 8901 13719
rect 14663 13685 14697 13719
rect 20275 13685 20309 13719
rect 29561 13685 29595 13719
rect 6193 13481 6227 13515
rect 8585 13481 8619 13515
rect 8953 13481 8987 13515
rect 9229 13481 9263 13515
rect 9505 13481 9539 13515
rect 9781 13481 9815 13515
rect 11437 13481 11471 13515
rect 11897 13481 11931 13515
rect 12265 13481 12299 13515
rect 14749 13481 14783 13515
rect 17969 13481 18003 13515
rect 18803 13481 18837 13515
rect 22391 13481 22425 13515
rect 24599 13481 24633 13515
rect 26157 13481 26191 13515
rect 28273 13481 28307 13515
rect 30021 13481 30055 13515
rect 30389 13481 30423 13515
rect 5641 13413 5675 13447
rect 15301 13413 15335 13447
rect 1225 13345 1259 13379
rect 3433 13345 3467 13379
rect 6009 13345 6043 13379
rect 6377 13345 6411 13379
rect 6653 13369 6687 13403
rect 9137 13345 9171 13379
rect 9413 13345 9447 13379
rect 9689 13345 9723 13379
rect 9965 13345 9999 13379
rect 10241 13345 10275 13379
rect 10517 13345 10551 13379
rect 10793 13345 10827 13379
rect 11161 13345 11195 13379
rect 11713 13345 11747 13379
rect 12173 13345 12207 13379
rect 12449 13345 12483 13379
rect 12868 13345 12902 13379
rect 14933 13345 14967 13379
rect 15025 13345 15059 13379
rect 15945 13345 15979 13379
rect 21833 13345 21867 13379
rect 21925 13345 21959 13379
rect 24041 13345 24075 13379
rect 26760 13345 26794 13379
rect 28641 13345 28675 13379
rect 28917 13345 28951 13379
rect 30573 13345 30607 13379
rect 1317 13277 1351 13311
rect 1644 13277 1678 13311
rect 1813 13295 1847 13329
rect 2053 13277 2087 13311
rect 3525 13277 3559 13311
rect 3852 13277 3886 13311
rect 3988 13279 4022 13313
rect 4261 13277 4295 13311
rect 6753 13277 6787 13311
rect 7072 13277 7106 13311
rect 7208 13277 7242 13311
rect 7481 13277 7515 13311
rect 12541 13277 12575 13311
rect 13047 13277 13081 13311
rect 13277 13277 13311 13311
rect 16129 13277 16163 13311
rect 16456 13277 16490 13311
rect 16592 13277 16626 13311
rect 16865 13277 16899 13311
rect 18337 13277 18371 13311
rect 18800 13277 18834 13311
rect 19073 13277 19107 13311
rect 22431 13277 22465 13311
rect 22661 13277 22695 13311
rect 24133 13277 24167 13311
rect 24596 13295 24630 13329
rect 24869 13277 24903 13311
rect 26433 13277 26467 13311
rect 26896 13277 26930 13311
rect 27169 13277 27203 13311
rect 11345 13209 11379 13243
rect 1041 13141 1075 13175
rect 5825 13141 5859 13175
rect 6469 13141 6503 13175
rect 10057 13141 10091 13175
rect 10333 13141 10367 13175
rect 10609 13141 10643 13175
rect 11989 13141 12023 13175
rect 14381 13141 14415 13175
rect 15761 13141 15795 13175
rect 20361 13141 20395 13175
rect 21649 13141 21683 13175
rect 3525 12937 3559 12971
rect 5917 12937 5951 12971
rect 8769 12937 8803 12971
rect 12541 12937 12575 12971
rect 18245 12937 18279 12971
rect 23121 12937 23155 12971
rect 25697 12937 25731 12971
rect 28733 12937 28767 12971
rect 29377 12937 29411 12971
rect 29653 12937 29687 12971
rect 29929 12937 29963 12971
rect 9045 12869 9079 12903
rect 30205 12869 30239 12903
rect 949 12801 983 12835
rect 1455 12801 1489 12835
rect 3065 12801 3099 12835
rect 4356 12801 4390 12835
rect 4629 12801 4663 12835
rect 6607 12799 6641 12833
rect 6837 12801 6871 12835
rect 10060 12801 10094 12835
rect 10333 12801 10367 12835
rect 12081 12801 12115 12835
rect 14016 12801 14050 12835
rect 16224 12801 16258 12835
rect 16497 12801 16531 12835
rect 19168 12801 19202 12835
rect 21376 12801 21410 12835
rect 24320 12801 24354 12835
rect 27205 12783 27239 12817
rect 1685 12733 1719 12767
rect 3433 12733 3467 12767
rect 3709 12733 3743 12767
rect 3893 12733 3927 12767
rect 6101 12733 6135 12767
rect 8401 12733 8435 12767
rect 8953 12733 8987 12767
rect 9229 12733 9263 12767
rect 9505 12733 9539 12767
rect 9597 12733 9631 12767
rect 9924 12733 9958 12767
rect 11713 12733 11747 12767
rect 11805 12733 11839 12767
rect 12357 12733 12391 12767
rect 12817 12733 12851 12767
rect 13093 12733 13127 12767
rect 13369 12733 13403 12767
rect 13553 12733 13587 12767
rect 14289 12733 14323 12767
rect 15761 12733 15795 12767
rect 16088 12733 16122 12767
rect 18153 12733 18187 12767
rect 18429 12733 18463 12767
rect 18705 12733 18739 12767
rect 19032 12733 19066 12767
rect 19441 12733 19475 12767
rect 20913 12733 20947 12767
rect 21649 12733 21683 12767
rect 23305 12733 23339 12767
rect 23581 12733 23615 12767
rect 23857 12733 23891 12767
rect 24593 12733 24627 12767
rect 26065 12733 26099 12767
rect 26709 12733 26743 12767
rect 27445 12733 27479 12767
rect 29561 12733 29595 12767
rect 29837 12733 29871 12767
rect 30113 12733 30147 12767
rect 30389 12733 30423 12767
rect 8217 12665 8251 12699
rect 20821 12665 20855 12699
rect 26341 12665 26375 12699
rect 29101 12665 29135 12699
rect 1415 12597 1449 12631
rect 3249 12597 3283 12631
rect 4359 12597 4393 12631
rect 6567 12597 6601 12631
rect 8585 12597 8619 12631
rect 9321 12597 9355 12631
rect 11989 12597 12023 12631
rect 12633 12597 12667 12631
rect 12909 12597 12943 12631
rect 13185 12597 13219 12631
rect 14019 12597 14053 12631
rect 15393 12597 15427 12631
rect 17601 12597 17635 12631
rect 17969 12597 18003 12631
rect 21379 12597 21413 12631
rect 22753 12597 22787 12631
rect 23397 12597 23431 12631
rect 24323 12597 24357 12631
rect 27175 12597 27209 12631
rect 29193 12597 29227 12631
rect 5825 12393 5859 12427
rect 6193 12393 6227 12427
rect 6935 12393 6969 12427
rect 8493 12393 8527 12427
rect 11253 12393 11287 12427
rect 13007 12393 13041 12427
rect 15301 12393 15335 12427
rect 16129 12393 16163 12427
rect 17423 12393 17457 12427
rect 18797 12393 18831 12427
rect 19717 12393 19751 12427
rect 20361 12393 20395 12427
rect 20913 12393 20947 12427
rect 21747 12393 21781 12427
rect 23121 12393 23155 12427
rect 23955 12393 23989 12427
rect 25329 12393 25363 12427
rect 26899 12393 26933 12427
rect 28273 12393 28307 12427
rect 30573 12393 30607 12427
rect 15025 12325 15059 12359
rect 26157 12325 26191 12359
rect 1225 12257 1259 12291
rect 1644 12257 1678 12291
rect 3433 12257 3467 12291
rect 4261 12257 4295 12291
rect 6009 12257 6043 12291
rect 6377 12257 6411 12291
rect 7205 12257 7239 12291
rect 9413 12257 9447 12291
rect 11161 12257 11195 12291
rect 11529 12257 11563 12291
rect 11805 12257 11839 12291
rect 12449 12257 12483 12291
rect 13277 12257 13311 12291
rect 14749 12257 14783 12291
rect 15485 12257 15519 12291
rect 15761 12257 15795 12291
rect 16313 12257 16347 12291
rect 16865 12257 16899 12291
rect 17693 12257 17727 12291
rect 19349 12257 19383 12291
rect 19625 12257 19659 12291
rect 19901 12257 19935 12291
rect 20545 12257 20579 12291
rect 20821 12257 20855 12291
rect 21097 12257 21131 12291
rect 21281 12257 21315 12291
rect 22017 12257 22051 12291
rect 24225 12257 24259 12291
rect 25789 12257 25823 12291
rect 28917 12257 28951 12291
rect 30389 12257 30423 12291
rect 1317 12189 1351 12223
rect 1780 12189 1814 12223
rect 2053 12189 2087 12223
rect 3525 12189 3559 12223
rect 3852 12189 3886 12223
rect 3988 12191 4022 12225
rect 6469 12189 6503 12223
rect 6932 12189 6966 12223
rect 8677 12189 8711 12223
rect 9004 12189 9038 12223
rect 9140 12191 9174 12225
rect 12541 12189 12575 12223
rect 13004 12207 13038 12241
rect 16957 12189 16991 12223
rect 17420 12191 17454 12225
rect 21744 12189 21778 12223
rect 23489 12189 23523 12223
rect 23952 12189 23986 12223
rect 26433 12189 26467 12223
rect 26896 12189 26930 12223
rect 27169 12189 27203 12223
rect 28641 12189 28675 12223
rect 11989 12121 12023 12155
rect 20637 12121 20671 12155
rect 1041 12053 1075 12087
rect 5549 12053 5583 12087
rect 10701 12053 10735 12087
rect 10977 12053 11011 12087
rect 11713 12053 11747 12087
rect 12265 12053 12299 12087
rect 14565 12053 14599 12087
rect 15577 12053 15611 12087
rect 16681 12053 16715 12087
rect 19165 12053 19199 12087
rect 19441 12053 19475 12087
rect 30021 12053 30055 12087
rect 2789 11849 2823 11883
rect 5825 11849 5859 11883
rect 15945 11849 15979 11883
rect 20729 11849 20763 11883
rect 22937 11849 22971 11883
rect 26249 11849 26283 11883
rect 28273 11849 28307 11883
rect 28641 11849 28675 11883
rect 30297 11849 30331 11883
rect 3249 11781 3283 11815
rect 12081 11781 12115 11815
rect 13369 11781 13403 11815
rect 16129 11781 16163 11815
rect 23213 11781 23247 11815
rect 29377 11781 29411 11815
rect 30389 11781 30423 11815
rect 1455 11713 1489 11747
rect 3801 11713 3835 11747
rect 4264 11713 4298 11747
rect 4537 11713 4571 11747
rect 6564 11713 6598 11747
rect 6837 11713 6871 11747
rect 8677 11713 8711 11747
rect 10060 11713 10094 11747
rect 10333 11713 10367 11747
rect 11805 11713 11839 11747
rect 14016 11695 14050 11729
rect 16911 11713 16945 11747
rect 18521 11713 18555 11747
rect 19168 11713 19202 11747
rect 21376 11713 21410 11747
rect 21649 11713 21683 11747
rect 24731 11713 24765 11747
rect 26896 11713 26930 11747
rect 949 11645 983 11679
rect 1685 11645 1719 11679
rect 3433 11645 3467 11679
rect 3709 11645 3743 11679
rect 6101 11645 6135 11679
rect 8585 11645 8619 11679
rect 9597 11645 9631 11679
rect 12265 11645 12299 11679
rect 12541 11645 12575 11679
rect 13001 11645 13035 11679
rect 13185 11645 13219 11679
rect 13553 11645 13587 11679
rect 14289 11645 14323 11679
rect 16313 11645 16347 11679
rect 16405 11645 16439 11679
rect 17141 11645 17175 11679
rect 18705 11645 18739 11679
rect 19441 11645 19475 11679
rect 20913 11645 20947 11679
rect 23397 11645 23431 11679
rect 23673 11645 23707 11679
rect 23857 11645 23891 11679
rect 24225 11645 24259 11679
rect 24961 11645 24995 11679
rect 26433 11645 26467 11679
rect 27169 11645 27203 11679
rect 28825 11645 28859 11679
rect 29101 11645 29135 11679
rect 29561 11645 29595 11679
rect 29837 11645 29871 11679
rect 30113 11645 30147 11679
rect 30573 11645 30607 11679
rect 8217 11577 8251 11611
rect 9137 11577 9171 11611
rect 1415 11509 1449 11543
rect 3525 11509 3559 11543
rect 4267 11509 4301 11543
rect 6567 11509 6601 11543
rect 8401 11509 8435 11543
rect 9413 11509 9447 11543
rect 10063 11509 10097 11543
rect 11621 11509 11655 11543
rect 12357 11509 12391 11543
rect 12817 11509 12851 11543
rect 14019 11509 14053 11543
rect 15393 11509 15427 11543
rect 16871 11509 16905 11543
rect 19171 11509 19205 11543
rect 21379 11509 21413 11543
rect 23489 11509 23523 11543
rect 24041 11509 24075 11543
rect 24691 11509 24725 11543
rect 26899 11509 26933 11543
rect 29193 11509 29227 11543
rect 29653 11509 29687 11543
rect 1317 11305 1351 11339
rect 1967 11305 2001 11339
rect 11529 11305 11563 11339
rect 13007 11305 13041 11339
rect 18889 11305 18923 11339
rect 23955 11305 23989 11339
rect 25329 11305 25363 11339
rect 27537 11305 27571 11339
rect 27813 11305 27847 11339
rect 29929 11305 29963 11339
rect 30481 11305 30515 11339
rect 3617 11237 3651 11271
rect 3985 11237 4019 11271
rect 5365 11237 5399 11271
rect 11897 11237 11931 11271
rect 15853 11237 15887 11271
rect 16313 11237 16347 11271
rect 19349 11237 19383 11271
rect 26709 11237 26743 11271
rect 27077 11237 27111 11271
rect 1041 11169 1075 11203
rect 1501 11169 1535 11203
rect 2237 11169 2271 11203
rect 3709 11169 3743 11203
rect 4445 11169 4479 11203
rect 4629 11169 4663 11203
rect 5089 11169 5123 11203
rect 5825 11169 5859 11203
rect 8217 11169 8251 11203
rect 9413 11169 9447 11203
rect 11161 11169 11195 11203
rect 11437 11169 11471 11203
rect 11713 11169 11747 11203
rect 12265 11169 12299 11203
rect 13277 11169 13311 11203
rect 14933 11169 14967 11203
rect 15209 11169 15243 11203
rect 17601 11169 17635 11203
rect 19073 11169 19107 11203
rect 24225 11169 24259 11203
rect 25789 11169 25823 11203
rect 26433 11169 26467 11203
rect 27721 11169 27755 11203
rect 27997 11169 28031 11203
rect 28416 11169 28450 11203
rect 28825 11169 28859 11203
rect 30297 11169 30331 11203
rect 1997 11119 2031 11153
rect 4905 11101 4939 11135
rect 6152 11101 6186 11135
rect 6288 11101 6322 11135
rect 6561 11101 6595 11135
rect 7941 11101 7975 11135
rect 8677 11101 8711 11135
rect 9004 11101 9038 11135
rect 9140 11103 9174 11137
rect 10793 11101 10827 11135
rect 12541 11101 12575 11135
rect 13004 11101 13038 11135
rect 16865 11101 16899 11135
rect 17192 11101 17226 11135
rect 17371 11101 17405 11135
rect 21281 11101 21315 11135
rect 21608 11101 21642 11135
rect 21777 11119 21811 11153
rect 22017 11101 22051 11135
rect 23489 11101 23523 11135
rect 23952 11101 23986 11135
rect 28089 11101 28123 11135
rect 28595 11101 28629 11135
rect 4261 11033 4295 11067
rect 11253 11033 11287 11067
rect 12081 11033 12115 11067
rect 12449 11033 12483 11067
rect 15025 11033 15059 11067
rect 23305 11033 23339 11067
rect 8401 10965 8435 10999
rect 10977 10965 11011 10999
rect 14381 10965 14415 10999
rect 14749 10965 14783 10999
rect 15485 10965 15519 10999
rect 25881 10965 25915 10999
rect 27169 10965 27203 10999
rect 23029 10761 23063 10795
rect 25881 10761 25915 10795
rect 30389 10761 30423 10795
rect 11621 10693 11655 10727
rect 13829 10693 13863 10727
rect 28457 10693 28491 10727
rect 29193 10693 29227 10727
rect 949 10625 983 10659
rect 1455 10625 1489 10659
rect 3712 10625 3746 10659
rect 6012 10625 6046 10659
rect 7665 10625 7699 10659
rect 8769 10625 8803 10659
rect 9924 10625 9958 10659
rect 10060 10625 10094 10659
rect 10333 10625 10367 10659
rect 13093 10625 13127 10659
rect 14248 10625 14282 10659
rect 14427 10625 14461 10659
rect 14657 10625 14691 10659
rect 16868 10625 16902 10659
rect 20683 10625 20717 10659
rect 24320 10625 24354 10659
rect 24593 10625 24627 10659
rect 26576 10625 26610 10659
rect 26712 10623 26746 10657
rect 1685 10557 1719 10591
rect 3249 10557 3283 10591
rect 3985 10557 4019 10591
rect 5549 10557 5583 10591
rect 5876 10557 5910 10591
rect 6285 10557 6319 10591
rect 8493 10557 8527 10591
rect 9045 10557 9079 10591
rect 9623 10557 9657 10591
rect 12909 10557 12943 10591
rect 13921 10557 13955 10591
rect 16405 10557 16439 10591
rect 16732 10557 16766 10591
rect 17141 10557 17175 10591
rect 18797 10557 18831 10591
rect 19165 10557 19199 10591
rect 20177 10557 20211 10591
rect 20913 10557 20947 10591
rect 22569 10557 22603 10591
rect 23213 10557 23247 10591
rect 23857 10557 23891 10591
rect 26249 10557 26283 10591
rect 26985 10557 27019 10591
rect 28641 10557 28675 10591
rect 29009 10557 29043 10591
rect 29377 10557 29411 10591
rect 29929 10557 29963 10591
rect 30205 10557 30239 10591
rect 30573 10557 30607 10591
rect 3065 10489 3099 10523
rect 5365 10489 5399 10523
rect 7849 10489 7883 10523
rect 11897 10489 11931 10523
rect 12449 10489 12483 10523
rect 12817 10489 12851 10523
rect 13645 10489 13679 10523
rect 18521 10489 18555 10523
rect 28365 10489 28399 10523
rect 1415 10421 1449 10455
rect 3715 10421 3749 10455
rect 7941 10421 7975 10455
rect 9229 10421 9263 10455
rect 11989 10421 12023 10455
rect 15761 10421 15795 10455
rect 20643 10421 20677 10455
rect 22017 10421 22051 10455
rect 22385 10421 22419 10455
rect 24323 10421 24357 10455
rect 29561 10421 29595 10455
rect 29745 10421 29779 10455
rect 30021 10421 30055 10455
rect 1507 10217 1541 10251
rect 3715 10217 3749 10251
rect 5457 10217 5491 10251
rect 9143 10217 9177 10251
rect 14295 10217 14329 10251
rect 17883 10217 17917 10251
rect 19257 10217 19291 10251
rect 20361 10217 20395 10251
rect 23305 10217 23339 10251
rect 26157 10217 26191 10251
rect 26899 10217 26933 10251
rect 16221 10149 16255 10183
rect 1041 10081 1075 10115
rect 3985 10081 4019 10115
rect 5641 10081 5675 10115
rect 5927 10081 5961 10115
rect 6193 10081 6227 10115
rect 8585 10081 8619 10115
rect 9413 10081 9447 10115
rect 13737 10081 13771 10115
rect 13829 10081 13863 10115
rect 16865 10081 16899 10115
rect 18153 10081 18187 10115
rect 19809 10081 19843 10115
rect 20545 10081 20579 10115
rect 20821 10081 20855 10115
rect 21097 10081 21131 10115
rect 21281 10081 21315 10115
rect 21608 10081 21642 10115
rect 22017 10081 22051 10115
rect 24460 10081 24494 10115
rect 28641 10081 28675 10115
rect 28917 10081 28951 10115
rect 30389 10081 30423 10115
rect 1537 10031 1571 10065
rect 1777 10013 1811 10047
rect 3249 10013 3283 10047
rect 3712 10013 3746 10047
rect 6469 10013 6503 10047
rect 6796 10013 6830 10047
rect 6975 10013 7009 10047
rect 7205 10013 7239 10047
rect 8677 10013 8711 10047
rect 9140 10031 9174 10065
rect 11161 10013 11195 10047
rect 11488 10013 11522 10047
rect 11624 10013 11658 10047
rect 11897 10013 11931 10047
rect 14292 10013 14326 10047
rect 14565 10013 14599 10047
rect 15945 10013 15979 10047
rect 17049 10013 17083 10047
rect 17417 10013 17451 10047
rect 17923 10013 17957 10047
rect 21787 10013 21821 10047
rect 24133 10013 24167 10047
rect 24639 10013 24673 10047
rect 24869 10013 24903 10047
rect 26433 10013 26467 10047
rect 26896 10013 26930 10047
rect 27169 10013 27203 10047
rect 20637 9945 20671 9979
rect 30481 9945 30515 9979
rect 3065 9877 3099 9911
rect 5273 9877 5307 9911
rect 10701 9877 10735 9911
rect 13001 9877 13035 9911
rect 13553 9877 13587 9911
rect 16497 9877 16531 9911
rect 19625 9877 19659 9911
rect 20913 9877 20947 9911
rect 28273 9877 28307 9911
rect 30021 9877 30055 9911
rect 5825 9673 5859 9707
rect 22753 9673 22787 9707
rect 26617 9673 26651 9707
rect 27997 9673 28031 9707
rect 10977 9605 11011 9639
rect 13553 9605 13587 9639
rect 16129 9605 16163 9639
rect 27445 9605 27479 9639
rect 27721 9605 27755 9639
rect 949 9537 983 9571
rect 1455 9537 1489 9571
rect 3804 9537 3838 9571
rect 5457 9537 5491 9571
rect 6101 9537 6135 9571
rect 6607 9537 6641 9571
rect 8953 9537 8987 9571
rect 9280 9537 9314 9571
rect 9459 9537 9493 9571
rect 11624 9537 11658 9571
rect 14335 9537 14369 9571
rect 16405 9537 16439 9571
rect 16868 9537 16902 9571
rect 19211 9537 19245 9571
rect 20821 9537 20855 9571
rect 21419 9537 21453 9571
rect 24593 9537 24627 9571
rect 25099 9537 25133 9571
rect 27261 9537 27295 9571
rect 1685 9469 1719 9503
rect 3341 9469 3375 9503
rect 4077 9469 4111 9503
rect 5733 9469 5767 9503
rect 6009 9469 6043 9503
rect 6837 9469 6871 9503
rect 8401 9469 8435 9503
rect 9689 9469 9723 9503
rect 11161 9469 11195 9503
rect 11488 9469 11522 9503
rect 11897 9469 11931 9503
rect 13737 9469 13771 9503
rect 13829 9469 13863 9503
rect 14565 9469 14599 9503
rect 16313 9469 16347 9503
rect 16732 9469 16766 9503
rect 17141 9469 17175 9503
rect 18705 9469 18739 9503
rect 19441 9469 19475 9503
rect 20913 9469 20947 9503
rect 21649 9469 21683 9503
rect 23673 9469 23707 9503
rect 24041 9469 24075 9503
rect 24317 9469 24351 9503
rect 24920 9469 24954 9503
rect 25329 9469 25363 9503
rect 27629 9469 27663 9503
rect 27905 9469 27939 9503
rect 28181 9469 28215 9503
rect 28457 9469 28491 9503
rect 8217 9401 8251 9435
rect 18521 9401 18555 9435
rect 26985 9401 27019 9435
rect 1415 9333 1449 9367
rect 2973 9333 3007 9367
rect 3807 9333 3841 9367
rect 5549 9333 5583 9367
rect 6567 9333 6601 9367
rect 8585 9333 8619 9367
rect 13001 9333 13035 9367
rect 14295 9333 14329 9367
rect 15669 9333 15703 9367
rect 19171 9333 19205 9367
rect 21379 9333 21413 9367
rect 23489 9333 23523 9367
rect 23857 9333 23891 9367
rect 24133 9333 24167 9367
rect 28273 9333 28307 9367
rect 3715 9129 3749 9163
rect 5273 9129 5307 9163
rect 7389 9129 7423 9163
rect 8131 9129 8165 9163
rect 9505 9129 9539 9163
rect 10057 9129 10091 9163
rect 10609 9129 10643 9163
rect 11627 9129 11661 9163
rect 17883 9129 17917 9163
rect 20177 9129 20211 9163
rect 21747 9129 21781 9163
rect 23121 9129 23155 9163
rect 23955 9129 23989 9163
rect 25329 9129 25363 9163
rect 25697 9129 25731 9163
rect 25973 9129 26007 9163
rect 30113 9129 30147 9163
rect 3157 9061 3191 9095
rect 17141 9061 17175 9095
rect 19533 9061 19567 9095
rect 20729 9061 20763 9095
rect 1368 8993 1402 9027
rect 1777 8993 1811 9027
rect 3985 8993 4019 9027
rect 5641 8993 5675 9027
rect 5825 8993 5859 9027
rect 6469 8993 6503 9027
rect 6929 8993 6963 9027
rect 7205 8993 7239 9027
rect 7573 8993 7607 9027
rect 7665 8993 7699 9027
rect 8401 8993 8435 9027
rect 10241 8993 10275 9027
rect 10517 8993 10551 9027
rect 10793 8993 10827 9027
rect 11161 8993 11195 9027
rect 11897 8993 11931 9027
rect 13645 8993 13679 9027
rect 14064 8993 14098 9027
rect 14473 8993 14507 9027
rect 16865 8993 16899 9027
rect 17417 8993 17451 9027
rect 19717 8993 19751 9027
rect 20361 8993 20395 9027
rect 22017 8993 22051 9027
rect 24225 8993 24259 9027
rect 25881 8993 25915 9027
rect 26157 8993 26191 9027
rect 26433 8993 26467 9027
rect 27169 8993 27203 9027
rect 28733 8993 28767 9027
rect 29009 8993 29043 9027
rect 1041 8925 1075 8959
rect 1547 8925 1581 8959
rect 3249 8925 3283 8959
rect 3712 8927 3746 8961
rect 6009 8925 6043 8959
rect 8128 8925 8162 8959
rect 11624 8927 11658 8961
rect 13737 8925 13771 8959
rect 14243 8925 14277 8959
rect 17923 8925 17957 8959
rect 18153 8925 18187 8959
rect 21005 8925 21039 8959
rect 21281 8925 21315 8959
rect 21787 8925 21821 8959
rect 23489 8925 23523 8959
rect 23995 8925 24029 8959
rect 26760 8925 26794 8959
rect 26896 8925 26930 8959
rect 6653 8857 6687 8891
rect 6745 8857 6779 8891
rect 19901 8857 19935 8891
rect 5457 8789 5491 8823
rect 7021 8789 7055 8823
rect 10333 8789 10367 8823
rect 13001 8789 13035 8823
rect 13461 8789 13495 8823
rect 15577 8789 15611 8823
rect 16313 8789 16347 8823
rect 16773 8789 16807 8823
rect 28273 8789 28307 8823
rect 5089 8585 5123 8619
rect 7389 8585 7423 8619
rect 8401 8585 8435 8619
rect 11713 8585 11747 8619
rect 11897 8585 11931 8619
rect 17969 8585 18003 8619
rect 18153 8585 18187 8619
rect 20545 8585 20579 8619
rect 21189 8585 21223 8619
rect 25881 8585 25915 8619
rect 8677 8517 8711 8551
rect 8953 8517 8987 8551
rect 13093 8517 13127 8551
rect 1455 8449 1489 8483
rect 3576 8449 3610 8483
rect 3712 8431 3746 8465
rect 6012 8449 6046 8483
rect 6285 8449 6319 8483
rect 10152 8449 10186 8483
rect 10425 8449 10459 8483
rect 12633 8449 12667 8483
rect 13737 8449 13771 8483
rect 14200 8449 14234 8483
rect 14473 8449 14507 8483
rect 15853 8449 15887 8483
rect 16408 8449 16442 8483
rect 19211 8449 19245 8483
rect 21557 8449 21591 8483
rect 22063 8447 22097 8481
rect 23673 8449 23707 8483
rect 24320 8449 24354 8483
rect 26341 8449 26375 8483
rect 26668 8449 26702 8483
rect 26847 8449 26881 8483
rect 949 8381 983 8415
rect 1685 8381 1719 8415
rect 3249 8381 3283 8415
rect 3985 8381 4019 8415
rect 5549 8381 5583 8415
rect 7757 8381 7791 8415
rect 8585 8381 8619 8415
rect 8861 8381 8895 8415
rect 9137 8381 9171 8415
rect 9597 8381 9631 8415
rect 9689 8381 9723 8415
rect 10016 8381 10050 8415
rect 12081 8381 12115 8415
rect 13001 8381 13035 8415
rect 13277 8381 13311 8415
rect 14064 8381 14098 8415
rect 15945 8381 15979 8415
rect 16681 8381 16715 8415
rect 18337 8381 18371 8415
rect 18705 8381 18739 8415
rect 19441 8381 19475 8415
rect 21465 8381 21499 8415
rect 22293 8381 22327 8415
rect 23857 8381 23891 8415
rect 24593 8381 24627 8415
rect 27077 8381 27111 8415
rect 28733 8381 28767 8415
rect 29101 8381 29135 8415
rect 30205 8381 30239 8415
rect 8033 8313 8067 8347
rect 12357 8313 12391 8347
rect 29653 8313 29687 8347
rect 1415 8245 1449 8279
rect 2789 8245 2823 8279
rect 6015 8245 6049 8279
rect 9413 8245 9447 8279
rect 12817 8245 12851 8279
rect 16411 8245 16445 8279
rect 19171 8245 19205 8279
rect 21281 8245 21315 8279
rect 22023 8245 22057 8279
rect 24323 8245 24357 8279
rect 28181 8245 28215 8279
rect 28549 8245 28583 8279
rect 29377 8245 29411 8279
rect 29745 8245 29779 8279
rect 30297 8245 30331 8279
rect 1691 8041 1725 8075
rect 8309 8041 8343 8075
rect 9143 8041 9177 8075
rect 12087 8041 12121 8075
rect 14295 8041 14329 8075
rect 16595 8041 16629 8075
rect 20177 8041 20211 8075
rect 23121 8041 23155 8075
rect 23955 8041 23989 8075
rect 25329 8041 25363 8075
rect 28187 8041 28221 8075
rect 29561 8041 29595 8075
rect 5917 7973 5951 8007
rect 1133 7905 1167 7939
rect 6285 7905 6319 7939
rect 7205 7905 7239 7939
rect 8677 7905 8711 7939
rect 11069 7905 11103 7939
rect 12357 7905 12391 7939
rect 16129 7905 16163 7939
rect 18664 7905 18698 7939
rect 20729 7905 20763 7939
rect 21097 7905 21131 7939
rect 22017 7905 22051 7939
rect 24225 7905 24259 7939
rect 25881 7905 25915 7939
rect 26157 7905 26191 7939
rect 26709 7905 26743 7939
rect 26985 7905 27019 7939
rect 27261 7905 27295 7939
rect 27629 7905 27663 7939
rect 28457 7905 28491 7939
rect 30113 7905 30147 7939
rect 1225 7837 1259 7871
rect 1731 7837 1765 7871
rect 1961 7837 1995 7871
rect 3525 7837 3559 7871
rect 3852 7837 3886 7871
rect 4031 7837 4065 7871
rect 4261 7837 4295 7871
rect 6469 7837 6503 7871
rect 6796 7837 6830 7871
rect 6965 7855 6999 7889
rect 9183 7837 9217 7871
rect 9413 7837 9447 7871
rect 11345 7837 11379 7871
rect 11621 7837 11655 7871
rect 12127 7837 12161 7871
rect 13829 7837 13863 7871
rect 14335 7837 14369 7871
rect 14565 7837 14599 7871
rect 16625 7855 16659 7889
rect 16865 7837 16899 7871
rect 18337 7837 18371 7871
rect 18843 7837 18877 7871
rect 19073 7837 19107 7871
rect 21281 7837 21315 7871
rect 21608 7837 21642 7871
rect 21787 7837 21821 7871
rect 23489 7837 23523 7871
rect 23995 7837 24029 7871
rect 27721 7837 27755 7871
rect 28200 7839 28234 7873
rect 15669 7769 15703 7803
rect 20545 7769 20579 7803
rect 26525 7769 26559 7803
rect 949 7701 983 7735
rect 3065 7701 3099 7735
rect 5549 7701 5583 7735
rect 10517 7701 10551 7735
rect 13461 7701 13495 7735
rect 17969 7701 18003 7735
rect 20913 7701 20947 7735
rect 25697 7701 25731 7735
rect 25973 7701 26007 7735
rect 26801 7701 26835 7735
rect 29929 7701 29963 7735
rect 2973 7497 3007 7531
rect 5825 7497 5859 7531
rect 13829 7497 13863 7531
rect 16957 7497 16991 7531
rect 18337 7497 18371 7531
rect 22753 7497 22787 7531
rect 25697 7497 25731 7531
rect 28733 7497 28767 7531
rect 5549 7429 5583 7463
rect 7941 7429 7975 7463
rect 8769 7429 8803 7463
rect 16589 7429 16623 7463
rect 17785 7429 17819 7463
rect 18061 7429 18095 7463
rect 20729 7429 20763 7463
rect 29285 7429 29319 7463
rect 1445 7343 1479 7377
rect 3341 7361 3375 7395
rect 3668 7361 3702 7395
rect 3847 7361 3881 7395
rect 6564 7361 6598 7395
rect 6837 7361 6871 7395
rect 9372 7361 9406 7395
rect 9551 7361 9585 7395
rect 11253 7361 11287 7395
rect 11759 7361 11793 7395
rect 14749 7361 14783 7395
rect 15076 7361 15110 7395
rect 15255 7361 15289 7395
rect 15485 7361 15519 7395
rect 19032 7361 19066 7395
rect 19211 7361 19245 7395
rect 20913 7361 20947 7395
rect 21419 7361 21453 7395
rect 24320 7361 24354 7395
rect 24593 7361 24627 7395
rect 27036 7361 27070 7395
rect 27215 7361 27249 7395
rect 949 7293 983 7327
rect 1685 7293 1719 7327
rect 4077 7293 4111 7327
rect 5733 7293 5767 7327
rect 6009 7293 6043 7327
rect 6101 7293 6135 7327
rect 8677 7293 8711 7327
rect 8953 7293 8987 7327
rect 9045 7293 9079 7327
rect 9781 7293 9815 7327
rect 11989 7293 12023 7327
rect 13645 7293 13679 7327
rect 14105 7293 14139 7327
rect 14197 7293 14231 7327
rect 14473 7293 14507 7327
rect 17141 7293 17175 7327
rect 17417 7293 17451 7327
rect 17693 7293 17727 7327
rect 17969 7293 18003 7327
rect 18245 7293 18279 7327
rect 18521 7293 18555 7327
rect 18705 7293 18739 7327
rect 19441 7293 19475 7327
rect 21649 7293 21683 7327
rect 23857 7293 23891 7327
rect 26065 7293 26099 7327
rect 26709 7293 26743 7327
rect 27445 7293 27479 7327
rect 29193 7293 29227 7327
rect 29469 7293 29503 7327
rect 23213 7225 23247 7259
rect 23581 7225 23615 7259
rect 26341 7225 26375 7259
rect 1415 7157 1449 7191
rect 5181 7157 5215 7191
rect 6567 7157 6601 7191
rect 8493 7157 8527 7191
rect 11069 7157 11103 7191
rect 11719 7157 11753 7191
rect 13093 7157 13127 7191
rect 13921 7157 13955 7191
rect 17233 7157 17267 7191
rect 17509 7157 17543 7191
rect 21379 7157 21413 7191
rect 24323 7157 24357 7191
rect 29009 7157 29043 7191
rect 1599 6953 1633 6987
rect 6101 6953 6135 6987
rect 6935 6953 6969 6987
rect 9143 6953 9177 6987
rect 10517 6953 10551 6987
rect 11437 6953 11471 6987
rect 11713 6953 11747 6987
rect 11989 6953 12023 6987
rect 12639 6953 12673 6987
rect 14841 6953 14875 6987
rect 15669 6953 15703 6987
rect 22299 6953 22333 6987
rect 24599 6953 24633 6987
rect 25973 6953 26007 6987
rect 28187 6953 28221 6987
rect 23949 6885 23983 6919
rect 1041 6817 1075 6851
rect 3249 6817 3283 6851
rect 3525 6817 3559 6851
rect 4261 6817 4295 6851
rect 6009 6817 6043 6851
rect 6285 6817 6319 6851
rect 7205 6817 7239 6851
rect 11161 6817 11195 6851
rect 11253 6817 11287 6851
rect 11529 6817 11563 6851
rect 11805 6817 11839 6851
rect 12173 6817 12207 6851
rect 12909 6817 12943 6851
rect 14749 6817 14783 6851
rect 15025 6817 15059 6851
rect 15209 6817 15243 6851
rect 15853 6817 15887 6851
rect 16497 6817 16531 6851
rect 19308 6817 19342 6851
rect 21833 6817 21867 6851
rect 24869 6817 24903 6851
rect 27261 6817 27295 6851
rect 27721 6817 27755 6851
rect 28457 6817 28491 6851
rect 1133 6749 1167 6783
rect 1639 6751 1673 6785
rect 1869 6749 1903 6783
rect 3852 6749 3886 6783
rect 4031 6749 4065 6783
rect 6469 6749 6503 6783
rect 6932 6749 6966 6783
rect 8677 6749 8711 6783
rect 9183 6749 9217 6783
rect 9413 6749 9447 6783
rect 12679 6749 12713 6783
rect 16773 6749 16807 6783
rect 17100 6749 17134 6783
rect 17236 6749 17270 6783
rect 17509 6749 17543 6783
rect 18981 6749 19015 6783
rect 19487 6749 19521 6783
rect 19717 6749 19751 6783
rect 21557 6749 21591 6783
rect 22339 6749 22373 6783
rect 22569 6749 22603 6783
rect 24133 6749 24167 6783
rect 24596 6749 24630 6783
rect 28227 6749 28261 6783
rect 5825 6681 5859 6715
rect 10977 6681 11011 6715
rect 14565 6681 14599 6715
rect 857 6613 891 6647
rect 5365 6613 5399 6647
rect 8309 6613 8343 6647
rect 14013 6613 14047 6647
rect 15485 6613 15519 6647
rect 16313 6613 16347 6647
rect 18797 6613 18831 6647
rect 21005 6613 21039 6647
rect 27353 6613 27387 6647
rect 29745 6613 29779 6647
rect 5825 6409 5859 6443
rect 8861 6409 8895 6443
rect 9137 6409 9171 6443
rect 9413 6409 9447 6443
rect 11345 6409 11379 6443
rect 11805 6409 11839 6443
rect 13185 6409 13219 6443
rect 16681 6409 16715 6443
rect 22293 6409 22327 6443
rect 26341 6409 26375 6443
rect 28549 6409 28583 6443
rect 5549 6341 5583 6375
rect 7941 6341 7975 6375
rect 12909 6341 12943 6375
rect 18245 6341 18279 6375
rect 1455 6273 1489 6307
rect 3668 6273 3702 6307
rect 3847 6273 3881 6307
rect 6607 6273 6641 6307
rect 6837 6273 6871 6307
rect 10011 6273 10045 6307
rect 14473 6273 14507 6307
rect 15120 6273 15154 6307
rect 15393 6273 15427 6307
rect 19349 6273 19383 6307
rect 20456 6273 20490 6307
rect 22109 6273 22143 6307
rect 24501 6273 24535 6307
rect 25007 6271 25041 6305
rect 25237 6273 25271 6307
rect 27172 6273 27206 6307
rect 949 6205 983 6239
rect 1685 6205 1719 6239
rect 3341 6205 3375 6239
rect 4077 6205 4111 6239
rect 5733 6205 5767 6239
rect 6009 6205 6043 6239
rect 6101 6205 6135 6239
rect 8585 6205 8619 6239
rect 8677 6205 8711 6239
rect 8953 6205 8987 6239
rect 9229 6205 9263 6239
rect 9505 6205 9539 6239
rect 10241 6205 10275 6239
rect 11989 6181 12023 6215
rect 12265 6205 12299 6239
rect 12541 6205 12575 6239
rect 12817 6205 12851 6239
rect 13093 6205 13127 6239
rect 13369 6205 13403 6239
rect 13737 6205 13771 6239
rect 14013 6205 14047 6239
rect 14657 6205 14691 6239
rect 16865 6205 16899 6239
rect 17601 6205 17635 6239
rect 17877 6205 17911 6239
rect 18153 6205 18187 6239
rect 18429 6205 18463 6239
rect 18889 6205 18923 6239
rect 19165 6205 19199 6239
rect 19901 6205 19935 6239
rect 19993 6205 20027 6239
rect 20729 6205 20763 6239
rect 22477 6205 22511 6239
rect 22753 6205 22787 6239
rect 23029 6205 23063 6239
rect 24133 6205 24167 6239
rect 24409 6205 24443 6239
rect 26709 6205 26743 6239
rect 27445 6205 27479 6239
rect 29193 6205 29227 6239
rect 14197 6137 14231 6171
rect 17141 6137 17175 6171
rect 1415 6069 1449 6103
rect 2973 6069 3007 6103
rect 5181 6069 5215 6103
rect 6567 6069 6601 6103
rect 8401 6069 8435 6103
rect 9971 6069 10005 6103
rect 12081 6069 12115 6103
rect 12357 6069 12391 6103
rect 12633 6069 12667 6103
rect 13553 6069 13587 6103
rect 13829 6069 13863 6103
rect 15123 6069 15157 6103
rect 17417 6069 17451 6103
rect 17693 6069 17727 6103
rect 17969 6069 18003 6103
rect 18705 6069 18739 6103
rect 19717 6069 19751 6103
rect 20459 6069 20493 6103
rect 22569 6069 22603 6103
rect 22845 6069 22879 6103
rect 23949 6069 23983 6103
rect 24225 6069 24259 6103
rect 24967 6069 25001 6103
rect 27175 6069 27209 6103
rect 29009 6069 29043 6103
rect 857 5865 891 5899
rect 4077 5865 4111 5899
rect 4445 5865 4479 5899
rect 5641 5865 5675 5899
rect 6377 5865 6411 5899
rect 16595 5865 16629 5899
rect 20361 5865 20395 5899
rect 21281 5865 21315 5899
rect 22391 5865 22425 5899
rect 29377 5865 29411 5899
rect 1041 5729 1075 5763
rect 1644 5729 1678 5763
rect 3985 5729 4019 5763
rect 4629 5729 4663 5763
rect 4905 5729 4939 5763
rect 5917 5729 5951 5763
rect 6285 5729 6319 5763
rect 6561 5729 6595 5763
rect 6837 5729 6871 5763
rect 7113 5729 7147 5763
rect 7389 5729 7423 5763
rect 7665 5729 7699 5763
rect 10241 5729 10275 5763
rect 10517 5729 10551 5763
rect 10793 5729 10827 5763
rect 11253 5729 11287 5763
rect 11345 5729 11379 5763
rect 12357 5729 12391 5763
rect 13737 5729 13771 5763
rect 14565 5729 14599 5763
rect 16865 5729 16899 5763
rect 19073 5729 19107 5763
rect 20729 5729 20763 5763
rect 21005 5729 21039 5763
rect 21465 5729 21499 5763
rect 21833 5729 21867 5763
rect 22661 5729 22695 5763
rect 24133 5729 24167 5763
rect 24460 5729 24494 5763
rect 24869 5729 24903 5763
rect 26617 5729 26651 5763
rect 26893 5729 26927 5763
rect 27169 5729 27203 5763
rect 27445 5729 27479 5763
rect 28273 5729 28307 5763
rect 1317 5661 1351 5695
rect 1813 5679 1847 5713
rect 2053 5661 2087 5695
rect 7849 5661 7883 5695
rect 8176 5661 8210 5695
rect 8355 5661 8389 5695
rect 8585 5661 8619 5695
rect 9965 5661 9999 5695
rect 11621 5661 11655 5695
rect 11948 5661 11982 5695
rect 12084 5661 12118 5695
rect 13829 5661 13863 5695
rect 14156 5661 14190 5695
rect 14292 5661 14326 5695
rect 16129 5661 16163 5695
rect 16635 5661 16669 5695
rect 18337 5661 18371 5695
rect 18664 5661 18698 5695
rect 18800 5661 18834 5695
rect 21925 5661 21959 5695
rect 22388 5661 22422 5695
rect 24041 5661 24075 5695
rect 24596 5661 24630 5695
rect 27537 5661 27571 5695
rect 27864 5661 27898 5695
rect 28000 5661 28034 5695
rect 4721 5593 4755 5627
rect 7481 5593 7515 5627
rect 10609 5593 10643 5627
rect 11529 5593 11563 5627
rect 20545 5593 20579 5627
rect 26433 5593 26467 5627
rect 3341 5525 3375 5559
rect 3801 5525 3835 5559
rect 5181 5525 5215 5559
rect 6653 5525 6687 5559
rect 6929 5525 6963 5559
rect 7205 5525 7239 5559
rect 10057 5525 10091 5559
rect 10333 5525 10367 5559
rect 11069 5525 11103 5559
rect 15853 5525 15887 5559
rect 18153 5525 18187 5559
rect 20821 5525 20855 5559
rect 21649 5525 21683 5559
rect 26157 5525 26191 5559
rect 26709 5525 26743 5559
rect 26985 5525 27019 5559
rect 27261 5525 27295 5559
rect 3249 5321 3283 5355
rect 15669 5321 15703 5355
rect 26065 5321 26099 5355
rect 29469 5321 29503 5355
rect 8125 5253 8159 5287
rect 28549 5253 28583 5287
rect 949 5185 983 5219
rect 1455 5185 1489 5219
rect 3525 5185 3559 5219
rect 3988 5185 4022 5219
rect 6101 5185 6135 5219
rect 6564 5185 6598 5219
rect 9508 5183 9542 5217
rect 9781 5185 9815 5219
rect 11161 5185 11195 5219
rect 11716 5185 11750 5219
rect 11989 5185 12023 5219
rect 13369 5185 13403 5219
rect 14108 5185 14142 5219
rect 16316 5185 16350 5219
rect 16589 5185 16623 5219
rect 19168 5185 19202 5219
rect 20821 5185 20855 5219
rect 21376 5185 21410 5219
rect 21649 5185 21683 5219
rect 24320 5185 24354 5219
rect 27172 5185 27206 5219
rect 27445 5185 27479 5219
rect 1685 5117 1719 5151
rect 3433 5117 3467 5151
rect 4261 5117 4295 5151
rect 6837 5117 6871 5151
rect 8593 5113 8627 5147
rect 8861 5117 8895 5151
rect 9045 5117 9079 5151
rect 11253 5117 11287 5151
rect 13645 5117 13679 5151
rect 13972 5117 14006 5151
rect 14381 5117 14415 5151
rect 15853 5117 15887 5151
rect 18061 5117 18095 5151
rect 18705 5117 18739 5151
rect 19441 5117 19475 5151
rect 20913 5117 20947 5151
rect 21240 5117 21274 5151
rect 23857 5117 23891 5151
rect 24593 5117 24627 5151
rect 26249 5117 26283 5151
rect 26709 5117 26743 5151
rect 29193 5117 29227 5151
rect 29285 5117 29319 5151
rect 3065 5049 3099 5083
rect 17969 5049 18003 5083
rect 18337 5049 18371 5083
rect 23305 5049 23339 5083
rect 1415 4981 1449 5015
rect 3991 4981 4025 5015
rect 5365 4981 5399 5015
rect 6567 4981 6601 5015
rect 8401 4981 8435 5015
rect 8677 4981 8711 5015
rect 9511 4981 9545 5015
rect 11719 4981 11753 5015
rect 16319 4981 16353 5015
rect 19171 4981 19205 5015
rect 22753 4981 22787 5015
rect 24323 4981 24357 5015
rect 25697 4981 25731 5015
rect 27175 4981 27209 5015
rect 29009 4981 29043 5015
rect 949 4777 983 4811
rect 3157 4777 3191 4811
rect 5549 4777 5583 4811
rect 6935 4777 6969 4811
rect 10701 4777 10735 4811
rect 12087 4777 12121 4811
rect 14295 4777 14329 4811
rect 16595 4777 16629 4811
rect 18153 4777 18187 4811
rect 18803 4777 18837 4811
rect 27077 4777 27111 4811
rect 28003 4777 28037 4811
rect 15945 4709 15979 4743
rect 1133 4641 1167 4675
rect 1317 4641 1351 4675
rect 1644 4641 1678 4675
rect 3525 4641 3559 4675
rect 5825 4641 5859 4675
rect 8585 4641 8619 4675
rect 9413 4641 9447 4675
rect 11161 4641 11195 4675
rect 12357 4641 12391 4675
rect 13737 4641 13771 4675
rect 14565 4641 14599 4675
rect 16865 4641 16899 4675
rect 19073 4641 19107 4675
rect 20729 4641 20763 4675
rect 21005 4641 21039 4675
rect 21281 4641 21315 4675
rect 21833 4641 21867 4675
rect 22569 4641 22603 4675
rect 23949 4641 23983 4675
rect 24777 4641 24811 4675
rect 26801 4641 26835 4675
rect 26893 4641 26927 4675
rect 27537 4641 27571 4675
rect 1813 4591 1847 4625
rect 2053 4573 2087 4607
rect 3852 4573 3886 4607
rect 4031 4573 4065 4607
rect 4261 4573 4295 4607
rect 6009 4573 6043 4607
rect 6469 4573 6503 4607
rect 6975 4573 7009 4607
rect 7205 4573 7239 4607
rect 8677 4573 8711 4607
rect 9004 4573 9038 4607
rect 9140 4573 9174 4607
rect 11621 4573 11655 4607
rect 12127 4573 12161 4607
rect 13829 4573 13863 4607
rect 14292 4573 14326 4607
rect 16129 4573 16163 4607
rect 16592 4573 16626 4607
rect 18337 4573 18371 4607
rect 18800 4573 18834 4607
rect 22160 4573 22194 4607
rect 22339 4573 22373 4607
rect 24041 4573 24075 4607
rect 24368 4573 24402 4607
rect 24504 4575 24538 4609
rect 28043 4573 28077 4607
rect 28273 4573 28307 4607
rect 20545 4505 20579 4539
rect 29377 4505 29411 4539
rect 11253 4437 11287 4471
rect 20361 4437 20395 4471
rect 20821 4437 20855 4471
rect 21465 4437 21499 4471
rect 26065 4437 26099 4471
rect 26617 4437 26651 4471
rect 11897 4233 11931 4267
rect 12541 4233 12575 4267
rect 18981 4233 19015 4267
rect 949 4097 983 4131
rect 1455 4097 1489 4131
rect 1685 4097 1719 4131
rect 3988 4097 4022 4131
rect 6380 4097 6414 4131
rect 8033 4097 8067 4131
rect 9505 4097 9539 4131
rect 10336 4097 10370 4131
rect 10609 4097 10643 4131
rect 13185 4097 13219 4131
rect 14156 4097 14190 4131
rect 14292 4095 14326 4129
rect 16911 4095 16945 4129
rect 17141 4097 17175 4131
rect 20364 4097 20398 4131
rect 20637 4097 20671 4131
rect 22017 4097 22051 4131
rect 22569 4097 22603 4131
rect 24031 4097 24065 4131
rect 24547 4097 24581 4131
rect 24777 4097 24811 4131
rect 26712 4097 26746 4131
rect 26985 4097 27019 4131
rect 3433 4029 3467 4063
rect 3525 4029 3559 4063
rect 4261 4029 4295 4063
rect 5917 4029 5951 4063
rect 6653 4029 6687 4063
rect 8585 4029 8619 4063
rect 8953 4029 8987 4063
rect 9229 4029 9263 4063
rect 9321 4029 9355 4063
rect 9873 4029 9907 4063
rect 10200 4029 10234 4063
rect 12265 4029 12299 4063
rect 12909 4029 12943 4063
rect 13737 4029 13771 4063
rect 13829 4029 13863 4063
rect 14565 4029 14599 4063
rect 16313 4029 16347 4063
rect 16405 4029 16439 4063
rect 19533 4029 19567 4063
rect 19801 4029 19835 4063
rect 19901 4029 19935 4063
rect 22293 4029 22327 4063
rect 23029 4029 23063 4063
rect 23305 4029 23339 4063
rect 23673 4029 23707 4063
rect 26249 4029 26283 4063
rect 12449 3961 12483 3995
rect 18889 3961 18923 3995
rect 1415 3893 1449 3927
rect 2789 3893 2823 3927
rect 3249 3893 3283 3927
rect 3991 3893 4025 3927
rect 5549 3893 5583 3927
rect 6383 3893 6417 3927
rect 8401 3893 8435 3927
rect 8769 3893 8803 3927
rect 9045 3893 9079 3927
rect 12081 3893 12115 3927
rect 13553 3893 13587 3927
rect 15853 3893 15887 3927
rect 16129 3893 16163 3927
rect 16871 3893 16905 3927
rect 18245 3893 18279 3927
rect 19349 3893 19383 3927
rect 19625 3893 19659 3927
rect 20367 3893 20401 3927
rect 22845 3893 22879 3927
rect 23121 3893 23155 3927
rect 23489 3893 23523 3927
rect 24507 3893 24541 3927
rect 26065 3893 26099 3927
rect 26715 3893 26749 3927
rect 28089 3893 28123 3927
rect 1041 3689 1075 3723
rect 1317 3689 1351 3723
rect 7757 3689 7791 3723
rect 14295 3689 14329 3723
rect 16595 3689 16629 3723
rect 18803 3689 18837 3723
rect 21747 3689 21781 3723
rect 23955 3689 23989 3723
rect 2881 3621 2915 3655
rect 10793 3621 10827 3655
rect 13737 3621 13771 3655
rect 20453 3621 20487 3655
rect 26985 3621 27019 3655
rect 27629 3621 27663 3655
rect 1225 3553 1259 3587
rect 1501 3553 1535 3587
rect 1777 3553 1811 3587
rect 2513 3553 2547 3587
rect 4261 3553 4295 3587
rect 6244 3553 6278 3587
rect 6653 3553 6687 3587
rect 8125 3553 8159 3587
rect 9413 3553 9447 3587
rect 11069 3553 11103 3587
rect 14565 3553 14599 3587
rect 15945 3553 15979 3587
rect 16865 3553 16899 3587
rect 18245 3553 18279 3587
rect 19073 3553 19107 3587
rect 20545 3553 20579 3587
rect 20821 3553 20855 3587
rect 22017 3553 22051 3587
rect 24225 3553 24259 3587
rect 25697 3553 25731 3587
rect 26617 3553 26651 3587
rect 26709 3553 26743 3587
rect 27353 3553 27387 3587
rect 27905 3553 27939 3587
rect 3249 3485 3283 3519
rect 3525 3485 3559 3519
rect 3852 3485 3886 3519
rect 3988 3485 4022 3519
rect 5641 3485 5675 3519
rect 5917 3485 5951 3519
rect 6423 3485 6457 3519
rect 8401 3485 8435 3519
rect 8677 3485 8711 3519
rect 9004 3485 9038 3519
rect 9183 3485 9217 3519
rect 11345 3485 11379 3519
rect 11621 3485 11655 3519
rect 11948 3485 11982 3519
rect 12084 3487 12118 3521
rect 12357 3485 12391 3519
rect 13829 3485 13863 3519
rect 14292 3485 14326 3519
rect 16129 3485 16163 3519
rect 16592 3487 16626 3521
rect 18337 3485 18371 3519
rect 18800 3485 18834 3519
rect 21281 3485 21315 3519
rect 21744 3485 21778 3519
rect 23489 3485 23523 3519
rect 23952 3485 23986 3519
rect 25881 3485 25915 3519
rect 28232 3485 28266 3519
rect 28411 3485 28445 3519
rect 28641 3485 28675 3519
rect 1593 3417 1627 3451
rect 29745 3417 29779 3451
rect 23305 3349 23339 3383
rect 25329 3349 25363 3383
rect 26433 3349 26467 3383
rect 5549 3145 5583 3179
rect 13277 3145 13311 3179
rect 22937 3077 22971 3111
rect 28641 3077 28675 3111
rect 949 3009 983 3043
rect 1445 2991 1479 3025
rect 3065 3009 3099 3043
rect 4215 3009 4249 3043
rect 6101 3009 6135 3043
rect 6564 2991 6598 3025
rect 8769 3009 8803 3043
rect 9508 3009 9542 3043
rect 9781 3009 9815 3043
rect 11161 3009 11195 3043
rect 11716 3009 11750 3043
rect 14151 3009 14185 3043
rect 16316 3009 16350 3043
rect 16589 3009 16623 3043
rect 17969 3009 18003 3043
rect 19168 3009 19202 3043
rect 20821 3009 20855 3043
rect 21376 3009 21410 3043
rect 24320 3009 24354 3043
rect 24593 3009 24627 3043
rect 26712 3009 26746 3043
rect 1685 2941 1719 2975
rect 3709 2941 3743 2975
rect 4445 2941 4479 2975
rect 6837 2941 6871 2975
rect 8217 2941 8251 2975
rect 9045 2941 9079 2975
rect 11253 2941 11287 2975
rect 11989 2941 12023 2975
rect 13645 2941 13679 2975
rect 14381 2941 14415 2975
rect 15853 2941 15887 2975
rect 18153 2941 18187 2975
rect 18705 2941 18739 2975
rect 19441 2941 19475 2975
rect 20913 2941 20947 2975
rect 21649 2941 21683 2975
rect 23581 2941 23615 2975
rect 23857 2941 23891 2975
rect 26249 2941 26283 2975
rect 26985 2941 27019 2975
rect 28457 2941 28491 2975
rect 8493 2873 8527 2907
rect 23213 2873 23247 2907
rect 1415 2805 1449 2839
rect 4175 2805 4209 2839
rect 6567 2805 6601 2839
rect 9511 2805 9545 2839
rect 11719 2805 11753 2839
rect 14111 2805 14145 2839
rect 15485 2805 15519 2839
rect 16319 2805 16353 2839
rect 18245 2805 18279 2839
rect 19171 2805 19205 2839
rect 21379 2805 21413 2839
rect 24323 2805 24357 2839
rect 25697 2805 25731 2839
rect 26715 2805 26749 2839
rect 28089 2805 28123 2839
rect 949 2601 983 2635
rect 6469 2601 6503 2635
rect 7481 2601 7515 2635
rect 8223 2601 8257 2635
rect 9781 2601 9815 2635
rect 10057 2601 10091 2635
rect 10333 2601 10367 2635
rect 10609 2601 10643 2635
rect 14203 2601 14237 2635
rect 16595 2601 16629 2635
rect 18803 2601 18837 2635
rect 20821 2601 20855 2635
rect 21747 2601 21781 2635
rect 25973 2601 26007 2635
rect 26617 2601 26651 2635
rect 27353 2601 27387 2635
rect 28089 2601 28123 2635
rect 30021 2601 30055 2635
rect 20729 2533 20763 2567
rect 26525 2533 26559 2567
rect 1133 2465 1167 2499
rect 1644 2465 1678 2499
rect 2053 2465 2087 2499
rect 3801 2465 3835 2499
rect 6193 2465 6227 2499
rect 6377 2465 6411 2499
rect 6837 2465 6871 2499
rect 7665 2465 7699 2499
rect 8493 2465 8527 2499
rect 10241 2465 10275 2499
rect 10517 2465 10551 2499
rect 10793 2465 10827 2499
rect 11069 2465 11103 2499
rect 13645 2465 13679 2499
rect 16129 2465 16163 2499
rect 16865 2465 16899 2499
rect 21281 2465 21315 2499
rect 23673 2465 23707 2499
rect 23949 2465 23983 2499
rect 24133 2465 24167 2499
rect 27261 2465 27295 2499
rect 27905 2465 27939 2499
rect 28181 2465 28215 2499
rect 28508 2465 28542 2499
rect 28917 2465 28951 2499
rect 1317 2397 1351 2431
rect 1823 2399 1857 2433
rect 7021 2397 7055 2431
rect 7757 2397 7791 2431
rect 8220 2397 8254 2431
rect 11529 2397 11563 2431
rect 11856 2397 11890 2431
rect 12035 2397 12069 2431
rect 12265 2397 12299 2431
rect 13737 2397 13771 2431
rect 14243 2399 14277 2433
rect 14473 2397 14507 2431
rect 16592 2397 16626 2431
rect 18337 2397 18371 2431
rect 18800 2397 18834 2431
rect 19073 2397 19107 2431
rect 20453 2397 20487 2431
rect 21777 2415 21811 2449
rect 22017 2397 22051 2431
rect 24460 2397 24494 2431
rect 24629 2415 24663 2449
rect 24869 2397 24903 2431
rect 28644 2397 28678 2431
rect 6009 2329 6043 2363
rect 23489 2329 23523 2363
rect 3341 2261 3375 2295
rect 11161 2261 11195 2295
rect 15761 2261 15795 2295
rect 18153 2261 18187 2295
rect 23121 2261 23155 2295
rect 23765 2261 23799 2295
rect 2973 2057 3007 2091
rect 5549 2057 5583 2091
rect 7849 2057 7883 2091
rect 17877 2057 17911 2091
rect 23397 2057 23431 2091
rect 28181 2057 28215 2091
rect 28733 2057 28767 2091
rect 3249 1989 3283 2023
rect 8033 1989 8067 2023
rect 18061 1989 18095 2023
rect 1445 1903 1479 1937
rect 1685 1921 1719 1955
rect 3525 1921 3559 1955
rect 3988 1919 4022 1953
rect 6152 1921 6186 1955
rect 6288 1919 6322 1953
rect 6561 1921 6595 1955
rect 9045 1921 9079 1955
rect 9508 1919 9542 1953
rect 9781 1921 9815 1955
rect 11161 1921 11195 1955
rect 11716 1921 11750 1955
rect 13369 1921 13403 1955
rect 14108 1921 14142 1955
rect 14381 1921 14415 1955
rect 15761 1921 15795 1955
rect 16316 1921 16350 1955
rect 16589 1921 16623 1955
rect 18705 1921 18739 1955
rect 19168 1921 19202 1955
rect 20821 1921 20855 1955
rect 21376 1921 21410 1955
rect 21649 1921 21683 1955
rect 24320 1921 24354 1955
rect 26804 1921 26838 1955
rect 27077 1921 27111 1955
rect 949 1853 983 1887
rect 3433 1853 3467 1887
rect 3852 1853 3886 1887
rect 4261 1853 4295 1887
rect 5825 1853 5859 1887
rect 8217 1853 8251 1887
rect 8677 1853 8711 1887
rect 8953 1853 8987 1887
rect 11253 1853 11287 1887
rect 11989 1853 12023 1887
rect 13645 1853 13679 1887
rect 13972 1853 14006 1887
rect 15853 1853 15887 1887
rect 18245 1853 18279 1887
rect 18521 1853 18555 1887
rect 19441 1853 19475 1887
rect 20939 1853 20973 1887
rect 23305 1853 23339 1887
rect 23581 1853 23615 1887
rect 23857 1853 23891 1887
rect 24593 1853 24627 1887
rect 26341 1853 26375 1887
rect 28549 1853 28583 1887
rect 29009 1853 29043 1887
rect 23029 1785 23063 1819
rect 1415 1717 1449 1751
rect 8493 1717 8527 1751
rect 8769 1717 8803 1751
rect 9511 1717 9545 1751
rect 11719 1717 11753 1751
rect 16319 1717 16353 1751
rect 18337 1717 18371 1751
rect 19171 1717 19205 1751
rect 21379 1717 21413 1751
rect 23121 1717 23155 1751
rect 24323 1717 24357 1751
rect 25697 1717 25731 1751
rect 26807 1717 26841 1751
rect 29193 1717 29227 1751
rect 857 1513 891 1547
rect 3341 1513 3375 1547
rect 3991 1513 4025 1547
rect 6935 1513 6969 1547
rect 8493 1513 8527 1547
rect 9143 1513 9177 1547
rect 10977 1513 11011 1547
rect 11253 1513 11287 1547
rect 11995 1513 12029 1547
rect 14203 1513 14237 1547
rect 15761 1513 15795 1547
rect 16595 1513 16629 1547
rect 18153 1513 18187 1547
rect 18803 1513 18837 1547
rect 21747 1513 21781 1547
rect 23305 1513 23339 1547
rect 26617 1513 26651 1547
rect 26893 1513 26927 1547
rect 27169 1513 27203 1547
rect 27445 1513 27479 1547
rect 28003 1513 28037 1547
rect 29377 1513 29411 1547
rect 10793 1445 10827 1479
rect 20453 1445 20487 1479
rect 1041 1377 1075 1411
rect 5825 1377 5859 1411
rect 9413 1377 9447 1411
rect 11161 1377 11195 1411
rect 11437 1377 11471 1411
rect 16129 1377 16163 1411
rect 20729 1377 20763 1411
rect 21005 1377 21039 1411
rect 23816 1377 23850 1411
rect 24225 1377 24259 1411
rect 25881 1377 25915 1411
rect 25973 1377 26007 1411
rect 26433 1377 26467 1411
rect 26709 1377 26743 1411
rect 26985 1377 27019 1411
rect 27261 1377 27295 1411
rect 27537 1377 27571 1411
rect 1317 1309 1351 1343
rect 1644 1309 1678 1343
rect 1823 1309 1857 1343
rect 2053 1309 2087 1343
rect 3525 1309 3559 1343
rect 4021 1311 4055 1345
rect 4261 1309 4295 1343
rect 6009 1309 6043 1343
rect 6469 1309 6503 1343
rect 6965 1327 6999 1361
rect 7205 1309 7239 1343
rect 8677 1309 8711 1343
rect 9140 1309 9174 1343
rect 11529 1309 11563 1343
rect 12035 1309 12069 1343
rect 12265 1309 12299 1343
rect 13737 1309 13771 1343
rect 14200 1309 14234 1343
rect 14473 1309 14507 1343
rect 16592 1309 16626 1343
rect 16865 1309 16899 1343
rect 18337 1309 18371 1343
rect 18800 1309 18834 1343
rect 19073 1309 19107 1343
rect 21281 1309 21315 1343
rect 21744 1327 21778 1361
rect 22017 1309 22051 1343
rect 23489 1309 23523 1343
rect 23952 1309 23986 1343
rect 28033 1327 28067 1361
rect 28273 1309 28307 1343
rect 5549 1241 5583 1275
rect 20545 1241 20579 1275
rect 20821 1241 20855 1275
rect 13369 1173 13403 1207
rect 25329 1173 25363 1207
rect 25697 1173 25731 1207
rect 26157 1173 26191 1207
rect 2973 969 3007 1003
rect 3525 969 3559 1003
rect 4169 969 4203 1003
rect 5181 969 5215 1003
rect 5457 969 5491 1003
rect 8125 969 8159 1003
rect 10701 969 10735 1003
rect 13277 969 13311 1003
rect 15761 969 15795 1003
rect 16129 969 16163 1003
rect 18705 969 18739 1003
rect 23397 969 23431 1003
rect 25973 969 26007 1003
rect 26433 969 26467 1003
rect 3617 901 3651 935
rect 8401 901 8435 935
rect 10977 901 11011 935
rect 15393 901 15427 935
rect 23857 901 23891 935
rect 28549 901 28583 935
rect 949 833 983 867
rect 1445 815 1479 849
rect 1685 833 1719 867
rect 6564 833 6598 867
rect 9183 833 9217 867
rect 11253 833 11287 867
rect 11759 831 11793 865
rect 13553 833 13587 867
rect 14059 833 14093 867
rect 16901 815 16935 849
rect 19487 833 19521 867
rect 21557 833 21591 867
rect 22063 833 22097 867
rect 22293 833 22327 867
rect 24639 833 24673 867
rect 27215 833 27249 867
rect 3801 765 3835 799
rect 5089 765 5123 799
rect 5365 765 5399 799
rect 5641 765 5675 799
rect 6009 765 6043 799
rect 6101 765 6135 799
rect 6837 765 6871 799
rect 8585 765 8619 799
rect 8677 765 8711 799
rect 9413 765 9447 799
rect 11161 765 11195 799
rect 11989 765 12023 799
rect 14289 765 14323 799
rect 15945 765 15979 799
rect 16313 765 16347 799
rect 16405 765 16439 799
rect 17141 765 17175 799
rect 18889 765 18923 799
rect 18981 765 19015 799
rect 19308 765 19342 799
rect 19717 765 19751 799
rect 21465 765 21499 799
rect 24041 765 24075 799
rect 24133 765 24167 799
rect 24869 765 24903 799
rect 26617 765 26651 799
rect 26709 765 26743 799
rect 27445 765 27479 799
rect 1415 629 1449 663
rect 4813 629 4847 663
rect 4905 629 4939 663
rect 5825 629 5859 663
rect 6567 629 6601 663
rect 9143 629 9177 663
rect 11719 629 11753 663
rect 14019 629 14053 663
rect 16871 629 16905 663
rect 18245 629 18279 663
rect 20821 629 20855 663
rect 21281 629 21315 663
rect 22023 629 22057 663
rect 24599 629 24633 663
rect 27175 629 27209 663
<< metal1 >>
rect 10962 22244 10968 22296
rect 11020 22284 11026 22296
rect 18874 22284 18880 22296
rect 11020 22256 18880 22284
rect 11020 22244 11026 22256
rect 18874 22244 18880 22256
rect 18932 22244 18938 22296
rect 24210 22244 24216 22296
rect 24268 22284 24274 22296
rect 25038 22284 25044 22296
rect 24268 22256 25044 22284
rect 24268 22244 24274 22256
rect 25038 22244 25044 22256
rect 25096 22284 25102 22296
rect 31202 22284 31208 22296
rect 25096 22256 31208 22284
rect 25096 22244 25102 22256
rect 31202 22244 31208 22256
rect 31260 22244 31266 22296
rect 9122 22176 9128 22228
rect 9180 22216 9186 22228
rect 15746 22216 15752 22228
rect 9180 22188 15752 22216
rect 9180 22176 9186 22188
rect 15746 22176 15752 22188
rect 15804 22176 15810 22228
rect 16758 22216 16764 22228
rect 15856 22188 16764 22216
rect 7558 22108 7564 22160
rect 7616 22148 7622 22160
rect 15856 22148 15884 22188
rect 16758 22176 16764 22188
rect 16816 22176 16822 22228
rect 16850 22176 16856 22228
rect 16908 22216 16914 22228
rect 27614 22216 27620 22228
rect 16908 22188 27620 22216
rect 16908 22176 16914 22188
rect 27614 22176 27620 22188
rect 27672 22176 27678 22228
rect 7616 22120 15884 22148
rect 7616 22108 7622 22120
rect 15930 22108 15936 22160
rect 15988 22148 15994 22160
rect 25866 22148 25872 22160
rect 15988 22120 25872 22148
rect 15988 22108 15994 22120
rect 25866 22108 25872 22120
rect 25924 22108 25930 22160
rect 10502 22040 10508 22092
rect 10560 22080 10566 22092
rect 16114 22080 16120 22092
rect 10560 22052 16120 22080
rect 10560 22040 10566 22052
rect 16114 22040 16120 22052
rect 16172 22040 16178 22092
rect 18690 22080 18696 22092
rect 17426 22052 18696 22080
rect 10134 22012 10140 22024
rect 5460 21984 10140 22012
rect 5460 21956 5488 21984
rect 10134 21972 10140 21984
rect 10192 21972 10198 22024
rect 10594 21972 10600 22024
rect 10652 22012 10658 22024
rect 15562 22012 15568 22024
rect 10652 21984 15568 22012
rect 10652 21972 10658 21984
rect 15562 21972 15568 21984
rect 15620 21972 15626 22024
rect 17426 22012 17454 22052
rect 18690 22040 18696 22052
rect 18748 22040 18754 22092
rect 19242 22040 19248 22092
rect 19300 22080 19306 22092
rect 24118 22080 24124 22092
rect 19300 22052 24124 22080
rect 19300 22040 19306 22052
rect 24118 22040 24124 22052
rect 24176 22080 24182 22092
rect 28718 22080 28724 22092
rect 24176 22052 28724 22080
rect 24176 22040 24182 22052
rect 28718 22040 28724 22052
rect 28776 22040 28782 22092
rect 30282 22012 30288 22024
rect 16040 21984 17454 22012
rect 17512 21984 30288 22012
rect 5442 21904 5448 21956
rect 5500 21904 5506 21956
rect 7742 21904 7748 21956
rect 7800 21944 7806 21956
rect 11422 21944 11428 21956
rect 7800 21916 11428 21944
rect 7800 21904 7806 21916
rect 11422 21904 11428 21916
rect 11480 21904 11486 21956
rect 4798 21836 4804 21888
rect 4856 21876 4862 21888
rect 10318 21876 10324 21888
rect 4856 21848 10324 21876
rect 4856 21836 4862 21848
rect 10318 21836 10324 21848
rect 10376 21836 10382 21888
rect 10410 21836 10416 21888
rect 10468 21876 10474 21888
rect 16040 21876 16068 21984
rect 17512 21888 17540 21984
rect 30282 21972 30288 21984
rect 30340 21972 30346 22024
rect 19720 21916 27844 21944
rect 19720 21888 19748 21916
rect 27816 21888 27844 21916
rect 10468 21848 16068 21876
rect 10468 21836 10474 21848
rect 17494 21836 17500 21888
rect 17552 21836 17558 21888
rect 19702 21836 19708 21888
rect 19760 21836 19766 21888
rect 20622 21836 20628 21888
rect 20680 21876 20686 21888
rect 23382 21876 23388 21888
rect 20680 21848 23388 21876
rect 20680 21836 20686 21848
rect 23382 21836 23388 21848
rect 23440 21836 23446 21888
rect 24578 21836 24584 21888
rect 24636 21876 24642 21888
rect 25958 21876 25964 21888
rect 24636 21848 25964 21876
rect 24636 21836 24642 21848
rect 25958 21836 25964 21848
rect 26016 21836 26022 21888
rect 27798 21836 27804 21888
rect 27856 21836 27862 21888
rect 552 21786 30912 21808
rect 552 21734 4193 21786
rect 4245 21734 4257 21786
rect 4309 21734 4321 21786
rect 4373 21734 4385 21786
rect 4437 21734 4449 21786
rect 4501 21734 11783 21786
rect 11835 21734 11847 21786
rect 11899 21734 11911 21786
rect 11963 21734 11975 21786
rect 12027 21734 12039 21786
rect 12091 21734 19373 21786
rect 19425 21734 19437 21786
rect 19489 21734 19501 21786
rect 19553 21734 19565 21786
rect 19617 21734 19629 21786
rect 19681 21734 26963 21786
rect 27015 21734 27027 21786
rect 27079 21734 27091 21786
rect 27143 21734 27155 21786
rect 27207 21734 27219 21786
rect 27271 21734 30912 21786
rect 552 21712 30912 21734
rect 7558 21672 7564 21684
rect 2746 21644 7564 21672
rect 1673 21539 1731 21545
rect 1418 21521 1624 21536
rect 1418 21490 1445 21521
rect 1433 21487 1445 21490
rect 1479 21508 1624 21521
rect 1479 21487 1491 21508
rect 1433 21481 1491 21487
rect 842 21428 848 21480
rect 900 21468 906 21480
rect 937 21471 995 21477
rect 937 21468 949 21471
rect 900 21440 949 21468
rect 900 21428 906 21440
rect 937 21437 949 21440
rect 983 21437 995 21471
rect 1596 21468 1624 21508
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 2746 21536 2774 21644
rect 7558 21632 7564 21644
rect 7616 21632 7622 21684
rect 8021 21675 8079 21681
rect 8021 21641 8033 21675
rect 8067 21672 8079 21675
rect 11698 21672 11704 21684
rect 8067 21644 11704 21672
rect 8067 21641 8079 21644
rect 8021 21635 8079 21641
rect 11698 21632 11704 21644
rect 11756 21632 11762 21684
rect 12526 21632 12532 21684
rect 12584 21672 12590 21684
rect 13725 21675 13783 21681
rect 13725 21672 13737 21675
rect 12584 21644 13737 21672
rect 12584 21632 12590 21644
rect 13725 21641 13737 21644
rect 13771 21641 13783 21675
rect 16850 21672 16856 21684
rect 13725 21635 13783 21641
rect 14292 21644 16856 21672
rect 1719 21508 2774 21536
rect 3053 21539 3111 21545
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 3053 21505 3065 21539
rect 3099 21536 3111 21539
rect 3700 21539 3758 21545
rect 3700 21536 3712 21539
rect 3099 21508 3712 21536
rect 3099 21505 3111 21508
rect 3053 21499 3111 21505
rect 3700 21505 3712 21508
rect 3746 21505 3758 21539
rect 6276 21539 6334 21545
rect 6276 21536 6288 21539
rect 3700 21499 3758 21505
rect 4080 21508 6288 21536
rect 4080 21480 4108 21508
rect 6276 21505 6288 21508
rect 6322 21505 6334 21539
rect 8662 21536 8668 21548
rect 6276 21499 6334 21505
rect 6472 21508 8668 21536
rect 2774 21468 2780 21480
rect 1596 21440 2780 21468
rect 937 21431 995 21437
rect 2774 21428 2780 21440
rect 2832 21428 2838 21480
rect 3234 21428 3240 21480
rect 3292 21428 3298 21480
rect 3973 21471 4031 21477
rect 3973 21468 3985 21471
rect 3344 21440 3985 21468
rect 2866 21360 2872 21412
rect 2924 21400 2930 21412
rect 3344 21400 3372 21440
rect 3973 21437 3985 21440
rect 4019 21437 4031 21471
rect 3973 21431 4031 21437
rect 4062 21428 4068 21480
rect 4120 21428 4126 21480
rect 5442 21428 5448 21480
rect 5500 21468 5506 21480
rect 5629 21471 5687 21477
rect 5629 21468 5641 21471
rect 5500 21440 5641 21468
rect 5500 21428 5506 21440
rect 5629 21437 5641 21440
rect 5675 21437 5687 21471
rect 5629 21431 5687 21437
rect 5813 21471 5871 21477
rect 5813 21437 5825 21471
rect 5859 21437 5871 21471
rect 5813 21431 5871 21437
rect 2924 21372 3372 21400
rect 2924 21360 2930 21372
rect 5350 21360 5356 21412
rect 5408 21360 5414 21412
rect 5718 21360 5724 21412
rect 5776 21400 5782 21412
rect 5828 21400 5856 21431
rect 6178 21428 6184 21480
rect 6236 21468 6242 21480
rect 6472 21468 6500 21508
rect 8662 21496 8668 21508
rect 8720 21545 8726 21548
rect 8720 21539 8774 21545
rect 8720 21505 8728 21539
rect 8762 21505 8774 21539
rect 8868 21521 8926 21527
rect 8868 21518 8880 21521
rect 8720 21499 8774 21505
rect 8720 21496 8726 21499
rect 8867 21487 8880 21518
rect 8914 21487 8926 21521
rect 9122 21496 9128 21548
rect 9180 21496 9186 21548
rect 9582 21496 9588 21548
rect 9640 21536 9646 21548
rect 9640 21508 10916 21536
rect 9640 21496 9646 21508
rect 8867 21484 8926 21487
rect 8823 21481 8926 21484
rect 6236 21440 6500 21468
rect 6549 21471 6607 21477
rect 6236 21428 6242 21440
rect 6549 21437 6561 21471
rect 6595 21468 6607 21471
rect 7374 21468 7380 21480
rect 6595 21440 7380 21468
rect 6595 21437 6607 21440
rect 6549 21431 6607 21437
rect 7374 21428 7380 21440
rect 7432 21428 7438 21480
rect 8205 21471 8263 21477
rect 8205 21437 8217 21471
rect 8251 21468 8263 21471
rect 8294 21468 8300 21480
rect 8251 21440 8300 21468
rect 8251 21437 8263 21440
rect 8205 21431 8263 21437
rect 8294 21428 8300 21440
rect 8352 21428 8358 21480
rect 8386 21428 8392 21480
rect 8444 21428 8450 21480
rect 8823 21468 8895 21481
rect 8496 21456 8895 21468
rect 8496 21440 8851 21456
rect 5776 21372 5856 21400
rect 5776 21360 5782 21372
rect 7282 21360 7288 21412
rect 7340 21400 7346 21412
rect 8496 21400 8524 21440
rect 9766 21428 9772 21480
rect 9824 21468 9830 21480
rect 10781 21471 10839 21477
rect 10781 21468 10793 21471
rect 9824 21440 10793 21468
rect 9824 21428 9830 21440
rect 10781 21437 10793 21440
rect 10827 21437 10839 21471
rect 10888 21468 10916 21508
rect 11054 21496 11060 21548
rect 11112 21536 11118 21548
rect 11612 21539 11670 21545
rect 11612 21536 11624 21539
rect 11112 21508 11624 21536
rect 11112 21496 11118 21508
rect 11612 21505 11624 21508
rect 11658 21505 11670 21539
rect 11612 21499 11670 21505
rect 11149 21471 11207 21477
rect 11149 21468 11161 21471
rect 10888 21440 11161 21468
rect 10781 21431 10839 21437
rect 11149 21437 11161 21440
rect 11195 21468 11207 21471
rect 11238 21468 11244 21480
rect 11195 21440 11244 21468
rect 11195 21437 11207 21440
rect 11149 21431 11207 21437
rect 11238 21428 11244 21440
rect 11296 21428 11302 21480
rect 11422 21428 11428 21480
rect 11480 21468 11486 21480
rect 14292 21477 14320 21644
rect 16850 21632 16856 21644
rect 16908 21632 16914 21684
rect 18874 21632 18880 21684
rect 18932 21632 18938 21684
rect 22112 21644 22968 21672
rect 15562 21564 15568 21616
rect 15620 21604 15626 21616
rect 22005 21607 22063 21613
rect 15620 21576 16896 21604
rect 15620 21564 15626 21576
rect 16301 21539 16359 21545
rect 16301 21536 16313 21539
rect 14384 21508 16313 21536
rect 11885 21471 11943 21477
rect 11885 21468 11897 21471
rect 11480 21440 11897 21468
rect 11480 21428 11486 21440
rect 11885 21437 11897 21440
rect 11931 21437 11943 21471
rect 14277 21471 14335 21477
rect 11885 21431 11943 21437
rect 12912 21440 13952 21468
rect 7340 21372 8524 21400
rect 10152 21372 11284 21400
rect 7340 21360 7346 21372
rect 1394 21292 1400 21344
rect 1452 21341 1458 21344
rect 1452 21295 1461 21341
rect 1452 21292 1458 21295
rect 3602 21292 3608 21344
rect 3660 21332 3666 21344
rect 3703 21335 3761 21341
rect 3703 21332 3715 21335
rect 3660 21304 3715 21332
rect 3660 21292 3666 21304
rect 3703 21301 3715 21304
rect 3749 21332 3761 21335
rect 3878 21332 3884 21344
rect 3749 21304 3884 21332
rect 3749 21301 3761 21304
rect 3703 21295 3761 21301
rect 3878 21292 3884 21304
rect 3936 21292 3942 21344
rect 5445 21335 5503 21341
rect 5445 21301 5457 21335
rect 5491 21332 5503 21335
rect 5902 21332 5908 21344
rect 5491 21304 5908 21332
rect 5491 21301 5503 21304
rect 5445 21295 5503 21301
rect 5902 21292 5908 21304
rect 5960 21292 5966 21344
rect 6086 21292 6092 21344
rect 6144 21332 6150 21344
rect 6279 21335 6337 21341
rect 6279 21332 6291 21335
rect 6144 21304 6291 21332
rect 6144 21292 6150 21304
rect 6279 21301 6291 21304
rect 6325 21301 6337 21335
rect 6279 21295 6337 21301
rect 6454 21292 6460 21344
rect 6512 21332 6518 21344
rect 7653 21335 7711 21341
rect 7653 21332 7665 21335
rect 6512 21304 7665 21332
rect 6512 21292 6518 21304
rect 7653 21301 7665 21304
rect 7699 21301 7711 21335
rect 7653 21295 7711 21301
rect 8662 21292 8668 21344
rect 8720 21332 8726 21344
rect 10152 21332 10180 21372
rect 8720 21304 10180 21332
rect 8720 21292 8726 21304
rect 10226 21292 10232 21344
rect 10284 21292 10290 21344
rect 10597 21335 10655 21341
rect 10597 21301 10609 21335
rect 10643 21332 10655 21335
rect 10962 21332 10968 21344
rect 10643 21304 10968 21332
rect 10643 21301 10655 21304
rect 10597 21295 10655 21301
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 11256 21332 11284 21372
rect 11606 21332 11612 21344
rect 11664 21341 11670 21344
rect 11256 21304 11612 21332
rect 11606 21292 11612 21304
rect 11664 21332 11673 21341
rect 12342 21332 12348 21344
rect 11664 21304 12348 21332
rect 11664 21295 11673 21304
rect 11664 21292 11670 21295
rect 12342 21292 12348 21304
rect 12400 21332 12406 21344
rect 12912 21332 12940 21440
rect 13633 21403 13691 21409
rect 13633 21369 13645 21403
rect 13679 21400 13691 21403
rect 13814 21400 13820 21412
rect 13679 21372 13820 21400
rect 13679 21369 13691 21372
rect 13633 21363 13691 21369
rect 13814 21360 13820 21372
rect 13872 21360 13878 21412
rect 13924 21400 13952 21440
rect 14277 21437 14289 21471
rect 14323 21437 14335 21471
rect 14277 21431 14335 21437
rect 14384 21400 14412 21508
rect 16301 21505 16313 21508
rect 16347 21505 16359 21539
rect 16868 21536 16896 21576
rect 22005 21573 22017 21607
rect 22051 21604 22063 21607
rect 22112 21604 22140 21644
rect 22051 21576 22140 21604
rect 22940 21604 22968 21644
rect 23382 21632 23388 21684
rect 23440 21632 23446 21684
rect 23676 21644 24440 21672
rect 23676 21604 23704 21644
rect 24210 21604 24216 21616
rect 22940 21576 23704 21604
rect 23768 21576 24216 21604
rect 22051 21573 22063 21576
rect 22005 21567 22063 21573
rect 17129 21539 17187 21545
rect 16868 21508 16988 21536
rect 16301 21499 16359 21505
rect 14553 21471 14611 21477
rect 14553 21437 14565 21471
rect 14599 21468 14611 21471
rect 14599 21440 16068 21468
rect 14599 21437 14611 21440
rect 14553 21431 14611 21437
rect 13924 21372 14412 21400
rect 15930 21360 15936 21412
rect 15988 21360 15994 21412
rect 12400 21304 12940 21332
rect 12400 21292 12406 21304
rect 12986 21292 12992 21344
rect 13044 21292 13050 21344
rect 14182 21292 14188 21344
rect 14240 21332 14246 21344
rect 15470 21332 15476 21344
rect 14240 21304 15476 21332
rect 14240 21292 14246 21304
rect 15470 21292 15476 21304
rect 15528 21292 15534 21344
rect 16040 21332 16068 21440
rect 16114 21428 16120 21480
rect 16172 21428 16178 21480
rect 16850 21428 16856 21480
rect 16908 21428 16914 21480
rect 16960 21468 16988 21508
rect 17129 21505 17141 21539
rect 17175 21536 17187 21539
rect 20809 21539 20867 21545
rect 20809 21536 20821 21539
rect 17175 21508 20821 21536
rect 17175 21505 17187 21508
rect 17129 21499 17187 21505
rect 20809 21505 20821 21508
rect 20855 21505 20867 21539
rect 20809 21499 20867 21505
rect 22094 21496 22100 21548
rect 22152 21536 22158 21548
rect 22398 21539 22456 21545
rect 22398 21536 22410 21539
rect 22152 21508 22410 21536
rect 22152 21496 22158 21508
rect 22398 21505 22410 21508
rect 22444 21505 22456 21539
rect 22398 21499 22456 21505
rect 22557 21539 22615 21545
rect 22557 21505 22569 21539
rect 22603 21536 22615 21539
rect 23768 21536 23796 21576
rect 24210 21564 24216 21576
rect 24268 21564 24274 21616
rect 24412 21548 24440 21644
rect 24486 21632 24492 21684
rect 24544 21672 24550 21684
rect 25685 21675 25743 21681
rect 25685 21672 25697 21675
rect 24544 21644 25697 21672
rect 24544 21632 24550 21644
rect 25685 21641 25697 21644
rect 25731 21641 25743 21675
rect 25685 21635 25743 21641
rect 25958 21632 25964 21684
rect 26016 21632 26022 21684
rect 27798 21632 27804 21684
rect 27856 21632 27862 21684
rect 29641 21675 29699 21681
rect 29641 21641 29653 21675
rect 29687 21672 29699 21675
rect 29687 21644 30604 21672
rect 29687 21641 29699 21644
rect 29641 21635 29699 21641
rect 22603 21508 23796 21536
rect 23845 21539 23903 21545
rect 22603 21505 22615 21508
rect 22557 21499 22615 21505
rect 23845 21505 23857 21539
rect 23891 21536 23903 21539
rect 23934 21536 23940 21548
rect 23891 21508 23940 21536
rect 23891 21505 23903 21508
rect 23845 21499 23903 21505
rect 23934 21496 23940 21508
rect 23992 21496 23998 21548
rect 24394 21496 24400 21548
rect 24452 21536 24458 21548
rect 24489 21539 24547 21545
rect 24489 21536 24501 21539
rect 24452 21508 24501 21536
rect 24452 21496 24458 21508
rect 24489 21505 24501 21508
rect 24535 21505 24547 21539
rect 24489 21499 24547 21505
rect 24765 21539 24823 21545
rect 24765 21505 24777 21539
rect 24811 21536 24823 21539
rect 25682 21536 25688 21548
rect 24811 21508 25688 21536
rect 24811 21505 24823 21508
rect 24765 21499 24823 21505
rect 25682 21496 25688 21508
rect 25740 21496 25746 21548
rect 25976 21536 26004 21632
rect 30576 21616 30604 21644
rect 30377 21607 30435 21613
rect 30377 21573 30389 21607
rect 30423 21573 30435 21607
rect 30377 21567 30435 21573
rect 26421 21539 26479 21545
rect 26421 21536 26433 21539
rect 25976 21508 26433 21536
rect 26421 21505 26433 21508
rect 26467 21505 26479 21539
rect 26421 21499 26479 21505
rect 26786 21496 26792 21548
rect 26844 21536 26850 21548
rect 30392 21536 30420 21567
rect 30558 21564 30564 21616
rect 30616 21564 30622 21616
rect 26844 21508 30420 21536
rect 26844 21496 26850 21508
rect 18785 21471 18843 21477
rect 18785 21468 18797 21471
rect 16960 21440 18797 21468
rect 18785 21437 18797 21440
rect 18831 21437 18843 21471
rect 18785 21431 18843 21437
rect 19242 21428 19248 21480
rect 19300 21468 19306 21480
rect 19429 21471 19487 21477
rect 19429 21468 19441 21471
rect 19300 21440 19441 21468
rect 19300 21428 19306 21440
rect 19429 21437 19441 21440
rect 19475 21437 19487 21471
rect 19429 21431 19487 21437
rect 19702 21428 19708 21480
rect 19760 21428 19766 21480
rect 21361 21471 21419 21477
rect 21361 21437 21373 21471
rect 21407 21437 21419 21471
rect 21361 21431 21419 21437
rect 18506 21360 18512 21412
rect 18564 21360 18570 21412
rect 21376 21344 21404 21431
rect 21450 21428 21456 21480
rect 21508 21468 21514 21480
rect 21545 21471 21603 21477
rect 21545 21468 21557 21471
rect 21508 21440 21557 21468
rect 21508 21428 21514 21440
rect 21545 21437 21557 21440
rect 21591 21437 21603 21471
rect 21545 21431 21603 21437
rect 22278 21428 22284 21480
rect 22336 21428 22342 21480
rect 23569 21471 23627 21477
rect 23569 21437 23581 21471
rect 23615 21468 23627 21471
rect 23658 21468 23664 21480
rect 23615 21440 23664 21468
rect 23615 21437 23627 21440
rect 23569 21431 23627 21437
rect 23658 21428 23664 21440
rect 23716 21428 23722 21480
rect 24029 21471 24087 21477
rect 24029 21437 24041 21471
rect 24075 21437 24087 21471
rect 24029 21431 24087 21437
rect 18598 21332 18604 21344
rect 16040 21304 18604 21332
rect 18598 21292 18604 21304
rect 18656 21292 18662 21344
rect 21358 21292 21364 21344
rect 21416 21292 21422 21344
rect 23014 21292 23020 21344
rect 23072 21332 23078 21344
rect 23201 21335 23259 21341
rect 23201 21332 23213 21335
rect 23072 21304 23213 21332
rect 23072 21292 23078 21304
rect 23201 21301 23213 21304
rect 23247 21301 23259 21335
rect 24044 21332 24072 21431
rect 24854 21428 24860 21480
rect 24912 21477 24918 21480
rect 24912 21471 24940 21477
rect 24928 21437 24940 21471
rect 24912 21431 24940 21437
rect 24912 21428 24918 21431
rect 25038 21428 25044 21480
rect 25096 21428 25102 21480
rect 25777 21471 25835 21477
rect 25777 21437 25789 21471
rect 25823 21468 25835 21471
rect 26326 21468 26332 21480
rect 25823 21440 26332 21468
rect 25823 21437 25835 21440
rect 25777 21431 25835 21437
rect 26326 21428 26332 21440
rect 26384 21428 26390 21480
rect 26697 21471 26755 21477
rect 26697 21437 26709 21471
rect 26743 21468 26755 21471
rect 27338 21468 27344 21480
rect 26743 21440 27344 21468
rect 26743 21437 26755 21440
rect 26697 21431 26755 21437
rect 27338 21428 27344 21440
rect 27396 21428 27402 21480
rect 27614 21428 27620 21480
rect 27672 21468 27678 21480
rect 28261 21471 28319 21477
rect 28261 21468 28273 21471
rect 27672 21440 28273 21468
rect 27672 21428 27678 21440
rect 28261 21437 28273 21440
rect 28307 21468 28319 21471
rect 28350 21468 28356 21480
rect 28307 21440 28356 21468
rect 28307 21437 28319 21440
rect 28261 21431 28319 21437
rect 28350 21428 28356 21440
rect 28408 21428 28414 21480
rect 29086 21428 29092 21480
rect 29144 21428 29150 21480
rect 29270 21428 29276 21480
rect 29328 21428 29334 21480
rect 29365 21471 29423 21477
rect 29365 21437 29377 21471
rect 29411 21468 29423 21471
rect 30561 21471 30619 21477
rect 29411 21440 29868 21468
rect 29411 21437 29423 21440
rect 29365 21431 29423 21437
rect 29840 21412 29868 21440
rect 30561 21437 30573 21471
rect 30607 21468 30619 21471
rect 31110 21468 31116 21480
rect 30607 21440 31116 21468
rect 30607 21437 30619 21440
rect 30561 21431 30619 21437
rect 31110 21428 31116 21440
rect 31168 21428 31174 21480
rect 26053 21403 26111 21409
rect 26053 21369 26065 21403
rect 26099 21369 26111 21403
rect 26053 21363 26111 21369
rect 25314 21332 25320 21344
rect 24044 21304 25320 21332
rect 23201 21295 23259 21301
rect 25314 21292 25320 21304
rect 25372 21292 25378 21344
rect 25774 21292 25780 21344
rect 25832 21332 25838 21344
rect 26068 21332 26096 21363
rect 29822 21360 29828 21412
rect 29880 21360 29886 21412
rect 29914 21360 29920 21412
rect 29972 21360 29978 21412
rect 25832 21304 26096 21332
rect 28537 21335 28595 21341
rect 25832 21292 25838 21304
rect 28537 21301 28549 21335
rect 28583 21332 28595 21335
rect 28718 21332 28724 21344
rect 28583 21304 28724 21332
rect 28583 21301 28595 21304
rect 28537 21295 28595 21301
rect 28718 21292 28724 21304
rect 28776 21292 28782 21344
rect 29730 21292 29736 21344
rect 29788 21332 29794 21344
rect 30009 21335 30067 21341
rect 30009 21332 30021 21335
rect 29788 21304 30021 21332
rect 29788 21292 29794 21304
rect 30009 21301 30021 21304
rect 30055 21301 30067 21335
rect 30009 21295 30067 21301
rect 552 21242 31072 21264
rect 552 21190 7988 21242
rect 8040 21190 8052 21242
rect 8104 21190 8116 21242
rect 8168 21190 8180 21242
rect 8232 21190 8244 21242
rect 8296 21190 15578 21242
rect 15630 21190 15642 21242
rect 15694 21190 15706 21242
rect 15758 21190 15770 21242
rect 15822 21190 15834 21242
rect 15886 21190 23168 21242
rect 23220 21190 23232 21242
rect 23284 21190 23296 21242
rect 23348 21190 23360 21242
rect 23412 21190 23424 21242
rect 23476 21190 30758 21242
rect 30810 21190 30822 21242
rect 30874 21190 30886 21242
rect 30938 21190 30950 21242
rect 31002 21190 31014 21242
rect 31066 21190 31072 21242
rect 552 21168 31072 21190
rect 1394 21088 1400 21140
rect 1452 21137 1458 21140
rect 1452 21091 1461 21137
rect 3602 21128 3608 21140
rect 3660 21137 3666 21140
rect 3569 21100 3608 21128
rect 1452 21088 1458 21091
rect 3602 21088 3608 21100
rect 3660 21091 3669 21137
rect 3660 21088 3666 21091
rect 5810 21088 5816 21140
rect 5868 21128 5874 21140
rect 6279 21131 6337 21137
rect 6279 21128 6291 21131
rect 5868 21100 6291 21128
rect 5868 21088 5874 21100
rect 6279 21097 6291 21100
rect 6325 21097 6337 21131
rect 6279 21091 6337 21097
rect 6546 21088 6552 21140
rect 6604 21128 6610 21140
rect 9953 21131 10011 21137
rect 9953 21128 9965 21131
rect 6604 21100 9965 21128
rect 6604 21088 6610 21100
rect 9953 21097 9965 21100
rect 9999 21097 10011 21131
rect 9953 21091 10011 21097
rect 10226 21088 10232 21140
rect 10284 21088 10290 21140
rect 14277 21131 14335 21137
rect 14277 21097 14289 21131
rect 14323 21128 14335 21131
rect 14458 21128 14464 21140
rect 14323 21100 14464 21128
rect 14323 21097 14335 21100
rect 14277 21091 14335 21097
rect 14458 21088 14464 21100
rect 14516 21088 14522 21140
rect 14737 21131 14795 21137
rect 14737 21097 14749 21131
rect 14783 21128 14795 21131
rect 14826 21128 14832 21140
rect 14783 21100 14832 21128
rect 14783 21097 14795 21100
rect 14737 21091 14795 21097
rect 14826 21088 14832 21100
rect 14884 21088 14890 21140
rect 15197 21131 15255 21137
rect 15197 21097 15209 21131
rect 15243 21128 15255 21131
rect 15378 21128 15384 21140
rect 15243 21100 15384 21128
rect 15243 21097 15255 21100
rect 15197 21091 15255 21097
rect 15378 21088 15384 21100
rect 15436 21088 15442 21140
rect 15654 21088 15660 21140
rect 15712 21088 15718 21140
rect 16574 21088 16580 21140
rect 16632 21128 16638 21140
rect 16632 21100 17080 21128
rect 16632 21088 16638 21100
rect 5261 21063 5319 21069
rect 5261 21029 5273 21063
rect 5307 21060 5319 21063
rect 5307 21032 5948 21060
rect 5307 21029 5319 21032
rect 5261 21023 5319 21029
rect 1670 20952 1676 21004
rect 1728 20952 1734 21004
rect 5353 20995 5411 21001
rect 5353 20961 5365 20995
rect 5399 20992 5411 20995
rect 5442 20992 5448 21004
rect 5399 20964 5448 20992
rect 5399 20961 5411 20964
rect 5353 20955 5411 20961
rect 5442 20952 5448 20964
rect 5500 20952 5506 21004
rect 5534 20952 5540 21004
rect 5592 20992 5598 21004
rect 5813 20995 5871 21001
rect 5813 20992 5825 20995
rect 5592 20964 5825 20992
rect 5592 20952 5598 20964
rect 5813 20961 5825 20964
rect 5859 20961 5871 20995
rect 5920 20992 5948 21032
rect 8754 20992 8760 21004
rect 5920 20964 6132 20992
rect 5813 20955 5871 20961
rect 934 20884 940 20936
rect 992 20884 998 20936
rect 1443 20927 1501 20933
rect 1443 20893 1455 20927
rect 1489 20924 1501 20927
rect 1854 20924 1860 20936
rect 1489 20896 1860 20924
rect 1489 20893 1501 20896
rect 1443 20887 1501 20893
rect 1854 20884 1860 20896
rect 1912 20884 1918 20936
rect 3145 20927 3203 20933
rect 3145 20893 3157 20927
rect 3191 20924 3203 20927
rect 3326 20924 3332 20936
rect 3191 20896 3332 20924
rect 3191 20893 3203 20896
rect 3145 20887 3203 20893
rect 3326 20884 3332 20896
rect 3384 20884 3390 20936
rect 3602 20884 3608 20936
rect 3660 20884 3666 20936
rect 3881 20927 3939 20933
rect 3881 20893 3893 20927
rect 3927 20924 3939 20927
rect 6104 20924 6132 20964
rect 8496 20964 8760 20992
rect 6276 20927 6334 20933
rect 6276 20924 6288 20927
rect 3927 20896 5764 20924
rect 6104 20896 6288 20924
rect 3927 20893 3939 20896
rect 3881 20887 3939 20893
rect 2958 20748 2964 20800
rect 3016 20748 3022 20800
rect 5534 20748 5540 20800
rect 5592 20748 5598 20800
rect 5736 20788 5764 20896
rect 6276 20893 6288 20896
rect 6322 20893 6334 20927
rect 6276 20887 6334 20893
rect 6549 20927 6607 20933
rect 6549 20893 6561 20927
rect 6595 20924 6607 20927
rect 6730 20924 6736 20936
rect 6595 20896 6736 20924
rect 6595 20893 6607 20896
rect 6549 20887 6607 20893
rect 6730 20884 6736 20896
rect 6788 20884 6794 20936
rect 8113 20927 8171 20933
rect 8113 20893 8125 20927
rect 8159 20893 8171 20927
rect 8113 20887 8171 20893
rect 7650 20788 7656 20800
rect 5736 20760 7656 20788
rect 7650 20748 7656 20760
rect 7708 20748 7714 20800
rect 7834 20748 7840 20800
rect 7892 20748 7898 20800
rect 8136 20788 8164 20887
rect 8386 20884 8392 20936
rect 8444 20933 8450 20936
rect 8496 20933 8524 20964
rect 8754 20952 8760 20964
rect 8812 20952 8818 21004
rect 9122 20952 9128 21004
rect 9180 20992 9186 21004
rect 10244 20992 10272 21088
rect 10410 21020 10416 21072
rect 10468 21020 10474 21072
rect 17052 21060 17080 21100
rect 17126 21088 17132 21140
rect 17184 21088 17190 21140
rect 17862 21128 17868 21140
rect 17236 21100 17868 21128
rect 17236 21060 17264 21100
rect 17862 21088 17868 21100
rect 17920 21088 17926 21140
rect 18598 21088 18604 21140
rect 18656 21088 18662 21140
rect 19242 21088 19248 21140
rect 19300 21088 19306 21140
rect 20809 21131 20867 21137
rect 20809 21097 20821 21131
rect 20855 21128 20867 21131
rect 21358 21128 21364 21140
rect 20855 21100 21364 21128
rect 20855 21097 20867 21100
rect 20809 21091 20867 21097
rect 21358 21088 21364 21100
rect 21416 21088 21422 21140
rect 22278 21088 22284 21140
rect 22336 21128 22342 21140
rect 23109 21131 23167 21137
rect 23109 21128 23121 21131
rect 22336 21100 23121 21128
rect 22336 21088 22342 21100
rect 23109 21097 23121 21100
rect 23155 21097 23167 21131
rect 23109 21091 23167 21097
rect 23382 21088 23388 21140
rect 23440 21128 23446 21140
rect 24762 21128 24768 21140
rect 23440 21100 24768 21128
rect 23440 21088 23446 21100
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 25314 21088 25320 21140
rect 25372 21088 25378 21140
rect 25685 21131 25743 21137
rect 25685 21097 25697 21131
rect 25731 21128 25743 21131
rect 29914 21128 29920 21140
rect 25731 21100 29920 21128
rect 25731 21097 25743 21100
rect 25685 21091 25743 21097
rect 29914 21088 29920 21100
rect 29972 21088 29978 21140
rect 19260 21060 19288 21088
rect 25130 21060 25136 21072
rect 17052 21032 17264 21060
rect 9180 20964 10272 20992
rect 9180 20952 9186 20964
rect 10318 20952 10324 21004
rect 10376 20992 10382 21004
rect 11701 20995 11759 21001
rect 11701 20992 11713 20995
rect 10376 20964 11713 20992
rect 10376 20952 10382 20964
rect 11701 20961 11713 20964
rect 11747 20961 11759 20995
rect 11701 20955 11759 20961
rect 12618 20952 12624 21004
rect 12676 20992 12682 21004
rect 13265 20995 13323 21001
rect 13265 20992 13277 20995
rect 12676 20964 13277 20992
rect 12676 20952 12682 20964
rect 13265 20961 13277 20964
rect 13311 20961 13323 20995
rect 13265 20955 13323 20961
rect 16114 20952 16120 21004
rect 16172 20992 16178 21004
rect 16301 20995 16359 21001
rect 16301 20992 16313 20995
rect 16172 20964 16313 20992
rect 16172 20952 16178 20964
rect 16301 20961 16313 20964
rect 16347 20961 16359 20995
rect 16301 20955 16359 20961
rect 16666 20952 16672 21004
rect 16724 20952 16730 21004
rect 17037 20995 17095 21001
rect 17037 20961 17049 20995
rect 17083 20992 17095 20995
rect 17236 20992 17264 21032
rect 18984 21032 19288 21060
rect 24978 21032 25136 21060
rect 17083 20964 17264 20992
rect 17083 20961 17095 20964
rect 17037 20955 17095 20961
rect 17494 20952 17500 21004
rect 17552 20952 17558 21004
rect 18984 20992 19012 21032
rect 25130 21020 25136 21032
rect 25188 21020 25194 21072
rect 26050 21020 26056 21072
rect 26108 21020 26114 21072
rect 20714 20992 20720 21004
rect 18892 20964 19012 20992
rect 20378 20964 20720 20992
rect 8662 20933 8668 20936
rect 8444 20927 8524 20933
rect 8444 20893 8452 20927
rect 8486 20896 8524 20927
rect 8619 20927 8668 20933
rect 8486 20893 8498 20896
rect 8444 20887 8498 20893
rect 8619 20893 8631 20927
rect 8665 20893 8668 20927
rect 8619 20887 8668 20893
rect 8444 20884 8450 20887
rect 8662 20884 8668 20887
rect 8720 20884 8726 20936
rect 8849 20927 8907 20933
rect 8849 20893 8861 20927
rect 8895 20924 8907 20927
rect 8938 20924 8944 20936
rect 8895 20896 8944 20924
rect 8895 20893 8907 20896
rect 8849 20887 8907 20893
rect 8938 20884 8944 20896
rect 8996 20884 9002 20936
rect 9030 20884 9036 20936
rect 9088 20924 9094 20936
rect 10965 20927 11023 20933
rect 10965 20924 10977 20927
rect 9088 20896 10977 20924
rect 9088 20884 9094 20896
rect 10965 20893 10977 20896
rect 11011 20893 11023 20927
rect 10965 20887 11023 20893
rect 11146 20884 11152 20936
rect 11204 20924 11210 20936
rect 11292 20927 11350 20933
rect 11292 20924 11304 20927
rect 11204 20896 11304 20924
rect 11204 20884 11210 20896
rect 11292 20893 11304 20896
rect 11338 20893 11350 20927
rect 11292 20887 11350 20893
rect 11422 20884 11428 20936
rect 11480 20884 11486 20936
rect 17221 20927 17279 20933
rect 17221 20893 17233 20927
rect 17267 20924 17279 20927
rect 18892 20924 18920 20964
rect 20714 20952 20720 20964
rect 20772 20952 20778 21004
rect 20993 20995 21051 21001
rect 20993 20961 21005 20995
rect 21039 20961 21051 20995
rect 23106 20992 23112 21004
rect 22678 20964 23112 20992
rect 20993 20955 21051 20961
rect 17267 20896 18920 20924
rect 18969 20927 19027 20933
rect 17267 20893 17279 20896
rect 17221 20887 17279 20893
rect 18969 20893 18981 20927
rect 19015 20893 19027 20927
rect 18969 20887 19027 20893
rect 19245 20927 19303 20933
rect 19245 20893 19257 20927
rect 19291 20924 19303 20927
rect 19702 20924 19708 20936
rect 19291 20896 19708 20924
rect 19291 20893 19303 20896
rect 19245 20887 19303 20893
rect 8478 20788 8484 20800
rect 8136 20760 8484 20788
rect 8478 20748 8484 20760
rect 8536 20788 8542 20800
rect 9582 20788 9588 20800
rect 8536 20760 9588 20788
rect 8536 20748 8542 20760
rect 9582 20748 9588 20760
rect 9640 20788 9646 20800
rect 10505 20791 10563 20797
rect 10505 20788 10517 20791
rect 9640 20760 10517 20788
rect 9640 20748 9646 20760
rect 10505 20757 10517 20760
rect 10551 20757 10563 20791
rect 10505 20751 10563 20757
rect 10778 20748 10784 20800
rect 10836 20788 10842 20800
rect 11422 20788 11428 20800
rect 10836 20760 11428 20788
rect 10836 20748 10842 20760
rect 11422 20748 11428 20760
rect 11480 20748 11486 20800
rect 12710 20748 12716 20800
rect 12768 20788 12774 20800
rect 12805 20791 12863 20797
rect 12805 20788 12817 20791
rect 12768 20760 12817 20788
rect 12768 20748 12774 20760
rect 12805 20757 12817 20760
rect 12851 20757 12863 20791
rect 12805 20751 12863 20757
rect 13170 20748 13176 20800
rect 13228 20788 13234 20800
rect 13357 20791 13415 20797
rect 13357 20788 13369 20791
rect 13228 20760 13369 20788
rect 13228 20748 13234 20760
rect 13357 20757 13369 20760
rect 13403 20757 13415 20791
rect 18984 20788 19012 20887
rect 19702 20884 19708 20896
rect 19760 20924 19766 20936
rect 21008 20924 21036 20955
rect 23106 20952 23112 20964
rect 23164 20952 23170 21004
rect 23293 20995 23351 21001
rect 23293 20961 23305 20995
rect 23339 20961 23351 20995
rect 23293 20955 23351 20961
rect 25501 20995 25559 21001
rect 25501 20961 25513 20995
rect 25547 20961 25559 20995
rect 25501 20955 25559 20961
rect 19760 20896 21036 20924
rect 19760 20884 19766 20896
rect 21266 20884 21272 20936
rect 21324 20884 21330 20936
rect 21545 20927 21603 20933
rect 21545 20893 21557 20927
rect 21591 20924 21603 20927
rect 23308 20924 23336 20955
rect 23477 20927 23535 20933
rect 23477 20924 23489 20927
rect 21591 20896 23489 20924
rect 21591 20893 21603 20896
rect 21545 20887 21603 20893
rect 23477 20893 23489 20896
rect 23523 20893 23535 20927
rect 23753 20927 23811 20933
rect 23753 20924 23765 20927
rect 23477 20887 23535 20893
rect 23584 20896 23765 20924
rect 21726 20788 21732 20800
rect 18984 20760 21732 20788
rect 13357 20751 13415 20757
rect 21726 20748 21732 20760
rect 21784 20748 21790 20800
rect 22186 20748 22192 20800
rect 22244 20788 22250 20800
rect 23584 20788 23612 20896
rect 23753 20893 23765 20896
rect 23799 20924 23811 20927
rect 25516 20924 25544 20955
rect 25590 20952 25596 21004
rect 25648 20992 25654 21004
rect 25869 20995 25927 21001
rect 25869 20992 25881 20995
rect 25648 20964 25881 20992
rect 25648 20952 25654 20964
rect 25869 20961 25881 20964
rect 25915 20961 25927 20995
rect 25869 20955 25927 20961
rect 26142 20952 26148 21004
rect 26200 20952 26206 21004
rect 26970 20952 26976 21004
rect 27028 20992 27034 21004
rect 28680 20995 28738 21001
rect 28680 20992 28692 20995
rect 27028 20964 28692 20992
rect 27028 20952 27034 20964
rect 28680 20961 28692 20964
rect 28726 20961 28738 20995
rect 28680 20955 28738 20961
rect 23799 20896 25544 20924
rect 23799 20893 23811 20896
rect 23753 20887 23811 20893
rect 26234 20884 26240 20936
rect 26292 20924 26298 20936
rect 26421 20927 26479 20933
rect 26421 20924 26433 20927
rect 26292 20896 26433 20924
rect 26292 20884 26298 20896
rect 26421 20893 26433 20896
rect 26467 20893 26479 20927
rect 26421 20887 26479 20893
rect 26697 20927 26755 20933
rect 26697 20893 26709 20927
rect 26743 20924 26755 20927
rect 27430 20924 27436 20936
rect 26743 20896 27436 20924
rect 26743 20893 26755 20896
rect 26697 20887 26755 20893
rect 27430 20884 27436 20896
rect 27488 20884 27494 20936
rect 27522 20884 27528 20936
rect 27580 20924 27586 20936
rect 28353 20927 28411 20933
rect 28353 20924 28365 20927
rect 27580 20896 28365 20924
rect 27580 20884 27586 20896
rect 28353 20893 28365 20896
rect 28399 20893 28411 20927
rect 28353 20887 28411 20893
rect 28859 20927 28917 20933
rect 28859 20893 28871 20927
rect 28905 20924 28917 20927
rect 28994 20924 29000 20936
rect 28905 20896 29000 20924
rect 28905 20893 28917 20896
rect 28859 20887 28917 20893
rect 28994 20884 29000 20896
rect 29052 20884 29058 20936
rect 29089 20927 29147 20933
rect 29089 20893 29101 20927
rect 29135 20924 29147 20927
rect 29822 20924 29828 20936
rect 29135 20896 29828 20924
rect 29135 20893 29147 20896
rect 29089 20887 29147 20893
rect 29822 20884 29828 20896
rect 29880 20884 29886 20936
rect 22244 20760 23612 20788
rect 27985 20791 28043 20797
rect 22244 20748 22250 20760
rect 27985 20757 27997 20791
rect 28031 20788 28043 20791
rect 28258 20788 28264 20800
rect 28031 20760 28264 20788
rect 28031 20757 28043 20760
rect 27985 20751 28043 20757
rect 28258 20748 28264 20760
rect 28316 20748 28322 20800
rect 28534 20748 28540 20800
rect 28592 20788 28598 20800
rect 30193 20791 30251 20797
rect 30193 20788 30205 20791
rect 28592 20760 30205 20788
rect 28592 20748 28598 20760
rect 30193 20757 30205 20760
rect 30239 20757 30251 20791
rect 30193 20751 30251 20757
rect 552 20698 30912 20720
rect 552 20646 4193 20698
rect 4245 20646 4257 20698
rect 4309 20646 4321 20698
rect 4373 20646 4385 20698
rect 4437 20646 4449 20698
rect 4501 20646 11783 20698
rect 11835 20646 11847 20698
rect 11899 20646 11911 20698
rect 11963 20646 11975 20698
rect 12027 20646 12039 20698
rect 12091 20646 19373 20698
rect 19425 20646 19437 20698
rect 19489 20646 19501 20698
rect 19553 20646 19565 20698
rect 19617 20646 19629 20698
rect 19681 20646 26963 20698
rect 27015 20646 27027 20698
rect 27079 20646 27091 20698
rect 27143 20646 27155 20698
rect 27207 20646 27219 20698
rect 27271 20646 30912 20698
rect 552 20624 30912 20646
rect 2961 20587 3019 20593
rect 952 20556 2774 20584
rect 842 20340 848 20392
rect 900 20380 906 20392
rect 952 20389 980 20556
rect 1302 20457 1308 20460
rect 1264 20451 1308 20457
rect 1264 20417 1276 20451
rect 1264 20411 1308 20417
rect 1302 20408 1308 20411
rect 1360 20408 1366 20460
rect 1578 20448 1584 20460
rect 1418 20433 1584 20448
rect 1418 20402 1445 20433
rect 1433 20399 1445 20402
rect 1479 20420 1584 20433
rect 1479 20399 1491 20420
rect 1578 20408 1584 20420
rect 1636 20408 1642 20460
rect 1670 20408 1676 20460
rect 1728 20408 1734 20460
rect 1433 20393 1491 20399
rect 937 20383 995 20389
rect 937 20380 949 20383
rect 900 20352 949 20380
rect 900 20340 906 20352
rect 937 20349 949 20352
rect 983 20349 995 20383
rect 2746 20380 2774 20556
rect 2961 20553 2973 20587
rect 3007 20584 3019 20587
rect 3602 20584 3608 20596
rect 3007 20556 3608 20584
rect 3007 20553 3019 20556
rect 2961 20547 3019 20553
rect 3602 20544 3608 20556
rect 3660 20544 3666 20596
rect 4706 20544 4712 20596
rect 4764 20584 4770 20596
rect 7929 20587 7987 20593
rect 7929 20584 7941 20587
rect 4764 20556 7941 20584
rect 4764 20544 4770 20556
rect 7929 20553 7941 20556
rect 7975 20553 7987 20587
rect 9122 20584 9128 20596
rect 7929 20547 7987 20553
rect 8036 20556 9128 20584
rect 4387 20451 4445 20457
rect 4387 20417 4399 20451
rect 4433 20448 4445 20451
rect 6270 20448 6276 20460
rect 4433 20420 6276 20448
rect 4433 20417 4445 20420
rect 4387 20411 4445 20417
rect 6270 20408 6276 20420
rect 6328 20408 6334 20460
rect 6638 20457 6644 20460
rect 6595 20451 6644 20457
rect 6595 20417 6607 20451
rect 6641 20417 6644 20451
rect 6595 20411 6644 20417
rect 6638 20408 6644 20411
rect 6696 20408 6702 20460
rect 6730 20408 6736 20460
rect 6788 20448 6794 20460
rect 8036 20448 8064 20556
rect 9122 20544 9128 20556
rect 9180 20544 9186 20596
rect 12986 20584 12992 20596
rect 10796 20556 12992 20584
rect 6788 20420 8064 20448
rect 8987 20451 9045 20457
rect 6788 20408 6794 20420
rect 8987 20417 8999 20451
rect 9033 20448 9045 20451
rect 10226 20448 10232 20460
rect 9033 20420 10232 20448
rect 9033 20417 9045 20420
rect 8987 20411 9045 20417
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 3329 20383 3387 20389
rect 3329 20380 3341 20383
rect 2746 20352 3341 20380
rect 937 20343 995 20349
rect 3329 20349 3341 20352
rect 3375 20380 3387 20383
rect 3418 20380 3424 20392
rect 3375 20352 3424 20380
rect 3375 20349 3387 20352
rect 3329 20343 3387 20349
rect 3418 20340 3424 20352
rect 3476 20340 3482 20392
rect 3881 20383 3939 20389
rect 3881 20349 3893 20383
rect 3927 20380 3939 20383
rect 4522 20380 4528 20392
rect 3927 20352 4528 20380
rect 3927 20349 3939 20352
rect 3881 20343 3939 20349
rect 4522 20340 4528 20352
rect 4580 20340 4586 20392
rect 4617 20383 4675 20389
rect 4617 20349 4629 20383
rect 4663 20380 4675 20383
rect 4890 20380 4896 20392
rect 4663 20352 4896 20380
rect 4663 20349 4675 20352
rect 4617 20343 4675 20349
rect 4890 20340 4896 20352
rect 4948 20340 4954 20392
rect 5718 20340 5724 20392
rect 5776 20380 5782 20392
rect 6089 20383 6147 20389
rect 6089 20380 6101 20383
rect 5776 20352 6101 20380
rect 5776 20340 5782 20352
rect 6089 20349 6101 20352
rect 6135 20349 6147 20383
rect 6089 20343 6147 20349
rect 6178 20340 6184 20392
rect 6236 20380 6242 20392
rect 6416 20383 6474 20389
rect 6416 20380 6428 20383
rect 6236 20352 6428 20380
rect 6236 20340 6242 20352
rect 6416 20349 6428 20352
rect 6462 20349 6474 20383
rect 6416 20343 6474 20349
rect 6825 20383 6883 20389
rect 6825 20349 6837 20383
rect 6871 20380 6883 20383
rect 6914 20380 6920 20392
rect 6871 20352 6920 20380
rect 6871 20349 6883 20352
rect 6825 20343 6883 20349
rect 6914 20340 6920 20352
rect 6972 20340 6978 20392
rect 7558 20340 7564 20392
rect 7616 20380 7622 20392
rect 8481 20383 8539 20389
rect 8481 20380 8493 20383
rect 7616 20352 8493 20380
rect 7616 20340 7622 20352
rect 8481 20349 8493 20352
rect 8527 20380 8539 20383
rect 8754 20380 8760 20392
rect 8527 20352 8760 20380
rect 8527 20349 8539 20352
rect 8481 20343 8539 20349
rect 8754 20340 8760 20352
rect 8812 20340 8818 20392
rect 9217 20383 9275 20389
rect 9217 20349 9229 20383
rect 9263 20380 9275 20383
rect 10686 20380 10692 20392
rect 9263 20352 10692 20380
rect 9263 20349 9275 20352
rect 9217 20343 9275 20349
rect 10686 20340 10692 20352
rect 10744 20340 10750 20392
rect 10796 20389 10824 20556
rect 12986 20544 12992 20556
rect 13044 20544 13050 20596
rect 13998 20544 14004 20596
rect 14056 20584 14062 20596
rect 16025 20587 16083 20593
rect 16025 20584 16037 20587
rect 14056 20556 16037 20584
rect 14056 20544 14062 20556
rect 16025 20553 16037 20556
rect 16071 20553 16083 20587
rect 16025 20547 16083 20553
rect 19061 20587 19119 20593
rect 19061 20553 19073 20587
rect 19107 20584 19119 20587
rect 21910 20584 21916 20596
rect 19107 20556 21916 20584
rect 19107 20553 19119 20556
rect 19061 20547 19119 20553
rect 21910 20544 21916 20556
rect 21968 20544 21974 20596
rect 23842 20544 23848 20596
rect 23900 20584 23906 20596
rect 25774 20584 25780 20596
rect 23900 20556 25780 20584
rect 23900 20544 23906 20556
rect 25774 20544 25780 20556
rect 25832 20544 25838 20596
rect 27522 20584 27528 20596
rect 26712 20556 27528 20584
rect 10870 20476 10876 20528
rect 10928 20516 10934 20528
rect 11057 20519 11115 20525
rect 11057 20516 11069 20519
rect 10928 20488 11069 20516
rect 10928 20476 10934 20488
rect 11057 20485 11069 20488
rect 11103 20485 11115 20519
rect 11057 20479 11115 20485
rect 20714 20476 20720 20528
rect 20772 20516 20778 20528
rect 21358 20516 21364 20528
rect 20772 20488 21364 20516
rect 20772 20476 20778 20488
rect 21358 20476 21364 20488
rect 21416 20476 21422 20528
rect 11704 20451 11762 20457
rect 11704 20448 11716 20451
rect 10888 20420 11716 20448
rect 10888 20392 10916 20420
rect 11704 20417 11716 20420
rect 11750 20417 11762 20451
rect 11704 20411 11762 20417
rect 14093 20451 14151 20457
rect 14093 20417 14105 20451
rect 14139 20448 14151 20451
rect 14182 20448 14188 20460
rect 14139 20420 14188 20448
rect 14139 20417 14151 20420
rect 14093 20411 14151 20417
rect 14182 20408 14188 20420
rect 14240 20448 14246 20460
rect 16117 20451 16175 20457
rect 16117 20448 16129 20451
rect 14240 20420 16129 20448
rect 14240 20408 14246 20420
rect 16117 20417 16129 20420
rect 16163 20417 16175 20451
rect 16117 20411 16175 20417
rect 18690 20408 18696 20460
rect 18748 20408 18754 20460
rect 19337 20451 19395 20457
rect 19337 20417 19349 20451
rect 19383 20448 19395 20451
rect 19702 20448 19708 20460
rect 19383 20420 19708 20448
rect 19383 20417 19395 20420
rect 19337 20411 19395 20417
rect 19702 20408 19708 20420
rect 19760 20408 19766 20460
rect 19978 20408 19984 20460
rect 20036 20448 20042 20460
rect 20732 20448 20760 20476
rect 26712 20460 26740 20556
rect 27522 20544 27528 20556
rect 27580 20544 27586 20596
rect 28166 20544 28172 20596
rect 28224 20584 28230 20596
rect 28350 20584 28356 20596
rect 28224 20556 28356 20584
rect 28224 20544 28230 20556
rect 28350 20544 28356 20556
rect 28408 20584 28414 20596
rect 30193 20587 30251 20593
rect 30193 20584 30205 20587
rect 28408 20556 30205 20584
rect 28408 20544 28414 20556
rect 30193 20553 30205 20556
rect 30239 20553 30251 20587
rect 30193 20547 30251 20553
rect 28902 20476 28908 20528
rect 28960 20516 28966 20528
rect 29454 20516 29460 20528
rect 28960 20488 29460 20516
rect 28960 20476 28966 20488
rect 29454 20476 29460 20488
rect 29512 20476 29518 20528
rect 20036 20420 20760 20448
rect 20036 20408 20042 20420
rect 10781 20383 10839 20389
rect 10781 20349 10793 20383
rect 10827 20349 10839 20383
rect 10781 20343 10839 20349
rect 10870 20340 10876 20392
rect 10928 20340 10934 20392
rect 11238 20340 11244 20392
rect 11296 20340 11302 20392
rect 11977 20383 12035 20389
rect 11977 20380 11989 20383
rect 11348 20352 11989 20380
rect 3694 20272 3700 20324
rect 3752 20272 3758 20324
rect 10597 20315 10655 20321
rect 10597 20281 10609 20315
rect 10643 20312 10655 20315
rect 11054 20312 11060 20324
rect 10643 20284 11060 20312
rect 10643 20281 10655 20284
rect 10597 20275 10655 20281
rect 11054 20272 11060 20284
rect 11112 20272 11118 20324
rect 4347 20247 4405 20253
rect 4347 20213 4359 20247
rect 4393 20244 4405 20247
rect 5810 20244 5816 20256
rect 4393 20216 5816 20244
rect 4393 20213 4405 20216
rect 4347 20207 4405 20213
rect 5810 20204 5816 20216
rect 5868 20204 5874 20256
rect 5905 20247 5963 20253
rect 5905 20213 5917 20247
rect 5951 20244 5963 20247
rect 7282 20244 7288 20256
rect 5951 20216 7288 20244
rect 5951 20213 5963 20216
rect 5905 20207 5963 20213
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 7466 20204 7472 20256
rect 7524 20244 7530 20256
rect 8947 20247 9005 20253
rect 8947 20244 8959 20247
rect 7524 20216 8959 20244
rect 7524 20204 7530 20216
rect 8947 20213 8959 20216
rect 8993 20244 9005 20247
rect 9122 20244 9128 20256
rect 8993 20216 9128 20244
rect 8993 20213 9005 20216
rect 8947 20207 9005 20213
rect 9122 20204 9128 20216
rect 9180 20204 9186 20256
rect 10502 20204 10508 20256
rect 10560 20244 10566 20256
rect 11348 20244 11376 20352
rect 11977 20349 11989 20352
rect 12023 20349 12035 20383
rect 11977 20343 12035 20349
rect 12066 20340 12072 20392
rect 12124 20380 12130 20392
rect 14277 20383 14335 20389
rect 14277 20380 14289 20383
rect 12124 20352 14289 20380
rect 12124 20340 12130 20352
rect 14277 20349 14289 20352
rect 14323 20349 14335 20383
rect 14277 20343 14335 20349
rect 16393 20383 16451 20389
rect 16393 20349 16405 20383
rect 16439 20380 16451 20383
rect 16666 20380 16672 20392
rect 16439 20352 16672 20380
rect 16439 20349 16451 20352
rect 16393 20343 16451 20349
rect 13817 20315 13875 20321
rect 13817 20281 13829 20315
rect 13863 20312 13875 20315
rect 13998 20312 14004 20324
rect 13863 20284 14004 20312
rect 13863 20281 13875 20284
rect 13817 20275 13875 20281
rect 13998 20272 14004 20284
rect 14056 20272 14062 20324
rect 14292 20312 14320 20343
rect 16666 20340 16672 20352
rect 16724 20340 16730 20392
rect 17957 20383 18015 20389
rect 17957 20349 17969 20383
rect 18003 20380 18015 20383
rect 18046 20380 18052 20392
rect 18003 20352 18052 20380
rect 18003 20349 18015 20352
rect 17957 20343 18015 20349
rect 18046 20340 18052 20352
rect 18104 20340 18110 20392
rect 18874 20340 18880 20392
rect 18932 20340 18938 20392
rect 20732 20366 20760 20420
rect 21821 20451 21879 20457
rect 21821 20417 21833 20451
rect 21867 20448 21879 20451
rect 24121 20451 24179 20457
rect 21867 20420 23612 20448
rect 21867 20417 21879 20420
rect 21821 20411 21879 20417
rect 21266 20380 21272 20392
rect 20916 20352 21272 20380
rect 14553 20315 14611 20321
rect 14292 20284 14504 20312
rect 14476 20256 14504 20284
rect 14553 20281 14565 20315
rect 14599 20312 14611 20315
rect 14826 20312 14832 20324
rect 14599 20284 14832 20312
rect 14599 20281 14611 20284
rect 14553 20275 14611 20281
rect 14826 20272 14832 20284
rect 14884 20272 14890 20324
rect 16114 20312 16120 20324
rect 15778 20284 16120 20312
rect 10560 20216 11376 20244
rect 10560 20204 10566 20216
rect 11606 20204 11612 20256
rect 11664 20244 11670 20256
rect 11707 20247 11765 20253
rect 11707 20244 11719 20247
rect 11664 20216 11719 20244
rect 11664 20204 11670 20216
rect 11707 20213 11719 20216
rect 11753 20213 11765 20247
rect 11707 20207 11765 20213
rect 13078 20204 13084 20256
rect 13136 20204 13142 20256
rect 14458 20204 14464 20256
rect 14516 20204 14522 20256
rect 15378 20204 15384 20256
rect 15436 20244 15442 20256
rect 15856 20244 15884 20284
rect 16114 20272 16120 20284
rect 16172 20272 16178 20324
rect 19613 20315 19671 20321
rect 19613 20281 19625 20315
rect 19659 20281 19671 20315
rect 19613 20275 19671 20281
rect 15436 20216 15884 20244
rect 15436 20204 15442 20216
rect 17494 20204 17500 20256
rect 17552 20204 17558 20256
rect 17862 20204 17868 20256
rect 17920 20244 17926 20256
rect 18049 20247 18107 20253
rect 18049 20244 18061 20247
rect 17920 20216 18061 20244
rect 17920 20204 17926 20216
rect 18049 20213 18061 20216
rect 18095 20213 18107 20247
rect 19628 20244 19656 20275
rect 20916 20244 20944 20352
rect 21266 20340 21272 20352
rect 21324 20380 21330 20392
rect 21361 20383 21419 20389
rect 21361 20380 21373 20383
rect 21324 20352 21373 20380
rect 21324 20340 21330 20352
rect 21361 20349 21373 20352
rect 21407 20349 21419 20383
rect 21361 20343 21419 20349
rect 21542 20340 21548 20392
rect 21600 20340 21606 20392
rect 23382 20389 23388 20392
rect 23364 20383 23388 20389
rect 23364 20349 23376 20383
rect 23364 20343 23388 20349
rect 23382 20340 23388 20343
rect 23440 20340 23446 20392
rect 23584 20389 23612 20420
rect 24121 20417 24133 20451
rect 24167 20448 24179 20451
rect 24167 20420 25912 20448
rect 24167 20417 24179 20420
rect 24121 20411 24179 20417
rect 23569 20383 23627 20389
rect 23569 20349 23581 20383
rect 23615 20380 23627 20383
rect 23845 20383 23903 20389
rect 23845 20380 23857 20383
rect 23615 20352 23857 20380
rect 23615 20349 23627 20352
rect 23569 20343 23627 20349
rect 23845 20349 23857 20352
rect 23891 20349 23903 20383
rect 23845 20343 23903 20349
rect 25130 20340 25136 20392
rect 25188 20380 25194 20392
rect 25884 20389 25912 20420
rect 26694 20408 26700 20460
rect 26752 20408 26758 20460
rect 26878 20408 26884 20460
rect 26936 20448 26942 20460
rect 27024 20451 27082 20457
rect 27024 20448 27036 20451
rect 26936 20420 27036 20448
rect 26936 20408 26942 20420
rect 27024 20417 27036 20420
rect 27070 20417 27082 20451
rect 27024 20411 27082 20417
rect 27203 20451 27261 20457
rect 27203 20417 27215 20451
rect 27249 20448 27261 20451
rect 27249 20420 29316 20448
rect 27249 20417 27261 20420
rect 27203 20411 27261 20417
rect 29288 20392 29316 20420
rect 25869 20383 25927 20389
rect 25188 20352 25254 20380
rect 25188 20340 25194 20352
rect 25869 20349 25881 20383
rect 25915 20349 25927 20383
rect 25869 20343 25927 20349
rect 27433 20383 27491 20389
rect 27433 20349 27445 20383
rect 27479 20380 27491 20383
rect 27479 20352 29040 20380
rect 27479 20349 27491 20352
rect 27433 20343 27491 20349
rect 22094 20312 22100 20324
rect 21192 20284 22100 20312
rect 21192 20253 21220 20284
rect 22094 20272 22100 20284
rect 22152 20272 22158 20324
rect 23106 20312 23112 20324
rect 23046 20284 23112 20312
rect 23106 20272 23112 20284
rect 23164 20312 23170 20324
rect 23750 20312 23756 20324
rect 23164 20284 23756 20312
rect 23164 20272 23170 20284
rect 23750 20272 23756 20284
rect 23808 20272 23814 20324
rect 26145 20315 26203 20321
rect 26145 20312 26157 20315
rect 25424 20284 26157 20312
rect 19628 20216 20944 20244
rect 21177 20247 21235 20253
rect 18049 20207 18107 20213
rect 21177 20213 21189 20247
rect 21223 20213 21235 20247
rect 21177 20207 21235 20213
rect 21358 20204 21364 20256
rect 21416 20244 21422 20256
rect 23124 20244 23152 20272
rect 21416 20216 23152 20244
rect 21416 20204 21422 20216
rect 24762 20204 24768 20256
rect 24820 20244 24826 20256
rect 25424 20244 25452 20284
rect 26145 20281 26157 20284
rect 26191 20281 26203 20315
rect 26145 20275 26203 20281
rect 24820 20216 25452 20244
rect 24820 20204 24826 20216
rect 25682 20204 25688 20256
rect 25740 20204 25746 20256
rect 26237 20247 26295 20253
rect 26237 20213 26249 20247
rect 26283 20244 26295 20247
rect 26326 20244 26332 20256
rect 26283 20216 26332 20244
rect 26283 20213 26295 20216
rect 26237 20207 26295 20213
rect 26326 20204 26332 20216
rect 26384 20204 26390 20256
rect 27522 20204 27528 20256
rect 27580 20244 27586 20256
rect 28537 20247 28595 20253
rect 28537 20244 28549 20247
rect 27580 20216 28549 20244
rect 27580 20204 27586 20216
rect 28537 20213 28549 20216
rect 28583 20213 28595 20247
rect 29012 20244 29040 20352
rect 29270 20340 29276 20392
rect 29328 20340 29334 20392
rect 29454 20340 29460 20392
rect 29512 20340 29518 20392
rect 29825 20383 29883 20389
rect 29825 20349 29837 20383
rect 29871 20380 29883 20383
rect 29914 20380 29920 20392
rect 29871 20352 29920 20380
rect 29871 20349 29883 20352
rect 29825 20343 29883 20349
rect 29914 20340 29920 20352
rect 29972 20340 29978 20392
rect 29086 20272 29092 20324
rect 29144 20272 29150 20324
rect 30098 20272 30104 20324
rect 30156 20272 30162 20324
rect 29454 20244 29460 20256
rect 29012 20216 29460 20244
rect 28537 20207 28595 20213
rect 29454 20204 29460 20216
rect 29512 20204 29518 20256
rect 29546 20204 29552 20256
rect 29604 20244 29610 20256
rect 29917 20247 29975 20253
rect 29917 20244 29929 20247
rect 29604 20216 29929 20244
rect 29604 20204 29610 20216
rect 29917 20213 29929 20216
rect 29963 20213 29975 20247
rect 29917 20207 29975 20213
rect 552 20154 31072 20176
rect 552 20102 7988 20154
rect 8040 20102 8052 20154
rect 8104 20102 8116 20154
rect 8168 20102 8180 20154
rect 8232 20102 8244 20154
rect 8296 20102 15578 20154
rect 15630 20102 15642 20154
rect 15694 20102 15706 20154
rect 15758 20102 15770 20154
rect 15822 20102 15834 20154
rect 15886 20102 23168 20154
rect 23220 20102 23232 20154
rect 23284 20102 23296 20154
rect 23348 20102 23360 20154
rect 23412 20102 23424 20154
rect 23476 20102 30758 20154
rect 30810 20102 30822 20154
rect 30874 20102 30886 20154
rect 30938 20102 30950 20154
rect 31002 20102 31014 20154
rect 31066 20102 31072 20154
rect 552 20080 31072 20102
rect 1302 20000 1308 20052
rect 1360 20040 1366 20052
rect 1403 20043 1461 20049
rect 1403 20040 1415 20043
rect 1360 20012 1415 20040
rect 1360 20000 1366 20012
rect 1403 20009 1415 20012
rect 1449 20040 1461 20043
rect 1762 20040 1768 20052
rect 1449 20012 1768 20040
rect 1449 20009 1461 20012
rect 1403 20003 1461 20009
rect 1762 20000 1768 20012
rect 1820 20000 1826 20052
rect 2961 20043 3019 20049
rect 2961 20009 2973 20043
rect 3007 20040 3019 20043
rect 4062 20040 4068 20052
rect 3007 20012 4068 20040
rect 3007 20009 3019 20012
rect 2961 20003 3019 20009
rect 4062 20000 4068 20012
rect 4120 20000 4126 20052
rect 5810 20000 5816 20052
rect 5868 20040 5874 20052
rect 6279 20043 6337 20049
rect 6279 20040 6291 20043
rect 5868 20012 6291 20040
rect 5868 20000 5874 20012
rect 6279 20009 6291 20012
rect 6325 20040 6337 20043
rect 7466 20040 7472 20052
rect 6325 20012 7472 20040
rect 6325 20009 6337 20012
rect 6279 20003 6337 20009
rect 7466 20000 7472 20012
rect 7524 20000 7530 20052
rect 13078 20040 13084 20052
rect 8128 20012 13084 20040
rect 5902 19972 5908 19984
rect 4908 19944 5908 19972
rect 3142 19904 3148 19916
rect 1596 19876 3148 19904
rect 1433 19857 1491 19863
rect 1433 19854 1445 19857
rect 842 19796 848 19848
rect 900 19836 906 19848
rect 937 19839 995 19845
rect 937 19836 949 19839
rect 900 19808 949 19836
rect 900 19796 906 19808
rect 937 19805 949 19808
rect 983 19805 995 19839
rect 1418 19823 1445 19854
rect 1479 19836 1491 19857
rect 1596 19836 1624 19876
rect 3142 19864 3148 19876
rect 3200 19864 3206 19916
rect 3421 19907 3479 19913
rect 3421 19873 3433 19907
rect 3467 19904 3479 19907
rect 3602 19904 3608 19916
rect 3467 19876 3608 19904
rect 3467 19873 3479 19876
rect 3421 19867 3479 19873
rect 3602 19864 3608 19876
rect 3660 19864 3666 19916
rect 3878 19913 3884 19916
rect 3840 19907 3884 19913
rect 3840 19873 3852 19907
rect 3936 19904 3942 19916
rect 4908 19904 4936 19944
rect 5902 19932 5908 19944
rect 5960 19932 5966 19984
rect 8128 19913 8156 20012
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 17494 20000 17500 20052
rect 17552 20000 17558 20052
rect 18874 20000 18880 20052
rect 18932 20040 18938 20052
rect 21266 20040 21272 20052
rect 18932 20012 21272 20040
rect 18932 20000 18938 20012
rect 21266 20000 21272 20012
rect 21324 20000 21330 20052
rect 21818 20000 21824 20052
rect 21876 20000 21882 20052
rect 23934 20000 23940 20052
rect 23992 20040 23998 20052
rect 24029 20043 24087 20049
rect 24029 20040 24041 20043
rect 23992 20012 24041 20040
rect 23992 20000 23998 20012
rect 24029 20009 24041 20012
rect 24075 20009 24087 20043
rect 25130 20040 25136 20052
rect 24029 20003 24087 20009
rect 24136 20012 25136 20040
rect 8386 19932 8392 19984
rect 8444 19932 8450 19984
rect 10594 19932 10600 19984
rect 10652 19932 10658 19984
rect 12066 19972 12072 19984
rect 11532 19944 12072 19972
rect 3936 19876 4936 19904
rect 5629 19907 5687 19913
rect 3840 19867 3884 19873
rect 3878 19864 3884 19867
rect 3936 19864 3942 19876
rect 5629 19873 5641 19907
rect 5675 19904 5687 19907
rect 8113 19907 8171 19913
rect 5675 19876 6224 19904
rect 5675 19873 5687 19876
rect 5629 19867 5687 19873
rect 1479 19823 1624 19836
rect 1418 19808 1624 19823
rect 937 19799 995 19805
rect 1670 19796 1676 19848
rect 1728 19796 1734 19848
rect 3326 19796 3332 19848
rect 3384 19836 3390 19848
rect 4062 19845 4068 19848
rect 3513 19839 3571 19845
rect 3513 19836 3525 19839
rect 3384 19808 3525 19836
rect 3384 19796 3390 19808
rect 3513 19805 3525 19808
rect 3559 19805 3571 19839
rect 3513 19799 3571 19805
rect 4019 19839 4068 19845
rect 4019 19805 4031 19839
rect 4065 19805 4068 19839
rect 4019 19799 4068 19805
rect 4062 19796 4068 19799
rect 4120 19796 4126 19848
rect 4249 19839 4307 19845
rect 4249 19805 4261 19839
rect 4295 19836 4307 19839
rect 5166 19836 5172 19848
rect 4295 19808 5172 19836
rect 4295 19805 4307 19808
rect 4249 19799 4307 19805
rect 5166 19796 5172 19808
rect 5224 19796 5230 19848
rect 5442 19796 5448 19848
rect 5500 19836 5506 19848
rect 5813 19839 5871 19845
rect 5813 19836 5825 19839
rect 5500 19808 5825 19836
rect 5500 19796 5506 19808
rect 5813 19805 5825 19808
rect 5859 19805 5871 19839
rect 6196 19838 6224 19876
rect 8113 19873 8125 19907
rect 8159 19873 8171 19907
rect 8404 19904 8432 19932
rect 8404 19876 8616 19904
rect 8113 19867 8171 19873
rect 6276 19841 6334 19847
rect 6276 19838 6288 19841
rect 6196 19810 6288 19838
rect 5813 19799 5871 19805
rect 6276 19807 6288 19810
rect 6322 19807 6334 19841
rect 6276 19801 6334 19807
rect 6454 19796 6460 19848
rect 6512 19836 6518 19848
rect 6549 19839 6607 19845
rect 6549 19836 6561 19839
rect 6512 19808 6561 19836
rect 6512 19796 6518 19808
rect 6549 19805 6561 19808
rect 6595 19805 6607 19839
rect 8386 19836 8392 19848
rect 6549 19799 6607 19805
rect 7760 19808 8392 19836
rect 3237 19703 3295 19709
rect 3237 19669 3249 19703
rect 3283 19700 3295 19703
rect 7760 19700 7788 19808
rect 8386 19796 8392 19808
rect 8444 19796 8450 19848
rect 8478 19796 8484 19848
rect 8536 19796 8542 19848
rect 8588 19836 8616 19876
rect 9030 19864 9036 19916
rect 9088 19904 9094 19916
rect 10965 19907 11023 19913
rect 10965 19904 10977 19907
rect 9088 19876 10977 19904
rect 9088 19864 9094 19876
rect 10965 19873 10977 19876
rect 11011 19873 11023 19907
rect 10965 19867 11023 19873
rect 11330 19864 11336 19916
rect 11388 19864 11394 19916
rect 11532 19913 11560 19944
rect 12066 19932 12072 19944
rect 12124 19932 12130 19984
rect 11517 19907 11575 19913
rect 11517 19873 11529 19907
rect 11563 19873 11575 19907
rect 11517 19867 11575 19873
rect 11609 19907 11667 19913
rect 11609 19873 11621 19907
rect 11655 19873 11667 19907
rect 11609 19867 11667 19873
rect 11701 19907 11759 19913
rect 11701 19873 11713 19907
rect 11747 19904 11759 19907
rect 11747 19876 14136 19904
rect 11747 19873 11759 19876
rect 11701 19867 11759 19873
rect 8808 19839 8866 19845
rect 8808 19836 8820 19839
rect 8588 19808 8820 19836
rect 8808 19805 8820 19808
rect 8854 19805 8866 19839
rect 8808 19799 8866 19805
rect 8938 19796 8944 19848
rect 8996 19836 9002 19848
rect 8996 19808 9041 19836
rect 8996 19796 9002 19808
rect 9214 19796 9220 19848
rect 9272 19796 9278 19848
rect 7837 19771 7895 19777
rect 7837 19737 7849 19771
rect 7883 19768 7895 19771
rect 11348 19768 11376 19864
rect 11624 19836 11652 19867
rect 11974 19836 11980 19848
rect 11624 19808 11980 19836
rect 11974 19796 11980 19808
rect 12032 19796 12038 19848
rect 12434 19845 12440 19848
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19805 12127 19839
rect 12069 19799 12127 19805
rect 12396 19839 12440 19845
rect 12396 19805 12408 19839
rect 12396 19799 12440 19805
rect 12084 19768 12112 19799
rect 12434 19796 12440 19799
rect 12492 19796 12498 19848
rect 12575 19839 12633 19845
rect 12575 19805 12587 19839
rect 12621 19836 12633 19839
rect 12710 19836 12716 19848
rect 12621 19808 12716 19836
rect 12621 19805 12633 19808
rect 12575 19799 12633 19805
rect 12710 19796 12716 19808
rect 12768 19796 12774 19848
rect 12802 19796 12808 19848
rect 12860 19796 12866 19848
rect 14108 19836 14136 19876
rect 14182 19864 14188 19916
rect 14240 19904 14246 19916
rect 14277 19907 14335 19913
rect 14277 19904 14289 19907
rect 14240 19876 14289 19904
rect 14240 19864 14246 19876
rect 14277 19873 14289 19876
rect 14323 19873 14335 19907
rect 14277 19867 14335 19873
rect 14553 19907 14611 19913
rect 14553 19873 14565 19907
rect 14599 19904 14611 19907
rect 15378 19904 15384 19916
rect 14599 19876 15384 19904
rect 14599 19873 14611 19876
rect 14553 19867 14611 19873
rect 14568 19836 14596 19867
rect 15378 19864 15384 19876
rect 15436 19864 15442 19916
rect 16393 19907 16451 19913
rect 16393 19873 16405 19907
rect 16439 19904 16451 19907
rect 17512 19904 17540 20000
rect 19889 19975 19947 19981
rect 19889 19941 19901 19975
rect 19935 19972 19947 19975
rect 20990 19972 20996 19984
rect 19935 19944 20996 19972
rect 19935 19941 19947 19944
rect 19889 19935 19947 19941
rect 20990 19932 20996 19944
rect 21048 19932 21054 19984
rect 21910 19932 21916 19984
rect 21968 19932 21974 19984
rect 23750 19972 23756 19984
rect 23690 19944 23756 19972
rect 23750 19932 23756 19944
rect 23808 19972 23814 19984
rect 24136 19972 24164 20012
rect 25130 20000 25136 20012
rect 25188 20000 25194 20052
rect 27338 20000 27344 20052
rect 27396 20040 27402 20052
rect 27801 20043 27859 20049
rect 27801 20040 27813 20043
rect 27396 20012 27813 20040
rect 27396 20000 27402 20012
rect 27801 20009 27813 20012
rect 27847 20009 27859 20043
rect 27801 20003 27859 20009
rect 23808 19944 24164 19972
rect 26053 19975 26111 19981
rect 23808 19932 23814 19944
rect 26053 19941 26065 19975
rect 26099 19972 26111 19975
rect 26099 19944 26556 19972
rect 26099 19941 26111 19944
rect 26053 19935 26111 19941
rect 16439 19876 17540 19904
rect 16439 19873 16451 19876
rect 16393 19867 16451 19873
rect 17954 19864 17960 19916
rect 18012 19904 18018 19916
rect 18141 19907 18199 19913
rect 18141 19904 18153 19907
rect 18012 19876 18153 19904
rect 18012 19864 18018 19876
rect 18141 19873 18153 19876
rect 18187 19873 18199 19907
rect 18141 19867 18199 19873
rect 20622 19864 20628 19916
rect 20680 19864 20686 19916
rect 20898 19864 20904 19916
rect 20956 19904 20962 19916
rect 21358 19904 21364 19916
rect 20956 19876 21364 19904
rect 20956 19864 20962 19876
rect 21358 19864 21364 19876
rect 21416 19864 21422 19916
rect 21450 19864 21456 19916
rect 21508 19864 21514 19916
rect 21542 19864 21548 19916
rect 21600 19864 21606 19916
rect 21928 19904 21956 19932
rect 22005 19907 22063 19913
rect 22005 19904 22017 19907
rect 21928 19876 22017 19904
rect 22005 19873 22017 19876
rect 22051 19873 22063 19907
rect 22005 19867 22063 19873
rect 22186 19864 22192 19916
rect 22244 19864 22250 19916
rect 24213 19907 24271 19913
rect 24213 19873 24225 19907
rect 24259 19873 24271 19907
rect 24673 19907 24731 19913
rect 24673 19904 24685 19907
rect 24213 19867 24271 19873
rect 24320 19876 24685 19904
rect 14108 19808 14596 19836
rect 15930 19796 15936 19848
rect 15988 19836 15994 19848
rect 16117 19839 16175 19845
rect 16117 19836 16129 19839
rect 15988 19808 16129 19836
rect 15988 19796 15994 19808
rect 16117 19805 16129 19808
rect 16163 19805 16175 19839
rect 16117 19799 16175 19805
rect 17218 19796 17224 19848
rect 17276 19836 17282 19848
rect 17862 19836 17868 19848
rect 17276 19808 17868 19836
rect 17276 19796 17282 19808
rect 17862 19796 17868 19808
rect 17920 19836 17926 19848
rect 18230 19836 18236 19848
rect 17920 19808 18236 19836
rect 17920 19796 17926 19808
rect 18230 19796 18236 19808
rect 18288 19796 18294 19848
rect 20993 19839 21051 19845
rect 20993 19805 21005 19839
rect 21039 19836 21051 19839
rect 21468 19836 21496 19864
rect 21039 19808 21496 19836
rect 21039 19805 21051 19808
rect 20993 19799 21051 19805
rect 7883 19740 8432 19768
rect 11348 19740 12112 19768
rect 21560 19768 21588 19864
rect 22465 19839 22523 19845
rect 22465 19836 22477 19839
rect 22296 19808 22477 19836
rect 22296 19768 22324 19808
rect 22465 19805 22477 19808
rect 22511 19836 22523 19839
rect 24228 19836 24256 19867
rect 22511 19808 24256 19836
rect 22511 19805 22523 19808
rect 22465 19799 22523 19805
rect 21560 19740 22324 19768
rect 7883 19737 7895 19740
rect 7837 19731 7895 19737
rect 3283 19672 7788 19700
rect 3283 19669 3295 19672
rect 3237 19663 3295 19669
rect 8294 19660 8300 19712
rect 8352 19660 8358 19712
rect 8404 19700 8432 19740
rect 23474 19728 23480 19780
rect 23532 19768 23538 19780
rect 24320 19768 24348 19876
rect 24673 19873 24685 19876
rect 24719 19873 24731 19907
rect 24673 19867 24731 19873
rect 26234 19864 26240 19916
rect 26292 19904 26298 19916
rect 26410 19907 26468 19913
rect 26410 19904 26422 19907
rect 26292 19876 26422 19904
rect 26292 19864 26298 19876
rect 26410 19873 26422 19876
rect 26456 19873 26468 19907
rect 26528 19904 26556 19944
rect 27890 19932 27896 19984
rect 27948 19972 27954 19984
rect 27948 19944 28488 19972
rect 27948 19932 27954 19944
rect 26697 19907 26755 19913
rect 26697 19904 26709 19907
rect 26528 19876 26709 19904
rect 26410 19867 26468 19873
rect 26697 19873 26709 19876
rect 26743 19873 26755 19907
rect 26697 19867 26755 19873
rect 28350 19864 28356 19916
rect 28408 19864 28414 19916
rect 28460 19904 28488 19944
rect 28460 19876 28948 19904
rect 24394 19796 24400 19848
rect 24452 19836 24458 19848
rect 24452 19808 25360 19836
rect 24452 19796 24458 19808
rect 23532 19740 24348 19768
rect 25332 19768 25360 19808
rect 25958 19796 25964 19848
rect 26016 19836 26022 19848
rect 26344 19836 26556 19838
rect 26016 19810 28304 19836
rect 26016 19808 26372 19810
rect 26528 19808 28304 19810
rect 26016 19796 26022 19808
rect 26418 19768 26424 19780
rect 25332 19740 26424 19768
rect 23532 19728 23538 19740
rect 26418 19728 26424 19740
rect 26476 19728 26482 19780
rect 28169 19771 28227 19777
rect 28169 19737 28181 19771
rect 28215 19737 28227 19771
rect 28169 19731 28227 19737
rect 8662 19700 8668 19712
rect 8404 19672 8668 19700
rect 8662 19660 8668 19672
rect 8720 19660 8726 19712
rect 11885 19703 11943 19709
rect 11885 19669 11897 19703
rect 11931 19700 11943 19703
rect 13722 19700 13728 19712
rect 11931 19672 13728 19700
rect 11931 19669 11943 19672
rect 11885 19663 11943 19669
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 13906 19660 13912 19712
rect 13964 19660 13970 19712
rect 15838 19660 15844 19712
rect 15896 19660 15902 19712
rect 17681 19703 17739 19709
rect 17681 19669 17693 19703
rect 17727 19700 17739 19703
rect 18138 19700 18144 19712
rect 17727 19672 18144 19700
rect 17727 19669 17739 19672
rect 17681 19663 17739 19669
rect 18138 19660 18144 19672
rect 18196 19660 18202 19712
rect 19150 19660 19156 19712
rect 19208 19700 19214 19712
rect 19245 19703 19303 19709
rect 19245 19700 19257 19703
rect 19208 19672 19257 19700
rect 19208 19660 19214 19672
rect 19245 19669 19257 19672
rect 19291 19669 19303 19703
rect 19245 19663 19303 19669
rect 21266 19660 21272 19712
rect 21324 19700 21330 19712
rect 21453 19703 21511 19709
rect 21453 19700 21465 19703
rect 21324 19672 21465 19700
rect 21324 19660 21330 19672
rect 21453 19669 21465 19672
rect 21499 19669 21511 19703
rect 21453 19663 21511 19669
rect 21542 19660 21548 19712
rect 21600 19700 21606 19712
rect 22646 19700 22652 19712
rect 21600 19672 22652 19700
rect 21600 19660 21606 19672
rect 22646 19660 22652 19672
rect 22704 19660 22710 19712
rect 23566 19660 23572 19712
rect 23624 19700 23630 19712
rect 28184 19700 28212 19731
rect 23624 19672 28212 19700
rect 28276 19700 28304 19808
rect 28442 19796 28448 19848
rect 28500 19796 28506 19848
rect 28810 19845 28816 19848
rect 28772 19839 28816 19845
rect 28772 19805 28784 19839
rect 28772 19799 28816 19805
rect 28810 19796 28816 19799
rect 28868 19796 28874 19848
rect 28920 19845 28948 19876
rect 28908 19839 28966 19845
rect 28908 19805 28920 19839
rect 28954 19805 28966 19839
rect 28908 19799 28966 19805
rect 29181 19839 29239 19845
rect 29181 19805 29193 19839
rect 29227 19836 29239 19839
rect 29638 19836 29644 19848
rect 29227 19808 29644 19836
rect 29227 19805 29239 19808
rect 29181 19799 29239 19805
rect 29638 19796 29644 19808
rect 29696 19796 29702 19848
rect 30285 19703 30343 19709
rect 30285 19700 30297 19703
rect 28276 19672 30297 19700
rect 23624 19660 23630 19672
rect 30285 19669 30297 19672
rect 30331 19669 30343 19703
rect 30285 19663 30343 19669
rect 552 19610 30912 19632
rect 552 19558 4193 19610
rect 4245 19558 4257 19610
rect 4309 19558 4321 19610
rect 4373 19558 4385 19610
rect 4437 19558 4449 19610
rect 4501 19558 11783 19610
rect 11835 19558 11847 19610
rect 11899 19558 11911 19610
rect 11963 19558 11975 19610
rect 12027 19558 12039 19610
rect 12091 19558 19373 19610
rect 19425 19558 19437 19610
rect 19489 19558 19501 19610
rect 19553 19558 19565 19610
rect 19617 19558 19629 19610
rect 19681 19558 26963 19610
rect 27015 19558 27027 19610
rect 27079 19558 27091 19610
rect 27143 19558 27155 19610
rect 27207 19558 27219 19610
rect 27271 19558 30912 19610
rect 552 19536 30912 19558
rect 2774 19456 2780 19508
rect 2832 19456 2838 19508
rect 3326 19456 3332 19508
rect 3384 19496 3390 19508
rect 4617 19499 4675 19505
rect 4617 19496 4629 19499
rect 3384 19468 4629 19496
rect 3384 19456 3390 19468
rect 4617 19465 4629 19468
rect 4663 19496 4675 19499
rect 5626 19496 5632 19508
rect 4663 19468 5632 19496
rect 4663 19465 4675 19468
rect 4617 19459 4675 19465
rect 5626 19456 5632 19468
rect 5684 19456 5690 19508
rect 5718 19456 5724 19508
rect 5776 19496 5782 19508
rect 5776 19468 6776 19496
rect 5776 19456 5782 19468
rect 5350 19388 5356 19440
rect 5408 19388 5414 19440
rect 1443 19363 1501 19369
rect 1443 19329 1455 19363
rect 1489 19360 1501 19363
rect 3050 19360 3056 19372
rect 1489 19332 3056 19360
rect 1489 19329 1501 19332
rect 1443 19323 1501 19329
rect 3050 19320 3056 19332
rect 3108 19320 3114 19372
rect 3878 19320 3884 19372
rect 3936 19320 3942 19372
rect 5368 19360 5396 19388
rect 5816 19363 5874 19369
rect 5816 19360 5828 19363
rect 5368 19332 5828 19360
rect 5816 19329 5828 19332
rect 5862 19329 5874 19363
rect 5816 19323 5874 19329
rect 5994 19320 6000 19372
rect 6052 19360 6058 19372
rect 6748 19360 6776 19468
rect 8294 19456 8300 19508
rect 8352 19496 8358 19508
rect 9582 19496 9588 19508
rect 8352 19468 9588 19496
rect 8352 19456 8358 19468
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 10226 19456 10232 19508
rect 10284 19456 10290 19508
rect 10686 19456 10692 19508
rect 10744 19496 10750 19508
rect 13446 19496 13452 19508
rect 10744 19468 13452 19496
rect 10744 19456 10750 19468
rect 13446 19456 13452 19468
rect 13504 19456 13510 19508
rect 13998 19456 14004 19508
rect 14056 19496 14062 19508
rect 14056 19468 15240 19496
rect 14056 19456 14062 19468
rect 6914 19388 6920 19440
rect 6972 19428 6978 19440
rect 6972 19400 8432 19428
rect 6972 19388 6978 19400
rect 6052 19332 6592 19360
rect 6748 19332 8340 19360
rect 6052 19320 6058 19332
rect 937 19295 995 19301
rect 937 19261 949 19295
rect 983 19292 995 19295
rect 1026 19292 1032 19304
rect 983 19264 1032 19292
rect 983 19261 995 19264
rect 937 19255 995 19261
rect 1026 19252 1032 19264
rect 1084 19252 1090 19304
rect 1673 19295 1731 19301
rect 1673 19261 1685 19295
rect 1719 19292 1731 19295
rect 2130 19292 2136 19304
rect 1719 19264 2136 19292
rect 1719 19261 1731 19264
rect 1673 19255 1731 19261
rect 2130 19252 2136 19264
rect 2188 19252 2194 19304
rect 3602 19252 3608 19304
rect 3660 19252 3666 19304
rect 3697 19295 3755 19301
rect 3697 19261 3709 19295
rect 3743 19261 3755 19295
rect 3697 19255 3755 19261
rect 4341 19295 4399 19301
rect 4341 19261 4353 19295
rect 4387 19292 4399 19295
rect 4522 19292 4528 19304
rect 4387 19264 4528 19292
rect 4387 19261 4399 19264
rect 4341 19255 4399 19261
rect 3712 19224 3740 19255
rect 4522 19252 4528 19264
rect 4580 19292 4586 19304
rect 5261 19295 5319 19301
rect 5261 19292 5273 19295
rect 4580 19264 5273 19292
rect 4580 19252 4586 19264
rect 5261 19261 5273 19264
rect 5307 19292 5319 19295
rect 5353 19295 5411 19301
rect 5353 19292 5365 19295
rect 5307 19264 5365 19292
rect 5307 19261 5319 19264
rect 5261 19255 5319 19261
rect 5353 19261 5365 19264
rect 5399 19292 5411 19295
rect 5442 19292 5448 19304
rect 5399 19264 5448 19292
rect 5399 19261 5411 19264
rect 5353 19255 5411 19261
rect 5442 19252 5448 19264
rect 5500 19252 5506 19304
rect 6089 19295 6147 19301
rect 6089 19261 6101 19295
rect 6135 19292 6147 19295
rect 6454 19292 6460 19304
rect 6135 19264 6460 19292
rect 6135 19261 6147 19264
rect 6089 19255 6147 19261
rect 6454 19252 6460 19264
rect 6512 19252 6518 19304
rect 6564 19292 6592 19332
rect 6564 19264 7239 19292
rect 3878 19224 3884 19236
rect 3712 19196 3884 19224
rect 3878 19184 3884 19196
rect 3936 19184 3942 19236
rect 4798 19224 4804 19236
rect 4356 19196 4804 19224
rect 1403 19159 1461 19165
rect 1403 19125 1415 19159
rect 1449 19156 1461 19159
rect 1762 19156 1768 19168
rect 1449 19128 1768 19156
rect 1449 19125 1461 19128
rect 1403 19119 1461 19125
rect 1762 19116 1768 19128
rect 1820 19116 1826 19168
rect 3421 19159 3479 19165
rect 3421 19125 3433 19159
rect 3467 19156 3479 19159
rect 4356 19156 4384 19196
rect 4798 19184 4804 19196
rect 4856 19184 4862 19236
rect 4893 19227 4951 19233
rect 4893 19193 4905 19227
rect 4939 19193 4951 19227
rect 7211 19224 7239 19264
rect 7282 19252 7288 19304
rect 7340 19292 7346 19304
rect 7745 19295 7803 19301
rect 7745 19292 7757 19295
rect 7340 19264 7757 19292
rect 7340 19252 7346 19264
rect 7745 19261 7757 19264
rect 7791 19261 7803 19295
rect 7745 19255 7803 19261
rect 7211 19196 7788 19224
rect 4893 19187 4951 19193
rect 3467 19128 4384 19156
rect 4908 19156 4936 19187
rect 5718 19156 5724 19168
rect 4908 19128 5724 19156
rect 3467 19125 3479 19128
rect 3421 19119 3479 19125
rect 5718 19116 5724 19128
rect 5776 19116 5782 19168
rect 5810 19116 5816 19168
rect 5868 19165 5874 19168
rect 5868 19119 5877 19165
rect 5868 19116 5874 19119
rect 6730 19116 6736 19168
rect 6788 19156 6794 19168
rect 7193 19159 7251 19165
rect 7193 19156 7205 19159
rect 6788 19128 7205 19156
rect 6788 19116 6794 19128
rect 7193 19125 7205 19128
rect 7239 19125 7251 19159
rect 7760 19156 7788 19196
rect 7834 19184 7840 19236
rect 7892 19224 7898 19236
rect 8021 19227 8079 19233
rect 8021 19224 8033 19227
rect 7892 19196 8033 19224
rect 7892 19184 7898 19196
rect 8021 19193 8033 19196
rect 8067 19193 8079 19227
rect 8312 19224 8340 19332
rect 8404 19301 8432 19400
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 8852 19363 8910 19369
rect 8852 19360 8864 19363
rect 8628 19332 8864 19360
rect 8628 19320 8634 19332
rect 8852 19329 8864 19332
rect 8898 19329 8910 19363
rect 8852 19323 8910 19329
rect 8938 19320 8944 19372
rect 8996 19360 9002 19372
rect 8996 19332 9536 19360
rect 8996 19320 9002 19332
rect 8389 19295 8447 19301
rect 8389 19261 8401 19295
rect 8435 19292 8447 19295
rect 8662 19292 8668 19304
rect 8435 19264 8668 19292
rect 8435 19261 8447 19264
rect 8389 19255 8447 19261
rect 8662 19252 8668 19264
rect 8720 19252 8726 19304
rect 9125 19295 9183 19301
rect 9125 19261 9137 19295
rect 9171 19292 9183 19295
rect 9398 19292 9404 19304
rect 9171 19264 9404 19292
rect 9171 19261 9183 19264
rect 9125 19255 9183 19261
rect 9398 19252 9404 19264
rect 9456 19252 9462 19304
rect 9508 19292 9536 19332
rect 11054 19320 11060 19372
rect 11112 19360 11118 19372
rect 11244 19363 11302 19369
rect 11244 19360 11256 19363
rect 11112 19332 11256 19360
rect 11112 19320 11118 19332
rect 11244 19329 11256 19332
rect 11290 19329 11302 19363
rect 11244 19323 11302 19329
rect 14182 19320 14188 19372
rect 14240 19320 14246 19372
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19360 14519 19363
rect 14826 19360 14832 19372
rect 14507 19332 14832 19360
rect 14507 19329 14519 19332
rect 14461 19323 14519 19329
rect 14826 19320 14832 19332
rect 14884 19320 14890 19372
rect 10781 19295 10839 19301
rect 10781 19292 10793 19295
rect 9508 19264 10793 19292
rect 10781 19261 10793 19264
rect 10827 19261 10839 19295
rect 11517 19295 11575 19301
rect 11517 19292 11529 19295
rect 10781 19255 10839 19261
rect 10888 19264 11529 19292
rect 8478 19224 8484 19236
rect 8312 19196 8484 19224
rect 8021 19187 8079 19193
rect 8478 19184 8484 19196
rect 8536 19184 8542 19236
rect 9950 19184 9956 19236
rect 10008 19224 10014 19236
rect 10888 19224 10916 19264
rect 11517 19261 11529 19264
rect 11563 19261 11575 19295
rect 11517 19255 11575 19261
rect 11974 19252 11980 19304
rect 12032 19292 12038 19304
rect 13173 19295 13231 19301
rect 13173 19292 13185 19295
rect 12032 19264 13185 19292
rect 12032 19252 12038 19264
rect 13173 19261 13185 19264
rect 13219 19292 13231 19295
rect 13262 19292 13268 19304
rect 13219 19264 13268 19292
rect 13219 19261 13231 19264
rect 13173 19255 13231 19261
rect 13262 19252 13268 19264
rect 13320 19252 13326 19304
rect 15212 19292 15240 19468
rect 16114 19456 16120 19508
rect 16172 19496 16178 19508
rect 22005 19499 22063 19505
rect 16172 19468 19656 19496
rect 16172 19456 16178 19468
rect 15838 19320 15844 19372
rect 15896 19360 15902 19372
rect 16209 19363 16267 19369
rect 16209 19360 16221 19363
rect 15896 19332 16221 19360
rect 15896 19320 15902 19332
rect 16209 19329 16221 19332
rect 16255 19329 16267 19363
rect 16209 19323 16267 19329
rect 17770 19320 17776 19372
rect 17828 19360 17834 19372
rect 18156 19369 18184 19468
rect 18141 19363 18199 19369
rect 17828 19332 18000 19360
rect 17828 19320 17834 19332
rect 15930 19292 15936 19304
rect 15212 19264 15936 19292
rect 15930 19252 15936 19264
rect 15988 19252 15994 19304
rect 17218 19292 17224 19304
rect 16040 19264 17224 19292
rect 10008 19196 10916 19224
rect 13725 19227 13783 19233
rect 10008 19184 10014 19196
rect 13725 19193 13737 19227
rect 13771 19193 13783 19227
rect 16040 19224 16068 19264
rect 17218 19252 17224 19264
rect 17276 19252 17282 19304
rect 17678 19252 17684 19304
rect 17736 19292 17742 19304
rect 17865 19295 17923 19301
rect 17865 19292 17877 19295
rect 17736 19264 17877 19292
rect 17736 19252 17742 19264
rect 17865 19261 17877 19264
rect 17911 19261 17923 19295
rect 17972 19292 18000 19332
rect 18141 19329 18153 19363
rect 18187 19329 18199 19363
rect 18141 19323 18199 19329
rect 18230 19320 18236 19372
rect 18288 19360 18294 19372
rect 18693 19363 18751 19369
rect 18693 19360 18705 19363
rect 18288 19332 18705 19360
rect 18288 19320 18294 19332
rect 18693 19329 18705 19332
rect 18739 19329 18751 19363
rect 19628 19360 19656 19468
rect 22005 19465 22017 19499
rect 22051 19496 22063 19499
rect 23474 19496 23480 19508
rect 22051 19468 23480 19496
rect 22051 19465 22063 19468
rect 22005 19459 22063 19465
rect 23474 19456 23480 19468
rect 23532 19456 23538 19508
rect 24394 19456 24400 19508
rect 24452 19456 24458 19508
rect 26510 19456 26516 19508
rect 26568 19496 26574 19508
rect 30098 19496 30104 19508
rect 26568 19468 30104 19496
rect 26568 19456 26574 19468
rect 30098 19456 30104 19468
rect 30156 19456 30162 19508
rect 21542 19388 21548 19440
rect 21600 19428 21606 19440
rect 22557 19431 22615 19437
rect 22557 19428 22569 19431
rect 21600 19400 22569 19428
rect 21600 19388 21606 19400
rect 22557 19397 22569 19400
rect 22603 19428 22615 19431
rect 24412 19428 24440 19456
rect 22603 19400 24440 19428
rect 22603 19397 22615 19400
rect 22557 19391 22615 19397
rect 19628 19332 22094 19360
rect 18693 19323 18751 19329
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17972 19264 18061 19292
rect 17865 19255 17923 19261
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18969 19295 19027 19301
rect 18969 19292 18981 19295
rect 18049 19255 18107 19261
rect 18800 19264 18981 19292
rect 13725 19187 13783 19193
rect 15672 19196 16068 19224
rect 17589 19227 17647 19233
rect 8855 19159 8913 19165
rect 8855 19156 8867 19159
rect 7760 19128 8867 19156
rect 7193 19119 7251 19125
rect 8855 19125 8867 19128
rect 8901 19156 8913 19159
rect 9122 19156 9128 19168
rect 8901 19128 9128 19156
rect 8901 19125 8913 19128
rect 8855 19119 8913 19125
rect 9122 19116 9128 19128
rect 9180 19116 9186 19168
rect 11146 19116 11152 19168
rect 11204 19156 11210 19168
rect 11247 19159 11305 19165
rect 11247 19156 11259 19159
rect 11204 19128 11259 19156
rect 11204 19116 11210 19128
rect 11247 19125 11259 19128
rect 11293 19125 11305 19159
rect 11247 19119 11305 19125
rect 11422 19116 11428 19168
rect 11480 19156 11486 19168
rect 12158 19156 12164 19168
rect 11480 19128 12164 19156
rect 11480 19116 11486 19128
rect 12158 19116 12164 19128
rect 12216 19116 12222 19168
rect 12526 19116 12532 19168
rect 12584 19156 12590 19168
rect 12621 19159 12679 19165
rect 12621 19156 12633 19159
rect 12584 19128 12633 19156
rect 12584 19116 12590 19128
rect 12621 19125 12633 19128
rect 12667 19125 12679 19159
rect 12621 19119 12679 19125
rect 12986 19116 12992 19168
rect 13044 19116 13050 19168
rect 13740 19156 13768 19187
rect 15672 19156 15700 19196
rect 17589 19193 17601 19227
rect 17635 19224 17647 19227
rect 18800 19224 18828 19264
rect 18969 19261 18981 19264
rect 19015 19261 19027 19295
rect 18969 19255 19027 19261
rect 20438 19252 20444 19304
rect 20496 19252 20502 19304
rect 20530 19252 20536 19304
rect 20588 19292 20594 19304
rect 20717 19295 20775 19301
rect 20717 19292 20729 19295
rect 20588 19264 20729 19292
rect 20588 19252 20594 19264
rect 20717 19261 20729 19264
rect 20763 19261 20775 19295
rect 22066 19292 22094 19332
rect 23566 19320 23572 19372
rect 23624 19320 23630 19372
rect 26694 19320 26700 19372
rect 26752 19320 26758 19372
rect 27203 19363 27261 19369
rect 27203 19329 27215 19363
rect 27249 19360 27261 19363
rect 27338 19360 27344 19372
rect 27249 19332 27344 19360
rect 27249 19329 27261 19332
rect 27203 19323 27261 19329
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 28902 19320 28908 19372
rect 28960 19360 28966 19372
rect 28997 19363 29055 19369
rect 28997 19360 29009 19363
rect 28960 19332 29009 19360
rect 28960 19320 28966 19332
rect 28997 19329 29009 19332
rect 29043 19329 29055 19363
rect 28997 19323 29055 19329
rect 22066 19264 22968 19292
rect 20717 19255 20775 19261
rect 17635 19196 18828 19224
rect 22281 19227 22339 19233
rect 17635 19193 17647 19196
rect 17589 19187 17647 19193
rect 22281 19193 22293 19227
rect 22327 19224 22339 19227
rect 22830 19224 22836 19236
rect 22327 19196 22836 19224
rect 22327 19193 22339 19196
rect 22281 19187 22339 19193
rect 22830 19184 22836 19196
rect 22888 19184 22894 19236
rect 22940 19224 22968 19264
rect 23014 19252 23020 19304
rect 23072 19292 23078 19304
rect 23293 19295 23351 19301
rect 23293 19292 23305 19295
rect 23072 19264 23305 19292
rect 23072 19252 23078 19264
rect 23293 19261 23305 19264
rect 23339 19261 23351 19295
rect 23293 19255 23351 19261
rect 23385 19295 23443 19301
rect 23385 19261 23397 19295
rect 23431 19292 23443 19295
rect 24486 19292 24492 19304
rect 23431 19264 24492 19292
rect 23431 19261 23443 19264
rect 23385 19255 23443 19261
rect 24486 19252 24492 19264
rect 24544 19252 24550 19304
rect 27062 19301 27068 19304
rect 27024 19295 27068 19301
rect 27024 19261 27036 19295
rect 27024 19255 27068 19261
rect 27062 19252 27068 19255
rect 27120 19252 27126 19304
rect 27433 19295 27491 19301
rect 27433 19261 27445 19295
rect 27479 19292 27491 19295
rect 29012 19292 29040 19323
rect 29273 19295 29331 19301
rect 27479 19264 28948 19292
rect 29012 19264 29224 19292
rect 27479 19261 27491 19264
rect 27433 19255 27491 19261
rect 23566 19224 23572 19236
rect 22940 19196 23572 19224
rect 23566 19184 23572 19196
rect 23624 19184 23630 19236
rect 24118 19184 24124 19236
rect 24176 19184 24182 19236
rect 24210 19184 24216 19236
rect 24268 19184 24274 19236
rect 26510 19184 26516 19236
rect 26568 19224 26574 19236
rect 28920 19224 28948 19264
rect 29086 19224 29092 19236
rect 26568 19196 26740 19224
rect 28920 19196 29092 19224
rect 26568 19184 26574 19196
rect 13740 19128 15700 19156
rect 15749 19159 15807 19165
rect 15749 19125 15761 19159
rect 15795 19156 15807 19159
rect 16022 19156 16028 19168
rect 15795 19128 16028 19156
rect 15795 19125 15807 19128
rect 15749 19119 15807 19125
rect 16022 19116 16028 19128
rect 16080 19116 16086 19168
rect 16298 19116 16304 19168
rect 16356 19156 16362 19168
rect 18325 19159 18383 19165
rect 18325 19156 18337 19159
rect 16356 19128 18337 19156
rect 16356 19116 16362 19128
rect 18325 19125 18337 19128
rect 18371 19125 18383 19159
rect 18325 19119 18383 19125
rect 20070 19116 20076 19168
rect 20128 19116 20134 19168
rect 22925 19159 22983 19165
rect 22925 19125 22937 19159
rect 22971 19156 22983 19159
rect 24228 19156 24256 19184
rect 22971 19128 24256 19156
rect 24397 19159 24455 19165
rect 22971 19125 22983 19128
rect 22925 19119 22983 19125
rect 24397 19125 24409 19159
rect 24443 19156 24455 19159
rect 24486 19156 24492 19168
rect 24443 19128 24492 19156
rect 24443 19125 24455 19128
rect 24397 19119 24455 19125
rect 24486 19116 24492 19128
rect 24544 19116 24550 19168
rect 24949 19159 25007 19165
rect 24949 19125 24961 19159
rect 24995 19156 25007 19159
rect 25130 19156 25136 19168
rect 24995 19128 25136 19156
rect 24995 19125 25007 19128
rect 24949 19119 25007 19125
rect 25130 19116 25136 19128
rect 25188 19116 25194 19168
rect 25409 19159 25467 19165
rect 25409 19125 25421 19159
rect 25455 19156 25467 19159
rect 25498 19156 25504 19168
rect 25455 19128 25504 19156
rect 25455 19125 25467 19128
rect 25409 19119 25467 19125
rect 25498 19116 25504 19128
rect 25556 19116 25562 19168
rect 25869 19159 25927 19165
rect 25869 19125 25881 19159
rect 25915 19156 25927 19159
rect 26050 19156 26056 19168
rect 25915 19128 26056 19156
rect 25915 19125 25927 19128
rect 25869 19119 25927 19125
rect 26050 19116 26056 19128
rect 26108 19116 26114 19168
rect 26329 19159 26387 19165
rect 26329 19125 26341 19159
rect 26375 19156 26387 19159
rect 26602 19156 26608 19168
rect 26375 19128 26608 19156
rect 26375 19125 26387 19128
rect 26329 19119 26387 19125
rect 26602 19116 26608 19128
rect 26660 19116 26666 19168
rect 26712 19156 26740 19196
rect 29086 19184 29092 19196
rect 29144 19184 29150 19236
rect 29196 19224 29224 19264
rect 29273 19261 29285 19295
rect 29319 19292 29331 19295
rect 29914 19292 29920 19304
rect 29319 19264 29920 19292
rect 29319 19261 29331 19264
rect 29273 19255 29331 19261
rect 29914 19252 29920 19264
rect 29972 19252 29978 19304
rect 29546 19224 29552 19236
rect 29196 19196 29552 19224
rect 29546 19184 29552 19196
rect 29604 19184 29610 19236
rect 30285 19227 30343 19233
rect 30285 19224 30297 19227
rect 30116 19196 30297 19224
rect 30116 19168 30144 19196
rect 30285 19193 30297 19196
rect 30331 19193 30343 19227
rect 30285 19187 30343 19193
rect 27706 19156 27712 19168
rect 26712 19128 27712 19156
rect 27706 19116 27712 19128
rect 27764 19116 27770 19168
rect 28534 19116 28540 19168
rect 28592 19116 28598 19168
rect 29917 19159 29975 19165
rect 29917 19125 29929 19159
rect 29963 19156 29975 19159
rect 30006 19156 30012 19168
rect 29963 19128 30012 19156
rect 29963 19125 29975 19128
rect 29917 19119 29975 19125
rect 30006 19116 30012 19128
rect 30064 19116 30070 19168
rect 30098 19116 30104 19168
rect 30156 19116 30162 19168
rect 30377 19159 30435 19165
rect 30377 19125 30389 19159
rect 30423 19156 30435 19159
rect 30650 19156 30656 19168
rect 30423 19128 30656 19156
rect 30423 19125 30435 19128
rect 30377 19119 30435 19125
rect 30650 19116 30656 19128
rect 30708 19116 30714 19168
rect 552 19066 31072 19088
rect 552 19014 7988 19066
rect 8040 19014 8052 19066
rect 8104 19014 8116 19066
rect 8168 19014 8180 19066
rect 8232 19014 8244 19066
rect 8296 19014 15578 19066
rect 15630 19014 15642 19066
rect 15694 19014 15706 19066
rect 15758 19014 15770 19066
rect 15822 19014 15834 19066
rect 15886 19014 23168 19066
rect 23220 19014 23232 19066
rect 23284 19014 23296 19066
rect 23348 19014 23360 19066
rect 23412 19014 23424 19066
rect 23476 19014 30758 19066
rect 30810 19014 30822 19066
rect 30874 19014 30886 19066
rect 30938 19014 30950 19066
rect 31002 19014 31014 19066
rect 31066 19014 31072 19066
rect 552 18992 31072 19014
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 1728 18924 2774 18952
rect 1728 18912 1734 18924
rect 2746 18884 2774 18924
rect 3142 18912 3148 18964
rect 3200 18912 3206 18964
rect 6822 18952 6828 18964
rect 5276 18924 6828 18952
rect 4157 18887 4215 18893
rect 4157 18884 4169 18887
rect 1136 18856 1348 18884
rect 2746 18856 4169 18884
rect 1136 18760 1164 18856
rect 1210 18776 1216 18828
rect 1268 18776 1274 18828
rect 1320 18825 1348 18856
rect 1305 18819 1363 18825
rect 1305 18785 1317 18819
rect 1351 18785 1363 18819
rect 2314 18816 2320 18828
rect 1305 18779 1363 18785
rect 1826 18788 2320 18816
rect 1118 18708 1124 18760
rect 1176 18708 1182 18760
rect 1826 18759 1854 18788
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 1632 18751 1690 18757
rect 1632 18748 1644 18751
rect 1320 18720 1644 18748
rect 1026 18572 1032 18624
rect 1084 18572 1090 18624
rect 1320 18612 1348 18720
rect 1632 18717 1644 18720
rect 1678 18717 1690 18751
rect 1632 18711 1690 18717
rect 1811 18753 1869 18759
rect 1811 18719 1823 18753
rect 1857 18719 1869 18753
rect 1811 18713 1869 18719
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18748 2099 18751
rect 2087 18720 2774 18748
rect 2087 18717 2099 18720
rect 2041 18711 2099 18717
rect 1762 18612 1768 18624
rect 1320 18584 1768 18612
rect 1762 18572 1768 18584
rect 1820 18572 1826 18624
rect 2746 18612 2774 18720
rect 3804 18680 3832 18856
rect 4157 18853 4169 18856
rect 4203 18853 4215 18887
rect 4157 18847 4215 18853
rect 4706 18844 4712 18896
rect 4764 18844 4770 18896
rect 5074 18844 5080 18896
rect 5132 18844 5138 18896
rect 5276 18893 5304 18924
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 8481 18955 8539 18961
rect 8481 18921 8493 18955
rect 8527 18952 8539 18955
rect 11974 18952 11980 18964
rect 8527 18924 11980 18952
rect 8527 18921 8539 18924
rect 8481 18915 8539 18921
rect 11974 18912 11980 18924
rect 12032 18912 12038 18964
rect 12342 18952 12348 18964
rect 12400 18961 12406 18964
rect 12309 18924 12348 18952
rect 12342 18912 12348 18924
rect 12400 18915 12409 18961
rect 12400 18912 12406 18915
rect 13814 18912 13820 18964
rect 13872 18952 13878 18964
rect 13909 18955 13967 18961
rect 13909 18952 13921 18955
rect 13872 18924 13921 18952
rect 13872 18912 13878 18924
rect 13909 18921 13921 18924
rect 13955 18921 13967 18955
rect 13909 18915 13967 18921
rect 16022 18912 16028 18964
rect 16080 18912 16086 18964
rect 17681 18955 17739 18961
rect 17681 18921 17693 18955
rect 17727 18952 17739 18955
rect 17954 18952 17960 18964
rect 17727 18924 17960 18952
rect 17727 18921 17739 18924
rect 17681 18915 17739 18921
rect 17954 18912 17960 18924
rect 18012 18912 18018 18964
rect 20622 18952 20628 18964
rect 20272 18924 20628 18952
rect 5261 18887 5319 18893
rect 5261 18853 5273 18887
rect 5307 18853 5319 18887
rect 5261 18847 5319 18853
rect 8113 18887 8171 18893
rect 8113 18853 8125 18887
rect 8159 18884 8171 18887
rect 8570 18884 8576 18896
rect 8159 18856 8576 18884
rect 8159 18853 8171 18856
rect 8113 18847 8171 18853
rect 8570 18844 8576 18856
rect 8628 18844 8634 18896
rect 10410 18844 10416 18896
rect 10468 18884 10474 18896
rect 10781 18887 10839 18893
rect 10468 18856 10640 18884
rect 10468 18844 10474 18856
rect 3878 18776 3884 18828
rect 3936 18776 3942 18828
rect 5902 18776 5908 18828
rect 5960 18816 5966 18828
rect 5997 18819 6055 18825
rect 5997 18816 6009 18819
rect 5960 18788 6009 18816
rect 5960 18776 5966 18788
rect 5997 18785 6009 18788
rect 6043 18785 6055 18819
rect 5997 18779 6055 18785
rect 6086 18776 6092 18828
rect 6144 18816 6150 18828
rect 6324 18819 6382 18825
rect 6324 18816 6336 18819
rect 6144 18788 6336 18816
rect 6144 18776 6150 18788
rect 6324 18785 6336 18788
rect 6370 18785 6382 18819
rect 6324 18779 6382 18785
rect 8389 18819 8447 18825
rect 8389 18785 8401 18819
rect 8435 18816 8447 18819
rect 8754 18816 8760 18828
rect 8435 18788 8760 18816
rect 8435 18785 8447 18788
rect 8389 18779 8447 18785
rect 8754 18776 8760 18788
rect 8812 18776 8818 18828
rect 9030 18825 9036 18828
rect 8992 18819 9036 18825
rect 8992 18785 9004 18819
rect 8992 18779 9036 18785
rect 9030 18776 9036 18779
rect 9088 18776 9094 18828
rect 10612 18816 10640 18856
rect 10781 18853 10793 18887
rect 10827 18884 10839 18887
rect 10870 18884 10876 18896
rect 10827 18856 10876 18884
rect 10827 18853 10839 18856
rect 10781 18847 10839 18853
rect 10870 18844 10876 18856
rect 10928 18844 10934 18896
rect 11348 18856 11928 18884
rect 11348 18828 11376 18856
rect 10965 18819 11023 18825
rect 10965 18816 10977 18819
rect 9324 18788 10548 18816
rect 10612 18788 10977 18816
rect 6104 18748 6132 18776
rect 5736 18720 6132 18748
rect 5736 18680 5764 18720
rect 6454 18708 6460 18760
rect 6512 18708 6518 18760
rect 6730 18708 6736 18760
rect 6788 18708 6794 18760
rect 8478 18748 8484 18760
rect 7392 18720 8484 18748
rect 3804 18652 5764 18680
rect 3786 18612 3792 18624
rect 2746 18584 3792 18612
rect 3786 18572 3792 18584
rect 3844 18572 3850 18624
rect 5537 18615 5595 18621
rect 5537 18581 5549 18615
rect 5583 18612 5595 18615
rect 7392 18612 7420 18720
rect 8478 18708 8484 18720
rect 8536 18708 8542 18760
rect 8570 18708 8576 18760
rect 8628 18748 8634 18760
rect 8665 18751 8723 18757
rect 8665 18748 8677 18751
rect 8628 18720 8677 18748
rect 8628 18708 8634 18720
rect 8665 18717 8677 18720
rect 8711 18717 8723 18751
rect 8665 18711 8723 18717
rect 9171 18751 9229 18757
rect 9171 18717 9183 18751
rect 9217 18748 9229 18751
rect 9324 18748 9352 18788
rect 10520 18760 10548 18788
rect 10965 18785 10977 18788
rect 11011 18785 11023 18819
rect 10965 18779 11023 18785
rect 11330 18776 11336 18828
rect 11388 18776 11394 18828
rect 11900 18825 11928 18856
rect 11517 18819 11575 18825
rect 11517 18785 11529 18819
rect 11563 18785 11575 18819
rect 11517 18779 11575 18785
rect 11885 18819 11943 18825
rect 11885 18785 11897 18819
rect 11931 18785 11943 18819
rect 12526 18816 12532 18828
rect 11885 18779 11943 18785
rect 12406 18788 12532 18816
rect 9217 18720 9352 18748
rect 9217 18717 9229 18720
rect 9171 18711 9229 18717
rect 9398 18708 9404 18760
rect 9456 18708 9462 18760
rect 9490 18708 9496 18760
rect 9548 18748 9554 18760
rect 9548 18720 10456 18748
rect 9548 18708 9554 18720
rect 8386 18640 8392 18692
rect 8444 18640 8450 18692
rect 10428 18680 10456 18720
rect 10502 18708 10508 18760
rect 10560 18708 10566 18760
rect 11146 18708 11152 18760
rect 11204 18708 11210 18760
rect 11532 18748 11560 18779
rect 12406 18759 12434 18788
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 12621 18819 12679 18825
rect 12621 18785 12633 18819
rect 12667 18816 12679 18819
rect 12986 18816 12992 18828
rect 12667 18788 12992 18816
rect 12667 18785 12679 18788
rect 12621 18779 12679 18785
rect 12986 18776 12992 18788
rect 13044 18776 13050 18828
rect 14550 18776 14556 18828
rect 14608 18776 14614 18828
rect 15930 18776 15936 18828
rect 15988 18776 15994 18828
rect 16040 18816 16068 18912
rect 16393 18819 16451 18825
rect 16393 18816 16405 18819
rect 16040 18788 16405 18816
rect 16393 18785 16405 18788
rect 16439 18785 16451 18819
rect 16393 18779 16451 18785
rect 17218 18776 17224 18828
rect 17276 18816 17282 18828
rect 17865 18819 17923 18825
rect 17865 18816 17877 18819
rect 17276 18788 17877 18816
rect 17276 18776 17282 18788
rect 17865 18785 17877 18788
rect 17911 18785 17923 18819
rect 17865 18779 17923 18785
rect 18138 18776 18144 18828
rect 18196 18776 18202 18828
rect 19886 18776 19892 18828
rect 19944 18776 19950 18828
rect 20272 18825 20300 18924
rect 20622 18912 20628 18924
rect 20680 18912 20686 18964
rect 22649 18955 22707 18961
rect 22649 18952 22661 18955
rect 20916 18924 22661 18952
rect 20916 18884 20944 18924
rect 22649 18921 22661 18924
rect 22695 18921 22707 18955
rect 22649 18915 22707 18921
rect 22830 18912 22836 18964
rect 22888 18912 22894 18964
rect 23293 18955 23351 18961
rect 23293 18921 23305 18955
rect 23339 18952 23351 18955
rect 23658 18952 23664 18964
rect 23339 18924 23664 18952
rect 23339 18921 23351 18924
rect 23293 18915 23351 18921
rect 23658 18912 23664 18924
rect 23716 18912 23722 18964
rect 23753 18955 23811 18961
rect 23753 18921 23765 18955
rect 23799 18952 23811 18955
rect 25222 18952 25228 18964
rect 23799 18924 25228 18952
rect 23799 18921 23811 18924
rect 23753 18915 23811 18921
rect 20640 18856 20944 18884
rect 22848 18884 22876 18912
rect 23768 18884 23796 18915
rect 25222 18912 25228 18924
rect 25280 18912 25286 18964
rect 25314 18912 25320 18964
rect 25372 18952 25378 18964
rect 28534 18952 28540 18964
rect 25372 18924 28540 18952
rect 25372 18912 25378 18924
rect 28534 18912 28540 18924
rect 28592 18912 28598 18964
rect 28810 18912 28816 18964
rect 28868 18952 28874 18964
rect 28911 18955 28969 18961
rect 28911 18952 28923 18955
rect 28868 18924 28923 18952
rect 28868 18912 28874 18924
rect 28911 18921 28923 18924
rect 28957 18921 28969 18955
rect 28911 18915 28969 18921
rect 29270 18912 29276 18964
rect 29328 18952 29334 18964
rect 30285 18955 30343 18961
rect 30285 18952 30297 18955
rect 29328 18924 30297 18952
rect 29328 18912 29334 18924
rect 30285 18921 30297 18924
rect 30331 18921 30343 18955
rect 30285 18915 30343 18921
rect 22848 18856 23796 18884
rect 20640 18828 20668 18856
rect 25590 18844 25596 18896
rect 25648 18884 25654 18896
rect 25648 18856 26648 18884
rect 28106 18870 28580 18884
rect 25648 18844 25654 18856
rect 20257 18819 20315 18825
rect 20257 18785 20269 18819
rect 20303 18785 20315 18819
rect 20257 18779 20315 18785
rect 20438 18776 20444 18828
rect 20496 18816 20502 18828
rect 20533 18819 20591 18825
rect 20533 18816 20545 18819
rect 20496 18788 20545 18816
rect 20496 18776 20502 18788
rect 20533 18785 20545 18788
rect 20579 18785 20591 18819
rect 20533 18779 20591 18785
rect 20622 18776 20628 18828
rect 20680 18776 20686 18828
rect 23017 18819 23075 18825
rect 23017 18816 23029 18819
rect 20916 18788 23029 18816
rect 12391 18753 12449 18759
rect 11532 18720 11928 18748
rect 11164 18680 11192 18708
rect 10428 18652 11192 18680
rect 11701 18683 11759 18689
rect 11701 18649 11713 18683
rect 11747 18680 11759 18683
rect 11790 18680 11796 18692
rect 11747 18652 11796 18680
rect 11747 18649 11759 18652
rect 11701 18643 11759 18649
rect 11790 18640 11796 18652
rect 11848 18640 11854 18692
rect 5583 18584 7420 18612
rect 8404 18612 8432 18640
rect 9398 18612 9404 18624
rect 8404 18584 9404 18612
rect 5583 18581 5595 18584
rect 5537 18575 5595 18581
rect 9398 18572 9404 18584
rect 9456 18572 9462 18624
rect 11900 18612 11928 18720
rect 12391 18719 12403 18753
rect 12437 18719 12449 18753
rect 12391 18713 12449 18719
rect 14277 18751 14335 18757
rect 14277 18717 14289 18751
rect 14323 18748 14335 18751
rect 15838 18748 15844 18760
rect 14323 18720 15844 18748
rect 14323 18717 14335 18720
rect 14277 18711 14335 18717
rect 15838 18708 15844 18720
rect 15896 18708 15902 18760
rect 15948 18748 15976 18776
rect 16117 18751 16175 18757
rect 16117 18748 16129 18751
rect 15948 18720 16129 18748
rect 16117 18717 16129 18720
rect 16163 18717 16175 18751
rect 19702 18748 19708 18760
rect 16117 18711 16175 18717
rect 18800 18720 19708 18748
rect 12618 18612 12624 18624
rect 11900 18584 12624 18612
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 15841 18615 15899 18621
rect 15841 18581 15853 18615
rect 15887 18612 15899 18615
rect 18800 18612 18828 18720
rect 19702 18708 19708 18720
rect 19760 18708 19766 18760
rect 19981 18751 20039 18757
rect 19981 18717 19993 18751
rect 20027 18748 20039 18751
rect 20916 18748 20944 18788
rect 23017 18785 23029 18788
rect 23063 18785 23075 18819
rect 23017 18779 23075 18785
rect 23661 18819 23719 18825
rect 23661 18785 23673 18819
rect 23707 18816 23719 18819
rect 23707 18788 24348 18816
rect 23707 18785 23719 18788
rect 23661 18779 23719 18785
rect 24320 18760 24348 18788
rect 24394 18776 24400 18828
rect 24452 18825 24458 18828
rect 24452 18819 24506 18825
rect 24452 18785 24460 18819
rect 24494 18785 24506 18819
rect 25958 18816 25964 18828
rect 24452 18779 24506 18785
rect 24780 18788 25964 18816
rect 24452 18776 24458 18779
rect 20027 18720 20944 18748
rect 20027 18717 20039 18720
rect 19981 18711 20039 18717
rect 21266 18708 21272 18760
rect 21324 18708 21330 18760
rect 21542 18708 21548 18760
rect 21600 18708 21606 18760
rect 24118 18708 24124 18760
rect 24176 18708 24182 18760
rect 24302 18708 24308 18760
rect 24360 18708 24366 18760
rect 24627 18751 24685 18757
rect 24627 18717 24639 18751
rect 24673 18748 24685 18751
rect 24780 18748 24808 18788
rect 25958 18776 25964 18788
rect 26016 18776 26022 18828
rect 26510 18776 26516 18828
rect 26568 18816 26574 18828
rect 26620 18825 26648 18856
rect 28092 18856 28580 18870
rect 26605 18819 26663 18825
rect 26605 18816 26617 18819
rect 26568 18788 26617 18816
rect 26568 18776 26574 18788
rect 26605 18785 26617 18788
rect 26651 18785 26663 18819
rect 26605 18779 26663 18785
rect 24673 18720 24808 18748
rect 24673 18717 24685 18720
rect 24627 18711 24685 18717
rect 24854 18708 24860 18760
rect 24912 18708 24918 18760
rect 25222 18708 25228 18760
rect 25280 18748 25286 18760
rect 26234 18748 26240 18760
rect 25280 18720 26240 18748
rect 25280 18708 25286 18720
rect 26234 18708 26240 18720
rect 26292 18708 26298 18760
rect 26881 18751 26939 18757
rect 26881 18748 26893 18751
rect 26712 18720 26893 18748
rect 18874 18640 18880 18692
rect 18932 18680 18938 18692
rect 18932 18652 19380 18680
rect 18932 18640 18938 18652
rect 15887 18584 18828 18612
rect 15887 18581 15899 18584
rect 15841 18575 15899 18581
rect 19058 18572 19064 18624
rect 19116 18612 19122 18624
rect 19245 18615 19303 18621
rect 19245 18612 19257 18615
rect 19116 18584 19257 18612
rect 19116 18572 19122 18584
rect 19245 18581 19257 18584
rect 19291 18581 19303 18615
rect 19352 18612 19380 18652
rect 20438 18640 20444 18692
rect 20496 18680 20502 18692
rect 21284 18680 21312 18708
rect 20496 18652 21312 18680
rect 23676 18652 23888 18680
rect 20496 18640 20502 18652
rect 20625 18615 20683 18621
rect 20625 18612 20637 18615
rect 19352 18584 20637 18612
rect 19245 18575 19303 18581
rect 20625 18581 20637 18584
rect 20671 18581 20683 18615
rect 20625 18575 20683 18581
rect 20990 18572 20996 18624
rect 21048 18612 21054 18624
rect 23676 18612 23704 18652
rect 21048 18584 23704 18612
rect 23860 18612 23888 18652
rect 25590 18640 25596 18692
rect 25648 18680 25654 18692
rect 26712 18680 26740 18720
rect 26881 18717 26893 18720
rect 26927 18748 26939 18751
rect 27614 18748 27620 18760
rect 26927 18720 27620 18748
rect 26927 18717 26939 18720
rect 26881 18711 26939 18717
rect 27614 18708 27620 18720
rect 27672 18708 27678 18760
rect 25648 18652 26740 18680
rect 25648 18640 25654 18652
rect 24762 18612 24768 18624
rect 23860 18584 24768 18612
rect 21048 18572 21054 18584
rect 24762 18572 24768 18584
rect 24820 18572 24826 18624
rect 24854 18572 24860 18624
rect 24912 18612 24918 18624
rect 25866 18612 25872 18624
rect 24912 18584 25872 18612
rect 24912 18572 24918 18584
rect 25866 18572 25872 18584
rect 25924 18572 25930 18624
rect 25958 18572 25964 18624
rect 26016 18572 26022 18624
rect 26050 18572 26056 18624
rect 26108 18612 26114 18624
rect 28092 18612 28120 18856
rect 28442 18776 28448 18828
rect 28500 18776 28506 18828
rect 28552 18816 28580 18856
rect 29270 18816 29276 18828
rect 28552 18788 29276 18816
rect 29270 18776 29276 18788
rect 29328 18816 29334 18828
rect 30006 18816 30012 18828
rect 29328 18788 30012 18816
rect 29328 18776 29334 18788
rect 30006 18776 30012 18788
rect 30064 18776 30070 18828
rect 28902 18708 28908 18760
rect 28960 18708 28966 18760
rect 29178 18708 29184 18760
rect 29236 18708 29242 18760
rect 26108 18584 28120 18612
rect 26108 18572 26114 18584
rect 28350 18572 28356 18624
rect 28408 18572 28414 18624
rect 552 18522 30912 18544
rect 552 18470 4193 18522
rect 4245 18470 4257 18522
rect 4309 18470 4321 18522
rect 4373 18470 4385 18522
rect 4437 18470 4449 18522
rect 4501 18470 11783 18522
rect 11835 18470 11847 18522
rect 11899 18470 11911 18522
rect 11963 18470 11975 18522
rect 12027 18470 12039 18522
rect 12091 18470 19373 18522
rect 19425 18470 19437 18522
rect 19489 18470 19501 18522
rect 19553 18470 19565 18522
rect 19617 18470 19629 18522
rect 19681 18470 26963 18522
rect 27015 18470 27027 18522
rect 27079 18470 27091 18522
rect 27143 18470 27155 18522
rect 27207 18470 27219 18522
rect 27271 18470 30912 18522
rect 552 18448 30912 18470
rect 1118 18368 1124 18420
rect 1176 18408 1182 18420
rect 2961 18411 3019 18417
rect 1176 18380 2912 18408
rect 1176 18368 1182 18380
rect 842 18232 848 18284
rect 900 18272 906 18284
rect 937 18275 995 18281
rect 937 18272 949 18275
rect 900 18244 949 18272
rect 900 18232 906 18244
rect 937 18241 949 18244
rect 983 18241 995 18275
rect 1673 18275 1731 18281
rect 1448 18263 1624 18272
rect 937 18235 995 18241
rect 1433 18257 1624 18263
rect 1433 18223 1445 18257
rect 1479 18244 1624 18257
rect 1479 18223 1491 18244
rect 1433 18217 1491 18223
rect 1596 18204 1624 18244
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 2682 18272 2688 18284
rect 1719 18244 2688 18272
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 2682 18232 2688 18244
rect 2740 18232 2746 18284
rect 2884 18272 2912 18380
rect 2961 18377 2973 18411
rect 3007 18408 3019 18411
rect 4062 18408 4068 18420
rect 3007 18380 4068 18408
rect 3007 18377 3019 18380
rect 2961 18371 3019 18377
rect 4062 18368 4068 18380
rect 4120 18368 4126 18420
rect 4154 18368 4160 18420
rect 4212 18408 4218 18420
rect 5905 18411 5963 18417
rect 4212 18380 5856 18408
rect 4212 18368 4218 18380
rect 3418 18300 3424 18352
rect 3476 18340 3482 18352
rect 3513 18343 3571 18349
rect 3513 18340 3525 18343
rect 3476 18312 3525 18340
rect 3476 18300 3482 18312
rect 3513 18309 3525 18312
rect 3559 18340 3571 18343
rect 3559 18312 3924 18340
rect 3559 18309 3571 18312
rect 3513 18303 3571 18309
rect 3896 18272 3924 18312
rect 4062 18272 4068 18284
rect 2884 18244 3740 18272
rect 3896 18244 4068 18272
rect 3712 18216 3740 18244
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 4387 18275 4445 18281
rect 4387 18241 4399 18275
rect 4433 18272 4445 18275
rect 4433 18244 5672 18272
rect 4433 18241 4445 18244
rect 4387 18235 4445 18241
rect 5644 18216 5672 18244
rect 1596 18176 3188 18204
rect 3160 18080 3188 18176
rect 3326 18164 3332 18216
rect 3384 18164 3390 18216
rect 3694 18164 3700 18216
rect 3752 18204 3758 18216
rect 3881 18207 3939 18213
rect 3881 18204 3893 18207
rect 3752 18176 3893 18204
rect 3752 18164 3758 18176
rect 3881 18173 3893 18176
rect 3927 18173 3939 18207
rect 3881 18167 3939 18173
rect 4614 18164 4620 18216
rect 4672 18164 4678 18216
rect 5626 18164 5632 18216
rect 5684 18164 5690 18216
rect 5828 18204 5856 18380
rect 5905 18377 5917 18411
rect 5951 18408 5963 18411
rect 6454 18408 6460 18420
rect 5951 18380 6460 18408
rect 5951 18377 5963 18380
rect 5905 18371 5963 18377
rect 6454 18368 6460 18380
rect 6512 18368 6518 18420
rect 9766 18408 9772 18420
rect 8220 18380 9772 18408
rect 8220 18352 8248 18380
rect 9766 18368 9772 18380
rect 9824 18368 9830 18420
rect 10597 18411 10655 18417
rect 10597 18377 10609 18411
rect 10643 18408 10655 18411
rect 11054 18408 11060 18420
rect 10643 18380 11060 18408
rect 10643 18377 10655 18380
rect 10597 18371 10655 18377
rect 11054 18368 11060 18380
rect 11112 18368 11118 18420
rect 13081 18411 13139 18417
rect 13081 18408 13093 18411
rect 11164 18380 13093 18408
rect 8202 18300 8208 18352
rect 8260 18300 8266 18352
rect 11164 18340 11192 18380
rect 13081 18377 13093 18380
rect 13127 18377 13139 18411
rect 13081 18371 13139 18377
rect 13354 18368 13360 18420
rect 13412 18408 13418 18420
rect 14093 18411 14151 18417
rect 14093 18408 14105 18411
rect 13412 18380 14105 18408
rect 13412 18368 13418 18380
rect 14093 18377 14105 18380
rect 14139 18377 14151 18411
rect 20070 18408 20076 18420
rect 14093 18371 14151 18377
rect 14200 18380 16344 18408
rect 11072 18312 11192 18340
rect 11072 18284 11100 18312
rect 13538 18300 13544 18352
rect 13596 18340 13602 18352
rect 14200 18340 14228 18380
rect 16316 18349 16344 18380
rect 18616 18380 20076 18408
rect 13596 18312 14228 18340
rect 16301 18343 16359 18349
rect 13596 18300 13602 18312
rect 16301 18309 16313 18343
rect 16347 18309 16359 18343
rect 16301 18303 16359 18309
rect 5994 18232 6000 18284
rect 6052 18272 6058 18284
rect 6552 18275 6610 18281
rect 6552 18272 6564 18275
rect 6052 18244 6564 18272
rect 6052 18232 6058 18244
rect 6552 18241 6564 18244
rect 6598 18241 6610 18275
rect 6552 18235 6610 18241
rect 9030 18232 9036 18284
rect 9088 18272 9094 18284
rect 9088 18244 9133 18272
rect 9088 18232 9094 18244
rect 11054 18232 11060 18284
rect 11112 18232 11118 18284
rect 11747 18275 11805 18281
rect 11747 18241 11759 18275
rect 11793 18272 11805 18275
rect 14924 18273 14982 18279
rect 11793 18244 14596 18272
rect 11793 18241 11805 18244
rect 11747 18235 11805 18241
rect 5902 18204 5908 18216
rect 5828 18176 5908 18204
rect 5902 18164 5908 18176
rect 5960 18204 5966 18216
rect 6089 18207 6147 18213
rect 6089 18204 6101 18207
rect 5960 18176 6101 18204
rect 5960 18164 5966 18176
rect 6089 18173 6101 18176
rect 6135 18173 6147 18207
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6089 18167 6147 18173
rect 6196 18176 6837 18204
rect 5350 18096 5356 18148
rect 5408 18136 5414 18148
rect 6196 18136 6224 18176
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 6825 18167 6883 18173
rect 8570 18164 8576 18216
rect 8628 18164 8634 18216
rect 9306 18164 9312 18216
rect 9364 18164 9370 18216
rect 10962 18164 10968 18216
rect 11020 18164 11026 18216
rect 11238 18164 11244 18216
rect 11296 18164 11302 18216
rect 11514 18164 11520 18216
rect 11572 18204 11578 18216
rect 11977 18207 12035 18213
rect 11977 18204 11989 18207
rect 11572 18176 11989 18204
rect 11572 18164 11578 18176
rect 11977 18173 11989 18176
rect 12023 18173 12035 18207
rect 11977 18167 12035 18173
rect 13814 18164 13820 18216
rect 13872 18164 13878 18216
rect 13906 18164 13912 18216
rect 13964 18204 13970 18216
rect 14001 18207 14059 18213
rect 14001 18204 14013 18207
rect 13964 18176 14013 18204
rect 13964 18164 13970 18176
rect 14001 18173 14013 18176
rect 14047 18173 14059 18207
rect 14001 18167 14059 18173
rect 14461 18207 14519 18213
rect 14461 18173 14473 18207
rect 14507 18173 14519 18207
rect 14568 18204 14596 18244
rect 14924 18239 14936 18273
rect 14970 18272 14982 18273
rect 15010 18272 15016 18284
rect 14970 18244 15016 18272
rect 14970 18239 14982 18244
rect 14924 18233 14982 18239
rect 15010 18232 15016 18244
rect 15068 18232 15074 18284
rect 15378 18272 15384 18284
rect 15120 18244 15384 18272
rect 15120 18204 15148 18244
rect 15378 18232 15384 18244
rect 15436 18232 15442 18284
rect 15838 18232 15844 18284
rect 15896 18272 15902 18284
rect 17034 18272 17040 18284
rect 15896 18244 17040 18272
rect 15896 18232 15902 18244
rect 17034 18232 17040 18244
rect 17092 18232 17098 18284
rect 17129 18275 17187 18281
rect 17129 18241 17141 18275
rect 17175 18272 17187 18275
rect 18616 18272 18644 18380
rect 20070 18368 20076 18380
rect 20128 18368 20134 18420
rect 20257 18411 20315 18417
rect 20257 18377 20269 18411
rect 20303 18408 20315 18411
rect 20530 18408 20536 18420
rect 20303 18380 20536 18408
rect 20303 18377 20315 18380
rect 20257 18371 20315 18377
rect 20530 18368 20536 18380
rect 20588 18368 20594 18420
rect 21174 18408 21180 18420
rect 20640 18380 21180 18408
rect 19702 18300 19708 18352
rect 19760 18340 19766 18352
rect 20640 18340 20668 18380
rect 21174 18368 21180 18380
rect 21232 18368 21238 18420
rect 21726 18368 21732 18420
rect 21784 18408 21790 18420
rect 23569 18411 23627 18417
rect 23569 18408 23581 18411
rect 21784 18380 23581 18408
rect 21784 18368 21790 18380
rect 23569 18377 23581 18380
rect 23615 18377 23627 18411
rect 23569 18371 23627 18377
rect 23845 18411 23903 18417
rect 23845 18377 23857 18411
rect 23891 18408 23903 18411
rect 26878 18408 26884 18420
rect 23891 18380 26884 18408
rect 23891 18377 23903 18380
rect 23845 18371 23903 18377
rect 26878 18368 26884 18380
rect 26936 18368 26942 18420
rect 28000 18380 29592 18408
rect 22833 18343 22891 18349
rect 22833 18340 22845 18343
rect 19760 18312 20668 18340
rect 22066 18312 22845 18340
rect 19760 18300 19766 18312
rect 17175 18244 18644 18272
rect 18693 18275 18751 18281
rect 17175 18241 17187 18244
rect 17129 18235 17187 18241
rect 18693 18241 18705 18275
rect 18739 18272 18751 18275
rect 18874 18272 18880 18284
rect 18739 18244 18880 18272
rect 18739 18241 18751 18244
rect 18693 18235 18751 18241
rect 14568 18176 15148 18204
rect 15197 18207 15255 18213
rect 14461 18167 14519 18173
rect 15197 18173 15209 18207
rect 15243 18204 15255 18207
rect 15286 18204 15292 18216
rect 15243 18176 15292 18204
rect 15243 18173 15255 18176
rect 15197 18167 15255 18173
rect 5408 18108 6224 18136
rect 8205 18139 8263 18145
rect 5408 18096 5414 18108
rect 8205 18105 8217 18139
rect 8251 18136 8263 18139
rect 8386 18136 8392 18148
rect 8251 18108 8392 18136
rect 8251 18105 8263 18108
rect 8205 18099 8263 18105
rect 8386 18096 8392 18108
rect 8444 18096 8450 18148
rect 11146 18096 11152 18148
rect 11204 18096 11210 18148
rect 13170 18096 13176 18148
rect 13228 18136 13234 18148
rect 13633 18139 13691 18145
rect 13633 18136 13645 18139
rect 13228 18108 13645 18136
rect 13228 18096 13234 18108
rect 13633 18105 13645 18108
rect 13679 18105 13691 18139
rect 13832 18136 13860 18164
rect 14476 18136 14504 18167
rect 15286 18164 15292 18176
rect 15344 18164 15350 18216
rect 16853 18207 16911 18213
rect 16853 18173 16865 18207
rect 16899 18204 16911 18207
rect 18046 18204 18052 18216
rect 16899 18176 18052 18204
rect 16899 18173 16911 18176
rect 16853 18167 16911 18173
rect 18046 18164 18052 18176
rect 18104 18204 18110 18216
rect 18708 18204 18736 18235
rect 18874 18232 18880 18244
rect 18932 18232 18938 18284
rect 18969 18275 19027 18281
rect 18969 18241 18981 18275
rect 19015 18272 19027 18275
rect 19058 18272 19064 18284
rect 19015 18244 19064 18272
rect 19015 18241 19027 18244
rect 18969 18235 19027 18241
rect 19058 18232 19064 18244
rect 19116 18232 19122 18284
rect 20806 18272 20812 18284
rect 19168 18244 20812 18272
rect 19168 18204 19196 18244
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 21131 18275 21189 18281
rect 21131 18241 21143 18275
rect 21177 18272 21189 18275
rect 21361 18275 21419 18281
rect 21177 18244 21312 18272
rect 21177 18241 21189 18244
rect 21131 18235 21189 18241
rect 18104 18176 18736 18204
rect 18800 18176 19196 18204
rect 20625 18207 20683 18213
rect 18104 18164 18110 18176
rect 18800 18136 18828 18176
rect 20625 18173 20637 18207
rect 20671 18204 20683 18207
rect 20714 18204 20720 18216
rect 20671 18176 20720 18204
rect 20671 18173 20683 18176
rect 20625 18167 20683 18173
rect 20714 18164 20720 18176
rect 20772 18164 20778 18216
rect 21284 18204 21312 18244
rect 21361 18241 21373 18275
rect 21407 18272 21419 18275
rect 22066 18272 22094 18312
rect 22833 18309 22845 18312
rect 22879 18309 22891 18343
rect 22833 18303 22891 18309
rect 24578 18300 24584 18352
rect 24636 18300 24642 18352
rect 27062 18340 27068 18352
rect 26252 18312 27068 18340
rect 26252 18284 26280 18312
rect 27062 18300 27068 18312
rect 27120 18300 27126 18352
rect 21407 18244 22094 18272
rect 21407 18241 21419 18244
rect 21361 18235 21419 18241
rect 22646 18232 22652 18284
rect 22704 18272 22710 18284
rect 22704 18244 23336 18272
rect 22704 18232 22710 18244
rect 21284 18176 22048 18204
rect 13832 18108 14504 18136
rect 17788 18108 18828 18136
rect 22020 18136 22048 18176
rect 22922 18164 22928 18216
rect 22980 18204 22986 18216
rect 23308 18213 23336 18244
rect 24486 18232 24492 18284
rect 24544 18272 24550 18284
rect 25038 18272 25044 18284
rect 24544 18244 25044 18272
rect 24544 18232 24550 18244
rect 25038 18232 25044 18244
rect 25096 18232 25102 18284
rect 25363 18275 25421 18281
rect 25363 18241 25375 18275
rect 25409 18272 25421 18275
rect 25958 18272 25964 18284
rect 25409 18244 25964 18272
rect 25409 18241 25421 18244
rect 25363 18235 25421 18241
rect 25958 18232 25964 18244
rect 26016 18232 26022 18284
rect 26234 18232 26240 18284
rect 26292 18232 26298 18284
rect 26510 18232 26516 18284
rect 26568 18272 26574 18284
rect 28000 18272 28028 18380
rect 29012 18281 29040 18380
rect 29564 18352 29592 18380
rect 29546 18300 29552 18352
rect 29604 18300 29610 18352
rect 26568 18244 28028 18272
rect 28997 18275 29055 18281
rect 26568 18232 26574 18244
rect 28997 18241 29009 18275
rect 29043 18241 29055 18275
rect 28997 18235 29055 18241
rect 23017 18207 23075 18213
rect 23017 18204 23029 18207
rect 22980 18176 23029 18204
rect 22980 18164 22986 18176
rect 23017 18173 23029 18176
rect 23063 18173 23075 18207
rect 23017 18167 23075 18173
rect 23293 18207 23351 18213
rect 23293 18173 23305 18207
rect 23339 18173 23351 18207
rect 23293 18167 23351 18173
rect 23658 18164 23664 18216
rect 23716 18204 23722 18216
rect 24029 18207 24087 18213
rect 24029 18204 24041 18207
rect 23716 18176 24041 18204
rect 23716 18164 23722 18176
rect 24029 18173 24041 18176
rect 24075 18173 24087 18207
rect 24029 18167 24087 18173
rect 24136 18176 24808 18204
rect 24136 18136 24164 18176
rect 24780 18148 24808 18176
rect 24854 18164 24860 18216
rect 24912 18164 24918 18216
rect 25498 18204 25504 18216
rect 24964 18176 25504 18204
rect 22020 18108 24164 18136
rect 13633 18099 13691 18105
rect 1403 18071 1461 18077
rect 1403 18037 1415 18071
rect 1449 18068 1461 18071
rect 1670 18068 1676 18080
rect 1449 18040 1676 18068
rect 1449 18037 1461 18040
rect 1403 18031 1461 18037
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 3142 18028 3148 18080
rect 3200 18028 3206 18080
rect 4347 18071 4405 18077
rect 4347 18037 4359 18071
rect 4393 18068 4405 18071
rect 4522 18068 4528 18080
rect 4393 18040 4528 18068
rect 4393 18037 4405 18040
rect 4347 18031 4405 18037
rect 4522 18028 4528 18040
rect 4580 18028 4586 18080
rect 6086 18028 6092 18080
rect 6144 18068 6150 18080
rect 6555 18071 6613 18077
rect 6555 18068 6567 18071
rect 6144 18040 6567 18068
rect 6144 18028 6150 18040
rect 6555 18037 6567 18040
rect 6601 18068 6613 18071
rect 6822 18068 6828 18080
rect 6601 18040 6828 18068
rect 6601 18037 6613 18040
rect 6555 18031 6613 18037
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 9030 18028 9036 18080
rect 9088 18077 9094 18080
rect 9088 18068 9097 18077
rect 9088 18040 9133 18068
rect 9088 18031 9097 18040
rect 9088 18028 9094 18031
rect 9582 18028 9588 18080
rect 9640 18068 9646 18080
rect 11330 18068 11336 18080
rect 9640 18040 11336 18068
rect 9640 18028 9646 18040
rect 11330 18028 11336 18040
rect 11388 18028 11394 18080
rect 11606 18028 11612 18080
rect 11664 18068 11670 18080
rect 11707 18071 11765 18077
rect 11707 18068 11719 18071
rect 11664 18040 11719 18068
rect 11664 18028 11670 18040
rect 11707 18037 11719 18040
rect 11753 18037 11765 18071
rect 11707 18031 11765 18037
rect 12066 18028 12072 18080
rect 12124 18068 12130 18080
rect 12710 18068 12716 18080
rect 12124 18040 12716 18068
rect 12124 18028 12130 18040
rect 12710 18028 12716 18040
rect 12768 18028 12774 18080
rect 12986 18028 12992 18080
rect 13044 18068 13050 18080
rect 13725 18071 13783 18077
rect 13725 18068 13737 18071
rect 13044 18040 13737 18068
rect 13044 18028 13050 18040
rect 13725 18037 13737 18040
rect 13771 18037 13783 18071
rect 13725 18031 13783 18037
rect 14274 18028 14280 18080
rect 14332 18068 14338 18080
rect 14927 18071 14985 18077
rect 14927 18068 14939 18071
rect 14332 18040 14939 18068
rect 14332 18028 14338 18040
rect 14927 18037 14939 18040
rect 14973 18037 14985 18071
rect 14927 18031 14985 18037
rect 15102 18028 15108 18080
rect 15160 18068 15166 18080
rect 17788 18068 17816 18108
rect 24394 18096 24400 18148
rect 24452 18096 24458 18148
rect 24762 18096 24768 18148
rect 24820 18096 24826 18148
rect 15160 18040 17816 18068
rect 18417 18071 18475 18077
rect 15160 18028 15166 18040
rect 18417 18037 18429 18071
rect 18463 18068 18475 18071
rect 19334 18068 19340 18080
rect 18463 18040 19340 18068
rect 18463 18037 18475 18040
rect 18417 18031 18475 18037
rect 19334 18028 19340 18040
rect 19392 18028 19398 18080
rect 21091 18071 21149 18077
rect 21091 18037 21103 18071
rect 21137 18068 21149 18071
rect 21450 18068 21456 18080
rect 21137 18040 21456 18068
rect 21137 18037 21149 18040
rect 21091 18031 21149 18037
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 21818 18028 21824 18080
rect 21876 18068 21882 18080
rect 22465 18071 22523 18077
rect 22465 18068 22477 18071
rect 21876 18040 22477 18068
rect 21876 18028 21882 18040
rect 22465 18037 22477 18040
rect 22511 18037 22523 18071
rect 22465 18031 22523 18037
rect 24026 18028 24032 18080
rect 24084 18068 24090 18080
rect 24964 18068 24992 18176
rect 25498 18164 25504 18176
rect 25556 18164 25562 18216
rect 25593 18207 25651 18213
rect 25593 18173 25605 18207
rect 25639 18204 25651 18207
rect 25639 18176 27016 18204
rect 25639 18173 25651 18176
rect 25593 18167 25651 18173
rect 24084 18040 24992 18068
rect 24084 18028 24090 18040
rect 25222 18028 25228 18080
rect 25280 18068 25286 18080
rect 25323 18071 25381 18077
rect 25323 18068 25335 18071
rect 25280 18040 25335 18068
rect 25280 18028 25286 18040
rect 25323 18037 25335 18040
rect 25369 18037 25381 18071
rect 25323 18031 25381 18037
rect 26694 18028 26700 18080
rect 26752 18028 26758 18080
rect 26988 18068 27016 18176
rect 27062 18164 27068 18216
rect 27120 18164 27126 18216
rect 27154 18164 27160 18216
rect 27212 18204 27218 18216
rect 27341 18207 27399 18213
rect 27341 18204 27353 18207
rect 27212 18176 27353 18204
rect 27212 18164 27218 18176
rect 27341 18173 27353 18176
rect 27387 18173 27399 18207
rect 27341 18167 27399 18173
rect 27614 18164 27620 18216
rect 27672 18204 27678 18216
rect 29273 18207 29331 18213
rect 29273 18204 29285 18207
rect 27672 18201 28954 18204
rect 29012 18201 29285 18204
rect 27672 18176 29285 18201
rect 27672 18164 27678 18176
rect 28926 18173 29040 18176
rect 29273 18173 29285 18176
rect 29319 18204 29331 18207
rect 30561 18207 30619 18213
rect 29319 18176 29960 18204
rect 29319 18173 29331 18176
rect 29273 18167 29331 18173
rect 29932 18148 29960 18176
rect 30561 18173 30573 18207
rect 30607 18204 30619 18207
rect 30607 18176 30696 18204
rect 30607 18173 30619 18176
rect 30561 18167 30619 18173
rect 29362 18136 29368 18148
rect 28368 18108 28994 18136
rect 28368 18068 28396 18108
rect 26988 18040 28396 18068
rect 28442 18028 28448 18080
rect 28500 18028 28506 18080
rect 28966 18068 28994 18108
rect 29104 18108 29368 18136
rect 29104 18068 29132 18108
rect 29362 18096 29368 18108
rect 29420 18096 29426 18148
rect 29914 18096 29920 18148
rect 29972 18096 29978 18148
rect 30668 18080 30696 18176
rect 28966 18040 29132 18068
rect 30098 18028 30104 18080
rect 30156 18028 30162 18080
rect 30190 18028 30196 18080
rect 30248 18068 30254 18080
rect 30285 18071 30343 18077
rect 30285 18068 30297 18071
rect 30248 18040 30297 18068
rect 30248 18028 30254 18040
rect 30285 18037 30297 18040
rect 30331 18037 30343 18071
rect 30285 18031 30343 18037
rect 30374 18028 30380 18080
rect 30432 18028 30438 18080
rect 30650 18028 30656 18080
rect 30708 18028 30714 18080
rect 552 17978 31072 18000
rect 552 17926 7988 17978
rect 8040 17926 8052 17978
rect 8104 17926 8116 17978
rect 8168 17926 8180 17978
rect 8232 17926 8244 17978
rect 8296 17926 15578 17978
rect 15630 17926 15642 17978
rect 15694 17926 15706 17978
rect 15758 17926 15770 17978
rect 15822 17926 15834 17978
rect 15886 17926 23168 17978
rect 23220 17926 23232 17978
rect 23284 17926 23296 17978
rect 23348 17926 23360 17978
rect 23412 17926 23424 17978
rect 23476 17926 30758 17978
rect 30810 17926 30822 17978
rect 30874 17926 30886 17978
rect 30938 17926 30950 17978
rect 31002 17926 31014 17978
rect 31066 17926 31072 17978
rect 552 17904 31072 17926
rect 1029 17867 1087 17873
rect 1029 17833 1041 17867
rect 1075 17864 1087 17867
rect 1075 17836 2774 17864
rect 1075 17833 1087 17836
rect 1029 17827 1087 17833
rect 1118 17756 1124 17808
rect 1176 17796 1182 17808
rect 2746 17796 2774 17836
rect 3142 17824 3148 17876
rect 3200 17824 3206 17876
rect 3979 17867 4037 17873
rect 3979 17833 3991 17867
rect 4025 17864 4037 17867
rect 4522 17864 4528 17876
rect 4025 17836 4528 17864
rect 4025 17833 4037 17836
rect 3979 17827 4037 17833
rect 4522 17824 4528 17836
rect 4580 17824 4586 17876
rect 6822 17824 6828 17876
rect 6880 17864 6886 17876
rect 6923 17867 6981 17873
rect 6923 17864 6935 17867
rect 6880 17836 6935 17864
rect 6880 17824 6886 17836
rect 6923 17833 6935 17836
rect 6969 17833 6981 17867
rect 12066 17864 12072 17876
rect 6923 17827 6981 17833
rect 8496 17836 12072 17864
rect 5629 17799 5687 17805
rect 1176 17768 1348 17796
rect 2746 17768 3372 17796
rect 1176 17756 1182 17768
rect 1320 17737 1348 17768
rect 1670 17737 1676 17740
rect 1213 17731 1271 17737
rect 1213 17697 1225 17731
rect 1259 17697 1271 17731
rect 1213 17691 1271 17697
rect 1305 17731 1363 17737
rect 1305 17697 1317 17731
rect 1351 17697 1363 17731
rect 1305 17691 1363 17697
rect 1632 17731 1676 17737
rect 1632 17697 1644 17731
rect 1632 17691 1676 17697
rect 1228 17524 1256 17691
rect 1670 17688 1676 17691
rect 1728 17688 1734 17740
rect 3142 17728 3148 17740
rect 1964 17700 3148 17728
rect 1801 17681 1859 17687
rect 1801 17647 1813 17681
rect 1847 17660 1859 17681
rect 1964 17660 1992 17700
rect 3142 17688 3148 17700
rect 3200 17688 3206 17740
rect 1847 17647 1992 17660
rect 1801 17641 1992 17647
rect 1826 17632 1992 17641
rect 2038 17620 2044 17672
rect 2096 17620 2102 17672
rect 3234 17524 3240 17536
rect 1228 17496 3240 17524
rect 3234 17484 3240 17496
rect 3292 17484 3298 17536
rect 3344 17524 3372 17768
rect 5629 17765 5641 17799
rect 5675 17796 5687 17799
rect 5994 17796 6000 17808
rect 5675 17768 6000 17796
rect 5675 17765 5687 17768
rect 5629 17759 5687 17765
rect 5994 17756 6000 17768
rect 6052 17756 6058 17808
rect 5905 17731 5963 17737
rect 4172 17700 5856 17728
rect 3513 17663 3571 17669
rect 3513 17629 3525 17663
rect 3559 17660 3571 17663
rect 3694 17660 3700 17672
rect 3559 17632 3700 17660
rect 3559 17629 3571 17632
rect 3513 17623 3571 17629
rect 3694 17620 3700 17632
rect 3752 17620 3758 17672
rect 4019 17663 4077 17669
rect 4019 17629 4031 17663
rect 4065 17660 4077 17663
rect 4172 17660 4200 17700
rect 5828 17672 5856 17700
rect 5905 17697 5917 17731
rect 5951 17728 5963 17731
rect 6546 17728 6552 17740
rect 5951 17700 6552 17728
rect 5951 17697 5963 17700
rect 5905 17691 5963 17697
rect 6546 17688 6552 17700
rect 6604 17688 6610 17740
rect 8496 17728 8524 17836
rect 12066 17824 12072 17836
rect 12124 17824 12130 17876
rect 12250 17824 12256 17876
rect 12308 17864 12314 17876
rect 12802 17864 12808 17876
rect 12308 17836 12808 17864
rect 12308 17824 12314 17836
rect 12802 17824 12808 17836
rect 12860 17824 12866 17876
rect 14274 17824 14280 17876
rect 14332 17873 14338 17876
rect 14332 17864 14341 17873
rect 14332 17836 14377 17864
rect 14332 17827 14341 17836
rect 14332 17824 14338 17827
rect 15378 17824 15384 17876
rect 15436 17864 15442 17876
rect 15657 17867 15715 17873
rect 15657 17864 15669 17867
rect 15436 17836 15669 17864
rect 15436 17824 15442 17836
rect 15657 17833 15669 17836
rect 15703 17833 15715 17867
rect 15657 17827 15715 17833
rect 16114 17824 16120 17876
rect 16172 17864 16178 17876
rect 16172 17836 16252 17864
rect 16172 17824 16178 17836
rect 10778 17756 10784 17808
rect 10836 17756 10842 17808
rect 15562 17756 15568 17808
rect 15620 17796 15626 17808
rect 16224 17805 16252 17836
rect 16574 17824 16580 17876
rect 16632 17864 16638 17876
rect 17037 17867 17095 17873
rect 17037 17864 17049 17867
rect 16632 17836 17049 17864
rect 16632 17824 16638 17836
rect 17037 17833 17049 17836
rect 17083 17833 17095 17867
rect 17770 17864 17776 17876
rect 17037 17827 17095 17833
rect 17236 17836 17776 17864
rect 16209 17799 16267 17805
rect 16209 17796 16221 17799
rect 15620 17768 16221 17796
rect 15620 17756 15626 17768
rect 16209 17765 16221 17768
rect 16255 17765 16267 17799
rect 16209 17759 16267 17765
rect 7208 17700 8524 17728
rect 8573 17731 8631 17737
rect 4065 17632 4200 17660
rect 4249 17663 4307 17669
rect 4065 17629 4077 17632
rect 4019 17623 4077 17629
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 5258 17660 5264 17672
rect 4295 17632 5264 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 5258 17620 5264 17632
rect 5316 17620 5322 17672
rect 5810 17620 5816 17672
rect 5868 17620 5874 17672
rect 6362 17620 6368 17672
rect 6420 17620 6426 17672
rect 6454 17620 6460 17672
rect 6512 17620 6518 17672
rect 6914 17620 6920 17672
rect 6972 17620 6978 17672
rect 7208 17669 7236 17700
rect 8573 17697 8585 17731
rect 8619 17728 8631 17731
rect 8619 17700 9171 17728
rect 8619 17697 8631 17700
rect 8573 17691 8631 17697
rect 7193 17663 7251 17669
rect 7193 17629 7205 17663
rect 7239 17629 7251 17663
rect 7193 17623 7251 17629
rect 8662 17620 8668 17672
rect 8720 17620 8726 17672
rect 9030 17669 9036 17672
rect 8992 17663 9036 17669
rect 8992 17629 9004 17663
rect 8992 17623 9036 17629
rect 9030 17620 9036 17623
rect 9088 17620 9094 17672
rect 9143 17671 9171 17700
rect 10318 17688 10324 17740
rect 10376 17728 10382 17740
rect 11606 17737 11612 17740
rect 11149 17731 11207 17737
rect 11149 17728 11161 17731
rect 10376 17700 11161 17728
rect 10376 17688 10382 17700
rect 11149 17697 11161 17700
rect 11195 17697 11207 17731
rect 11149 17691 11207 17697
rect 11568 17731 11612 17737
rect 11568 17697 11580 17731
rect 11568 17691 11612 17697
rect 9128 17665 9186 17671
rect 9128 17631 9140 17665
rect 9174 17631 9186 17665
rect 9128 17625 9186 17631
rect 9398 17620 9404 17672
rect 9456 17620 9462 17672
rect 6380 17592 6408 17620
rect 4908 17564 6408 17592
rect 4908 17524 4936 17564
rect 3344 17496 4936 17524
rect 6181 17527 6239 17533
rect 6181 17493 6193 17527
rect 6227 17524 6239 17527
rect 9858 17524 9864 17536
rect 6227 17496 9864 17524
rect 6227 17493 6239 17496
rect 6181 17487 6239 17493
rect 9858 17484 9864 17496
rect 9916 17484 9922 17536
rect 10962 17484 10968 17536
rect 11020 17484 11026 17536
rect 11164 17524 11192 17691
rect 11606 17688 11612 17691
rect 11664 17688 11670 17740
rect 11762 17700 13032 17728
rect 11238 17620 11244 17672
rect 11296 17620 11302 17672
rect 11762 17671 11790 17700
rect 11747 17665 11805 17671
rect 11747 17631 11759 17665
rect 11793 17631 11805 17665
rect 11747 17625 11805 17631
rect 11882 17620 11888 17672
rect 11940 17660 11946 17672
rect 11977 17663 12035 17669
rect 11977 17660 11989 17663
rect 11940 17632 11989 17660
rect 11940 17620 11946 17632
rect 11977 17629 11989 17632
rect 12023 17629 12035 17663
rect 11977 17623 12035 17629
rect 12066 17620 12072 17672
rect 12124 17660 12130 17672
rect 12894 17660 12900 17672
rect 12124 17632 12900 17660
rect 12124 17620 12130 17632
rect 12894 17620 12900 17632
rect 12952 17620 12958 17672
rect 13004 17660 13032 17700
rect 13262 17688 13268 17740
rect 13320 17728 13326 17740
rect 13449 17731 13507 17737
rect 13449 17728 13461 17731
rect 13320 17700 13461 17728
rect 13320 17688 13326 17700
rect 13449 17697 13461 17700
rect 13495 17697 13507 17731
rect 16114 17728 16120 17740
rect 13449 17691 13507 17697
rect 14476 17700 16120 17728
rect 13004 17632 13768 17660
rect 12986 17524 12992 17536
rect 11164 17496 12992 17524
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 13078 17484 13084 17536
rect 13136 17484 13142 17536
rect 13630 17484 13636 17536
rect 13688 17484 13694 17536
rect 13740 17524 13768 17632
rect 13814 17620 13820 17672
rect 13872 17620 13878 17672
rect 14323 17663 14381 17669
rect 14323 17629 14335 17663
rect 14369 17660 14381 17663
rect 14476 17660 14504 17700
rect 16114 17688 16120 17700
rect 16172 17688 16178 17740
rect 16574 17688 16580 17740
rect 16632 17688 16638 17740
rect 16945 17731 17003 17737
rect 16945 17697 16957 17731
rect 16991 17728 17003 17731
rect 17236 17728 17264 17836
rect 17770 17824 17776 17836
rect 17828 17824 17834 17876
rect 21634 17864 21640 17876
rect 19260 17836 21640 17864
rect 19260 17728 19288 17836
rect 21634 17824 21640 17836
rect 21692 17824 21698 17876
rect 23014 17824 23020 17876
rect 23072 17864 23078 17876
rect 24578 17864 24584 17876
rect 23072 17836 24584 17864
rect 23072 17824 23078 17836
rect 24578 17824 24584 17836
rect 24636 17824 24642 17876
rect 24762 17824 24768 17876
rect 24820 17864 24826 17876
rect 25961 17867 26019 17873
rect 25961 17864 25973 17867
rect 24820 17836 25973 17864
rect 24820 17824 24826 17836
rect 25961 17833 25973 17836
rect 26007 17833 26019 17867
rect 25961 17827 26019 17833
rect 27430 17824 27436 17876
rect 27488 17864 27494 17876
rect 27801 17867 27859 17873
rect 27801 17864 27813 17867
rect 27488 17836 27813 17864
rect 27488 17824 27494 17836
rect 27801 17833 27813 17836
rect 27847 17833 27859 17867
rect 28810 17864 28816 17876
rect 28868 17873 28874 17876
rect 27801 17827 27859 17833
rect 27908 17836 28816 17864
rect 23584 17768 24164 17796
rect 16991 17700 17264 17728
rect 17788 17700 19288 17728
rect 16991 17697 17003 17700
rect 16945 17691 17003 17697
rect 14369 17632 14504 17660
rect 14553 17663 14611 17669
rect 14369 17629 14381 17632
rect 14323 17623 14381 17629
rect 14553 17629 14565 17663
rect 14599 17660 14611 17663
rect 16666 17660 16672 17672
rect 14599 17632 16672 17660
rect 14599 17629 14611 17632
rect 14553 17623 14611 17629
rect 16666 17620 16672 17632
rect 16724 17620 16730 17672
rect 17034 17620 17040 17672
rect 17092 17660 17098 17672
rect 17494 17669 17500 17672
rect 17129 17663 17187 17669
rect 17129 17660 17141 17663
rect 17092 17632 17141 17660
rect 17092 17620 17098 17632
rect 17129 17629 17141 17632
rect 17175 17629 17187 17663
rect 17129 17623 17187 17629
rect 17456 17663 17500 17669
rect 17456 17629 17468 17663
rect 17456 17623 17500 17629
rect 17494 17620 17500 17623
rect 17552 17620 17558 17672
rect 17635 17663 17693 17669
rect 17635 17629 17647 17663
rect 17681 17660 17693 17663
rect 17788 17660 17816 17700
rect 19334 17688 19340 17740
rect 19392 17728 19398 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 19392 17700 19717 17728
rect 19392 17688 19398 17700
rect 19705 17697 19717 17700
rect 19751 17697 19763 17731
rect 19705 17691 19763 17697
rect 21085 17731 21143 17737
rect 21085 17697 21097 17731
rect 21131 17728 21143 17731
rect 23584 17728 23612 17768
rect 21131 17700 23612 17728
rect 21131 17697 21143 17700
rect 21085 17691 21143 17697
rect 23658 17688 23664 17740
rect 23716 17688 23722 17740
rect 23750 17688 23756 17740
rect 23808 17728 23814 17740
rect 24029 17731 24087 17737
rect 24029 17728 24041 17731
rect 23808 17700 24041 17728
rect 23808 17688 23814 17700
rect 24029 17697 24041 17700
rect 24075 17697 24087 17731
rect 24136 17728 24164 17768
rect 26697 17731 26755 17737
rect 26697 17728 26709 17731
rect 24136 17700 26709 17728
rect 24029 17691 24087 17697
rect 26697 17697 26709 17700
rect 26743 17697 26755 17731
rect 26697 17691 26755 17697
rect 17681 17632 17816 17660
rect 17681 17629 17693 17632
rect 17635 17623 17693 17629
rect 17862 17620 17868 17672
rect 17920 17620 17926 17672
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17660 19487 17663
rect 20438 17660 20444 17672
rect 19475 17632 20444 17660
rect 19475 17629 19487 17632
rect 19429 17623 19487 17629
rect 20438 17620 20444 17632
rect 20496 17620 20502 17672
rect 20714 17620 20720 17672
rect 20772 17660 20778 17672
rect 21269 17663 21327 17669
rect 21269 17660 21281 17663
rect 20772 17632 21281 17660
rect 20772 17620 20778 17632
rect 21269 17629 21281 17632
rect 21315 17629 21327 17663
rect 21269 17623 21327 17629
rect 15470 17524 15476 17536
rect 13740 17496 15476 17524
rect 15470 17484 15476 17496
rect 15528 17484 15534 17536
rect 17586 17484 17592 17536
rect 17644 17524 17650 17536
rect 18969 17527 19027 17533
rect 18969 17524 18981 17527
rect 17644 17496 18981 17524
rect 17644 17484 17650 17496
rect 18969 17493 18981 17496
rect 19015 17493 19027 17527
rect 21284 17524 21312 17623
rect 21450 17620 21456 17672
rect 21508 17660 21514 17672
rect 21596 17663 21654 17669
rect 21596 17660 21608 17663
rect 21508 17632 21608 17660
rect 21508 17620 21514 17632
rect 21596 17629 21608 17632
rect 21642 17629 21654 17663
rect 21596 17623 21654 17629
rect 21775 17663 21833 17669
rect 21775 17629 21787 17663
rect 21821 17660 21833 17663
rect 21910 17660 21916 17672
rect 21821 17632 21916 17660
rect 21821 17629 21833 17632
rect 21775 17623 21833 17629
rect 21910 17620 21916 17632
rect 21968 17620 21974 17672
rect 22005 17663 22063 17669
rect 22005 17629 22017 17663
rect 22051 17660 22063 17663
rect 22051 17632 23520 17660
rect 22051 17629 22063 17632
rect 22005 17623 22063 17629
rect 23492 17601 23520 17632
rect 23566 17620 23572 17672
rect 23624 17660 23630 17672
rect 24486 17669 24492 17672
rect 24121 17663 24179 17669
rect 24121 17660 24133 17663
rect 23624 17632 24133 17660
rect 23624 17620 23630 17632
rect 24121 17629 24133 17632
rect 24167 17629 24179 17663
rect 24121 17623 24179 17629
rect 24448 17663 24492 17669
rect 24448 17629 24460 17663
rect 24448 17623 24492 17629
rect 24486 17620 24492 17623
rect 24544 17620 24550 17672
rect 24584 17665 24642 17671
rect 24584 17631 24596 17665
rect 24630 17660 24642 17665
rect 24670 17660 24676 17672
rect 24630 17632 24676 17660
rect 24630 17631 24642 17632
rect 24584 17625 24642 17631
rect 24670 17620 24676 17632
rect 24728 17620 24734 17672
rect 24854 17620 24860 17672
rect 24912 17620 24918 17672
rect 25038 17620 25044 17672
rect 25096 17660 25102 17672
rect 25096 17632 25544 17660
rect 25096 17620 25102 17632
rect 23477 17595 23535 17601
rect 23477 17561 23489 17595
rect 23523 17561 23535 17595
rect 25516 17592 25544 17632
rect 26418 17620 26424 17672
rect 26476 17620 26482 17672
rect 27338 17620 27344 17672
rect 27396 17660 27402 17672
rect 27908 17660 27936 17836
rect 28810 17824 28816 17836
rect 28868 17864 28877 17873
rect 28868 17836 28913 17864
rect 28868 17827 28877 17836
rect 28868 17824 28874 17827
rect 28994 17824 29000 17876
rect 29052 17864 29058 17876
rect 30193 17867 30251 17873
rect 30193 17864 30205 17867
rect 29052 17836 30205 17864
rect 29052 17824 29058 17836
rect 30193 17833 30205 17836
rect 30239 17833 30251 17867
rect 30193 17827 30251 17833
rect 29012 17700 29960 17728
rect 27396 17632 27936 17660
rect 28353 17663 28411 17669
rect 27396 17620 27402 17632
rect 28353 17629 28365 17663
rect 28399 17660 28411 17663
rect 28534 17660 28540 17672
rect 28399 17632 28540 17660
rect 28399 17629 28411 17632
rect 28353 17623 28411 17629
rect 28534 17620 28540 17632
rect 28592 17620 28598 17672
rect 28859 17663 28917 17669
rect 28859 17629 28871 17663
rect 28905 17660 28917 17663
rect 29012 17660 29040 17700
rect 29932 17672 29960 17700
rect 28905 17632 29040 17660
rect 29089 17663 29147 17669
rect 28905 17629 28917 17632
rect 28859 17623 28917 17629
rect 29089 17629 29101 17663
rect 29135 17660 29147 17663
rect 29730 17660 29736 17672
rect 29135 17632 29736 17660
rect 29135 17629 29147 17632
rect 29089 17623 29147 17629
rect 29730 17620 29736 17632
rect 29788 17620 29794 17672
rect 29914 17620 29920 17672
rect 29972 17620 29978 17672
rect 25516 17564 26464 17592
rect 23477 17555 23535 17561
rect 26436 17536 26464 17564
rect 22002 17524 22008 17536
rect 21284 17496 22008 17524
rect 18969 17487 19027 17493
rect 22002 17484 22008 17496
rect 22060 17484 22066 17536
rect 22738 17484 22744 17536
rect 22796 17524 22802 17536
rect 23109 17527 23167 17533
rect 23109 17524 23121 17527
rect 22796 17496 23121 17524
rect 22796 17484 22802 17496
rect 23109 17493 23121 17496
rect 23155 17493 23167 17527
rect 23109 17487 23167 17493
rect 23845 17527 23903 17533
rect 23845 17493 23857 17527
rect 23891 17524 23903 17527
rect 25498 17524 25504 17536
rect 23891 17496 25504 17524
rect 23891 17493 23903 17496
rect 23845 17487 23903 17493
rect 25498 17484 25504 17496
rect 25556 17484 25562 17536
rect 26418 17484 26424 17536
rect 26476 17484 26482 17536
rect 29270 17484 29276 17536
rect 29328 17524 29334 17536
rect 30098 17524 30104 17536
rect 29328 17496 30104 17524
rect 29328 17484 29334 17496
rect 30098 17484 30104 17496
rect 30156 17484 30162 17536
rect 552 17434 30912 17456
rect 552 17382 4193 17434
rect 4245 17382 4257 17434
rect 4309 17382 4321 17434
rect 4373 17382 4385 17434
rect 4437 17382 4449 17434
rect 4501 17382 11783 17434
rect 11835 17382 11847 17434
rect 11899 17382 11911 17434
rect 11963 17382 11975 17434
rect 12027 17382 12039 17434
rect 12091 17382 19373 17434
rect 19425 17382 19437 17434
rect 19489 17382 19501 17434
rect 19553 17382 19565 17434
rect 19617 17382 19629 17434
rect 19681 17382 26963 17434
rect 27015 17382 27027 17434
rect 27079 17382 27091 17434
rect 27143 17382 27155 17434
rect 27207 17382 27219 17434
rect 27271 17382 30912 17434
rect 552 17360 30912 17382
rect 1578 17280 1584 17332
rect 1636 17320 1642 17332
rect 2777 17323 2835 17329
rect 2777 17320 2789 17323
rect 1636 17292 2789 17320
rect 1636 17280 1642 17292
rect 2777 17289 2789 17292
rect 2823 17289 2835 17323
rect 2777 17283 2835 17289
rect 3234 17280 3240 17332
rect 3292 17320 3298 17332
rect 5905 17323 5963 17329
rect 3292 17292 5856 17320
rect 3292 17280 3298 17292
rect 3694 17212 3700 17264
rect 3752 17212 3758 17264
rect 937 17187 995 17193
rect 937 17153 949 17187
rect 983 17184 995 17187
rect 1118 17184 1124 17196
rect 983 17156 1124 17184
rect 983 17153 995 17156
rect 937 17147 995 17153
rect 1118 17144 1124 17156
rect 1176 17144 1182 17196
rect 1443 17187 1501 17193
rect 1443 17153 1455 17187
rect 1489 17184 1501 17187
rect 2774 17184 2780 17196
rect 1489 17156 2780 17184
rect 1489 17153 1501 17156
rect 1443 17147 1501 17153
rect 2774 17144 2780 17156
rect 2832 17144 2838 17196
rect 3712 17184 3740 17212
rect 3881 17187 3939 17193
rect 3881 17184 3893 17187
rect 3712 17156 3893 17184
rect 3881 17153 3893 17156
rect 3927 17184 3939 17187
rect 4062 17184 4068 17196
rect 3927 17156 4068 17184
rect 3927 17153 3939 17156
rect 3881 17147 3939 17153
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 4387 17187 4445 17193
rect 4387 17153 4399 17187
rect 4433 17184 4445 17187
rect 5534 17184 5540 17196
rect 4433 17156 5540 17184
rect 4433 17153 4445 17156
rect 4387 17147 4445 17153
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17116 1731 17119
rect 2406 17116 2412 17128
rect 1719 17088 2412 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 2406 17076 2412 17088
rect 2464 17076 2470 17128
rect 3234 17076 3240 17128
rect 3292 17076 3298 17128
rect 4617 17119 4675 17125
rect 4617 17085 4629 17119
rect 4663 17116 4675 17119
rect 5074 17116 5080 17128
rect 4663 17088 5080 17116
rect 4663 17085 4675 17088
rect 4617 17079 4675 17085
rect 5074 17076 5080 17088
rect 5132 17076 5138 17128
rect 5828 17116 5856 17292
rect 5905 17289 5917 17323
rect 5951 17320 5963 17323
rect 6914 17320 6920 17332
rect 5951 17292 6920 17320
rect 5951 17289 5963 17292
rect 5905 17283 5963 17289
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 8113 17323 8171 17329
rect 8113 17289 8125 17323
rect 8159 17320 8171 17323
rect 8478 17320 8484 17332
rect 8159 17292 8484 17320
rect 8159 17289 8171 17292
rect 8113 17283 8171 17289
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 10226 17320 10232 17332
rect 8588 17292 10232 17320
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 6089 17187 6147 17193
rect 6089 17184 6101 17187
rect 5960 17156 6101 17184
rect 5960 17144 5966 17156
rect 6089 17153 6101 17156
rect 6135 17184 6147 17187
rect 6454 17184 6460 17196
rect 6135 17156 6460 17184
rect 6135 17153 6147 17156
rect 6089 17147 6147 17153
rect 6454 17144 6460 17156
rect 6512 17144 6518 17196
rect 6546 17144 6552 17196
rect 6604 17184 6610 17196
rect 6825 17187 6883 17193
rect 6604 17156 6649 17184
rect 6604 17144 6610 17156
rect 6825 17153 6837 17187
rect 6871 17184 6883 17187
rect 8386 17184 8392 17196
rect 6871 17156 8392 17184
rect 6871 17153 6883 17156
rect 6825 17147 6883 17153
rect 8386 17144 8392 17156
rect 8444 17144 8450 17196
rect 7466 17116 7472 17128
rect 5828 17088 7472 17116
rect 7466 17076 7472 17088
rect 7524 17076 7530 17128
rect 8588 17125 8616 17292
rect 10226 17280 10232 17292
rect 10284 17280 10290 17332
rect 10502 17280 10508 17332
rect 10560 17280 10566 17332
rect 11514 17320 11520 17332
rect 10612 17292 11520 17320
rect 8662 17144 8668 17196
rect 8720 17144 8726 17196
rect 9030 17193 9036 17196
rect 8992 17187 9036 17193
rect 8992 17153 9004 17187
rect 8992 17147 9036 17153
rect 9030 17144 9036 17147
rect 9088 17144 9094 17196
rect 9122 17144 9128 17196
rect 9180 17191 9186 17196
rect 9180 17185 9229 17191
rect 9180 17151 9183 17185
rect 9217 17151 9229 17185
rect 9180 17145 9229 17151
rect 9401 17187 9459 17193
rect 9401 17153 9413 17187
rect 9447 17184 9459 17187
rect 9582 17184 9588 17196
rect 9447 17156 9588 17184
rect 9447 17153 9459 17156
rect 9401 17147 9459 17153
rect 9180 17144 9186 17145
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17085 8631 17119
rect 10612 17116 10640 17292
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 11698 17280 11704 17332
rect 11756 17320 11762 17332
rect 13725 17323 13783 17329
rect 13725 17320 13737 17323
rect 11756 17292 13737 17320
rect 11756 17280 11762 17292
rect 13725 17289 13737 17292
rect 13771 17289 13783 17323
rect 13725 17283 13783 17289
rect 15194 17280 15200 17332
rect 15252 17320 15258 17332
rect 15565 17323 15623 17329
rect 15565 17320 15577 17323
rect 15252 17292 15577 17320
rect 15252 17280 15258 17292
rect 15565 17289 15577 17292
rect 15611 17289 15623 17323
rect 18233 17323 18291 17329
rect 18233 17320 18245 17323
rect 15565 17283 15623 17289
rect 16040 17292 18245 17320
rect 13262 17212 13268 17264
rect 13320 17252 13326 17264
rect 14093 17255 14151 17261
rect 14093 17252 14105 17255
rect 13320 17224 14105 17252
rect 13320 17212 13326 17224
rect 14093 17221 14105 17224
rect 14139 17221 14151 17255
rect 14093 17215 14151 17221
rect 14458 17212 14464 17264
rect 14516 17212 14522 17264
rect 15378 17212 15384 17264
rect 15436 17252 15442 17264
rect 15933 17255 15991 17261
rect 15933 17252 15945 17255
rect 15436 17224 15945 17252
rect 15436 17212 15442 17224
rect 15933 17221 15945 17224
rect 15979 17221 15991 17255
rect 15933 17215 15991 17221
rect 11790 17191 11796 17196
rect 11747 17185 11796 17191
rect 11747 17151 11759 17185
rect 11793 17151 11796 17185
rect 11747 17145 11796 17151
rect 11790 17144 11796 17145
rect 11848 17144 11854 17196
rect 8573 17079 8631 17085
rect 8772 17088 10640 17116
rect 3513 17051 3571 17057
rect 3513 17017 3525 17051
rect 3559 17017 3571 17051
rect 3513 17011 3571 17017
rect 1403 16983 1461 16989
rect 1403 16949 1415 16983
rect 1449 16980 1461 16983
rect 1762 16980 1768 16992
rect 1449 16952 1768 16980
rect 1449 16949 1461 16952
rect 1403 16943 1461 16949
rect 1762 16940 1768 16952
rect 1820 16980 1826 16992
rect 3528 16980 3556 17011
rect 4347 16983 4405 16989
rect 4347 16980 4359 16983
rect 1820 16952 4359 16980
rect 1820 16940 1826 16952
rect 4347 16949 4359 16952
rect 4393 16980 4405 16983
rect 4522 16980 4528 16992
rect 4393 16952 4528 16980
rect 4393 16949 4405 16952
rect 4347 16943 4405 16949
rect 4522 16940 4528 16952
rect 4580 16980 4586 16992
rect 4982 16980 4988 16992
rect 4580 16952 4988 16980
rect 4580 16940 4586 16952
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 6555 16983 6613 16989
rect 6555 16949 6567 16983
rect 6601 16980 6613 16983
rect 6822 16980 6828 16992
rect 6601 16952 6828 16980
rect 6601 16949 6613 16952
rect 6555 16943 6613 16949
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 8389 16983 8447 16989
rect 8389 16949 8401 16983
rect 8435 16980 8447 16983
rect 8772 16980 8800 17088
rect 10962 17076 10968 17128
rect 11020 17076 11026 17128
rect 11238 17076 11244 17128
rect 11296 17076 11302 17128
rect 11974 17076 11980 17128
rect 12032 17076 12038 17128
rect 13633 17119 13691 17125
rect 13633 17085 13645 17119
rect 13679 17116 13691 17119
rect 13998 17116 14004 17128
rect 13679 17112 13768 17116
rect 13924 17112 14004 17116
rect 13679 17088 14004 17112
rect 13679 17085 13691 17088
rect 13633 17079 13691 17085
rect 13740 17084 13952 17088
rect 13998 17076 14004 17088
rect 14056 17076 14062 17128
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 14476 17125 14504 17212
rect 16040 17184 16068 17292
rect 18233 17289 18245 17292
rect 18279 17289 18291 17323
rect 18233 17283 18291 17289
rect 20257 17323 20315 17329
rect 20257 17289 20269 17323
rect 20303 17320 20315 17323
rect 21542 17320 21548 17332
rect 20303 17292 21548 17320
rect 20303 17289 20315 17292
rect 20257 17283 20315 17289
rect 21542 17280 21548 17292
rect 21600 17280 21606 17332
rect 22094 17280 22100 17332
rect 22152 17320 22158 17332
rect 22152 17292 26740 17320
rect 22152 17280 22158 17292
rect 23385 17255 23443 17261
rect 23385 17252 23397 17255
rect 22066 17224 23397 17252
rect 15028 17156 16068 17184
rect 16899 17187 16957 17193
rect 15028 17128 15056 17156
rect 16899 17153 16911 17187
rect 16945 17184 16957 17187
rect 18969 17187 19027 17193
rect 16945 17156 18920 17184
rect 16945 17153 16957 17156
rect 16899 17147 16957 17153
rect 14277 17119 14335 17125
rect 14277 17116 14289 17119
rect 14148 17088 14289 17116
rect 14148 17076 14154 17088
rect 14277 17085 14289 17088
rect 14323 17085 14335 17119
rect 14461 17119 14519 17125
rect 14461 17116 14473 17119
rect 14277 17079 14335 17085
rect 14384 17088 14473 17116
rect 10134 17008 10140 17060
rect 10192 17048 10198 17060
rect 10778 17048 10784 17060
rect 10192 17020 10784 17048
rect 10192 17008 10198 17020
rect 10778 17008 10784 17020
rect 10836 17048 10842 17060
rect 11149 17051 11207 17057
rect 11149 17048 11161 17051
rect 10836 17020 11161 17048
rect 10836 17008 10842 17020
rect 11149 17017 11161 17020
rect 11195 17017 11207 17051
rect 14384 17048 14412 17088
rect 14461 17085 14473 17088
rect 14507 17085 14519 17119
rect 14461 17079 14519 17085
rect 14737 17119 14795 17125
rect 14737 17085 14749 17119
rect 14783 17085 14795 17119
rect 14737 17079 14795 17085
rect 11149 17011 11207 17017
rect 12642 17020 14412 17048
rect 8435 16952 8800 16980
rect 8435 16949 8447 16952
rect 8389 16943 8447 16949
rect 9490 16940 9496 16992
rect 9548 16980 9554 16992
rect 11054 16980 11060 16992
rect 9548 16952 11060 16980
rect 9548 16940 9554 16952
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 11606 16940 11612 16992
rect 11664 16980 11670 16992
rect 11707 16983 11765 16989
rect 11707 16980 11719 16983
rect 11664 16952 11719 16980
rect 11664 16940 11670 16952
rect 11707 16949 11719 16952
rect 11753 16949 11765 16983
rect 11707 16943 11765 16949
rect 12066 16940 12072 16992
rect 12124 16980 12130 16992
rect 12642 16980 12670 17020
rect 14642 17008 14648 17060
rect 14700 17048 14706 17060
rect 14752 17048 14780 17079
rect 15010 17076 15016 17128
rect 15068 17076 15074 17128
rect 15841 17119 15899 17125
rect 15841 17116 15853 17119
rect 15120 17088 15853 17116
rect 14700 17020 14780 17048
rect 14700 17008 14706 17020
rect 14918 17008 14924 17060
rect 14976 17048 14982 17060
rect 15120 17048 15148 17088
rect 15841 17085 15853 17088
rect 15887 17116 15899 17119
rect 15930 17116 15936 17128
rect 15887 17088 15936 17116
rect 15887 17085 15899 17088
rect 15841 17079 15899 17085
rect 15930 17076 15936 17088
rect 15988 17076 15994 17128
rect 16117 17119 16175 17125
rect 16117 17085 16129 17119
rect 16163 17085 16175 17119
rect 16117 17079 16175 17085
rect 16393 17119 16451 17125
rect 16393 17085 16405 17119
rect 16439 17116 16451 17119
rect 17034 17116 17040 17128
rect 16439 17088 17040 17116
rect 16439 17085 16451 17088
rect 16393 17079 16451 17085
rect 14976 17020 15148 17048
rect 14976 17008 14982 17020
rect 15194 17008 15200 17060
rect 15252 17048 15258 17060
rect 16132 17048 16160 17079
rect 17034 17076 17040 17088
rect 17092 17076 17098 17128
rect 17126 17076 17132 17128
rect 17184 17076 17190 17128
rect 18693 17119 18751 17125
rect 18693 17085 18705 17119
rect 18739 17116 18751 17119
rect 18782 17116 18788 17128
rect 18739 17088 18788 17116
rect 18739 17085 18751 17088
rect 18693 17079 18751 17085
rect 18782 17076 18788 17088
rect 18840 17076 18846 17128
rect 18892 17116 18920 17156
rect 18969 17153 18981 17187
rect 19015 17184 19027 17187
rect 19150 17184 19156 17196
rect 19015 17156 19156 17184
rect 19015 17153 19027 17156
rect 18969 17147 19027 17153
rect 19150 17144 19156 17156
rect 19208 17144 19214 17196
rect 21131 17187 21189 17193
rect 20548 17156 21036 17184
rect 20548 17116 20576 17156
rect 18892 17088 20576 17116
rect 20625 17119 20683 17125
rect 20625 17085 20637 17119
rect 20671 17116 20683 17119
rect 20714 17116 20720 17128
rect 20671 17088 20720 17116
rect 20671 17085 20683 17088
rect 20625 17079 20683 17085
rect 16482 17048 16488 17060
rect 15252 17020 15700 17048
rect 16132 17020 16488 17048
rect 15252 17008 15258 17020
rect 12124 16952 12670 16980
rect 12124 16940 12130 16952
rect 12710 16940 12716 16992
rect 12768 16980 12774 16992
rect 13081 16983 13139 16989
rect 13081 16980 13093 16983
rect 12768 16952 13093 16980
rect 12768 16940 12774 16952
rect 13081 16949 13093 16952
rect 13127 16949 13139 16983
rect 13081 16943 13139 16949
rect 13262 16940 13268 16992
rect 13320 16980 13326 16992
rect 15381 16983 15439 16989
rect 15381 16980 15393 16983
rect 13320 16952 15393 16980
rect 13320 16940 13326 16952
rect 15381 16949 15393 16952
rect 15427 16980 15439 16983
rect 15562 16980 15568 16992
rect 15427 16952 15568 16980
rect 15427 16949 15439 16952
rect 15381 16943 15439 16949
rect 15562 16940 15568 16952
rect 15620 16940 15626 16992
rect 15672 16989 15700 17020
rect 16482 17008 16488 17020
rect 16540 17008 16546 17060
rect 20640 17048 20668 17079
rect 20714 17076 20720 17088
rect 20772 17076 20778 17128
rect 21008 17116 21036 17156
rect 21131 17153 21143 17187
rect 21177 17184 21189 17187
rect 21266 17184 21272 17196
rect 21177 17156 21272 17184
rect 21177 17153 21189 17156
rect 21131 17147 21189 17153
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 21361 17187 21419 17193
rect 21361 17153 21373 17187
rect 21407 17184 21419 17187
rect 22066 17184 22094 17224
rect 23385 17221 23397 17224
rect 23431 17221 23443 17255
rect 23385 17215 23443 17221
rect 23658 17212 23664 17264
rect 23716 17252 23722 17264
rect 24118 17252 24124 17264
rect 23716 17224 24124 17252
rect 23716 17212 23722 17224
rect 24118 17212 24124 17224
rect 24176 17212 24182 17264
rect 24210 17212 24216 17264
rect 24268 17252 24274 17264
rect 24670 17252 24676 17264
rect 24268 17224 24676 17252
rect 24268 17212 24274 17224
rect 21407 17156 22094 17184
rect 21407 17153 21419 17156
rect 21361 17147 21419 17153
rect 22278 17144 22284 17196
rect 22336 17144 22342 17196
rect 23014 17144 23020 17196
rect 23072 17184 23078 17196
rect 23750 17184 23756 17196
rect 23072 17156 23756 17184
rect 23072 17144 23078 17156
rect 23750 17144 23756 17156
rect 23808 17184 23814 17196
rect 23808 17156 24072 17184
rect 23808 17144 23814 17156
rect 21818 17116 21824 17128
rect 21008 17088 21824 17116
rect 21818 17076 21824 17088
rect 21876 17076 21882 17128
rect 22002 17076 22008 17128
rect 22060 17076 22066 17128
rect 22296 17116 22324 17144
rect 23569 17119 23627 17125
rect 23569 17116 23581 17119
rect 22296 17088 23581 17116
rect 23569 17085 23581 17088
rect 23615 17116 23627 17119
rect 23658 17116 23664 17128
rect 23615 17088 23664 17116
rect 23615 17085 23627 17088
rect 23569 17079 23627 17085
rect 23658 17076 23664 17088
rect 23716 17076 23722 17128
rect 24044 17125 24072 17156
rect 24320 17125 24348 17224
rect 24670 17212 24676 17224
rect 24728 17212 24734 17264
rect 26712 17261 26740 17292
rect 28966 17292 29960 17320
rect 26697 17255 26755 17261
rect 26697 17221 26709 17255
rect 26743 17221 26755 17255
rect 26697 17215 26755 17221
rect 28350 17212 28356 17264
rect 28408 17252 28414 17264
rect 28966 17252 28994 17292
rect 28408 17224 28994 17252
rect 28408 17212 28414 17224
rect 29546 17212 29552 17264
rect 29604 17212 29610 17264
rect 24486 17144 24492 17196
rect 24544 17184 24550 17196
rect 25222 17193 25228 17196
rect 24581 17187 24639 17193
rect 24581 17184 24593 17187
rect 24544 17156 24593 17184
rect 24544 17144 24550 17156
rect 24581 17153 24593 17156
rect 24627 17184 24639 17187
rect 25184 17187 25228 17193
rect 25184 17184 25196 17187
rect 24627 17156 25196 17184
rect 24627 17153 24639 17156
rect 24581 17147 24639 17153
rect 25184 17153 25196 17156
rect 25184 17147 25228 17153
rect 25222 17144 25228 17147
rect 25280 17144 25286 17196
rect 25314 17144 25320 17196
rect 25372 17184 25378 17196
rect 25372 17156 25417 17184
rect 25372 17144 25378 17156
rect 25498 17144 25504 17196
rect 25556 17184 25562 17196
rect 25593 17187 25651 17193
rect 25593 17184 25605 17187
rect 25556 17156 25605 17184
rect 25556 17144 25562 17156
rect 25593 17153 25605 17156
rect 25639 17153 25651 17187
rect 25593 17147 25651 17153
rect 27341 17187 27399 17193
rect 27341 17153 27353 17187
rect 27387 17184 27399 17187
rect 28442 17184 28448 17196
rect 27387 17156 28448 17184
rect 27387 17153 27399 17156
rect 27341 17147 27399 17153
rect 28442 17144 28448 17156
rect 28500 17144 28506 17196
rect 24029 17119 24087 17125
rect 24029 17085 24041 17119
rect 24075 17085 24087 17119
rect 24029 17079 24087 17085
rect 24305 17119 24363 17125
rect 24305 17085 24317 17119
rect 24351 17085 24363 17119
rect 24854 17116 24860 17128
rect 24305 17079 24363 17085
rect 24412 17088 24860 17116
rect 19904 17020 20668 17048
rect 22020 17048 22048 17076
rect 22925 17051 22983 17057
rect 22925 17048 22937 17051
rect 22020 17020 22937 17048
rect 19904 16992 19932 17020
rect 22925 17017 22937 17020
rect 22971 17017 22983 17051
rect 24412 17048 24440 17088
rect 24854 17076 24860 17088
rect 24912 17076 24918 17128
rect 26418 17076 26424 17128
rect 26476 17116 26482 17128
rect 29564 17125 29592 17212
rect 27065 17119 27123 17125
rect 27065 17116 27077 17119
rect 26476 17088 27077 17116
rect 26476 17076 26482 17088
rect 27065 17085 27077 17088
rect 27111 17116 27123 17119
rect 29549 17119 29607 17125
rect 27111 17088 28028 17116
rect 27111 17085 27123 17088
rect 27065 17079 27123 17085
rect 22925 17011 22983 17017
rect 23584 17020 24440 17048
rect 28000 17048 28028 17088
rect 29549 17085 29561 17119
rect 29595 17085 29607 17119
rect 29549 17079 29607 17085
rect 29825 17119 29883 17125
rect 29825 17085 29837 17119
rect 29871 17085 29883 17119
rect 29932 17116 29960 17292
rect 30101 17119 30159 17125
rect 30101 17116 30113 17119
rect 29932 17088 30113 17116
rect 29825 17079 29883 17085
rect 30101 17085 30113 17088
rect 30147 17085 30159 17119
rect 30101 17079 30159 17085
rect 28000 17020 28672 17048
rect 23584 16992 23612 17020
rect 28644 16992 28672 17020
rect 28718 17008 28724 17060
rect 28776 17008 28782 17060
rect 29089 17051 29147 17057
rect 29089 17017 29101 17051
rect 29135 17017 29147 17051
rect 29840 17048 29868 17079
rect 30006 17048 30012 17060
rect 29840 17020 30012 17048
rect 29089 17011 29147 17017
rect 15657 16983 15715 16989
rect 15657 16949 15669 16983
rect 15703 16949 15715 16983
rect 15657 16943 15715 16949
rect 16859 16983 16917 16989
rect 16859 16949 16871 16983
rect 16905 16980 16917 16983
rect 17494 16980 17500 16992
rect 16905 16952 17500 16980
rect 16905 16949 16917 16952
rect 16859 16943 16917 16949
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 19886 16940 19892 16992
rect 19944 16940 19950 16992
rect 21091 16983 21149 16989
rect 21091 16949 21103 16983
rect 21137 16980 21149 16983
rect 21450 16980 21456 16992
rect 21137 16952 21456 16980
rect 21137 16949 21149 16952
rect 21091 16943 21149 16949
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 21818 16940 21824 16992
rect 21876 16980 21882 16992
rect 22002 16980 22008 16992
rect 21876 16952 22008 16980
rect 21876 16940 21882 16952
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 22462 16940 22468 16992
rect 22520 16940 22526 16992
rect 23201 16983 23259 16989
rect 23201 16949 23213 16983
rect 23247 16980 23259 16983
rect 23566 16980 23572 16992
rect 23247 16952 23572 16980
rect 23247 16949 23259 16952
rect 23201 16943 23259 16949
rect 23566 16940 23572 16952
rect 23624 16940 23630 16992
rect 23842 16940 23848 16992
rect 23900 16940 23906 16992
rect 25590 16940 25596 16992
rect 25648 16980 25654 16992
rect 27982 16980 27988 16992
rect 25648 16952 27988 16980
rect 25648 16940 25654 16952
rect 27982 16940 27988 16952
rect 28040 16940 28046 16992
rect 28626 16940 28632 16992
rect 28684 16940 28690 16992
rect 29104 16980 29132 17011
rect 30006 17008 30012 17020
rect 30064 17008 30070 17060
rect 29270 16980 29276 16992
rect 29104 16952 29276 16980
rect 29270 16940 29276 16952
rect 29328 16940 29334 16992
rect 29546 16940 29552 16992
rect 29604 16980 29610 16992
rect 29917 16983 29975 16989
rect 29917 16980 29929 16983
rect 29604 16952 29929 16980
rect 29604 16940 29610 16952
rect 29917 16949 29929 16952
rect 29963 16949 29975 16983
rect 29917 16943 29975 16949
rect 30374 16940 30380 16992
rect 30432 16940 30438 16992
rect 552 16890 31072 16912
rect 552 16838 7988 16890
rect 8040 16838 8052 16890
rect 8104 16838 8116 16890
rect 8168 16838 8180 16890
rect 8232 16838 8244 16890
rect 8296 16838 15578 16890
rect 15630 16838 15642 16890
rect 15694 16838 15706 16890
rect 15758 16838 15770 16890
rect 15822 16838 15834 16890
rect 15886 16838 23168 16890
rect 23220 16838 23232 16890
rect 23284 16838 23296 16890
rect 23348 16838 23360 16890
rect 23412 16838 23424 16890
rect 23476 16838 30758 16890
rect 30810 16838 30822 16890
rect 30874 16838 30886 16890
rect 30938 16838 30950 16890
rect 31002 16838 31014 16890
rect 31066 16838 31072 16890
rect 552 16816 31072 16838
rect 937 16779 995 16785
rect 937 16745 949 16779
rect 983 16745 995 16779
rect 937 16739 995 16745
rect 952 16708 980 16739
rect 1026 16736 1032 16788
rect 1084 16776 1090 16788
rect 1854 16776 1860 16788
rect 1084 16748 1860 16776
rect 1084 16736 1090 16748
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 3050 16736 3056 16788
rect 3108 16736 3114 16788
rect 6546 16736 6552 16788
rect 6604 16776 6610 16788
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 6604 16748 7665 16776
rect 6604 16736 6610 16748
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 7653 16739 7711 16745
rect 8021 16779 8079 16785
rect 8021 16745 8033 16779
rect 8067 16776 8079 16779
rect 9950 16776 9956 16788
rect 8067 16748 9956 16776
rect 8067 16745 8079 16748
rect 8021 16739 8079 16745
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 10870 16736 10876 16788
rect 10928 16736 10934 16788
rect 11882 16776 11888 16788
rect 11164 16748 11888 16776
rect 1302 16708 1308 16720
rect 952 16680 1308 16708
rect 1302 16668 1308 16680
rect 1360 16668 1366 16720
rect 5626 16668 5632 16720
rect 5684 16668 5690 16720
rect 7374 16668 7380 16720
rect 7432 16708 7438 16720
rect 7834 16708 7840 16720
rect 7432 16680 7840 16708
rect 7432 16668 7438 16680
rect 7834 16668 7840 16680
rect 7892 16668 7898 16720
rect 8128 16680 8524 16708
rect 1118 16600 1124 16652
rect 1176 16600 1182 16652
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 4249 16643 4307 16649
rect 4120 16612 4200 16640
rect 4120 16600 4126 16612
rect 1709 16593 1767 16599
rect 1709 16590 1721 16593
rect 1210 16532 1216 16584
rect 1268 16532 1274 16584
rect 1578 16581 1584 16584
rect 1540 16575 1584 16581
rect 1540 16541 1552 16575
rect 1540 16535 1584 16541
rect 1578 16532 1584 16535
rect 1636 16532 1642 16584
rect 1688 16559 1721 16590
rect 1755 16584 1767 16593
rect 1755 16559 1768 16584
rect 1688 16544 1768 16559
rect 1762 16532 1768 16544
rect 1820 16532 1826 16584
rect 1854 16532 1860 16584
rect 1912 16572 1918 16584
rect 1949 16575 2007 16581
rect 1949 16572 1961 16575
rect 1912 16544 1961 16572
rect 1912 16532 1918 16544
rect 1949 16541 1961 16544
rect 1995 16541 2007 16575
rect 1949 16535 2007 16541
rect 3510 16532 3516 16584
rect 3568 16532 3574 16584
rect 3878 16581 3884 16584
rect 3840 16575 3884 16581
rect 3840 16541 3852 16575
rect 3840 16535 3884 16541
rect 3878 16532 3884 16535
rect 3936 16532 3942 16584
rect 3970 16532 3976 16584
rect 4028 16572 4034 16584
rect 4172 16572 4200 16612
rect 4249 16609 4261 16643
rect 4295 16640 4307 16643
rect 4706 16640 4712 16652
rect 4295 16612 4712 16640
rect 4295 16609 4307 16612
rect 4249 16603 4307 16609
rect 4706 16600 4712 16612
rect 4764 16600 4770 16652
rect 4982 16600 4988 16652
rect 5040 16640 5046 16652
rect 6140 16643 6198 16649
rect 6140 16640 6152 16643
rect 5040 16612 6152 16640
rect 5040 16600 5046 16612
rect 6140 16609 6152 16612
rect 6186 16609 6198 16643
rect 6140 16603 6198 16609
rect 6546 16600 6552 16652
rect 6604 16600 6610 16652
rect 7466 16600 7472 16652
rect 7524 16640 7530 16652
rect 8128 16640 8156 16680
rect 8496 16649 8524 16680
rect 7524 16612 8156 16640
rect 8205 16643 8263 16649
rect 7524 16600 7530 16612
rect 8205 16609 8217 16643
rect 8251 16609 8263 16643
rect 8205 16603 8263 16609
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16609 8539 16643
rect 8481 16603 8539 16609
rect 8573 16643 8631 16649
rect 8573 16609 8585 16643
rect 8619 16640 8631 16643
rect 8662 16640 8668 16652
rect 8619 16612 8668 16640
rect 8619 16609 8631 16612
rect 8573 16603 8631 16609
rect 6362 16583 6368 16584
rect 5813 16575 5871 16581
rect 5813 16572 5825 16575
rect 4028 16544 4073 16572
rect 4172 16544 5825 16572
rect 4028 16532 4034 16544
rect 5813 16541 5825 16544
rect 5859 16541 5871 16575
rect 5813 16535 5871 16541
rect 6319 16577 6368 16583
rect 6319 16543 6331 16577
rect 6365 16543 6368 16577
rect 6319 16537 6368 16543
rect 6362 16532 6368 16537
rect 6420 16532 6426 16584
rect 7006 16532 7012 16584
rect 7064 16572 7070 16584
rect 8110 16572 8116 16584
rect 7064 16544 8116 16572
rect 7064 16532 7070 16544
rect 8110 16532 8116 16544
rect 8168 16532 8174 16584
rect 8220 16504 8248 16603
rect 8496 16572 8524 16603
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 9214 16640 9220 16652
rect 8772 16612 9220 16640
rect 8772 16572 8800 16612
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 9309 16643 9367 16649
rect 9309 16609 9321 16643
rect 9355 16640 9367 16643
rect 9950 16640 9956 16652
rect 9355 16612 9956 16640
rect 9355 16609 9367 16612
rect 9309 16603 9367 16609
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 10888 16640 10916 16736
rect 11164 16717 11192 16748
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12894 16736 12900 16788
rect 12952 16776 12958 16788
rect 13449 16779 13507 16785
rect 13449 16776 13461 16779
rect 12952 16748 13461 16776
rect 12952 16736 12958 16748
rect 13449 16745 13461 16748
rect 13495 16745 13507 16779
rect 13449 16739 13507 16745
rect 15194 16736 15200 16788
rect 15252 16736 15258 16788
rect 15470 16736 15476 16788
rect 15528 16776 15534 16788
rect 15657 16779 15715 16785
rect 15657 16776 15669 16779
rect 15528 16748 15669 16776
rect 15528 16736 15534 16748
rect 15657 16745 15669 16748
rect 15703 16745 15715 16779
rect 15657 16739 15715 16745
rect 15930 16736 15936 16788
rect 15988 16776 15994 16788
rect 16301 16779 16359 16785
rect 16301 16776 16313 16779
rect 15988 16748 16313 16776
rect 15988 16736 15994 16748
rect 16301 16745 16313 16748
rect 16347 16745 16359 16779
rect 16301 16739 16359 16745
rect 16666 16736 16672 16788
rect 16724 16736 16730 16788
rect 18969 16779 19027 16785
rect 18969 16776 18981 16779
rect 16776 16748 18981 16776
rect 11149 16711 11207 16717
rect 11149 16677 11161 16711
rect 11195 16677 11207 16711
rect 11149 16671 11207 16677
rect 11330 16668 11336 16720
rect 11388 16708 11394 16720
rect 12434 16708 12440 16720
rect 11388 16680 12440 16708
rect 11388 16668 11394 16680
rect 12434 16668 12440 16680
rect 12492 16708 12498 16720
rect 12492 16680 13676 16708
rect 12492 16668 12498 16680
rect 11974 16640 11980 16652
rect 10888 16612 11980 16640
rect 11974 16600 11980 16612
rect 12032 16600 12038 16652
rect 12066 16600 12072 16652
rect 12124 16600 12130 16652
rect 12342 16600 12348 16652
rect 12400 16640 12406 16652
rect 12986 16640 12992 16652
rect 12400 16612 12992 16640
rect 12400 16600 12406 16612
rect 12986 16600 12992 16612
rect 13044 16600 13050 16652
rect 13173 16643 13231 16649
rect 13173 16609 13185 16643
rect 13219 16640 13231 16643
rect 13262 16640 13268 16652
rect 13219 16612 13268 16640
rect 13219 16609 13231 16612
rect 13173 16603 13231 16609
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 13648 16649 13676 16680
rect 13633 16643 13691 16649
rect 13633 16609 13645 16643
rect 13679 16609 13691 16643
rect 13633 16603 13691 16609
rect 14553 16643 14611 16649
rect 14553 16609 14565 16643
rect 14599 16640 14611 16643
rect 15212 16640 15240 16736
rect 16114 16668 16120 16720
rect 16172 16708 16178 16720
rect 16776 16708 16804 16748
rect 18969 16745 18981 16748
rect 19015 16745 19027 16779
rect 22462 16776 22468 16788
rect 18969 16739 19027 16745
rect 19536 16748 22468 16776
rect 16172 16680 16804 16708
rect 16172 16668 16178 16680
rect 14599 16612 15240 16640
rect 14599 16609 14611 16612
rect 14553 16603 14611 16609
rect 15562 16600 15568 16652
rect 15620 16640 15626 16652
rect 16209 16643 16267 16649
rect 16209 16640 16221 16643
rect 15620 16612 16221 16640
rect 15620 16600 15626 16612
rect 16209 16609 16221 16612
rect 16255 16640 16267 16643
rect 16298 16640 16304 16652
rect 16255 16612 16304 16640
rect 16255 16609 16267 16612
rect 16209 16603 16267 16609
rect 16298 16600 16304 16612
rect 16356 16600 16362 16652
rect 16850 16640 16856 16652
rect 16684 16612 16856 16640
rect 8938 16581 8944 16584
rect 8496 16544 8800 16572
rect 8900 16575 8944 16581
rect 8900 16541 8912 16575
rect 8900 16535 8944 16541
rect 8938 16532 8944 16535
rect 8996 16532 9002 16584
rect 9079 16577 9137 16583
rect 9079 16543 9091 16577
rect 9125 16572 9137 16577
rect 9490 16572 9496 16584
rect 9125 16544 9496 16572
rect 9125 16543 9137 16544
rect 9079 16537 9137 16543
rect 9490 16532 9496 16544
rect 9548 16532 9554 16584
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 10042 16572 10048 16584
rect 9732 16544 10048 16572
rect 9732 16532 9738 16544
rect 10042 16532 10048 16544
rect 10100 16572 10106 16584
rect 11425 16575 11483 16581
rect 11425 16572 11437 16575
rect 10100 16544 11437 16572
rect 10100 16532 10106 16544
rect 11425 16541 11437 16544
rect 11471 16572 11483 16575
rect 11698 16572 11704 16584
rect 11471 16544 11704 16572
rect 11471 16541 11483 16544
rect 11425 16535 11483 16541
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 13814 16532 13820 16584
rect 13872 16581 13878 16584
rect 14182 16581 14188 16584
rect 13872 16572 13883 16581
rect 14144 16575 14188 16581
rect 13872 16544 13917 16572
rect 13872 16535 13883 16544
rect 14144 16541 14156 16575
rect 14144 16535 14188 16541
rect 13872 16532 13878 16535
rect 14182 16532 14188 16535
rect 14240 16532 14246 16584
rect 14323 16575 14381 16581
rect 14323 16541 14335 16575
rect 14369 16572 14381 16575
rect 15010 16572 15016 16584
rect 14369 16544 15016 16572
rect 14369 16541 14381 16544
rect 14323 16535 14381 16541
rect 15010 16532 15016 16544
rect 15068 16532 15074 16584
rect 16684 16516 16712 16612
rect 16850 16600 16856 16612
rect 16908 16600 16914 16652
rect 17034 16600 17040 16652
rect 17092 16640 17098 16652
rect 17129 16643 17187 16649
rect 17129 16640 17141 16643
rect 17092 16612 17141 16640
rect 17092 16600 17098 16612
rect 17129 16609 17141 16612
rect 17175 16640 17187 16643
rect 17218 16640 17224 16652
rect 17175 16612 17224 16640
rect 17175 16609 17187 16612
rect 17129 16603 17187 16609
rect 17218 16600 17224 16612
rect 17276 16600 17282 16652
rect 19536 16640 19564 16748
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 22646 16736 22652 16788
rect 22704 16776 22710 16788
rect 23109 16779 23167 16785
rect 23109 16776 23121 16779
rect 22704 16748 23121 16776
rect 22704 16736 22710 16748
rect 23109 16745 23121 16748
rect 23155 16745 23167 16779
rect 23842 16776 23848 16788
rect 23109 16739 23167 16745
rect 23216 16748 23848 16776
rect 21082 16668 21088 16720
rect 21140 16668 21146 16720
rect 17788 16612 19564 16640
rect 19705 16643 19763 16649
rect 17625 16593 17683 16599
rect 17494 16581 17500 16584
rect 17456 16575 17500 16581
rect 17456 16541 17468 16575
rect 17456 16535 17500 16541
rect 17494 16532 17500 16535
rect 17552 16532 17558 16584
rect 17625 16559 17637 16593
rect 17671 16572 17683 16593
rect 17788 16572 17816 16612
rect 19705 16609 19717 16643
rect 19751 16640 19763 16643
rect 20622 16640 20628 16652
rect 19751 16612 20628 16640
rect 19751 16609 19763 16612
rect 19705 16603 19763 16609
rect 20622 16600 20628 16612
rect 20680 16600 20686 16652
rect 20898 16640 20904 16652
rect 20732 16612 20904 16640
rect 17671 16559 17816 16572
rect 17625 16553 17816 16559
rect 17640 16544 17816 16553
rect 17865 16575 17923 16581
rect 17865 16541 17877 16575
rect 17911 16572 17923 16575
rect 18046 16572 18052 16584
rect 17911 16544 18052 16572
rect 17911 16541 17923 16544
rect 17865 16535 17923 16541
rect 18046 16532 18052 16544
rect 18104 16532 18110 16584
rect 19429 16575 19487 16581
rect 19429 16541 19441 16575
rect 19475 16572 19487 16575
rect 20732 16572 20760 16612
rect 20898 16600 20904 16612
rect 20956 16600 20962 16652
rect 22005 16643 22063 16649
rect 22005 16609 22017 16643
rect 22051 16640 22063 16643
rect 23216 16640 23244 16748
rect 23842 16736 23848 16748
rect 23900 16736 23906 16788
rect 23943 16779 24001 16785
rect 23943 16745 23955 16779
rect 23989 16776 24001 16779
rect 24210 16776 24216 16788
rect 23989 16748 24216 16776
rect 23989 16745 24001 16748
rect 23943 16739 24001 16745
rect 24210 16736 24216 16748
rect 24268 16776 24274 16788
rect 24486 16776 24492 16788
rect 24268 16748 24492 16776
rect 24268 16736 24274 16748
rect 24486 16736 24492 16748
rect 24544 16736 24550 16788
rect 24872 16748 27844 16776
rect 24213 16643 24271 16649
rect 24213 16640 24225 16643
rect 22051 16612 23244 16640
rect 23676 16612 24225 16640
rect 22051 16609 22063 16612
rect 22005 16603 22063 16609
rect 21765 16593 21823 16599
rect 19475 16544 20760 16572
rect 19475 16541 19487 16544
rect 19429 16535 19487 16541
rect 21266 16532 21272 16584
rect 21324 16532 21330 16584
rect 21450 16532 21456 16584
rect 21508 16572 21514 16584
rect 21596 16575 21654 16581
rect 21596 16572 21608 16575
rect 21508 16544 21608 16572
rect 21508 16532 21514 16544
rect 21596 16541 21608 16544
rect 21642 16541 21654 16575
rect 21765 16559 21777 16593
rect 21811 16584 21823 16593
rect 23676 16584 23704 16612
rect 24213 16609 24225 16612
rect 24259 16609 24271 16643
rect 24872 16640 24900 16748
rect 24946 16668 24952 16720
rect 25004 16668 25010 16720
rect 25222 16668 25228 16720
rect 25280 16708 25286 16720
rect 25280 16680 25912 16708
rect 25280 16668 25286 16680
rect 24213 16603 24271 16609
rect 24320 16612 24900 16640
rect 24964 16640 24992 16668
rect 25777 16643 25835 16649
rect 25777 16640 25789 16643
rect 24964 16612 25789 16640
rect 21811 16559 21824 16584
rect 21765 16553 21824 16559
rect 21790 16544 21824 16553
rect 21596 16535 21654 16541
rect 21818 16532 21824 16544
rect 21876 16532 21882 16584
rect 21910 16532 21916 16584
rect 21968 16572 21974 16584
rect 22370 16572 22376 16584
rect 21968 16544 22376 16572
rect 21968 16532 21974 16544
rect 22370 16532 22376 16544
rect 22428 16572 22434 16584
rect 23014 16572 23020 16584
rect 22428 16544 23020 16572
rect 22428 16532 22434 16544
rect 23014 16532 23020 16544
rect 23072 16532 23078 16584
rect 23474 16532 23480 16584
rect 23532 16532 23538 16584
rect 23658 16532 23664 16584
rect 23716 16532 23722 16584
rect 23956 16577 24014 16583
rect 23956 16543 23968 16577
rect 24002 16572 24014 16577
rect 24320 16572 24348 16612
rect 25777 16609 25789 16612
rect 25823 16609 25835 16643
rect 25884 16640 25912 16680
rect 27816 16652 27844 16748
rect 27982 16736 27988 16788
rect 28040 16776 28046 16788
rect 28261 16779 28319 16785
rect 28261 16776 28273 16779
rect 28040 16748 28273 16776
rect 28040 16736 28046 16748
rect 28261 16745 28273 16748
rect 28307 16745 28319 16779
rect 28261 16739 28319 16745
rect 29362 16736 29368 16788
rect 29420 16776 29426 16788
rect 30377 16779 30435 16785
rect 30377 16776 30389 16779
rect 29420 16748 30389 16776
rect 29420 16736 29426 16748
rect 30377 16745 30389 16748
rect 30423 16745 30435 16779
rect 30377 16739 30435 16745
rect 30282 16668 30288 16720
rect 30340 16668 30346 16720
rect 26748 16643 26806 16649
rect 26748 16640 26760 16643
rect 25884 16612 26760 16640
rect 25777 16603 25835 16609
rect 26748 16609 26760 16612
rect 26794 16609 26806 16643
rect 27522 16640 27528 16652
rect 26748 16603 26806 16609
rect 26899 16612 27528 16640
rect 24002 16544 24348 16572
rect 24002 16543 24014 16544
rect 23956 16537 24014 16543
rect 25682 16532 25688 16584
rect 25740 16532 25746 16584
rect 25792 16572 25820 16603
rect 26899 16583 26927 16612
rect 27522 16600 27528 16612
rect 27580 16600 27586 16652
rect 27798 16600 27804 16652
rect 27856 16600 27862 16652
rect 28258 16600 28264 16652
rect 28316 16640 28322 16652
rect 28905 16643 28963 16649
rect 28905 16640 28917 16643
rect 28316 16612 28917 16640
rect 28316 16600 28322 16612
rect 28905 16609 28917 16612
rect 28951 16609 28963 16643
rect 28905 16603 28963 16609
rect 30098 16600 30104 16652
rect 30156 16640 30162 16652
rect 30466 16640 30472 16652
rect 30156 16612 30472 16640
rect 30156 16600 30162 16612
rect 30466 16600 30472 16612
rect 30524 16640 30530 16652
rect 30561 16643 30619 16649
rect 30561 16640 30573 16643
rect 30524 16612 30573 16640
rect 30524 16600 30530 16612
rect 30561 16609 30573 16612
rect 30607 16609 30619 16643
rect 30561 16603 30619 16609
rect 26421 16575 26479 16581
rect 26421 16572 26433 16575
rect 25792 16544 26433 16572
rect 26421 16541 26433 16544
rect 26467 16541 26479 16575
rect 26421 16535 26479 16541
rect 26884 16577 26942 16583
rect 26884 16543 26896 16577
rect 26930 16543 26942 16577
rect 26884 16537 26942 16543
rect 26970 16532 26976 16584
rect 27028 16572 27034 16584
rect 27157 16575 27215 16581
rect 27157 16572 27169 16575
rect 27028 16544 27169 16572
rect 27028 16532 27034 16544
rect 27157 16541 27169 16544
rect 27203 16541 27215 16575
rect 27157 16535 27215 16541
rect 28626 16532 28632 16584
rect 28684 16532 28690 16584
rect 8478 16504 8484 16516
rect 8220 16476 8484 16504
rect 8478 16464 8484 16476
rect 8536 16464 8542 16516
rect 16022 16464 16028 16516
rect 16080 16504 16086 16516
rect 16390 16504 16396 16516
rect 16080 16476 16396 16504
rect 16080 16464 16086 16476
rect 16390 16464 16396 16476
rect 16448 16464 16454 16516
rect 16666 16464 16672 16516
rect 16724 16464 16730 16516
rect 25700 16504 25728 16532
rect 25958 16504 25964 16516
rect 18892 16476 19472 16504
rect 2038 16396 2044 16448
rect 2096 16436 2102 16448
rect 3786 16436 3792 16448
rect 2096 16408 3792 16436
rect 2096 16396 2102 16408
rect 3786 16396 3792 16408
rect 3844 16396 3850 16448
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 7190 16436 7196 16448
rect 4120 16408 7196 16436
rect 4120 16396 4126 16408
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 8297 16439 8355 16445
rect 8297 16405 8309 16439
rect 8343 16436 8355 16439
rect 9214 16436 9220 16448
rect 8343 16408 9220 16436
rect 8343 16405 8355 16408
rect 8297 16399 8355 16405
rect 9214 16396 9220 16408
rect 9272 16396 9278 16448
rect 10410 16396 10416 16448
rect 10468 16396 10474 16448
rect 10962 16396 10968 16448
rect 11020 16436 11026 16448
rect 12434 16436 12440 16448
rect 11020 16408 12440 16436
rect 11020 16396 11026 16408
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 13354 16396 13360 16448
rect 13412 16396 13418 16448
rect 14458 16396 14464 16448
rect 14516 16436 14522 16448
rect 17586 16436 17592 16448
rect 14516 16408 17592 16436
rect 14516 16396 14522 16408
rect 17586 16396 17592 16408
rect 17644 16396 17650 16448
rect 17678 16396 17684 16448
rect 17736 16436 17742 16448
rect 18892 16436 18920 16476
rect 17736 16408 18920 16436
rect 19444 16436 19472 16476
rect 20732 16476 20944 16504
rect 25700 16476 25964 16504
rect 20732 16436 20760 16476
rect 19444 16408 20760 16436
rect 20916 16436 20944 16476
rect 25958 16464 25964 16476
rect 26016 16464 26022 16516
rect 22922 16436 22928 16448
rect 20916 16408 22928 16436
rect 17736 16396 17742 16408
rect 22922 16396 22928 16408
rect 22980 16396 22986 16448
rect 23014 16396 23020 16448
rect 23072 16436 23078 16448
rect 25317 16439 25375 16445
rect 25317 16436 25329 16439
rect 23072 16408 25329 16436
rect 23072 16396 23078 16408
rect 25317 16405 25329 16408
rect 25363 16405 25375 16439
rect 25317 16399 25375 16405
rect 26694 16396 26700 16448
rect 26752 16436 26758 16448
rect 28074 16436 28080 16448
rect 26752 16408 28080 16436
rect 26752 16396 26758 16408
rect 28074 16396 28080 16408
rect 28132 16436 28138 16448
rect 30098 16436 30104 16448
rect 28132 16408 30104 16436
rect 28132 16396 28138 16408
rect 30098 16396 30104 16408
rect 30156 16396 30162 16448
rect 552 16346 30912 16368
rect 552 16294 4193 16346
rect 4245 16294 4257 16346
rect 4309 16294 4321 16346
rect 4373 16294 4385 16346
rect 4437 16294 4449 16346
rect 4501 16294 11783 16346
rect 11835 16294 11847 16346
rect 11899 16294 11911 16346
rect 11963 16294 11975 16346
rect 12027 16294 12039 16346
rect 12091 16294 19373 16346
rect 19425 16294 19437 16346
rect 19489 16294 19501 16346
rect 19553 16294 19565 16346
rect 19617 16294 19629 16346
rect 19681 16294 26963 16346
rect 27015 16294 27027 16346
rect 27079 16294 27091 16346
rect 27143 16294 27155 16346
rect 27207 16294 27219 16346
rect 27271 16294 30912 16346
rect 552 16272 30912 16294
rect 2314 16192 2320 16244
rect 2372 16232 2378 16244
rect 2777 16235 2835 16241
rect 2777 16232 2789 16235
rect 2372 16204 2789 16232
rect 2372 16192 2378 16204
rect 2777 16201 2789 16204
rect 2823 16201 2835 16235
rect 5626 16232 5632 16244
rect 2777 16195 2835 16201
rect 3252 16204 5632 16232
rect 842 16056 848 16108
rect 900 16096 906 16108
rect 1443 16099 1501 16105
rect 900 16068 1348 16096
rect 900 16056 906 16068
rect 937 16031 995 16037
rect 937 15997 949 16031
rect 983 15997 995 16031
rect 1320 16028 1348 16068
rect 1443 16065 1455 16099
rect 1489 16096 1501 16099
rect 3252 16096 3280 16204
rect 5626 16192 5632 16204
rect 5684 16192 5690 16244
rect 7929 16235 7987 16241
rect 7929 16232 7941 16235
rect 6104 16204 7941 16232
rect 3694 16164 3700 16176
rect 1489 16068 3280 16096
rect 3344 16136 3700 16164
rect 1489 16065 1501 16068
rect 1443 16059 1501 16065
rect 3344 16037 3372 16136
rect 3694 16124 3700 16136
rect 3752 16124 3758 16176
rect 3786 16124 3792 16176
rect 3844 16124 3850 16176
rect 5810 16124 5816 16176
rect 5868 16124 5874 16176
rect 3804 16096 3832 16124
rect 4295 16099 4353 16105
rect 3804 16068 4200 16096
rect 1673 16031 1731 16037
rect 1673 16028 1685 16031
rect 1320 16000 1685 16028
rect 937 15991 995 15997
rect 1673 15997 1685 16000
rect 1719 15997 1731 16031
rect 1673 15991 1731 15997
rect 3329 16031 3387 16037
rect 3329 15997 3341 16031
rect 3375 15997 3387 16031
rect 3789 16031 3847 16037
rect 3789 16028 3801 16031
rect 3329 15991 3387 15997
rect 3620 16000 3801 16028
rect 952 15892 980 15991
rect 1302 15892 1308 15904
rect 952 15864 1308 15892
rect 1302 15852 1308 15864
rect 1360 15852 1366 15904
rect 1403 15895 1461 15901
rect 1403 15861 1415 15895
rect 1449 15892 1461 15895
rect 1578 15892 1584 15904
rect 1449 15864 1584 15892
rect 1449 15861 1461 15864
rect 1403 15855 1461 15861
rect 1578 15852 1584 15864
rect 1636 15852 1642 15904
rect 3510 15852 3516 15904
rect 3568 15892 3574 15904
rect 3620 15901 3648 16000
rect 3789 15997 3801 16000
rect 3835 15997 3847 16031
rect 4172 16028 4200 16068
rect 4295 16065 4307 16099
rect 4341 16096 4353 16099
rect 6104 16096 6132 16204
rect 7929 16201 7941 16204
rect 7975 16201 7987 16235
rect 7929 16195 7987 16201
rect 8110 16192 8116 16244
rect 8168 16232 8174 16244
rect 10502 16232 10508 16244
rect 8168 16204 10508 16232
rect 8168 16192 8174 16204
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 13081 16235 13139 16241
rect 13081 16232 13093 16235
rect 10980 16204 13093 16232
rect 6454 16105 6460 16108
rect 4341 16068 6132 16096
rect 6416 16099 6460 16105
rect 4341 16065 4353 16068
rect 4295 16059 4353 16065
rect 6416 16065 6428 16099
rect 6416 16059 6460 16065
rect 6454 16056 6460 16059
rect 6512 16056 6518 16108
rect 6595 16097 6653 16103
rect 6595 16063 6607 16097
rect 6641 16096 6653 16097
rect 8478 16096 8484 16108
rect 6641 16068 8484 16096
rect 6641 16063 6653 16068
rect 6595 16057 6653 16063
rect 8478 16056 8484 16068
rect 8536 16056 8542 16108
rect 9069 16081 9127 16087
rect 9069 16047 9081 16081
rect 9115 16047 9127 16081
rect 9214 16056 9220 16108
rect 9272 16096 9278 16108
rect 9309 16099 9367 16105
rect 9309 16096 9321 16099
rect 9272 16068 9321 16096
rect 9272 16056 9278 16068
rect 9309 16065 9321 16068
rect 9355 16065 9367 16099
rect 9309 16059 9367 16065
rect 9069 16044 9127 16047
rect 9069 16041 9168 16044
rect 4430 16028 4436 16040
rect 4172 16000 4436 16028
rect 3789 15991 3847 15997
rect 4430 15988 4436 16000
rect 4488 15988 4494 16040
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 16028 4583 16031
rect 4982 16028 4988 16040
rect 4571 16000 4988 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 4982 15988 4988 16000
rect 5040 15988 5046 16040
rect 6086 15988 6092 16040
rect 6144 15988 6150 16040
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6196 16000 6837 16028
rect 5442 15920 5448 15972
rect 5500 15960 5506 15972
rect 6196 15960 6224 16000
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 6825 15991 6883 15997
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 16028 8631 16031
rect 8662 16028 8668 16040
rect 8619 16000 8668 16028
rect 8619 15997 8631 16000
rect 8573 15991 8631 15997
rect 8662 15988 8668 16000
rect 8720 15988 8726 16040
rect 8938 16037 8944 16040
rect 8900 16031 8944 16037
rect 8900 15997 8912 16031
rect 8900 15991 8944 15997
rect 8938 15988 8944 15991
rect 8996 15988 9002 16040
rect 9084 16028 9168 16041
rect 10980 16028 11008 16204
rect 13081 16201 13093 16204
rect 13127 16201 13139 16235
rect 13081 16195 13139 16201
rect 13446 16192 13452 16244
rect 13504 16232 13510 16244
rect 14093 16235 14151 16241
rect 14093 16232 14105 16235
rect 13504 16204 14105 16232
rect 13504 16192 13510 16204
rect 14093 16201 14105 16204
rect 14139 16201 14151 16235
rect 14093 16195 14151 16201
rect 14461 16235 14519 16241
rect 14461 16201 14473 16235
rect 14507 16232 14519 16235
rect 15286 16232 15292 16244
rect 14507 16204 15292 16232
rect 14507 16201 14519 16204
rect 14461 16195 14519 16201
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 16666 16232 16672 16244
rect 15528 16204 16672 16232
rect 15528 16192 15534 16204
rect 16666 16192 16672 16204
rect 16724 16192 16730 16244
rect 17126 16192 17132 16244
rect 17184 16232 17190 16244
rect 17497 16235 17555 16241
rect 17497 16232 17509 16235
rect 17184 16204 17509 16232
rect 17184 16192 17190 16204
rect 17497 16201 17509 16204
rect 17543 16201 17555 16235
rect 17497 16195 17555 16201
rect 17773 16235 17831 16241
rect 17773 16201 17785 16235
rect 17819 16232 17831 16235
rect 17862 16232 17868 16244
rect 17819 16204 17868 16232
rect 17819 16201 17831 16204
rect 17773 16195 17831 16201
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 18417 16235 18475 16241
rect 18417 16201 18429 16235
rect 18463 16232 18475 16235
rect 19886 16232 19892 16244
rect 18463 16204 19892 16232
rect 18463 16201 18475 16204
rect 18417 16195 18475 16201
rect 19886 16192 19892 16204
rect 19944 16192 19950 16244
rect 22738 16232 22744 16244
rect 20640 16204 22744 16232
rect 16298 16124 16304 16176
rect 16356 16164 16362 16176
rect 17221 16167 17279 16173
rect 16356 16136 16988 16164
rect 16356 16124 16362 16136
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11606 16105 11612 16108
rect 11568 16099 11612 16105
rect 11112 16068 11192 16096
rect 11112 16056 11118 16068
rect 11164 16037 11192 16068
rect 11568 16065 11580 16099
rect 11568 16059 11612 16065
rect 11606 16056 11612 16059
rect 11664 16056 11670 16108
rect 11747 16099 11805 16105
rect 11747 16065 11759 16099
rect 11793 16096 11805 16099
rect 13538 16096 13544 16108
rect 11793 16068 13544 16096
rect 11793 16065 11805 16068
rect 11747 16059 11805 16065
rect 13538 16056 13544 16068
rect 13596 16056 13602 16108
rect 14737 16099 14795 16105
rect 14737 16096 14749 16099
rect 13832 16068 14749 16096
rect 13832 16040 13860 16068
rect 14737 16065 14749 16068
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 15243 16099 15301 16105
rect 15243 16065 15255 16099
rect 15289 16096 15301 16099
rect 15289 16068 16528 16096
rect 15289 16065 15301 16068
rect 15243 16059 15301 16065
rect 9084 16016 11008 16028
rect 9140 16000 11008 16016
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 15997 11207 16031
rect 11149 15991 11207 15997
rect 11238 15988 11244 16040
rect 11296 15988 11302 16040
rect 11977 16031 12035 16037
rect 11977 16028 11989 16031
rect 11348 16000 11989 16028
rect 10686 15960 10692 15972
rect 5500 15932 6224 15960
rect 10336 15932 10692 15960
rect 5500 15920 5506 15932
rect 3605 15895 3663 15901
rect 3605 15892 3617 15895
rect 3568 15864 3617 15892
rect 3568 15852 3574 15864
rect 3605 15861 3617 15864
rect 3651 15861 3663 15895
rect 3605 15855 3663 15861
rect 3878 15852 3884 15904
rect 3936 15892 3942 15904
rect 4255 15895 4313 15901
rect 4255 15892 4267 15895
rect 3936 15864 4267 15892
rect 3936 15852 3942 15864
rect 4255 15861 4267 15864
rect 4301 15861 4313 15895
rect 4255 15855 4313 15861
rect 4430 15852 4436 15904
rect 4488 15892 4494 15904
rect 10336 15892 10364 15932
rect 10686 15920 10692 15932
rect 10744 15920 10750 15972
rect 4488 15864 10364 15892
rect 4488 15852 4494 15864
rect 10410 15852 10416 15904
rect 10468 15852 10474 15904
rect 10965 15895 11023 15901
rect 10965 15861 10977 15895
rect 11011 15892 11023 15895
rect 11348 15892 11376 16000
rect 11977 15997 11989 16000
rect 12023 15997 12035 16031
rect 11977 15991 12035 15997
rect 13814 15988 13820 16040
rect 13872 15988 13878 16040
rect 13906 15988 13912 16040
rect 13964 16028 13970 16040
rect 14277 16031 14335 16037
rect 14277 16028 14289 16031
rect 13964 16000 14289 16028
rect 13964 15988 13970 16000
rect 14277 15997 14289 16000
rect 14323 15997 14335 16031
rect 14277 15991 14335 15997
rect 14645 16031 14703 16037
rect 14645 15997 14657 16031
rect 14691 16028 14703 16031
rect 15473 16031 15531 16037
rect 14691 16000 14780 16028
rect 14691 15997 14703 16000
rect 14645 15991 14703 15997
rect 13538 15920 13544 15972
rect 13596 15960 13602 15972
rect 13633 15963 13691 15969
rect 13633 15960 13645 15963
rect 13596 15932 13645 15960
rect 13596 15920 13602 15932
rect 13633 15929 13645 15932
rect 13679 15929 13691 15963
rect 13633 15923 13691 15929
rect 13998 15920 14004 15972
rect 14056 15960 14062 15972
rect 14752 15960 14780 16000
rect 15473 15997 15485 16031
rect 15519 16028 15531 16031
rect 16114 16028 16120 16040
rect 15519 16000 16120 16028
rect 15519 15997 15531 16000
rect 15473 15991 15531 15997
rect 16114 15988 16120 16000
rect 16172 15988 16178 16040
rect 14056 15932 14780 15960
rect 16500 15960 16528 16068
rect 16960 16040 16988 16136
rect 17221 16133 17233 16167
rect 17267 16133 17279 16167
rect 17221 16127 17279 16133
rect 17236 16096 17264 16127
rect 19199 16099 19257 16105
rect 17236 16068 18828 16096
rect 16942 15988 16948 16040
rect 17000 15988 17006 16040
rect 17405 16031 17463 16037
rect 17405 15997 17417 16031
rect 17451 16028 17463 16031
rect 17586 16028 17592 16040
rect 17451 16000 17592 16028
rect 17451 15997 17463 16000
rect 17405 15991 17463 15997
rect 17586 15988 17592 16000
rect 17644 15988 17650 16040
rect 17678 15988 17684 16040
rect 17736 15988 17742 16040
rect 17957 16031 18015 16037
rect 17957 15997 17969 16031
rect 18003 16028 18015 16031
rect 18598 16028 18604 16040
rect 18003 16000 18604 16028
rect 18003 15997 18015 16000
rect 17957 15991 18015 15997
rect 18598 15988 18604 16000
rect 18656 15988 18662 16040
rect 18693 16031 18751 16037
rect 18693 15997 18705 16031
rect 18739 15997 18751 16031
rect 18800 16028 18828 16068
rect 19199 16065 19211 16099
rect 19245 16096 19257 16099
rect 20640 16096 20668 16204
rect 22738 16192 22744 16204
rect 22796 16192 22802 16244
rect 22922 16192 22928 16244
rect 22980 16232 22986 16244
rect 22980 16204 25728 16232
rect 22980 16192 22986 16204
rect 25700 16173 25728 16204
rect 25866 16192 25872 16244
rect 25924 16232 25930 16244
rect 28994 16232 29000 16244
rect 25924 16204 29000 16232
rect 25924 16192 25930 16204
rect 28994 16192 29000 16204
rect 29052 16192 29058 16244
rect 29564 16204 30420 16232
rect 25685 16167 25743 16173
rect 25685 16133 25697 16167
rect 25731 16133 25743 16167
rect 25685 16127 25743 16133
rect 27706 16124 27712 16176
rect 27764 16164 27770 16176
rect 28442 16164 28448 16176
rect 27764 16136 28448 16164
rect 27764 16124 27770 16136
rect 28442 16124 28448 16136
rect 28500 16124 28506 16176
rect 19245 16068 20668 16096
rect 19245 16065 19257 16068
rect 19199 16059 19257 16065
rect 20806 16056 20812 16108
rect 20864 16056 20870 16108
rect 21818 16096 21824 16108
rect 20916 16068 21824 16096
rect 20916 16037 20944 16068
rect 21818 16056 21824 16068
rect 21876 16056 21882 16108
rect 22002 16056 22008 16108
rect 22060 16105 22066 16108
rect 24210 16105 24216 16108
rect 22060 16099 22109 16105
rect 22060 16065 22063 16099
rect 22097 16096 22109 16099
rect 24172 16099 24216 16105
rect 22097 16068 22153 16096
rect 22204 16068 23999 16096
rect 22097 16065 22109 16068
rect 22060 16059 22109 16065
rect 22060 16056 22066 16059
rect 19429 16031 19487 16037
rect 19429 16028 19441 16031
rect 18800 16000 19441 16028
rect 18693 15991 18751 15997
rect 19429 15997 19441 16000
rect 19475 15997 19487 16031
rect 19429 15991 19487 15997
rect 20901 16031 20959 16037
rect 20901 15997 20913 16031
rect 20947 15997 20959 16031
rect 20901 15991 20959 15997
rect 21545 16031 21603 16037
rect 21545 15997 21557 16031
rect 21591 16028 21603 16031
rect 22204 16028 22232 16068
rect 21591 16000 22232 16028
rect 21591 15997 21603 16000
rect 21545 15991 21603 15997
rect 17862 15960 17868 15972
rect 16500 15932 17868 15960
rect 14056 15920 14062 15932
rect 14752 15904 14780 15932
rect 17862 15920 17868 15932
rect 17920 15920 17926 15972
rect 18141 15963 18199 15969
rect 18141 15929 18153 15963
rect 18187 15960 18199 15963
rect 18708 15960 18736 15991
rect 22278 15988 22284 16040
rect 22336 15988 22342 16040
rect 23474 15988 23480 16040
rect 23532 16028 23538 16040
rect 23842 16028 23848 16040
rect 23532 16000 23848 16028
rect 23532 15988 23538 16000
rect 23842 15988 23848 16000
rect 23900 15988 23906 16040
rect 18187 15932 18736 15960
rect 21177 15963 21235 15969
rect 18187 15929 18199 15932
rect 18141 15923 18199 15929
rect 21177 15929 21189 15963
rect 21223 15960 21235 15963
rect 21450 15960 21456 15972
rect 21223 15932 21456 15960
rect 21223 15929 21235 15932
rect 21177 15923 21235 15929
rect 11011 15864 11376 15892
rect 11011 15861 11023 15864
rect 10965 15855 11023 15861
rect 11514 15852 11520 15904
rect 11572 15892 11578 15904
rect 13078 15892 13084 15904
rect 11572 15864 13084 15892
rect 11572 15852 11578 15864
rect 13078 15852 13084 15864
rect 13136 15852 13142 15904
rect 13722 15852 13728 15904
rect 13780 15852 13786 15904
rect 14734 15852 14740 15904
rect 14792 15852 14798 15904
rect 14826 15852 14832 15904
rect 14884 15892 14890 15904
rect 15203 15895 15261 15901
rect 15203 15892 15215 15895
rect 14884 15864 15215 15892
rect 14884 15852 14890 15864
rect 15203 15861 15215 15864
rect 15249 15861 15261 15895
rect 15203 15855 15261 15861
rect 16574 15852 16580 15904
rect 16632 15852 16638 15904
rect 17126 15852 17132 15904
rect 17184 15852 17190 15904
rect 17218 15852 17224 15904
rect 17276 15892 17282 15904
rect 18156 15892 18184 15923
rect 21450 15920 21456 15932
rect 21508 15920 21514 15972
rect 23661 15963 23719 15969
rect 23661 15929 23673 15963
rect 23707 15960 23719 15963
rect 23750 15960 23756 15972
rect 23707 15932 23756 15960
rect 23707 15929 23719 15932
rect 23661 15923 23719 15929
rect 23750 15920 23756 15932
rect 23808 15920 23814 15972
rect 17276 15864 18184 15892
rect 17276 15852 17282 15864
rect 18966 15852 18972 15904
rect 19024 15892 19030 15904
rect 19159 15895 19217 15901
rect 19159 15892 19171 15895
rect 19024 15864 19171 15892
rect 19024 15852 19030 15864
rect 19159 15861 19171 15864
rect 19205 15861 19217 15895
rect 19159 15855 19217 15861
rect 19518 15852 19524 15904
rect 19576 15892 19582 15904
rect 21910 15892 21916 15904
rect 19576 15864 21916 15892
rect 19576 15852 19582 15864
rect 21910 15852 21916 15864
rect 21968 15852 21974 15904
rect 22011 15895 22069 15901
rect 22011 15861 22023 15895
rect 22057 15892 22069 15895
rect 22646 15892 22652 15904
rect 22057 15864 22652 15892
rect 22057 15861 22069 15864
rect 22011 15855 22069 15861
rect 22646 15852 22652 15864
rect 22704 15852 22710 15904
rect 23971 15892 23999 16068
rect 24172 16065 24184 16099
rect 24172 16059 24216 16065
rect 24210 16056 24216 16059
rect 24268 16056 24274 16108
rect 24308 16097 24366 16103
rect 24308 16063 24320 16097
rect 24354 16063 24366 16097
rect 24308 16057 24366 16063
rect 24323 16028 24351 16057
rect 24394 16056 24400 16108
rect 24452 16096 24458 16108
rect 24581 16099 24639 16105
rect 24581 16096 24593 16099
rect 24452 16068 24593 16096
rect 24452 16056 24458 16068
rect 24581 16065 24593 16068
rect 24627 16065 24639 16099
rect 24581 16059 24639 16065
rect 25866 16056 25872 16108
rect 25924 16056 25930 16108
rect 25958 16056 25964 16108
rect 26016 16096 26022 16108
rect 26053 16099 26111 16105
rect 26053 16096 26065 16099
rect 26016 16068 26065 16096
rect 26016 16056 26022 16068
rect 26053 16065 26065 16068
rect 26099 16065 26111 16099
rect 26516 16099 26574 16105
rect 26516 16096 26528 16099
rect 26053 16059 26111 16065
rect 26344 16068 26528 16096
rect 24486 16028 24492 16040
rect 24323 16000 24492 16028
rect 24486 15988 24492 16000
rect 24544 15988 24550 16040
rect 25884 16028 25912 16056
rect 26344 16040 26372 16068
rect 26516 16065 26528 16068
rect 26562 16065 26574 16099
rect 26516 16059 26574 16065
rect 26789 16099 26847 16105
rect 26789 16065 26801 16099
rect 26835 16096 26847 16099
rect 29564 16096 29592 16204
rect 30006 16164 30012 16176
rect 26835 16094 29390 16096
rect 29472 16094 29592 16096
rect 26835 16068 29592 16094
rect 29748 16136 30012 16164
rect 26835 16065 26847 16068
rect 29362 16066 29500 16068
rect 26789 16059 26847 16065
rect 25884 16000 26188 16028
rect 25958 15920 25964 15972
rect 26016 15920 26022 15972
rect 25976 15892 26004 15920
rect 23971 15864 26004 15892
rect 26160 15892 26188 16000
rect 26326 15988 26332 16040
rect 26384 15988 26390 16040
rect 28721 16031 28779 16037
rect 28721 16028 28733 16031
rect 27540 16000 28733 16028
rect 27540 15904 27568 16000
rect 28721 15997 28733 16000
rect 28767 15997 28779 16031
rect 28721 15991 28779 15997
rect 27706 15920 27712 15972
rect 27764 15960 27770 15972
rect 28353 15963 28411 15969
rect 28353 15960 28365 15963
rect 27764 15932 28365 15960
rect 27764 15920 27770 15932
rect 28353 15929 28365 15932
rect 28399 15929 28411 15963
rect 28736 15960 28764 15991
rect 29086 15988 29092 16040
rect 29144 15988 29150 16040
rect 29178 15988 29184 16040
rect 29236 15988 29242 16040
rect 29365 16031 29423 16037
rect 29365 15997 29377 16031
rect 29411 16006 29423 16031
rect 29748 16006 29776 16136
rect 30006 16124 30012 16136
rect 30064 16124 30070 16176
rect 30392 16173 30420 16204
rect 30377 16167 30435 16173
rect 30377 16133 30389 16167
rect 30423 16133 30435 16167
rect 30377 16127 30435 16133
rect 30006 16038 30012 16040
rect 29840 16037 30012 16038
rect 29411 15997 29776 16006
rect 29365 15991 29776 15997
rect 29835 16031 30012 16037
rect 29835 15997 29847 16031
rect 29881 16010 30012 16031
rect 29881 15997 29893 16010
rect 29835 15991 29893 15997
rect 29380 15978 29776 15991
rect 30006 15988 30012 16010
rect 30064 15988 30070 16040
rect 30561 16031 30619 16037
rect 30561 15997 30573 16031
rect 30607 15997 30619 16031
rect 30561 15991 30619 15997
rect 28994 15960 29000 15972
rect 28736 15932 29000 15960
rect 28353 15923 28411 15929
rect 28994 15920 29000 15932
rect 29052 15920 29058 15972
rect 30098 15920 30104 15972
rect 30156 15920 30162 15972
rect 26519 15895 26577 15901
rect 26519 15892 26531 15895
rect 26160 15864 26531 15892
rect 26519 15861 26531 15864
rect 26565 15892 26577 15895
rect 26694 15892 26700 15904
rect 26565 15864 26700 15892
rect 26565 15861 26577 15864
rect 26519 15855 26577 15861
rect 26694 15852 26700 15864
rect 26752 15852 26758 15904
rect 27522 15852 27528 15904
rect 27580 15852 27586 15904
rect 27890 15852 27896 15904
rect 27948 15852 27954 15904
rect 29362 15852 29368 15904
rect 29420 15892 29426 15904
rect 29641 15895 29699 15901
rect 29641 15892 29653 15895
rect 29420 15864 29653 15892
rect 29420 15852 29426 15864
rect 29641 15861 29653 15864
rect 29687 15861 29699 15895
rect 30576 15892 30604 15991
rect 30576 15864 31156 15892
rect 29641 15855 29699 15861
rect 552 15802 31072 15824
rect 552 15750 7988 15802
rect 8040 15750 8052 15802
rect 8104 15750 8116 15802
rect 8168 15750 8180 15802
rect 8232 15750 8244 15802
rect 8296 15750 15578 15802
rect 15630 15750 15642 15802
rect 15694 15750 15706 15802
rect 15758 15750 15770 15802
rect 15822 15750 15834 15802
rect 15886 15750 23168 15802
rect 23220 15750 23232 15802
rect 23284 15750 23296 15802
rect 23348 15750 23360 15802
rect 23412 15750 23424 15802
rect 23476 15750 30758 15802
rect 30810 15750 30822 15802
rect 30874 15750 30886 15802
rect 30938 15750 30950 15802
rect 31002 15750 31014 15802
rect 31066 15750 31072 15802
rect 552 15728 31072 15750
rect 3050 15688 3056 15700
rect 1228 15660 3056 15688
rect 1228 15561 1256 15660
rect 3050 15648 3056 15660
rect 3108 15648 3114 15700
rect 3142 15648 3148 15700
rect 3200 15648 3206 15700
rect 5534 15648 5540 15700
rect 5592 15648 5598 15700
rect 10410 15688 10416 15700
rect 5828 15660 10416 15688
rect 1213 15555 1271 15561
rect 1213 15521 1225 15555
rect 1259 15521 1271 15555
rect 4249 15555 4307 15561
rect 1213 15515 1271 15521
rect 1964 15524 4200 15552
rect 1801 15505 1859 15511
rect 1670 15493 1676 15496
rect 1305 15487 1363 15493
rect 1305 15453 1317 15487
rect 1351 15453 1363 15487
rect 1305 15447 1363 15453
rect 1632 15487 1676 15493
rect 1632 15453 1644 15487
rect 1632 15447 1676 15453
rect 1320 15360 1348 15447
rect 1670 15444 1676 15447
rect 1728 15444 1734 15496
rect 1801 15471 1813 15505
rect 1847 15484 1859 15505
rect 1964 15484 1992 15524
rect 1847 15471 1992 15484
rect 1801 15465 1992 15471
rect 1826 15456 1992 15465
rect 2038 15444 2044 15496
rect 2096 15444 2102 15496
rect 3510 15444 3516 15496
rect 3568 15444 3574 15496
rect 3878 15493 3884 15496
rect 3840 15487 3884 15493
rect 3840 15453 3852 15487
rect 3840 15447 3884 15453
rect 3878 15444 3884 15447
rect 3936 15444 3942 15496
rect 3976 15489 4034 15495
rect 3976 15455 3988 15489
rect 4022 15484 4034 15489
rect 4062 15484 4068 15496
rect 4022 15456 4068 15484
rect 4022 15455 4034 15456
rect 3976 15449 4034 15455
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 4172 15484 4200 15524
rect 4249 15521 4261 15555
rect 4295 15552 4307 15555
rect 4522 15552 4528 15564
rect 4295 15524 4528 15552
rect 4295 15521 4307 15524
rect 4249 15515 4307 15521
rect 4522 15512 4528 15524
rect 4580 15512 4586 15564
rect 5828 15484 5856 15660
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 11514 15688 11520 15700
rect 10980 15660 11520 15688
rect 5905 15555 5963 15561
rect 5905 15521 5917 15555
rect 5951 15521 5963 15555
rect 5905 15515 5963 15521
rect 4172 15456 5856 15484
rect 1026 15308 1032 15360
rect 1084 15308 1090 15360
rect 1302 15308 1308 15360
rect 1360 15348 1366 15360
rect 3528 15348 3556 15444
rect 3786 15348 3792 15360
rect 1360 15320 3792 15348
rect 1360 15308 1366 15320
rect 3786 15308 3792 15320
rect 3844 15348 3850 15360
rect 5920 15348 5948 15515
rect 6454 15512 6460 15564
rect 6512 15552 6518 15564
rect 6692 15555 6750 15561
rect 6692 15552 6704 15555
rect 6512 15524 6704 15552
rect 6512 15512 6518 15524
rect 6692 15521 6704 15524
rect 6738 15521 6750 15555
rect 8294 15552 8300 15564
rect 6692 15515 6750 15521
rect 7024 15524 8300 15552
rect 6828 15505 6886 15511
rect 6365 15487 6423 15493
rect 6365 15484 6377 15487
rect 6196 15456 6377 15484
rect 6196 15360 6224 15456
rect 6365 15453 6377 15456
rect 6411 15453 6423 15487
rect 6828 15471 6840 15505
rect 6874 15484 6886 15505
rect 7024 15484 7052 15524
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 8662 15512 8668 15564
rect 8720 15512 8726 15564
rect 10980 15552 11008 15660
rect 11514 15648 11520 15660
rect 11572 15648 11578 15700
rect 11606 15648 11612 15700
rect 11664 15688 11670 15700
rect 12075 15691 12133 15697
rect 12075 15688 12087 15691
rect 11664 15660 12087 15688
rect 11664 15648 11670 15660
rect 12075 15657 12087 15660
rect 12121 15657 12133 15691
rect 12075 15651 12133 15657
rect 13446 15648 13452 15700
rect 13504 15648 13510 15700
rect 16574 15688 16580 15700
rect 13556 15660 16580 15688
rect 9232 15524 11008 15552
rect 11057 15555 11115 15561
rect 6874 15471 7052 15484
rect 6828 15465 7052 15471
rect 6843 15456 7052 15465
rect 6365 15447 6423 15453
rect 7098 15444 7104 15496
rect 7156 15444 7162 15496
rect 8202 15444 8208 15496
rect 8260 15484 8266 15496
rect 8573 15487 8631 15493
rect 8573 15484 8585 15487
rect 8260 15456 8585 15484
rect 8260 15444 8266 15456
rect 8573 15453 8585 15456
rect 8619 15484 8631 15487
rect 8680 15484 8708 15512
rect 9069 15505 9127 15511
rect 8938 15493 8944 15496
rect 8619 15456 8708 15484
rect 8900 15487 8944 15493
rect 8619 15453 8631 15456
rect 8573 15447 8631 15453
rect 8900 15453 8912 15487
rect 8900 15447 8944 15453
rect 3844 15320 5948 15348
rect 3844 15308 3850 15320
rect 6178 15308 6184 15360
rect 6236 15308 6242 15360
rect 6270 15308 6276 15360
rect 6328 15348 6334 15360
rect 8205 15351 8263 15357
rect 8205 15348 8217 15351
rect 6328 15320 8217 15348
rect 6328 15308 6334 15320
rect 8205 15317 8217 15320
rect 8251 15317 8263 15351
rect 8588 15348 8616 15447
rect 8938 15444 8944 15447
rect 8996 15444 9002 15496
rect 9069 15471 9081 15505
rect 9115 15484 9127 15505
rect 9232 15484 9260 15524
rect 11057 15521 11069 15555
rect 11103 15521 11115 15555
rect 13556 15552 13584 15660
rect 16574 15648 16580 15660
rect 16632 15648 16638 15700
rect 16942 15648 16948 15700
rect 17000 15648 17006 15700
rect 17034 15648 17040 15700
rect 17092 15688 17098 15700
rect 17129 15691 17187 15697
rect 17129 15688 17141 15691
rect 17092 15660 17141 15688
rect 17092 15648 17098 15660
rect 17129 15657 17141 15660
rect 17175 15657 17187 15691
rect 17129 15651 17187 15657
rect 17586 15648 17592 15700
rect 17644 15688 17650 15700
rect 20714 15688 20720 15700
rect 17644 15660 20720 15688
rect 17644 15648 17650 15660
rect 20714 15648 20720 15660
rect 20772 15648 20778 15700
rect 20993 15691 21051 15697
rect 20993 15657 21005 15691
rect 21039 15688 21051 15691
rect 22830 15688 22836 15700
rect 21039 15660 22836 15688
rect 21039 15657 21051 15660
rect 20993 15651 21051 15657
rect 22830 15648 22836 15660
rect 22888 15648 22894 15700
rect 23014 15648 23020 15700
rect 23072 15648 23078 15700
rect 23943 15691 24001 15697
rect 23943 15657 23955 15691
rect 23989 15688 24001 15691
rect 24210 15688 24216 15700
rect 23989 15660 24216 15688
rect 23989 15657 24001 15660
rect 23943 15651 24001 15657
rect 24210 15648 24216 15660
rect 24268 15648 24274 15700
rect 24486 15648 24492 15700
rect 24544 15688 24550 15700
rect 28261 15691 28319 15697
rect 28261 15688 28273 15691
rect 24544 15660 28273 15688
rect 24544 15648 24550 15660
rect 28261 15657 28273 15660
rect 28307 15657 28319 15691
rect 28261 15651 28319 15657
rect 30377 15691 30435 15697
rect 30377 15657 30389 15691
rect 30423 15657 30435 15691
rect 30377 15651 30435 15657
rect 15930 15580 15936 15632
rect 15988 15580 15994 15632
rect 14182 15561 14188 15564
rect 11057 15515 11115 15521
rect 12268 15524 13584 15552
rect 14144 15555 14188 15561
rect 9115 15471 9260 15484
rect 9069 15465 9260 15471
rect 9084 15456 9260 15465
rect 9306 15444 9312 15496
rect 9364 15444 9370 15496
rect 11072 15416 11100 15515
rect 11609 15487 11667 15493
rect 11609 15453 11621 15487
rect 11655 15453 11667 15487
rect 11609 15447 11667 15453
rect 12115 15487 12173 15493
rect 12115 15453 12127 15487
rect 12161 15484 12173 15487
rect 12268 15484 12296 15524
rect 14144 15521 14156 15555
rect 14240 15552 14246 15564
rect 14826 15552 14832 15564
rect 14240 15524 14832 15552
rect 14144 15515 14188 15521
rect 14182 15512 14188 15515
rect 14240 15512 14246 15524
rect 14826 15512 14832 15524
rect 14884 15512 14890 15564
rect 16960 15561 16988 15648
rect 19518 15620 19524 15632
rect 19306 15592 19524 15620
rect 16117 15555 16175 15561
rect 16117 15552 16129 15555
rect 16040 15524 16129 15552
rect 16040 15496 16068 15524
rect 16117 15521 16129 15524
rect 16163 15552 16175 15555
rect 16669 15555 16727 15561
rect 16669 15552 16681 15555
rect 16163 15524 16681 15552
rect 16163 15521 16175 15524
rect 16117 15515 16175 15521
rect 16669 15521 16681 15524
rect 16715 15521 16727 15555
rect 16669 15515 16727 15521
rect 16945 15555 17003 15561
rect 16945 15521 16957 15555
rect 16991 15521 17003 15555
rect 17494 15552 17500 15564
rect 16945 15515 17003 15521
rect 17144 15524 17500 15552
rect 12161 15456 12296 15484
rect 12161 15453 12173 15456
rect 12115 15447 12173 15453
rect 9968 15388 11100 15416
rect 9968 15348 9996 15388
rect 11238 15376 11244 15428
rect 11296 15416 11302 15428
rect 11624 15416 11652 15447
rect 12342 15444 12348 15496
rect 12400 15444 12406 15496
rect 13814 15444 13820 15496
rect 13872 15444 13878 15496
rect 14323 15487 14381 15493
rect 14323 15453 14335 15487
rect 14369 15484 14381 15487
rect 14458 15484 14464 15496
rect 14369 15456 14464 15484
rect 14369 15453 14381 15456
rect 14323 15447 14381 15453
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 14553 15487 14611 15493
rect 14553 15453 14565 15487
rect 14599 15484 14611 15487
rect 15378 15484 15384 15496
rect 14599 15456 15384 15484
rect 14599 15453 14611 15456
rect 14553 15447 14611 15453
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 16022 15444 16028 15496
rect 16080 15444 16086 15496
rect 16393 15487 16451 15493
rect 16393 15453 16405 15487
rect 16439 15453 16451 15487
rect 16393 15447 16451 15453
rect 16408 15416 16436 15447
rect 16758 15444 16764 15496
rect 16816 15484 16822 15496
rect 17144 15484 17172 15524
rect 17494 15512 17500 15524
rect 17552 15561 17558 15564
rect 17552 15555 17606 15561
rect 17552 15521 17560 15555
rect 17594 15521 17606 15555
rect 17552 15515 17606 15521
rect 17880 15524 18092 15552
rect 17552 15512 17558 15515
rect 16816 15456 17172 15484
rect 16816 15444 16822 15456
rect 17218 15444 17224 15496
rect 17276 15444 17282 15496
rect 17727 15487 17785 15493
rect 17727 15453 17739 15487
rect 17773 15484 17785 15487
rect 17880 15484 17908 15524
rect 17773 15456 17908 15484
rect 17773 15453 17785 15456
rect 17727 15447 17785 15453
rect 17954 15444 17960 15496
rect 18012 15444 18018 15496
rect 18064 15484 18092 15524
rect 18598 15512 18604 15564
rect 18656 15552 18662 15564
rect 19306 15552 19334 15592
rect 19518 15580 19524 15592
rect 19576 15580 19582 15632
rect 18656 15524 19334 15552
rect 18656 15512 18662 15524
rect 19702 15512 19708 15564
rect 19760 15512 19766 15564
rect 19794 15512 19800 15564
rect 19852 15552 19858 15564
rect 21358 15552 21364 15564
rect 19852 15524 21364 15552
rect 19852 15512 19858 15524
rect 21358 15512 21364 15524
rect 21416 15512 21422 15564
rect 23032 15552 23060 15648
rect 26234 15580 26240 15632
rect 26292 15580 26298 15632
rect 29730 15580 29736 15632
rect 29788 15620 29794 15632
rect 30392 15620 30420 15651
rect 31128 15620 31156 15864
rect 29788 15592 30420 15620
rect 30484 15592 31156 15620
rect 29788 15580 29794 15592
rect 21790 15524 23060 15552
rect 18064 15456 19380 15484
rect 11296 15388 11652 15416
rect 15212 15388 16436 15416
rect 11296 15376 11302 15388
rect 8588 15320 9996 15348
rect 8205 15311 8263 15317
rect 10410 15308 10416 15360
rect 10468 15308 10474 15360
rect 10502 15308 10508 15360
rect 10560 15348 10566 15360
rect 15212 15348 15240 15388
rect 16850 15376 16856 15428
rect 16908 15376 16914 15428
rect 17236 15416 17264 15444
rect 17052 15388 17264 15416
rect 10560 15320 15240 15348
rect 10560 15308 10566 15320
rect 15562 15308 15568 15360
rect 15620 15348 15626 15360
rect 16301 15351 16359 15357
rect 16301 15348 16313 15351
rect 15620 15320 16313 15348
rect 15620 15308 15626 15320
rect 16301 15317 16313 15320
rect 16347 15348 16359 15351
rect 16390 15348 16396 15360
rect 16347 15320 16396 15348
rect 16347 15317 16359 15320
rect 16301 15311 16359 15317
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 16574 15308 16580 15360
rect 16632 15348 16638 15360
rect 17052 15348 17080 15388
rect 16632 15320 17080 15348
rect 16632 15308 16638 15320
rect 19058 15308 19064 15360
rect 19116 15308 19122 15360
rect 19352 15348 19380 15456
rect 19426 15444 19432 15496
rect 19484 15444 19490 15496
rect 21266 15444 21272 15496
rect 21324 15444 21330 15496
rect 21450 15444 21456 15496
rect 21508 15484 21514 15496
rect 21790 15493 21818 15524
rect 23750 15512 23756 15564
rect 23808 15552 23814 15564
rect 23808 15524 23983 15552
rect 23808 15512 23814 15524
rect 21596 15487 21654 15493
rect 21596 15484 21608 15487
rect 21508 15456 21608 15484
rect 21508 15444 21514 15456
rect 21596 15453 21608 15456
rect 21642 15453 21654 15487
rect 21596 15447 21654 15453
rect 21775 15487 21833 15493
rect 21775 15453 21787 15487
rect 21821 15453 21833 15487
rect 21775 15447 21833 15453
rect 21910 15444 21916 15496
rect 21968 15493 21974 15496
rect 21968 15487 22017 15493
rect 21968 15453 21971 15487
rect 22005 15453 22017 15487
rect 21968 15447 22017 15453
rect 23477 15487 23535 15493
rect 23477 15453 23489 15487
rect 23523 15484 23535 15487
rect 23842 15484 23848 15496
rect 23523 15456 23848 15484
rect 23523 15453 23535 15456
rect 23477 15447 23535 15453
rect 21968 15444 21974 15447
rect 23842 15444 23848 15456
rect 23900 15444 23906 15496
rect 23955 15495 23983 15524
rect 24670 15512 24676 15564
rect 24728 15552 24734 15564
rect 25866 15552 25872 15564
rect 24728 15524 25872 15552
rect 24728 15512 24734 15524
rect 25866 15512 25872 15524
rect 25924 15512 25930 15564
rect 25958 15512 25964 15564
rect 26016 15552 26022 15564
rect 26421 15555 26479 15561
rect 26421 15552 26433 15555
rect 26016 15524 26433 15552
rect 26016 15512 26022 15524
rect 26421 15521 26433 15524
rect 26467 15521 26479 15555
rect 26421 15515 26479 15521
rect 23940 15489 23998 15495
rect 23940 15455 23952 15489
rect 23986 15455 23998 15489
rect 23940 15449 23998 15455
rect 24210 15444 24216 15496
rect 24268 15444 24274 15496
rect 19702 15348 19708 15360
rect 19352 15320 19708 15348
rect 19702 15308 19708 15320
rect 19760 15308 19766 15360
rect 19794 15308 19800 15360
rect 19852 15348 19858 15360
rect 23109 15351 23167 15357
rect 23109 15348 23121 15351
rect 19852 15320 23121 15348
rect 19852 15308 19858 15320
rect 23109 15317 23121 15320
rect 23155 15317 23167 15351
rect 23109 15311 23167 15317
rect 23658 15308 23664 15360
rect 23716 15348 23722 15360
rect 25317 15351 25375 15357
rect 25317 15348 25329 15351
rect 23716 15320 25329 15348
rect 23716 15308 23722 15320
rect 25317 15317 25329 15320
rect 25363 15317 25375 15351
rect 26436 15348 26464 15515
rect 26694 15512 26700 15564
rect 26752 15561 26758 15564
rect 26752 15555 26806 15561
rect 26752 15521 26760 15555
rect 26794 15521 26806 15555
rect 26752 15515 26806 15521
rect 26752 15512 26758 15515
rect 26970 15512 26976 15564
rect 27028 15552 27034 15564
rect 27157 15555 27215 15561
rect 27157 15552 27169 15555
rect 27028 15524 27169 15552
rect 27028 15512 27034 15524
rect 27157 15521 27169 15524
rect 27203 15521 27215 15555
rect 27157 15515 27215 15521
rect 28718 15512 28724 15564
rect 28776 15552 28782 15564
rect 28905 15555 28963 15561
rect 28905 15552 28917 15555
rect 28776 15524 28917 15552
rect 28776 15512 28782 15524
rect 28905 15521 28917 15524
rect 28951 15521 28963 15555
rect 28905 15515 28963 15521
rect 28994 15512 29000 15564
rect 29052 15552 29058 15564
rect 30484 15552 30512 15592
rect 29052 15524 30512 15552
rect 30561 15555 30619 15561
rect 29052 15512 29058 15524
rect 30561 15521 30573 15555
rect 30607 15552 30619 15555
rect 30607 15524 30696 15552
rect 30607 15521 30619 15524
rect 30561 15515 30619 15521
rect 30668 15496 30696 15524
rect 26878 15444 26884 15496
rect 26936 15444 26942 15496
rect 28629 15487 28687 15493
rect 28629 15453 28641 15487
rect 28675 15484 28687 15487
rect 28810 15484 28816 15496
rect 28675 15456 28816 15484
rect 28675 15453 28687 15456
rect 28629 15447 28687 15453
rect 28810 15444 28816 15456
rect 28868 15444 28874 15496
rect 29362 15444 29368 15496
rect 29420 15484 29426 15496
rect 30282 15484 30288 15496
rect 29420 15456 30288 15484
rect 29420 15444 29426 15456
rect 30282 15444 30288 15456
rect 30340 15444 30346 15496
rect 30650 15444 30656 15496
rect 30708 15444 30714 15496
rect 28810 15348 28816 15360
rect 26436 15320 28816 15348
rect 25317 15311 25375 15317
rect 28810 15308 28816 15320
rect 28868 15308 28874 15360
rect 30006 15308 30012 15360
rect 30064 15308 30070 15360
rect 552 15258 30912 15280
rect 552 15206 4193 15258
rect 4245 15206 4257 15258
rect 4309 15206 4321 15258
rect 4373 15206 4385 15258
rect 4437 15206 4449 15258
rect 4501 15206 11783 15258
rect 11835 15206 11847 15258
rect 11899 15206 11911 15258
rect 11963 15206 11975 15258
rect 12027 15206 12039 15258
rect 12091 15206 19373 15258
rect 19425 15206 19437 15258
rect 19489 15206 19501 15258
rect 19553 15206 19565 15258
rect 19617 15206 19629 15258
rect 19681 15206 26963 15258
rect 27015 15206 27027 15258
rect 27079 15206 27091 15258
rect 27143 15206 27155 15258
rect 27207 15206 27219 15258
rect 27271 15206 30912 15258
rect 552 15184 30912 15206
rect 2774 15104 2780 15156
rect 2832 15104 2838 15156
rect 5813 15147 5871 15153
rect 3712 15116 5212 15144
rect 2498 15036 2504 15088
rect 2556 15076 2562 15088
rect 3510 15076 3516 15088
rect 2556 15048 3516 15076
rect 2556 15036 2562 15048
rect 3510 15036 3516 15048
rect 3568 15036 3574 15088
rect 937 15011 995 15017
rect 937 14977 949 15011
rect 983 15008 995 15011
rect 1302 15008 1308 15020
rect 983 14980 1308 15008
rect 983 14977 995 14980
rect 937 14971 995 14977
rect 1302 14968 1308 14980
rect 1360 14968 1366 15020
rect 1443 15011 1501 15017
rect 1443 14977 1455 15011
rect 1489 15008 1501 15011
rect 2130 15008 2136 15020
rect 1489 14980 2136 15008
rect 1489 14977 1501 14980
rect 1443 14971 1501 14977
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 1673 14943 1731 14949
rect 1673 14909 1685 14943
rect 1719 14940 1731 14943
rect 1762 14940 1768 14952
rect 1719 14912 1768 14940
rect 1719 14909 1731 14912
rect 1673 14903 1731 14909
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 3234 14900 3240 14952
rect 3292 14940 3298 14952
rect 3712 14940 3740 15116
rect 5184 15076 5212 15116
rect 5813 15113 5825 15147
rect 5859 15144 5871 15147
rect 6362 15144 6368 15156
rect 5859 15116 6368 15144
rect 5859 15113 5871 15116
rect 5813 15107 5871 15113
rect 6362 15104 6368 15116
rect 6420 15104 6426 15156
rect 6730 15104 6736 15156
rect 6788 15144 6794 15156
rect 7929 15147 7987 15153
rect 7929 15144 7941 15147
rect 6788 15116 7941 15144
rect 6788 15104 6794 15116
rect 7929 15113 7941 15116
rect 7975 15113 7987 15147
rect 10502 15144 10508 15156
rect 7929 15107 7987 15113
rect 8128 15116 10508 15144
rect 6086 15076 6092 15088
rect 5184 15048 6092 15076
rect 6086 15036 6092 15048
rect 6144 15036 6150 15088
rect 3786 14968 3792 15020
rect 3844 14968 3850 15020
rect 4295 15011 4353 15017
rect 4295 14977 4307 15011
rect 4341 15008 4353 15011
rect 6270 15008 6276 15020
rect 4341 14980 6276 15008
rect 4341 14977 4353 14980
rect 4295 14971 4353 14977
rect 6270 14968 6276 14980
rect 6328 14968 6334 15020
rect 6595 15011 6653 15017
rect 6595 14977 6607 15011
rect 6641 15008 6653 15011
rect 8128 15008 8156 15116
rect 10502 15104 10508 15116
rect 10560 15104 10566 15156
rect 13722 15144 13728 15156
rect 11262 15116 13728 15144
rect 10134 15036 10140 15088
rect 10192 15076 10198 15088
rect 10413 15079 10471 15085
rect 10413 15076 10425 15079
rect 10192 15048 10425 15076
rect 10192 15036 10198 15048
rect 10413 15045 10425 15048
rect 10459 15045 10471 15079
rect 10413 15039 10471 15045
rect 10594 15036 10600 15088
rect 10652 15076 10658 15088
rect 10965 15079 11023 15085
rect 10965 15076 10977 15079
rect 10652 15048 10977 15076
rect 10652 15036 10658 15048
rect 10965 15045 10977 15048
rect 11011 15045 11023 15079
rect 10965 15039 11023 15045
rect 6641 14980 8156 15008
rect 6641 14977 6653 14980
rect 6595 14971 6653 14977
rect 8202 14968 8208 15020
rect 8260 15008 8266 15020
rect 8573 15011 8631 15017
rect 8573 15008 8585 15011
rect 8260 14980 8585 15008
rect 8260 14968 8266 14980
rect 8573 14977 8585 14980
rect 8619 14977 8631 15011
rect 8573 14971 8631 14977
rect 9048 14993 9996 15008
rect 9048 14962 9081 14993
rect 9069 14959 9081 14962
rect 9115 14980 9996 14993
rect 9115 14959 9127 14980
rect 9069 14953 9127 14959
rect 3292 14912 3740 14940
rect 3292 14900 3298 14912
rect 3878 14900 3884 14952
rect 3936 14940 3942 14952
rect 4116 14943 4174 14949
rect 4116 14940 4128 14943
rect 3936 14912 4128 14940
rect 3936 14900 3942 14912
rect 4116 14909 4128 14912
rect 4162 14909 4174 14943
rect 4116 14903 4174 14909
rect 4522 14900 4528 14952
rect 4580 14900 4586 14952
rect 6089 14943 6147 14949
rect 6089 14909 6101 14943
rect 6135 14909 6147 14943
rect 6089 14903 6147 14909
rect 3513 14875 3571 14881
rect 3513 14872 3525 14875
rect 2746 14844 3525 14872
rect 1403 14807 1461 14813
rect 1403 14773 1415 14807
rect 1449 14804 1461 14807
rect 1670 14804 1676 14816
rect 1449 14776 1676 14804
rect 1449 14773 1461 14776
rect 1403 14767 1461 14773
rect 1670 14764 1676 14776
rect 1728 14804 1734 14816
rect 2746 14804 2774 14844
rect 3513 14841 3525 14844
rect 3559 14872 3571 14875
rect 3896 14872 3924 14900
rect 3559 14844 3924 14872
rect 3559 14841 3571 14844
rect 3513 14835 3571 14841
rect 6104 14816 6132 14903
rect 6362 14900 6368 14952
rect 6420 14940 6426 14952
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6420 14912 6837 14940
rect 6420 14900 6426 14912
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 9309 14943 9367 14949
rect 9309 14909 9321 14943
rect 9355 14940 9367 14943
rect 9674 14940 9680 14952
rect 9355 14912 9680 14940
rect 9355 14909 9367 14912
rect 9309 14903 9367 14909
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 9968 14940 9996 14980
rect 10226 14968 10232 15020
rect 10284 15008 10290 15020
rect 11262 15008 11290 15116
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 16025 15147 16083 15153
rect 16025 15144 16037 15147
rect 13883 15116 16037 15144
rect 11606 15017 11612 15020
rect 10284 14980 11290 15008
rect 11568 15011 11612 15017
rect 10284 14968 10290 14980
rect 11568 14977 11580 15011
rect 11568 14971 11612 14977
rect 11606 14968 11612 14971
rect 11664 14968 11670 15020
rect 11747 15011 11805 15017
rect 11747 14977 11759 15011
rect 11793 15008 11805 15011
rect 11882 15008 11888 15020
rect 11793 14980 11888 15008
rect 11793 14977 11805 14980
rect 11747 14971 11805 14977
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 11974 14966 11980 15018
rect 12032 14966 12038 15018
rect 12066 14968 12072 15020
rect 12124 15008 12130 15020
rect 13883 15008 13911 15116
rect 16025 15113 16037 15116
rect 16071 15113 16083 15147
rect 16025 15107 16083 15113
rect 18046 15104 18052 15156
rect 18104 15144 18110 15156
rect 19245 15147 19303 15153
rect 19245 15144 19257 15147
rect 18104 15116 19257 15144
rect 18104 15104 18110 15116
rect 19245 15113 19257 15116
rect 19291 15113 19303 15147
rect 19245 15107 19303 15113
rect 19521 15147 19579 15153
rect 19521 15113 19533 15147
rect 19567 15144 19579 15147
rect 21910 15144 21916 15156
rect 19567 15116 21916 15144
rect 19567 15113 19579 15116
rect 19521 15107 19579 15113
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 22189 15147 22247 15153
rect 22189 15113 22201 15147
rect 22235 15144 22247 15147
rect 23017 15147 23075 15153
rect 22235 15116 22968 15144
rect 22235 15113 22247 15116
rect 22189 15107 22247 15113
rect 17862 15036 17868 15088
rect 17920 15076 17926 15088
rect 18233 15079 18291 15085
rect 18233 15076 18245 15079
rect 17920 15048 18245 15076
rect 17920 15036 17926 15048
rect 18233 15045 18245 15048
rect 18279 15045 18291 15079
rect 18233 15039 18291 15045
rect 22462 15036 22468 15088
rect 22520 15036 22526 15088
rect 22940 15076 22968 15116
rect 23017 15113 23029 15147
rect 23063 15144 23075 15147
rect 24210 15144 24216 15156
rect 23063 15116 24216 15144
rect 23063 15113 23075 15116
rect 23017 15107 23075 15113
rect 24210 15104 24216 15116
rect 24268 15104 24274 15156
rect 24946 15104 24952 15156
rect 25004 15144 25010 15156
rect 27522 15144 27528 15156
rect 25004 15116 27528 15144
rect 25004 15104 25010 15116
rect 27522 15104 27528 15116
rect 27580 15104 27586 15156
rect 27798 15104 27804 15156
rect 27856 15144 27862 15156
rect 27893 15147 27951 15153
rect 27893 15144 27905 15147
rect 27856 15116 27905 15144
rect 27856 15104 27862 15116
rect 27893 15113 27905 15116
rect 27939 15113 27951 15147
rect 30098 15144 30104 15156
rect 27893 15107 27951 15113
rect 28276 15116 30104 15144
rect 23566 15076 23572 15088
rect 22940 15048 23572 15076
rect 23566 15036 23572 15048
rect 23624 15036 23630 15088
rect 26050 15076 26056 15088
rect 25884 15048 26056 15076
rect 12124 14980 13911 15008
rect 14691 15011 14749 15017
rect 12124 14968 12130 14980
rect 14691 14977 14703 15011
rect 14737 15008 14749 15011
rect 16393 15011 16451 15017
rect 14737 14980 15608 15008
rect 14737 14977 14749 14980
rect 14691 14971 14749 14977
rect 10870 14940 10876 14952
rect 9968 14912 10876 14940
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 11146 14900 11152 14952
rect 11204 14900 11210 14952
rect 11238 14900 11244 14952
rect 11296 14940 11302 14952
rect 13633 14943 13691 14949
rect 13633 14940 13645 14943
rect 11296 14936 11928 14940
rect 12084 14936 13645 14940
rect 11296 14912 13645 14936
rect 11296 14900 11302 14912
rect 11900 14908 12112 14912
rect 13633 14909 13645 14912
rect 13679 14909 13691 14943
rect 13633 14903 13691 14909
rect 13814 14900 13820 14952
rect 13872 14940 13878 14952
rect 14185 14943 14243 14949
rect 14185 14940 14197 14943
rect 13872 14912 14197 14940
rect 13872 14900 13878 14912
rect 14185 14909 14197 14912
rect 14231 14909 14243 14943
rect 14921 14943 14979 14949
rect 14921 14940 14933 14943
rect 14185 14903 14243 14909
rect 14292 14912 14933 14940
rect 14292 14872 14320 14912
rect 14921 14909 14933 14912
rect 14967 14909 14979 14943
rect 14921 14903 14979 14909
rect 10336 14844 11100 14872
rect 1728 14776 2774 14804
rect 1728 14764 1734 14776
rect 3602 14764 3608 14816
rect 3660 14804 3666 14816
rect 4614 14804 4620 14816
rect 3660 14776 4620 14804
rect 3660 14764 3666 14776
rect 4614 14764 4620 14776
rect 4672 14804 4678 14816
rect 5534 14804 5540 14816
rect 4672 14776 5540 14804
rect 4672 14764 4678 14776
rect 5534 14764 5540 14776
rect 5592 14804 5598 14816
rect 5902 14804 5908 14816
rect 5592 14776 5908 14804
rect 5592 14764 5598 14776
rect 5902 14764 5908 14776
rect 5960 14764 5966 14816
rect 6086 14764 6092 14816
rect 6144 14764 6150 14816
rect 6454 14764 6460 14816
rect 6512 14804 6518 14816
rect 6555 14807 6613 14813
rect 6555 14804 6567 14807
rect 6512 14776 6567 14804
rect 6512 14764 6518 14776
rect 6555 14773 6567 14776
rect 6601 14804 6613 14807
rect 8938 14804 8944 14816
rect 6601 14776 8944 14804
rect 6601 14773 6613 14776
rect 6555 14767 6613 14773
rect 8938 14764 8944 14776
rect 8996 14804 9002 14816
rect 9039 14807 9097 14813
rect 9039 14804 9051 14807
rect 8996 14776 9051 14804
rect 8996 14764 9002 14776
rect 9039 14773 9051 14776
rect 9085 14773 9097 14807
rect 9039 14767 9097 14773
rect 9766 14764 9772 14816
rect 9824 14804 9830 14816
rect 10336 14804 10364 14844
rect 9824 14776 10364 14804
rect 11072 14804 11100 14844
rect 13648 14844 14320 14872
rect 13648 14816 13676 14844
rect 13081 14807 13139 14813
rect 13081 14804 13093 14807
rect 11072 14776 13093 14804
rect 9824 14764 9830 14776
rect 13081 14773 13093 14776
rect 13127 14773 13139 14807
rect 13081 14767 13139 14773
rect 13630 14764 13636 14816
rect 13688 14764 13694 14816
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 13909 14807 13967 14813
rect 13909 14804 13921 14807
rect 13872 14776 13921 14804
rect 13872 14764 13878 14776
rect 13909 14773 13921 14776
rect 13955 14773 13967 14807
rect 13909 14767 13967 14773
rect 14651 14807 14709 14813
rect 14651 14773 14663 14807
rect 14697 14804 14709 14807
rect 14826 14804 14832 14816
rect 14697 14776 14832 14804
rect 14697 14773 14709 14776
rect 14651 14767 14709 14773
rect 14826 14764 14832 14776
rect 14884 14764 14890 14816
rect 15580 14804 15608 14980
rect 16393 14977 16405 15011
rect 16439 15008 16451 15011
rect 16574 15008 16580 15020
rect 16439 14980 16580 15008
rect 16439 14977 16451 14980
rect 16393 14971 16451 14977
rect 16574 14968 16580 14980
rect 16632 14968 16638 15020
rect 16899 15011 16957 15017
rect 16899 14977 16911 15011
rect 16945 15008 16957 15011
rect 19794 15008 19800 15020
rect 16945 14980 19800 15008
rect 16945 14977 16957 14980
rect 16899 14971 16957 14977
rect 19794 14968 19800 14980
rect 19852 14968 19858 15020
rect 19886 14968 19892 15020
rect 19944 14968 19950 15020
rect 20395 15011 20453 15017
rect 20395 14977 20407 15011
rect 20441 15008 20453 15011
rect 20530 15008 20536 15020
rect 20441 14980 20536 15008
rect 20441 14977 20453 14980
rect 20395 14971 20453 14977
rect 20530 14968 20536 14980
rect 20588 14968 20594 15020
rect 20622 14968 20628 15020
rect 20680 14968 20686 15020
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 20772 14980 22692 15008
rect 20772 14968 20778 14980
rect 17129 14943 17187 14949
rect 17129 14909 17141 14943
rect 17175 14940 17187 14943
rect 17175 14912 18552 14940
rect 17175 14909 17187 14912
rect 17129 14903 17187 14909
rect 18524 14872 18552 14912
rect 18690 14900 18696 14952
rect 18748 14900 18754 14952
rect 19429 14943 19487 14949
rect 19429 14909 19441 14943
rect 19475 14909 19487 14943
rect 19429 14903 19487 14909
rect 18874 14872 18880 14884
rect 18524 14844 18880 14872
rect 18874 14832 18880 14844
rect 18932 14832 18938 14884
rect 18966 14832 18972 14884
rect 19024 14832 19030 14884
rect 19444 14872 19472 14903
rect 19702 14900 19708 14952
rect 19760 14940 19766 14952
rect 22664 14949 22692 14980
rect 22830 14968 22836 15020
rect 22888 15008 22894 15020
rect 22888 14980 22968 15008
rect 22888 14968 22894 14980
rect 22940 14949 22968 14980
rect 23750 14968 23756 15020
rect 23808 14968 23814 15020
rect 24210 15017 24216 15020
rect 24172 15011 24216 15017
rect 24172 14977 24184 15011
rect 24172 14971 24216 14977
rect 24210 14968 24216 14971
rect 24268 14968 24274 15020
rect 24341 15011 24399 15017
rect 24341 14977 24353 15011
rect 24387 15008 24399 15011
rect 25884 15008 25912 15048
rect 26050 15036 26056 15048
rect 26108 15036 26114 15088
rect 24387 14980 25912 15008
rect 24387 14977 24399 14980
rect 24341 14971 24399 14977
rect 25958 14968 25964 15020
rect 26016 14968 26022 15020
rect 26516 15011 26574 15017
rect 26516 15008 26528 15011
rect 26160 14980 26528 15008
rect 22373 14943 22431 14949
rect 22373 14940 22385 14943
rect 19760 14912 22385 14940
rect 19760 14900 19766 14912
rect 22373 14909 22385 14912
rect 22419 14909 22431 14943
rect 22373 14903 22431 14909
rect 22649 14943 22707 14949
rect 22649 14909 22661 14943
rect 22695 14940 22707 14943
rect 22925 14943 22983 14949
rect 22695 14912 22876 14940
rect 22695 14909 22707 14912
rect 22649 14903 22707 14909
rect 19978 14872 19984 14884
rect 19444 14844 19984 14872
rect 19978 14832 19984 14844
rect 20036 14832 20042 14884
rect 22388 14872 22416 14903
rect 22848 14872 22876 14912
rect 22925 14909 22937 14943
rect 22971 14909 22983 14943
rect 22925 14903 22983 14909
rect 23198 14900 23204 14952
rect 23256 14900 23262 14952
rect 23661 14943 23719 14949
rect 23661 14940 23673 14943
rect 23308 14912 23673 14940
rect 23014 14872 23020 14884
rect 22388 14844 22692 14872
rect 22848 14844 23020 14872
rect 16390 14804 16396 14816
rect 15580 14776 16396 14804
rect 16390 14764 16396 14776
rect 16448 14764 16454 14816
rect 16758 14764 16764 14816
rect 16816 14804 16822 14816
rect 16859 14807 16917 14813
rect 16859 14804 16871 14807
rect 16816 14776 16871 14804
rect 16816 14764 16822 14776
rect 16859 14773 16871 14776
rect 16905 14804 16917 14807
rect 18984 14804 19012 14832
rect 22664 14816 22692 14844
rect 23014 14832 23020 14844
rect 23072 14872 23078 14884
rect 23308 14872 23336 14912
rect 23661 14909 23673 14912
rect 23707 14940 23719 14943
rect 23768 14940 23796 14968
rect 23707 14912 23796 14940
rect 23707 14909 23719 14912
rect 23661 14903 23719 14909
rect 23842 14900 23848 14952
rect 23900 14900 23906 14952
rect 24581 14943 24639 14949
rect 24581 14940 24593 14943
rect 23952 14936 24164 14940
rect 24320 14936 24593 14940
rect 23952 14912 24593 14936
rect 23952 14872 23980 14912
rect 24136 14908 24348 14912
rect 24581 14909 24593 14912
rect 24627 14909 24639 14943
rect 25976 14940 26004 14968
rect 26053 14943 26111 14949
rect 26053 14940 26065 14943
rect 25976 14912 26065 14940
rect 24581 14903 24639 14909
rect 26053 14909 26065 14912
rect 26099 14909 26111 14943
rect 26053 14903 26111 14909
rect 23072 14844 23336 14872
rect 23400 14844 23980 14872
rect 23072 14832 23078 14844
rect 16905 14776 19012 14804
rect 16905 14773 16917 14776
rect 16859 14767 16917 14773
rect 20254 14764 20260 14816
rect 20312 14804 20318 14816
rect 20355 14807 20413 14813
rect 20355 14804 20367 14807
rect 20312 14776 20367 14804
rect 20312 14764 20318 14776
rect 20355 14773 20367 14776
rect 20401 14804 20413 14807
rect 21450 14804 21456 14816
rect 20401 14776 21456 14804
rect 20401 14773 20413 14776
rect 20355 14767 20413 14773
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 21726 14764 21732 14816
rect 21784 14764 21790 14816
rect 22646 14764 22652 14816
rect 22704 14764 22710 14816
rect 22741 14807 22799 14813
rect 22741 14773 22753 14807
rect 22787 14804 22799 14807
rect 23400 14804 23428 14844
rect 22787 14776 23428 14804
rect 23477 14807 23535 14813
rect 22787 14773 22799 14776
rect 22741 14767 22799 14773
rect 23477 14773 23489 14807
rect 23523 14804 23535 14807
rect 24210 14804 24216 14816
rect 23523 14776 24216 14804
rect 23523 14773 23535 14776
rect 23477 14767 23535 14773
rect 24210 14764 24216 14776
rect 24268 14764 24274 14816
rect 25682 14764 25688 14816
rect 25740 14764 25746 14816
rect 26050 14764 26056 14816
rect 26108 14804 26114 14816
rect 26160 14804 26188 14980
rect 26516 14977 26528 14980
rect 26562 14977 26574 15011
rect 26516 14971 26574 14977
rect 26602 14968 26608 15020
rect 26660 15008 26666 15020
rect 28166 15008 28172 15020
rect 26660 14980 28172 15008
rect 26660 14968 26666 14980
rect 28166 14968 28172 14980
rect 28224 14968 28230 15020
rect 26789 14943 26847 14949
rect 26789 14909 26801 14943
rect 26835 14940 26847 14943
rect 28276 14940 28304 15116
rect 30098 15104 30104 15116
rect 30156 15104 30162 15156
rect 29733 15079 29791 15085
rect 29733 15076 29745 15079
rect 26835 14912 28304 14940
rect 28368 15048 29745 15076
rect 26835 14909 26847 14912
rect 26789 14903 26847 14909
rect 27982 14832 27988 14884
rect 28040 14872 28046 14884
rect 28368 14881 28396 15048
rect 29733 15045 29745 15048
rect 29779 15045 29791 15079
rect 29733 15039 29791 15045
rect 28534 14968 28540 15020
rect 28592 15008 28598 15020
rect 29365 15011 29423 15017
rect 29365 15008 29377 15011
rect 28592 14980 29377 15008
rect 28592 14968 28598 14980
rect 29365 14977 29377 14980
rect 29411 14977 29423 15011
rect 29365 14971 29423 14977
rect 28353 14875 28411 14881
rect 28353 14872 28365 14875
rect 28040 14844 28365 14872
rect 28040 14832 28046 14844
rect 28353 14841 28365 14844
rect 28399 14841 28411 14875
rect 28353 14835 28411 14841
rect 26108 14776 26188 14804
rect 26519 14807 26577 14813
rect 26108 14764 26114 14776
rect 26519 14773 26531 14807
rect 26565 14804 26577 14807
rect 26694 14804 26700 14816
rect 26565 14776 26700 14804
rect 26565 14773 26577 14776
rect 26519 14767 26577 14773
rect 26694 14764 26700 14776
rect 26752 14764 26758 14816
rect 26786 14764 26792 14816
rect 26844 14804 26850 14816
rect 27522 14804 27528 14816
rect 26844 14776 27528 14804
rect 26844 14764 26850 14776
rect 27522 14764 27528 14776
rect 27580 14804 27586 14816
rect 28552 14804 28580 14968
rect 28718 14900 28724 14952
rect 28776 14940 28782 14952
rect 28776 14912 29500 14940
rect 28776 14900 28782 14912
rect 28810 14832 28816 14884
rect 28868 14872 28874 14884
rect 29089 14875 29147 14881
rect 29089 14872 29101 14875
rect 28868 14844 29101 14872
rect 28868 14832 28874 14844
rect 29089 14841 29101 14844
rect 29135 14841 29147 14875
rect 29472 14872 29500 14912
rect 29546 14900 29552 14952
rect 29604 14900 29610 14952
rect 29730 14872 29736 14884
rect 29472 14844 29736 14872
rect 29089 14835 29147 14841
rect 29730 14832 29736 14844
rect 29788 14832 29794 14884
rect 30193 14875 30251 14881
rect 30193 14841 30205 14875
rect 30239 14841 30251 14875
rect 30193 14835 30251 14841
rect 27580 14776 28580 14804
rect 27580 14764 27586 14776
rect 29270 14764 29276 14816
rect 29328 14804 29334 14816
rect 30208 14804 30236 14835
rect 29328 14776 30236 14804
rect 30469 14807 30527 14813
rect 29328 14764 29334 14776
rect 30469 14773 30481 14807
rect 30515 14804 30527 14807
rect 31110 14804 31116 14816
rect 30515 14776 31116 14804
rect 30515 14773 30527 14776
rect 30469 14767 30527 14773
rect 31110 14764 31116 14776
rect 31168 14764 31174 14816
rect 552 14714 31072 14736
rect 552 14662 7988 14714
rect 8040 14662 8052 14714
rect 8104 14662 8116 14714
rect 8168 14662 8180 14714
rect 8232 14662 8244 14714
rect 8296 14662 15578 14714
rect 15630 14662 15642 14714
rect 15694 14662 15706 14714
rect 15758 14662 15770 14714
rect 15822 14662 15834 14714
rect 15886 14662 23168 14714
rect 23220 14662 23232 14714
rect 23284 14662 23296 14714
rect 23348 14662 23360 14714
rect 23412 14662 23424 14714
rect 23476 14662 30758 14714
rect 30810 14662 30822 14714
rect 30874 14662 30886 14714
rect 30938 14662 30950 14714
rect 31002 14662 31014 14714
rect 31066 14662 31072 14714
rect 552 14640 31072 14662
rect 2498 14600 2504 14612
rect 1412 14572 2504 14600
rect 1412 14473 1440 14572
rect 2498 14560 2504 14572
rect 2556 14560 2562 14612
rect 2590 14560 2596 14612
rect 2648 14600 2654 14612
rect 2648 14572 3280 14600
rect 2648 14560 2654 14572
rect 3050 14492 3056 14544
rect 3108 14492 3114 14544
rect 3252 14532 3280 14572
rect 3418 14560 3424 14612
rect 3476 14600 3482 14612
rect 3973 14603 4031 14609
rect 3973 14600 3985 14603
rect 3476 14572 3985 14600
rect 3476 14560 3482 14572
rect 3973 14569 3985 14572
rect 4019 14569 4031 14603
rect 3973 14563 4031 14569
rect 4430 14560 4436 14612
rect 4488 14560 4494 14612
rect 4522 14560 4528 14612
rect 4580 14600 4586 14612
rect 4709 14603 4767 14609
rect 4709 14600 4721 14603
rect 4580 14572 4721 14600
rect 4580 14560 4586 14572
rect 4709 14569 4721 14572
rect 4755 14569 4767 14603
rect 4709 14563 4767 14569
rect 4982 14560 4988 14612
rect 5040 14560 5046 14612
rect 5442 14560 5448 14612
rect 5500 14560 5506 14612
rect 6089 14603 6147 14609
rect 6089 14569 6101 14603
rect 6135 14600 6147 14603
rect 6135 14572 6319 14600
rect 6135 14569 6147 14572
rect 6089 14563 6147 14569
rect 6291 14532 6319 14572
rect 6362 14560 6368 14612
rect 6420 14560 6426 14612
rect 7098 14600 7104 14612
rect 6610 14572 7104 14600
rect 6610 14532 6638 14572
rect 7098 14560 7104 14572
rect 7156 14560 7162 14612
rect 7282 14560 7288 14612
rect 7340 14600 7346 14612
rect 7340 14572 8892 14600
rect 7340 14560 7346 14572
rect 3252 14504 4752 14532
rect 1121 14467 1179 14473
rect 1121 14433 1133 14467
rect 1167 14464 1179 14467
rect 1397 14467 1455 14473
rect 1397 14464 1409 14467
rect 1167 14436 1409 14464
rect 1167 14433 1179 14436
rect 1121 14427 1179 14433
rect 1397 14433 1409 14436
rect 1443 14433 1455 14467
rect 1397 14427 1455 14433
rect 1486 14424 1492 14476
rect 1544 14424 1550 14476
rect 2590 14464 2596 14476
rect 1596 14436 2596 14464
rect 1596 14396 1624 14436
rect 2590 14424 2596 14436
rect 2648 14424 2654 14476
rect 3068 14464 3096 14492
rect 4724 14476 4752 14504
rect 4908 14504 6132 14532
rect 6291 14504 6638 14532
rect 3881 14467 3939 14473
rect 3881 14464 3893 14467
rect 3068 14436 3893 14464
rect 3881 14433 3893 14436
rect 3927 14433 3939 14467
rect 3881 14427 3939 14433
rect 4157 14467 4215 14473
rect 4157 14433 4169 14467
rect 4203 14464 4215 14467
rect 4430 14464 4436 14476
rect 4203 14436 4436 14464
rect 4203 14433 4215 14436
rect 4157 14427 4215 14433
rect 952 14368 1624 14396
rect 952 14337 980 14368
rect 1670 14356 1676 14408
rect 1728 14396 1734 14408
rect 2038 14407 2044 14408
rect 1816 14399 1874 14405
rect 1816 14396 1828 14399
rect 1728 14368 1828 14396
rect 1728 14356 1734 14368
rect 1816 14365 1828 14368
rect 1862 14365 1874 14399
rect 1816 14359 1874 14365
rect 1995 14401 2044 14407
rect 1995 14367 2007 14401
rect 2041 14367 2044 14401
rect 1995 14361 2044 14367
rect 2038 14356 2044 14361
rect 2096 14356 2102 14408
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 3142 14396 3148 14408
rect 2271 14368 3148 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 3142 14356 3148 14368
rect 3200 14356 3206 14408
rect 3605 14399 3663 14405
rect 3605 14365 3617 14399
rect 3651 14396 3663 14399
rect 3786 14396 3792 14408
rect 3651 14368 3792 14396
rect 3651 14365 3663 14368
rect 3605 14359 3663 14365
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 3896 14396 3924 14427
rect 4430 14424 4436 14436
rect 4488 14424 4494 14476
rect 4614 14424 4620 14476
rect 4672 14424 4678 14476
rect 4706 14424 4712 14476
rect 4764 14424 4770 14476
rect 4908 14473 4936 14504
rect 4893 14467 4951 14473
rect 4893 14433 4905 14467
rect 4939 14433 4951 14467
rect 4893 14427 4951 14433
rect 4982 14424 4988 14476
rect 5040 14464 5046 14476
rect 5169 14467 5227 14473
rect 5169 14464 5181 14467
rect 5040 14436 5181 14464
rect 5040 14424 5046 14436
rect 5169 14433 5181 14436
rect 5215 14464 5227 14467
rect 5629 14467 5687 14473
rect 5629 14464 5641 14467
rect 5215 14436 5641 14464
rect 5215 14433 5227 14436
rect 5169 14427 5227 14433
rect 5629 14433 5641 14436
rect 5675 14433 5687 14467
rect 5629 14427 5687 14433
rect 5350 14396 5356 14408
rect 3896 14368 5356 14396
rect 5350 14356 5356 14368
rect 5408 14356 5414 14408
rect 5644 14396 5672 14427
rect 5902 14424 5908 14476
rect 5960 14464 5966 14476
rect 5997 14467 6055 14473
rect 5997 14464 6009 14467
rect 5960 14436 6009 14464
rect 5960 14424 5966 14436
rect 5997 14433 6009 14436
rect 6043 14433 6055 14467
rect 6104 14464 6132 14504
rect 6270 14464 6276 14476
rect 6104 14436 6276 14464
rect 5997 14427 6055 14433
rect 6270 14424 6276 14436
rect 6328 14424 6334 14476
rect 6362 14424 6368 14476
rect 6420 14464 6426 14476
rect 6549 14467 6607 14473
rect 6549 14464 6561 14467
rect 6420 14436 6561 14464
rect 6420 14424 6426 14436
rect 6549 14433 6561 14436
rect 6595 14433 6607 14467
rect 6549 14427 6607 14433
rect 6638 14424 6644 14476
rect 6696 14424 6702 14476
rect 8864 14473 8892 14572
rect 8938 14560 8944 14612
rect 8996 14560 9002 14612
rect 9030 14560 9036 14612
rect 9088 14560 9094 14612
rect 9306 14560 9312 14612
rect 9364 14600 9370 14612
rect 9401 14603 9459 14609
rect 9401 14600 9413 14603
rect 9364 14572 9413 14600
rect 9364 14560 9370 14572
rect 9401 14569 9413 14572
rect 9447 14569 9459 14603
rect 9401 14563 9459 14569
rect 9674 14560 9680 14612
rect 9732 14560 9738 14612
rect 9950 14560 9956 14612
rect 10008 14560 10014 14612
rect 10042 14560 10048 14612
rect 10100 14560 10106 14612
rect 10321 14603 10379 14609
rect 10321 14569 10333 14603
rect 10367 14600 10379 14603
rect 11974 14600 11980 14612
rect 10367 14572 11980 14600
rect 10367 14569 10379 14572
rect 10321 14563 10379 14569
rect 11974 14560 11980 14572
rect 12032 14560 12038 14612
rect 13446 14560 13452 14612
rect 13504 14560 13510 14612
rect 14283 14603 14341 14609
rect 14283 14569 14295 14603
rect 14329 14600 14341 14603
rect 14826 14600 14832 14612
rect 14329 14572 14832 14600
rect 14329 14569 14341 14572
rect 14283 14563 14341 14569
rect 14826 14560 14832 14572
rect 14884 14560 14890 14612
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 16853 14603 16911 14609
rect 16853 14600 16865 14603
rect 14976 14572 16865 14600
rect 14976 14560 14982 14572
rect 16853 14569 16865 14572
rect 16899 14569 16911 14603
rect 16853 14563 16911 14569
rect 18322 14560 18328 14612
rect 18380 14600 18386 14612
rect 20073 14603 20131 14609
rect 20073 14600 20085 14603
rect 18380 14572 20085 14600
rect 18380 14560 18386 14572
rect 20073 14569 20085 14572
rect 20119 14569 20131 14603
rect 20073 14563 20131 14569
rect 20257 14603 20315 14609
rect 20257 14569 20269 14603
rect 20303 14600 20315 14603
rect 20622 14600 20628 14612
rect 20303 14572 20628 14600
rect 20303 14569 20315 14572
rect 20257 14563 20315 14569
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 21726 14600 21732 14612
rect 20824 14572 21732 14600
rect 8849 14467 8907 14473
rect 6748 14436 8432 14464
rect 6748 14396 6776 14436
rect 7006 14405 7012 14408
rect 5644 14368 6776 14396
rect 6968 14399 7012 14405
rect 6968 14365 6980 14399
rect 6968 14359 7012 14365
rect 7006 14356 7012 14359
rect 7064 14356 7070 14408
rect 7147 14399 7205 14405
rect 7147 14365 7159 14399
rect 7193 14396 7205 14399
rect 7282 14396 7288 14408
rect 7193 14368 7288 14396
rect 7193 14365 7205 14368
rect 7147 14359 7205 14365
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 7374 14356 7380 14408
rect 7432 14356 7438 14408
rect 7558 14356 7564 14408
rect 7616 14396 7622 14408
rect 7616 14368 8340 14396
rect 7616 14356 7622 14368
rect 937 14331 995 14337
rect 937 14297 949 14331
rect 983 14297 995 14331
rect 4706 14328 4712 14340
rect 937 14291 995 14297
rect 3436 14300 4712 14328
rect 1213 14263 1271 14269
rect 1213 14229 1225 14263
rect 1259 14260 1271 14263
rect 3436 14260 3464 14300
rect 4706 14288 4712 14300
rect 4764 14288 4770 14340
rect 5718 14288 5724 14340
rect 5776 14328 5782 14340
rect 6362 14328 6368 14340
rect 5776 14300 6368 14328
rect 5776 14288 5782 14300
rect 6362 14288 6368 14300
rect 6420 14288 6426 14340
rect 1259 14232 3464 14260
rect 3697 14263 3755 14269
rect 1259 14229 1271 14232
rect 1213 14223 1271 14229
rect 3697 14229 3709 14263
rect 3743 14260 3755 14263
rect 4798 14260 4804 14272
rect 3743 14232 4804 14260
rect 3743 14229 3755 14232
rect 3697 14223 3755 14229
rect 4798 14220 4804 14232
rect 4856 14220 4862 14272
rect 5810 14220 5816 14272
rect 5868 14220 5874 14272
rect 5994 14220 6000 14272
rect 6052 14260 6058 14272
rect 6638 14260 6644 14272
rect 6052 14232 6644 14260
rect 6052 14220 6058 14232
rect 6638 14220 6644 14232
rect 6696 14220 6702 14272
rect 8312 14260 8340 14368
rect 8404 14340 8432 14436
rect 8849 14433 8861 14467
rect 8895 14433 8907 14467
rect 8956 14464 8984 14560
rect 9048 14532 9076 14560
rect 10060 14532 10088 14560
rect 10962 14532 10968 14544
rect 9048 14504 9628 14532
rect 9324 14476 9352 14504
rect 9125 14467 9183 14473
rect 9125 14464 9137 14467
rect 8956 14436 9137 14464
rect 8849 14427 8907 14433
rect 9125 14433 9137 14436
rect 9171 14433 9183 14467
rect 9125 14427 9183 14433
rect 8864 14396 8892 14427
rect 9306 14424 9312 14476
rect 9364 14424 9370 14476
rect 9600 14473 9628 14504
rect 10060 14504 10968 14532
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14433 9643 14467
rect 9585 14427 9643 14433
rect 9861 14467 9919 14473
rect 9861 14433 9873 14467
rect 9907 14464 9919 14467
rect 9950 14464 9956 14476
rect 9907 14436 9956 14464
rect 9907 14433 9919 14436
rect 9861 14427 9919 14433
rect 9950 14424 9956 14436
rect 10008 14464 10014 14476
rect 10060 14464 10088 14504
rect 10962 14492 10968 14504
rect 11020 14492 11026 14544
rect 11333 14535 11391 14541
rect 11333 14501 11345 14535
rect 11379 14532 11391 14535
rect 11514 14532 11520 14544
rect 11379 14504 11520 14532
rect 11379 14501 11391 14504
rect 11333 14495 11391 14501
rect 11514 14492 11520 14504
rect 11572 14532 11578 14544
rect 11572 14504 11744 14532
rect 11572 14492 11578 14504
rect 10008 14436 10088 14464
rect 10137 14467 10195 14473
rect 10008 14424 10014 14436
rect 10137 14433 10149 14467
rect 10183 14464 10195 14467
rect 10226 14464 10232 14476
rect 10183 14436 10232 14464
rect 10183 14433 10195 14436
rect 10137 14427 10195 14433
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 10318 14424 10324 14476
rect 10376 14464 10382 14476
rect 10505 14467 10563 14473
rect 10505 14464 10517 14467
rect 10376 14436 10517 14464
rect 10376 14424 10382 14436
rect 10505 14433 10517 14436
rect 10551 14433 10563 14467
rect 10505 14427 10563 14433
rect 10778 14424 10784 14476
rect 10836 14424 10842 14476
rect 11057 14467 11115 14473
rect 11057 14433 11069 14467
rect 11103 14433 11115 14467
rect 11057 14427 11115 14433
rect 11072 14396 11100 14427
rect 11238 14424 11244 14476
rect 11296 14464 11302 14476
rect 11609 14467 11667 14473
rect 11609 14464 11621 14467
rect 11296 14436 11621 14464
rect 11296 14424 11302 14436
rect 11609 14433 11621 14436
rect 11655 14433 11667 14467
rect 11716 14464 11744 14504
rect 19536 14504 20484 14532
rect 11936 14467 11994 14473
rect 11936 14464 11948 14467
rect 11716 14436 11948 14464
rect 11609 14427 11667 14433
rect 11936 14433 11948 14436
rect 11982 14433 11994 14467
rect 15933 14467 15991 14473
rect 15933 14464 15945 14467
rect 11936 14427 11994 14433
rect 12120 14436 15945 14464
rect 11790 14396 11796 14408
rect 8864 14368 11796 14396
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 12120 14407 12148 14436
rect 15933 14433 15945 14436
rect 15979 14433 15991 14467
rect 16209 14467 16267 14473
rect 16209 14464 16221 14467
rect 15933 14427 15991 14433
rect 16040 14436 16221 14464
rect 12105 14401 12163 14407
rect 12105 14367 12117 14401
rect 12151 14367 12163 14401
rect 12105 14361 12163 14367
rect 12250 14356 12256 14408
rect 12308 14405 12314 14408
rect 12308 14399 12357 14405
rect 12308 14365 12311 14399
rect 12345 14365 12357 14399
rect 12308 14359 12357 14365
rect 12308 14356 12314 14359
rect 13814 14356 13820 14408
rect 13872 14356 13878 14408
rect 14323 14399 14381 14405
rect 14323 14365 14335 14399
rect 14369 14396 14381 14399
rect 14458 14396 14464 14408
rect 14369 14368 14464 14396
rect 14369 14365 14381 14368
rect 14323 14359 14381 14365
rect 14458 14356 14464 14368
rect 14516 14356 14522 14408
rect 14550 14356 14556 14408
rect 14608 14356 14614 14408
rect 14642 14356 14648 14408
rect 14700 14396 14706 14408
rect 15378 14396 15384 14408
rect 14700 14368 15384 14396
rect 14700 14356 14706 14368
rect 15378 14356 15384 14368
rect 15436 14356 15442 14408
rect 8386 14288 8392 14340
rect 8444 14288 8450 14340
rect 10134 14328 10140 14340
rect 8496 14300 10140 14328
rect 8496 14260 8524 14300
rect 10134 14288 10140 14300
rect 10192 14288 10198 14340
rect 10870 14288 10876 14340
rect 10928 14288 10934 14340
rect 8312 14232 8524 14260
rect 8665 14263 8723 14269
rect 8665 14229 8677 14263
rect 8711 14260 8723 14263
rect 10042 14260 10048 14272
rect 8711 14232 10048 14260
rect 8711 14229 8723 14232
rect 8665 14223 8723 14229
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 10226 14220 10232 14272
rect 10284 14260 10290 14272
rect 10410 14260 10416 14272
rect 10284 14232 10416 14260
rect 10284 14220 10290 14232
rect 10410 14220 10416 14232
rect 10468 14220 10474 14272
rect 10594 14220 10600 14272
rect 10652 14220 10658 14272
rect 10888 14260 10916 14288
rect 12710 14260 12716 14272
rect 10888 14232 12716 14260
rect 12710 14220 12716 14232
rect 12768 14220 12774 14272
rect 13832 14260 13860 14356
rect 14182 14260 14188 14272
rect 13832 14232 14188 14260
rect 14182 14220 14188 14232
rect 14240 14260 14246 14272
rect 16040 14260 16068 14436
rect 16209 14433 16221 14436
rect 16255 14433 16267 14467
rect 16209 14427 16267 14433
rect 16666 14424 16672 14476
rect 16724 14424 16730 14476
rect 16758 14424 16764 14476
rect 16816 14464 16822 14476
rect 19536 14473 19564 14504
rect 17456 14467 17514 14473
rect 17456 14464 17468 14467
rect 16816 14436 17468 14464
rect 16816 14424 16822 14436
rect 17456 14433 17468 14436
rect 17502 14433 17514 14467
rect 19521 14467 19579 14473
rect 17456 14427 17514 14433
rect 17788 14436 19472 14464
rect 17129 14399 17187 14405
rect 17129 14396 17141 14399
rect 16592 14368 17141 14396
rect 16592 14272 16620 14368
rect 17129 14365 17141 14368
rect 17175 14365 17187 14399
rect 17129 14359 17187 14365
rect 17635 14399 17693 14405
rect 17635 14365 17647 14399
rect 17681 14396 17693 14399
rect 17788 14396 17816 14436
rect 17681 14368 17816 14396
rect 17865 14399 17923 14405
rect 17681 14365 17693 14368
rect 17635 14359 17693 14365
rect 17865 14365 17877 14399
rect 17911 14396 17923 14399
rect 19444 14396 19472 14436
rect 19521 14433 19533 14467
rect 19567 14433 19579 14467
rect 19521 14427 19579 14433
rect 19797 14467 19855 14473
rect 19797 14433 19809 14467
rect 19843 14464 19855 14467
rect 20162 14464 20168 14476
rect 19843 14436 20168 14464
rect 19843 14433 19855 14436
rect 19797 14427 19855 14433
rect 20162 14424 20168 14436
rect 20220 14424 20226 14476
rect 20456 14473 20484 14504
rect 20441 14467 20499 14473
rect 20441 14433 20453 14467
rect 20487 14464 20499 14467
rect 20530 14464 20536 14476
rect 20487 14436 20536 14464
rect 20487 14433 20499 14436
rect 20441 14427 20499 14433
rect 20530 14424 20536 14436
rect 20588 14424 20594 14476
rect 20714 14464 20720 14476
rect 20772 14473 20778 14476
rect 20683 14436 20720 14464
rect 20714 14424 20720 14436
rect 20772 14427 20783 14473
rect 20772 14424 20778 14427
rect 20824 14396 20852 14572
rect 21726 14560 21732 14572
rect 21784 14560 21790 14612
rect 22646 14560 22652 14612
rect 22704 14600 22710 14612
rect 23658 14600 23664 14612
rect 22704 14572 23664 14600
rect 22704 14560 22710 14572
rect 23658 14560 23664 14572
rect 23716 14560 23722 14612
rect 23753 14603 23811 14609
rect 23753 14569 23765 14603
rect 23799 14569 23811 14603
rect 23753 14563 23811 14569
rect 23768 14532 23796 14563
rect 23842 14560 23848 14612
rect 23900 14600 23906 14612
rect 24026 14600 24032 14612
rect 23900 14572 24032 14600
rect 23900 14560 23906 14572
rect 24026 14560 24032 14572
rect 24084 14560 24090 14612
rect 24394 14560 24400 14612
rect 24452 14600 24458 14612
rect 24495 14603 24553 14609
rect 24495 14600 24507 14603
rect 24452 14572 24507 14600
rect 24452 14560 24458 14572
rect 24495 14569 24507 14572
rect 24541 14600 24553 14603
rect 24541 14572 25452 14600
rect 24541 14569 24553 14572
rect 24495 14563 24553 14569
rect 25424 14532 25452 14572
rect 26050 14560 26056 14612
rect 26108 14560 26114 14612
rect 27338 14600 27344 14612
rect 26896 14572 27344 14600
rect 26786 14532 26792 14544
rect 17911 14368 19380 14396
rect 19444 14368 20852 14396
rect 21008 14504 21312 14532
rect 23768 14504 24164 14532
rect 25424 14504 26792 14532
rect 17911 14365 17923 14368
rect 17865 14359 17923 14365
rect 18966 14288 18972 14340
rect 19024 14288 19030 14340
rect 19352 14337 19380 14368
rect 19337 14331 19395 14337
rect 19337 14297 19349 14331
rect 19383 14297 19395 14331
rect 20533 14331 20591 14337
rect 19337 14291 19395 14297
rect 19444 14300 19932 14328
rect 14240 14232 16068 14260
rect 16485 14263 16543 14269
rect 14240 14220 14246 14232
rect 16485 14229 16497 14263
rect 16531 14260 16543 14263
rect 16574 14260 16580 14272
rect 16531 14232 16580 14260
rect 16531 14229 16543 14232
rect 16485 14223 16543 14229
rect 16574 14220 16580 14232
rect 16632 14220 16638 14272
rect 18690 14220 18696 14272
rect 18748 14260 18754 14272
rect 19444 14260 19472 14300
rect 18748 14232 19472 14260
rect 19613 14263 19671 14269
rect 18748 14220 18754 14232
rect 19613 14229 19625 14263
rect 19659 14260 19671 14263
rect 19794 14260 19800 14272
rect 19659 14232 19800 14260
rect 19659 14229 19671 14232
rect 19613 14223 19671 14229
rect 19794 14220 19800 14232
rect 19852 14220 19858 14272
rect 19904 14260 19932 14300
rect 20533 14297 20545 14331
rect 20579 14328 20591 14331
rect 21008 14328 21036 14504
rect 21085 14467 21143 14473
rect 21085 14433 21097 14467
rect 21131 14433 21143 14467
rect 21284 14464 21312 14504
rect 22005 14467 22063 14473
rect 22005 14464 22017 14467
rect 21284 14436 22017 14464
rect 21085 14427 21143 14433
rect 22005 14433 22017 14436
rect 22051 14433 22063 14467
rect 22005 14427 22063 14433
rect 20579 14300 21036 14328
rect 20579 14297 20591 14300
rect 20533 14291 20591 14297
rect 20806 14260 20812 14272
rect 19904 14232 20812 14260
rect 20806 14220 20812 14232
rect 20864 14220 20870 14272
rect 20901 14263 20959 14269
rect 20901 14229 20913 14263
rect 20947 14260 20959 14263
rect 20990 14260 20996 14272
rect 20947 14232 20996 14260
rect 20947 14229 20959 14232
rect 20901 14223 20959 14229
rect 20990 14220 20996 14232
rect 21048 14220 21054 14272
rect 21100 14260 21128 14427
rect 22094 14424 22100 14476
rect 22152 14464 22158 14476
rect 22830 14464 22836 14476
rect 22152 14436 22836 14464
rect 22152 14424 22158 14436
rect 22830 14424 22836 14436
rect 22888 14464 22894 14476
rect 23658 14464 23664 14476
rect 22888 14436 23664 14464
rect 22888 14424 22894 14436
rect 23658 14424 23664 14436
rect 23716 14424 23722 14476
rect 23750 14424 23756 14476
rect 23808 14464 23814 14476
rect 23937 14467 23995 14473
rect 23937 14464 23949 14467
rect 23808 14436 23949 14464
rect 23808 14424 23814 14436
rect 23937 14433 23949 14436
rect 23983 14433 23995 14467
rect 24136 14464 24164 14504
rect 26786 14492 26792 14504
rect 26844 14532 26850 14544
rect 26896 14541 26924 14572
rect 27338 14560 27344 14572
rect 27396 14560 27402 14612
rect 28543 14603 28601 14609
rect 28543 14569 28555 14603
rect 28589 14600 28601 14603
rect 28718 14600 28724 14612
rect 28589 14572 28724 14600
rect 28589 14569 28601 14572
rect 28543 14563 28601 14569
rect 28718 14560 28724 14572
rect 28776 14560 28782 14612
rect 29914 14560 29920 14612
rect 29972 14560 29978 14612
rect 26881 14535 26939 14541
rect 26881 14532 26893 14535
rect 26844 14504 26893 14532
rect 26844 14492 26850 14504
rect 26881 14501 26893 14504
rect 26927 14501 26939 14535
rect 26881 14495 26939 14501
rect 27522 14492 27528 14544
rect 27580 14492 27586 14544
rect 27724 14504 28212 14532
rect 24765 14467 24823 14473
rect 24765 14464 24777 14467
rect 24136 14436 24777 14464
rect 23937 14427 23995 14433
rect 24765 14433 24777 14436
rect 24811 14433 24823 14467
rect 24765 14427 24823 14433
rect 24854 14424 24860 14476
rect 24912 14464 24918 14476
rect 26418 14464 26424 14476
rect 24912 14436 26424 14464
rect 24912 14424 24918 14436
rect 26418 14424 26424 14436
rect 26476 14464 26482 14476
rect 26605 14467 26663 14473
rect 26605 14464 26617 14467
rect 26476 14436 26617 14464
rect 26476 14424 26482 14436
rect 26605 14433 26617 14436
rect 26651 14433 26663 14467
rect 26605 14427 26663 14433
rect 27062 14424 27068 14476
rect 27120 14464 27126 14476
rect 27341 14467 27399 14473
rect 27341 14464 27353 14467
rect 27120 14436 27353 14464
rect 27120 14424 27126 14436
rect 27341 14433 27353 14436
rect 27387 14464 27399 14467
rect 27724 14464 27752 14504
rect 27387 14436 27752 14464
rect 28077 14467 28135 14473
rect 27387 14433 27399 14436
rect 27341 14427 27399 14433
rect 28077 14433 28089 14467
rect 28123 14433 28135 14467
rect 28184 14464 28212 14504
rect 28184 14436 28994 14464
rect 28077 14427 28135 14433
rect 21266 14356 21272 14408
rect 21324 14356 21330 14408
rect 21450 14356 21456 14408
rect 21508 14396 21514 14408
rect 21596 14399 21654 14405
rect 21596 14396 21608 14399
rect 21508 14368 21608 14396
rect 21508 14356 21514 14368
rect 21596 14365 21608 14368
rect 21642 14365 21654 14399
rect 21596 14359 21654 14365
rect 21775 14399 21833 14405
rect 21775 14365 21787 14399
rect 21821 14396 21833 14399
rect 22922 14396 22928 14408
rect 21821 14368 22928 14396
rect 21821 14365 21833 14368
rect 21775 14359 21833 14365
rect 22922 14356 22928 14368
rect 22980 14356 22986 14408
rect 24026 14356 24032 14408
rect 24084 14356 24090 14408
rect 24486 14356 24492 14408
rect 24544 14396 24550 14408
rect 24544 14368 24589 14396
rect 24544 14356 24550 14368
rect 23934 14328 23940 14340
rect 23124 14300 23940 14328
rect 23124 14260 23152 14300
rect 23934 14288 23940 14300
rect 23992 14288 23998 14340
rect 27801 14331 27859 14337
rect 27801 14328 27813 14331
rect 26528 14300 27813 14328
rect 26528 14272 26556 14300
rect 27801 14297 27813 14300
rect 27847 14328 27859 14331
rect 28092 14328 28120 14427
rect 28583 14399 28641 14405
rect 28583 14365 28595 14399
rect 28629 14396 28641 14399
rect 28718 14396 28724 14408
rect 28629 14368 28724 14396
rect 28629 14365 28641 14368
rect 28583 14359 28641 14365
rect 28718 14356 28724 14368
rect 28776 14356 28782 14408
rect 28810 14356 28816 14408
rect 28868 14356 28874 14408
rect 28966 14396 28994 14436
rect 29914 14424 29920 14476
rect 29972 14464 29978 14476
rect 30285 14467 30343 14473
rect 30285 14464 30297 14467
rect 29972 14436 30297 14464
rect 29972 14424 29978 14436
rect 30285 14433 30297 14436
rect 30331 14464 30343 14467
rect 30558 14464 30564 14476
rect 30331 14436 30564 14464
rect 30331 14433 30343 14436
rect 30285 14427 30343 14433
rect 30558 14424 30564 14436
rect 30616 14424 30622 14476
rect 31110 14424 31116 14476
rect 31168 14424 31174 14476
rect 31128 14396 31156 14424
rect 28966 14368 31156 14396
rect 27847 14300 28120 14328
rect 27847 14297 27859 14300
rect 27801 14291 27859 14297
rect 29914 14288 29920 14340
rect 29972 14328 29978 14340
rect 29972 14300 30604 14328
rect 29972 14288 29978 14300
rect 30576 14272 30604 14300
rect 21100 14232 23152 14260
rect 23290 14220 23296 14272
rect 23348 14220 23354 14272
rect 23477 14263 23535 14269
rect 23477 14229 23489 14263
rect 23523 14260 23535 14263
rect 24670 14260 24676 14272
rect 23523 14232 24676 14260
rect 23523 14229 23535 14232
rect 23477 14223 23535 14229
rect 24670 14220 24676 14232
rect 24728 14220 24734 14272
rect 26510 14220 26516 14272
rect 26568 14220 26574 14272
rect 27157 14263 27215 14269
rect 27157 14229 27169 14263
rect 27203 14260 27215 14263
rect 27338 14260 27344 14272
rect 27203 14232 27344 14260
rect 27203 14229 27215 14232
rect 27157 14223 27215 14229
rect 27338 14220 27344 14232
rect 27396 14220 27402 14272
rect 27706 14220 27712 14272
rect 27764 14260 27770 14272
rect 30469 14263 30527 14269
rect 30469 14260 30481 14263
rect 27764 14232 30481 14260
rect 27764 14220 27770 14232
rect 30469 14229 30481 14232
rect 30515 14229 30527 14263
rect 30469 14223 30527 14229
rect 30558 14220 30564 14272
rect 30616 14220 30622 14272
rect 552 14170 30912 14192
rect 552 14118 4193 14170
rect 4245 14118 4257 14170
rect 4309 14118 4321 14170
rect 4373 14118 4385 14170
rect 4437 14118 4449 14170
rect 4501 14118 11783 14170
rect 11835 14118 11847 14170
rect 11899 14118 11911 14170
rect 11963 14118 11975 14170
rect 12027 14118 12039 14170
rect 12091 14118 19373 14170
rect 19425 14118 19437 14170
rect 19489 14118 19501 14170
rect 19553 14118 19565 14170
rect 19617 14118 19629 14170
rect 19681 14118 26963 14170
rect 27015 14118 27027 14170
rect 27079 14118 27091 14170
rect 27143 14118 27155 14170
rect 27207 14118 27219 14170
rect 27271 14118 30912 14170
rect 552 14096 30912 14118
rect 1118 14016 1124 14068
rect 1176 14056 1182 14068
rect 4982 14056 4988 14068
rect 1176 14028 4988 14056
rect 1176 14016 1182 14028
rect 934 13880 940 13932
rect 992 13880 998 13932
rect 1302 13929 1308 13932
rect 1264 13923 1308 13929
rect 1264 13889 1276 13923
rect 1264 13883 1308 13889
rect 1302 13880 1308 13883
rect 1360 13880 1366 13932
rect 2314 13920 2320 13932
rect 1418 13905 2320 13920
rect 1418 13874 1445 13905
rect 1433 13871 1445 13874
rect 1479 13892 2320 13905
rect 1479 13871 1491 13892
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 1433 13865 1491 13871
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 2590 13852 2596 13864
rect 1719 13824 2596 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 3050 13812 3056 13864
rect 3108 13812 3114 13864
rect 3712 13861 3740 14028
rect 4982 14016 4988 14028
rect 5040 14016 5046 14068
rect 5810 14016 5816 14068
rect 5868 14016 5874 14068
rect 7190 14016 7196 14068
rect 7248 14056 7254 14068
rect 7929 14059 7987 14065
rect 7929 14056 7941 14059
rect 7248 14028 7941 14056
rect 7248 14016 7254 14028
rect 7929 14025 7941 14028
rect 7975 14025 7987 14059
rect 9766 14056 9772 14068
rect 7929 14019 7987 14025
rect 8404 14028 9772 14056
rect 3786 13948 3792 14000
rect 3844 13948 3850 14000
rect 3804 13920 3832 13948
rect 4252 13923 4310 13929
rect 4252 13920 4264 13923
rect 3804 13892 4264 13920
rect 4252 13889 4264 13892
rect 4298 13889 4310 13923
rect 4614 13920 4620 13932
rect 4252 13883 4310 13889
rect 4448 13892 4620 13920
rect 3421 13855 3479 13861
rect 3421 13821 3433 13855
rect 3467 13852 3479 13855
rect 3697 13855 3755 13861
rect 3697 13852 3709 13855
rect 3467 13824 3709 13852
rect 3467 13821 3479 13824
rect 3421 13815 3479 13821
rect 3697 13821 3709 13824
rect 3743 13821 3755 13855
rect 3697 13815 3755 13821
rect 3786 13812 3792 13864
rect 3844 13812 3850 13864
rect 4448 13852 4476 13892
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 4706 13880 4712 13932
rect 4764 13880 4770 13932
rect 5828 13920 5856 14016
rect 6595 13923 6653 13929
rect 5828 13892 6408 13920
rect 3896 13824 4476 13852
rect 4525 13855 4583 13861
rect 3896 13784 3924 13824
rect 4525 13821 4537 13855
rect 4571 13852 4583 13855
rect 4724 13852 4752 13880
rect 4571 13824 4752 13852
rect 4571 13821 4583 13824
rect 4525 13815 4583 13821
rect 5902 13812 5908 13864
rect 5960 13812 5966 13864
rect 6086 13812 6092 13864
rect 6144 13812 6150 13864
rect 6380 13852 6408 13892
rect 6595 13889 6607 13923
rect 6641 13920 6653 13923
rect 8404 13920 8432 14028
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 10134 14016 10140 14068
rect 10192 14016 10198 14068
rect 10502 14016 10508 14068
rect 10560 14056 10566 14068
rect 13081 14059 13139 14065
rect 13081 14056 13093 14059
rect 10560 14028 13093 14056
rect 10560 14016 10566 14028
rect 13081 14025 13093 14028
rect 13127 14025 13139 14059
rect 13081 14019 13139 14025
rect 13630 14016 13636 14068
rect 13688 14016 13694 14068
rect 13832 14028 16068 14056
rect 10152 13988 10180 14016
rect 10873 13991 10931 13997
rect 10873 13988 10885 13991
rect 10152 13960 10885 13988
rect 10873 13957 10885 13960
rect 10919 13957 10931 13991
rect 10873 13951 10931 13957
rect 8852 13923 8910 13929
rect 8852 13920 8864 13923
rect 6641 13892 8432 13920
rect 8772 13892 8864 13920
rect 6641 13889 6653 13892
rect 6595 13883 6653 13889
rect 8772 13864 8800 13892
rect 8852 13889 8864 13892
rect 8898 13889 8910 13923
rect 8852 13883 8910 13889
rect 8938 13880 8944 13932
rect 8996 13920 9002 13932
rect 9306 13920 9312 13932
rect 8996 13892 9312 13920
rect 8996 13880 9002 13892
rect 9306 13880 9312 13892
rect 9364 13880 9370 13932
rect 10134 13880 10140 13932
rect 10192 13920 10198 13932
rect 10505 13923 10563 13929
rect 10505 13920 10517 13923
rect 10192 13892 10517 13920
rect 10192 13880 10198 13892
rect 10505 13889 10517 13892
rect 10551 13889 10563 13923
rect 10505 13883 10563 13889
rect 10594 13880 10600 13932
rect 10652 13920 10658 13932
rect 11606 13929 11612 13932
rect 11568 13923 11612 13929
rect 10652 13892 11376 13920
rect 10652 13880 10658 13892
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6380 13824 6837 13852
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 7558 13812 7564 13864
rect 7616 13852 7622 13864
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 7616 13824 8401 13852
rect 7616 13812 7622 13824
rect 8389 13821 8401 13824
rect 8435 13821 8447 13855
rect 8389 13815 8447 13821
rect 8754 13812 8760 13864
rect 8812 13812 8818 13864
rect 9125 13855 9183 13861
rect 9125 13821 9137 13855
rect 9171 13852 9183 13855
rect 10870 13852 10876 13864
rect 9171 13824 10876 13852
rect 9171 13821 9183 13824
rect 9125 13815 9183 13821
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 10962 13812 10968 13864
rect 11020 13852 11026 13864
rect 11057 13855 11115 13861
rect 11057 13852 11069 13855
rect 11020 13824 11069 13852
rect 11020 13812 11026 13824
rect 11057 13821 11069 13824
rect 11103 13821 11115 13855
rect 11057 13815 11115 13821
rect 11238 13812 11244 13864
rect 11296 13812 11302 13864
rect 11348 13852 11376 13892
rect 11568 13889 11580 13923
rect 11568 13883 11612 13889
rect 11606 13880 11612 13883
rect 11664 13880 11670 13932
rect 11747 13923 11805 13929
rect 11747 13889 11759 13923
rect 11793 13920 11805 13923
rect 13832 13920 13860 14028
rect 16040 13997 16068 14028
rect 16390 14016 16396 14068
rect 16448 14056 16454 14068
rect 18233 14059 18291 14065
rect 18233 14056 18245 14059
rect 16448 14028 18245 14056
rect 16448 14016 16454 14028
rect 18233 14025 18245 14028
rect 18279 14025 18291 14059
rect 23290 14056 23296 14068
rect 18233 14019 18291 14025
rect 18800 14028 23296 14056
rect 13909 13991 13967 13997
rect 13909 13957 13921 13991
rect 13955 13957 13967 13991
rect 13909 13951 13967 13957
rect 16025 13991 16083 13997
rect 16025 13957 16037 13991
rect 16071 13957 16083 13991
rect 16025 13951 16083 13957
rect 18693 13991 18751 13997
rect 18693 13957 18705 13991
rect 18739 13957 18751 13991
rect 18693 13951 18751 13957
rect 11793 13892 13860 13920
rect 13924 13920 13952 13951
rect 14691 13923 14749 13929
rect 13924 13892 14504 13920
rect 11793 13889 11805 13892
rect 11747 13883 11805 13889
rect 11977 13855 12035 13861
rect 11977 13852 11989 13855
rect 11348 13824 11989 13852
rect 11977 13821 11989 13824
rect 12023 13821 12035 13855
rect 11977 13815 12035 13821
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 14090 13812 14096 13864
rect 14148 13812 14154 13864
rect 14182 13812 14188 13864
rect 14240 13812 14246 13864
rect 14476 13852 14504 13892
rect 14691 13889 14703 13923
rect 14737 13920 14749 13923
rect 15102 13920 15108 13932
rect 14737 13892 15108 13920
rect 14737 13889 14749 13892
rect 14691 13883 14749 13889
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 16393 13923 16451 13929
rect 16393 13889 16405 13923
rect 16439 13920 16451 13923
rect 16574 13920 16580 13932
rect 16439 13892 16580 13920
rect 16439 13889 16451 13892
rect 16393 13883 16451 13889
rect 16574 13880 16580 13892
rect 16632 13880 16638 13932
rect 16758 13929 16764 13932
rect 16720 13923 16764 13929
rect 16720 13889 16732 13923
rect 16720 13883 16764 13889
rect 16758 13880 16764 13883
rect 16816 13880 16822 13932
rect 16899 13923 16957 13929
rect 16899 13889 16911 13923
rect 16945 13920 16957 13923
rect 17129 13923 17187 13929
rect 16945 13892 17080 13920
rect 16945 13889 16957 13892
rect 16899 13883 16957 13889
rect 14921 13855 14979 13861
rect 14921 13852 14933 13855
rect 14476 13824 14933 13852
rect 14921 13821 14933 13824
rect 14967 13821 14979 13855
rect 17052 13852 17080 13892
rect 17129 13889 17141 13923
rect 17175 13920 17187 13923
rect 18708 13920 18736 13951
rect 17175 13892 18736 13920
rect 17175 13889 17187 13892
rect 17129 13883 17187 13889
rect 18800 13852 18828 14028
rect 23290 14016 23296 14028
rect 23348 14016 23354 14068
rect 23569 14059 23627 14065
rect 23569 14025 23581 14059
rect 23615 14056 23627 14059
rect 23842 14056 23848 14068
rect 23615 14028 23848 14056
rect 23615 14025 23627 14028
rect 23569 14019 23627 14025
rect 23842 14016 23848 14028
rect 23900 14016 23906 14068
rect 24026 14016 24032 14068
rect 24084 14056 24090 14068
rect 24084 14028 25452 14056
rect 24084 14016 24090 14028
rect 18874 13948 18880 14000
rect 18932 13988 18938 14000
rect 18969 13991 19027 13997
rect 18969 13988 18981 13991
rect 18932 13960 18981 13988
rect 18932 13948 18938 13960
rect 18969 13957 18981 13960
rect 19015 13957 19027 13991
rect 18969 13951 19027 13957
rect 19150 13948 19156 14000
rect 19208 13948 19214 14000
rect 19794 13948 19800 14000
rect 19852 13948 19858 14000
rect 21358 13948 21364 14000
rect 21416 13988 21422 14000
rect 21637 13991 21695 13997
rect 21637 13988 21649 13991
rect 21416 13960 21649 13988
rect 21416 13948 21422 13960
rect 21637 13957 21649 13960
rect 21683 13957 21695 13991
rect 21637 13951 21695 13957
rect 21750 13960 21956 13988
rect 17052 13824 18828 13852
rect 18877 13855 18935 13861
rect 14921 13815 14979 13821
rect 18877 13821 18889 13855
rect 18923 13852 18935 13855
rect 18966 13852 18972 13864
rect 18923 13824 18972 13852
rect 18923 13821 18935 13824
rect 18877 13815 18935 13821
rect 18966 13812 18972 13824
rect 19024 13812 19030 13864
rect 19168 13861 19196 13948
rect 19426 13880 19432 13932
rect 19484 13880 19490 13932
rect 19812 13920 19840 13948
rect 20303 13923 20361 13929
rect 19812 13892 20116 13920
rect 19153 13855 19211 13861
rect 19153 13821 19165 13855
rect 19199 13821 19211 13855
rect 19153 13815 19211 13821
rect 19797 13855 19855 13861
rect 19797 13821 19809 13855
rect 19843 13852 19855 13855
rect 19886 13852 19892 13864
rect 19843 13824 19892 13852
rect 19843 13821 19855 13824
rect 19797 13815 19855 13821
rect 19886 13812 19892 13824
rect 19944 13812 19950 13864
rect 20088 13852 20116 13892
rect 20303 13889 20315 13923
rect 20349 13920 20361 13923
rect 20622 13920 20628 13932
rect 20349 13892 20628 13920
rect 20349 13889 20361 13892
rect 20303 13883 20361 13889
rect 20622 13880 20628 13892
rect 20680 13880 20686 13932
rect 21174 13880 21180 13932
rect 21232 13920 21238 13932
rect 21750 13920 21778 13960
rect 21232 13892 21778 13920
rect 21232 13880 21238 13892
rect 21818 13880 21824 13932
rect 21876 13880 21882 13932
rect 21928 13920 21956 13960
rect 22281 13923 22339 13929
rect 22281 13920 22293 13923
rect 21928 13892 22293 13920
rect 22281 13889 22293 13892
rect 22327 13889 22339 13923
rect 23842 13920 23848 13932
rect 22281 13883 22339 13889
rect 22940 13892 23848 13920
rect 20533 13855 20591 13861
rect 20533 13852 20545 13855
rect 20088 13824 20545 13852
rect 20533 13821 20545 13824
rect 20579 13821 20591 13855
rect 20533 13815 20591 13821
rect 20806 13812 20812 13864
rect 20864 13852 20870 13864
rect 21836 13852 21864 13880
rect 22005 13855 22063 13861
rect 22005 13852 22017 13855
rect 20864 13824 21778 13852
rect 21836 13824 22017 13852
rect 20864 13812 20870 13824
rect 3528 13756 3924 13784
rect 7484 13756 8064 13784
rect 3234 13676 3240 13728
rect 3292 13676 3298 13728
rect 3528 13725 3556 13756
rect 3513 13719 3571 13725
rect 3513 13685 3525 13719
rect 3559 13685 3571 13719
rect 3513 13679 3571 13685
rect 3878 13676 3884 13728
rect 3936 13716 3942 13728
rect 4255 13719 4313 13725
rect 4255 13716 4267 13719
rect 3936 13688 4267 13716
rect 3936 13676 3942 13688
rect 4255 13685 4267 13688
rect 4301 13685 4313 13719
rect 4255 13679 4313 13685
rect 6454 13676 6460 13728
rect 6512 13716 6518 13728
rect 6555 13719 6613 13725
rect 6555 13716 6567 13719
rect 6512 13688 6567 13716
rect 6512 13676 6518 13688
rect 6555 13685 6567 13688
rect 6601 13685 6613 13719
rect 6555 13679 6613 13685
rect 7190 13676 7196 13728
rect 7248 13716 7254 13728
rect 7484 13716 7512 13756
rect 7248 13688 7512 13716
rect 8036 13716 8064 13756
rect 9858 13744 9864 13796
rect 9916 13784 9922 13796
rect 10597 13787 10655 13793
rect 10597 13784 10609 13787
rect 9916 13756 10609 13784
rect 9916 13744 9922 13756
rect 10597 13753 10609 13756
rect 10643 13753 10655 13787
rect 10597 13747 10655 13753
rect 10686 13744 10692 13796
rect 10744 13784 10750 13796
rect 10744 13756 11376 13784
rect 10744 13744 10750 13756
rect 8855 13719 8913 13725
rect 8855 13716 8867 13719
rect 8036 13688 8867 13716
rect 7248 13676 7254 13688
rect 8855 13685 8867 13688
rect 8901 13685 8913 13719
rect 8855 13679 8913 13685
rect 9122 13676 9128 13728
rect 9180 13716 9186 13728
rect 11238 13716 11244 13728
rect 9180 13688 11244 13716
rect 9180 13676 9186 13688
rect 11238 13676 11244 13688
rect 11296 13676 11302 13728
rect 11348 13716 11376 13756
rect 15930 13744 15936 13796
rect 15988 13784 15994 13796
rect 16206 13784 16212 13796
rect 15988 13756 16212 13784
rect 15988 13744 15994 13756
rect 16206 13744 16212 13756
rect 16264 13744 16270 13796
rect 21750 13784 21778 13824
rect 22005 13821 22017 13824
rect 22051 13821 22063 13855
rect 22940 13852 22968 13892
rect 23842 13880 23848 13892
rect 23900 13880 23906 13932
rect 24044 13929 24072 14016
rect 24394 13929 24400 13932
rect 24029 13923 24087 13929
rect 24029 13889 24041 13923
rect 24075 13889 24087 13923
rect 24029 13883 24087 13889
rect 24356 13923 24400 13929
rect 24356 13889 24368 13923
rect 24356 13883 24400 13889
rect 24394 13880 24400 13883
rect 24452 13880 24458 13932
rect 24578 13927 24584 13932
rect 24535 13921 24584 13927
rect 24535 13887 24547 13921
rect 24581 13887 24584 13921
rect 24535 13881 24584 13887
rect 24578 13880 24584 13881
rect 24636 13880 24642 13932
rect 24670 13880 24676 13932
rect 24728 13920 24734 13932
rect 24765 13923 24823 13929
rect 24765 13920 24777 13923
rect 24728 13892 24777 13920
rect 24728 13880 24734 13892
rect 24765 13889 24777 13892
rect 24811 13889 24823 13923
rect 24765 13883 24823 13889
rect 24946 13880 24952 13932
rect 25004 13880 25010 13932
rect 25424 13920 25452 14028
rect 25866 14016 25872 14068
rect 25924 14016 25930 14068
rect 26053 14059 26111 14065
rect 26053 14025 26065 14059
rect 26099 14056 26111 14059
rect 26326 14056 26332 14068
rect 26099 14028 26332 14056
rect 26099 14025 26111 14028
rect 26053 14019 26111 14025
rect 26326 14016 26332 14028
rect 26384 14016 26390 14068
rect 27430 14016 27436 14068
rect 27488 14056 27494 14068
rect 28537 14059 28595 14065
rect 28537 14056 28549 14059
rect 27488 14028 28549 14056
rect 27488 14016 27494 14028
rect 28537 14025 28549 14028
rect 28583 14025 28595 14059
rect 30101 14059 30159 14065
rect 28537 14019 28595 14025
rect 28644 14028 29592 14056
rect 25884 13988 25912 14016
rect 26605 13991 26663 13997
rect 26605 13988 26617 13991
rect 25884 13960 26617 13988
rect 26605 13957 26617 13960
rect 26651 13957 26663 13991
rect 26605 13951 26663 13957
rect 28166 13948 28172 14000
rect 28224 13988 28230 14000
rect 28644 13988 28672 14028
rect 28224 13960 28672 13988
rect 28224 13948 28230 13960
rect 28994 13948 29000 14000
rect 29052 13988 29058 14000
rect 29270 13988 29276 14000
rect 29052 13960 29276 13988
rect 29052 13948 29058 13960
rect 29270 13948 29276 13960
rect 29328 13948 29334 14000
rect 26694 13920 26700 13932
rect 25424 13892 26700 13920
rect 26694 13880 26700 13892
rect 26752 13880 26758 13932
rect 27203 13923 27261 13929
rect 27203 13889 27215 13923
rect 27249 13920 27261 13923
rect 27433 13923 27491 13929
rect 27249 13892 27384 13920
rect 27249 13889 27261 13892
rect 27203 13883 27261 13889
rect 22005 13815 22063 13821
rect 22112 13824 22968 13852
rect 22112 13784 22140 13824
rect 23658 13812 23664 13864
rect 23716 13852 23722 13864
rect 24964 13852 24992 13880
rect 23716 13824 24992 13852
rect 26421 13855 26479 13861
rect 23716 13812 23722 13824
rect 26421 13821 26433 13855
rect 26467 13821 26479 13855
rect 26421 13815 26479 13821
rect 26436 13784 26464 13815
rect 26786 13812 26792 13864
rect 26844 13852 26850 13864
rect 27024 13855 27082 13861
rect 27024 13852 27036 13855
rect 26844 13824 27036 13852
rect 26844 13812 26850 13824
rect 27024 13821 27036 13824
rect 27070 13821 27082 13855
rect 27356 13852 27384 13892
rect 27433 13889 27445 13923
rect 27479 13920 27491 13923
rect 29564 13920 29592 14028
rect 30101 14025 30113 14059
rect 30147 14056 30159 14059
rect 30466 14056 30472 14068
rect 30147 14028 30472 14056
rect 30147 14025 30159 14028
rect 30101 14019 30159 14025
rect 30466 14016 30472 14028
rect 30524 14016 30530 14068
rect 30282 13948 30288 14000
rect 30340 13948 30346 14000
rect 27479 13892 29316 13920
rect 29564 13892 29684 13920
rect 27479 13889 27491 13892
rect 27433 13883 27491 13889
rect 29288 13864 29316 13892
rect 29656 13868 29684 13892
rect 30374 13880 30380 13932
rect 30432 13880 30438 13932
rect 27356 13824 28304 13852
rect 27024 13815 27082 13821
rect 26602 13784 26608 13796
rect 21750 13756 22140 13784
rect 23308 13756 24164 13784
rect 26436 13756 26608 13784
rect 11882 13716 11888 13728
rect 11348 13688 11888 13716
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 14651 13719 14709 13725
rect 14651 13685 14663 13719
rect 14697 13716 14709 13719
rect 14826 13716 14832 13728
rect 14697 13688 14832 13716
rect 14697 13685 14709 13688
rect 14651 13679 14709 13685
rect 14826 13676 14832 13688
rect 14884 13676 14890 13728
rect 20254 13676 20260 13728
rect 20312 13725 20318 13728
rect 20312 13679 20321 13725
rect 20312 13676 20318 13679
rect 20990 13676 20996 13728
rect 21048 13716 21054 13728
rect 23308 13716 23336 13756
rect 21048 13688 23336 13716
rect 24136 13716 24164 13756
rect 26602 13744 26608 13756
rect 26660 13744 26666 13796
rect 28276 13728 28304 13824
rect 28994 13812 29000 13864
rect 29052 13852 29058 13864
rect 29089 13855 29147 13861
rect 29089 13852 29101 13855
rect 29052 13824 29101 13852
rect 29052 13812 29058 13824
rect 29089 13821 29101 13824
rect 29135 13852 29147 13855
rect 29178 13852 29184 13864
rect 29135 13824 29184 13852
rect 29135 13821 29147 13824
rect 29089 13815 29147 13821
rect 29178 13812 29184 13824
rect 29236 13812 29242 13864
rect 29270 13812 29276 13864
rect 29328 13812 29334 13864
rect 29362 13812 29368 13864
rect 29420 13852 29426 13864
rect 29656 13852 29776 13868
rect 29825 13855 29883 13861
rect 29825 13852 29837 13855
rect 29420 13824 29500 13852
rect 29656 13840 29837 13852
rect 29748 13824 29837 13840
rect 29420 13812 29426 13824
rect 28534 13744 28540 13796
rect 28592 13784 28598 13796
rect 29472 13793 29500 13824
rect 29825 13821 29837 13824
rect 29871 13821 29883 13855
rect 30392 13852 30420 13880
rect 30469 13855 30527 13861
rect 30469 13852 30481 13855
rect 30392 13824 30481 13852
rect 29825 13815 29883 13821
rect 30469 13821 30481 13824
rect 30515 13821 30527 13855
rect 30469 13815 30527 13821
rect 29457 13787 29515 13793
rect 29457 13784 29469 13787
rect 28592 13756 29469 13784
rect 28592 13744 28598 13756
rect 29457 13753 29469 13756
rect 29503 13753 29515 13787
rect 29457 13747 29515 13753
rect 27706 13716 27712 13728
rect 24136 13688 27712 13716
rect 21048 13676 21054 13688
rect 27706 13676 27712 13688
rect 27764 13676 27770 13728
rect 28258 13676 28264 13728
rect 28316 13676 28322 13728
rect 28626 13676 28632 13728
rect 28684 13716 28690 13728
rect 29549 13719 29607 13725
rect 29549 13716 29561 13719
rect 28684 13688 29561 13716
rect 28684 13676 28690 13688
rect 29549 13685 29561 13688
rect 29595 13716 29607 13719
rect 30558 13716 30564 13728
rect 29595 13688 30564 13716
rect 29595 13685 29607 13688
rect 29549 13679 29607 13685
rect 30558 13676 30564 13688
rect 30616 13676 30622 13728
rect 552 13626 31072 13648
rect 552 13574 7988 13626
rect 8040 13574 8052 13626
rect 8104 13574 8116 13626
rect 8168 13574 8180 13626
rect 8232 13574 8244 13626
rect 8296 13574 15578 13626
rect 15630 13574 15642 13626
rect 15694 13574 15706 13626
rect 15758 13574 15770 13626
rect 15822 13574 15834 13626
rect 15886 13574 23168 13626
rect 23220 13574 23232 13626
rect 23284 13574 23296 13626
rect 23348 13574 23360 13626
rect 23412 13574 23424 13626
rect 23476 13574 30758 13626
rect 30810 13574 30822 13626
rect 30874 13574 30886 13626
rect 30938 13574 30950 13626
rect 31002 13574 31014 13626
rect 31066 13574 31072 13626
rect 552 13552 31072 13574
rect 750 13472 756 13524
rect 808 13512 814 13524
rect 1762 13512 1768 13524
rect 808 13484 1768 13512
rect 808 13472 814 13484
rect 1762 13472 1768 13484
rect 1820 13472 1826 13524
rect 5258 13512 5264 13524
rect 2746 13484 5264 13512
rect 1118 13404 1124 13456
rect 1176 13404 1182 13456
rect 1136 13376 1164 13404
rect 1213 13379 1271 13385
rect 1213 13376 1225 13379
rect 1136 13348 1225 13376
rect 1213 13345 1225 13348
rect 1259 13345 1271 13379
rect 1213 13339 1271 13345
rect 1801 13329 1859 13335
rect 1302 13268 1308 13320
rect 1360 13308 1366 13320
rect 1486 13308 1492 13320
rect 1360 13280 1492 13308
rect 1360 13268 1366 13280
rect 1486 13268 1492 13280
rect 1544 13268 1550 13320
rect 1670 13317 1676 13320
rect 1632 13311 1676 13317
rect 1632 13277 1644 13311
rect 1632 13271 1676 13277
rect 1670 13268 1676 13271
rect 1728 13268 1734 13320
rect 1801 13295 1813 13329
rect 1847 13308 1859 13329
rect 1946 13308 1952 13320
rect 1847 13295 1952 13308
rect 1801 13289 1952 13295
rect 1826 13280 1952 13289
rect 1946 13268 1952 13280
rect 2004 13268 2010 13320
rect 2038 13268 2044 13320
rect 2096 13268 2102 13320
rect 1029 13175 1087 13181
rect 1029 13141 1041 13175
rect 1075 13172 1087 13175
rect 2746 13172 2774 13484
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 5350 13472 5356 13524
rect 5408 13512 5414 13524
rect 6086 13512 6092 13524
rect 5408 13484 6092 13512
rect 5408 13472 5414 13484
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 6181 13515 6239 13521
rect 6181 13481 6193 13515
rect 6227 13512 6239 13515
rect 7374 13512 7380 13524
rect 6227 13484 7380 13512
rect 6227 13481 6239 13484
rect 6181 13475 6239 13481
rect 7374 13472 7380 13484
rect 7432 13472 7438 13524
rect 8570 13472 8576 13524
rect 8628 13472 8634 13524
rect 8662 13472 8668 13524
rect 8720 13472 8726 13524
rect 8938 13472 8944 13524
rect 8996 13472 9002 13524
rect 9214 13472 9220 13524
rect 9272 13472 9278 13524
rect 9398 13472 9404 13524
rect 9456 13512 9462 13524
rect 9493 13515 9551 13521
rect 9493 13512 9505 13515
rect 9456 13484 9505 13512
rect 9456 13472 9462 13484
rect 9493 13481 9505 13484
rect 9539 13481 9551 13515
rect 9493 13475 9551 13481
rect 9582 13472 9588 13524
rect 9640 13512 9646 13524
rect 9769 13515 9827 13521
rect 9769 13512 9781 13515
rect 9640 13484 9781 13512
rect 9640 13472 9646 13484
rect 9769 13481 9781 13484
rect 9815 13481 9827 13515
rect 9769 13475 9827 13481
rect 11146 13472 11152 13524
rect 11204 13472 11210 13524
rect 11422 13472 11428 13524
rect 11480 13472 11486 13524
rect 11882 13472 11888 13524
rect 11940 13472 11946 13524
rect 12158 13472 12164 13524
rect 12216 13512 12222 13524
rect 12253 13515 12311 13521
rect 12253 13512 12265 13515
rect 12216 13484 12265 13512
rect 12216 13472 12222 13484
rect 12253 13481 12265 13484
rect 12299 13481 12311 13515
rect 12526 13512 12532 13524
rect 12253 13475 12311 13481
rect 12452 13484 12532 13512
rect 5629 13447 5687 13453
rect 5629 13413 5641 13447
rect 5675 13444 5687 13447
rect 6270 13444 6276 13456
rect 5675 13416 6276 13444
rect 5675 13413 5687 13416
rect 5629 13407 5687 13413
rect 6270 13404 6276 13416
rect 6328 13404 6334 13456
rect 8680 13444 8708 13472
rect 11164 13444 11192 13472
rect 11606 13444 11612 13456
rect 8680 13416 9444 13444
rect 6641 13403 6699 13409
rect 6641 13400 6653 13403
rect 3421 13379 3479 13385
rect 3421 13345 3433 13379
rect 3467 13376 3479 13379
rect 5997 13379 6055 13385
rect 3467 13348 4019 13376
rect 3467 13345 3479 13348
rect 3421 13339 3479 13345
rect 3878 13317 3884 13320
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13277 3571 13311
rect 3513 13271 3571 13277
rect 3840 13311 3884 13317
rect 3840 13277 3852 13311
rect 3840 13271 3884 13277
rect 1075 13144 2774 13172
rect 3528 13172 3556 13271
rect 3878 13268 3884 13271
rect 3936 13268 3942 13320
rect 3991 13319 4019 13348
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 6362 13376 6368 13388
rect 6043 13348 6368 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 3976 13313 4034 13319
rect 3976 13279 3988 13313
rect 4022 13279 4034 13313
rect 3976 13273 4034 13279
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13308 4307 13311
rect 5810 13308 5816 13320
rect 4295 13280 5816 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 4982 13200 4988 13252
rect 5040 13240 5046 13252
rect 6012 13240 6040 13339
rect 6362 13336 6368 13348
rect 6420 13336 6426 13388
rect 6567 13380 6653 13400
rect 6475 13376 6653 13380
rect 6472 13372 6653 13376
rect 6472 13352 6595 13372
rect 6641 13369 6653 13372
rect 6687 13369 6699 13403
rect 6641 13363 6699 13369
rect 9125 13379 9183 13385
rect 6472 13348 6503 13352
rect 6086 13268 6092 13320
rect 6144 13308 6150 13320
rect 6472 13308 6500 13348
rect 9125 13345 9137 13379
rect 9171 13376 9183 13379
rect 9306 13376 9312 13388
rect 9171 13348 9312 13376
rect 9171 13345 9183 13348
rect 9125 13339 9183 13345
rect 9306 13336 9312 13348
rect 9364 13336 9370 13388
rect 9416 13385 9444 13416
rect 9968 13416 11612 13444
rect 9401 13379 9459 13385
rect 9401 13345 9413 13379
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 9674 13336 9680 13388
rect 9732 13336 9738 13388
rect 9858 13336 9864 13388
rect 9916 13376 9922 13388
rect 9968 13385 9996 13416
rect 11606 13404 11612 13416
rect 11664 13404 11670 13456
rect 9953 13379 10011 13385
rect 9953 13376 9965 13379
rect 9916 13348 9965 13376
rect 9916 13336 9922 13348
rect 9953 13345 9965 13348
rect 9999 13345 10011 13379
rect 9953 13339 10011 13345
rect 10226 13336 10232 13388
rect 10284 13336 10290 13388
rect 10318 13336 10324 13388
rect 10376 13376 10382 13388
rect 10505 13379 10563 13385
rect 10505 13376 10517 13379
rect 10376 13348 10517 13376
rect 10376 13336 10382 13348
rect 10505 13345 10517 13348
rect 10551 13345 10563 13379
rect 10505 13339 10563 13345
rect 10778 13336 10784 13388
rect 10836 13336 10842 13388
rect 11054 13336 11060 13388
rect 11112 13376 11118 13388
rect 11149 13379 11207 13385
rect 11149 13376 11161 13379
rect 11112 13348 11161 13376
rect 11112 13336 11118 13348
rect 11149 13345 11161 13348
rect 11195 13376 11207 13379
rect 11422 13376 11428 13388
rect 11195 13348 11428 13376
rect 11195 13345 11207 13348
rect 11149 13339 11207 13345
rect 11422 13336 11428 13348
rect 11480 13376 11486 13388
rect 12452 13385 12480 13484
rect 12526 13472 12532 13484
rect 12584 13512 12590 13524
rect 13262 13512 13268 13524
rect 12584 13484 13268 13512
rect 12584 13472 12590 13484
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 14550 13472 14556 13524
rect 14608 13512 14614 13524
rect 14737 13515 14795 13521
rect 14737 13512 14749 13515
rect 14608 13484 14749 13512
rect 14608 13472 14614 13484
rect 14737 13481 14749 13484
rect 14783 13481 14795 13515
rect 14737 13475 14795 13481
rect 14826 13472 14832 13524
rect 14884 13472 14890 13524
rect 15102 13472 15108 13524
rect 15160 13512 15166 13524
rect 17957 13515 18015 13521
rect 17957 13512 17969 13515
rect 15160 13484 17969 13512
rect 15160 13472 15166 13484
rect 17957 13481 17969 13484
rect 18003 13481 18015 13515
rect 17957 13475 18015 13481
rect 18791 13515 18849 13521
rect 18791 13481 18803 13515
rect 18837 13512 18849 13515
rect 19150 13512 19156 13524
rect 18837 13484 19156 13512
rect 18837 13481 18849 13484
rect 18791 13475 18849 13481
rect 19150 13472 19156 13484
rect 19208 13472 19214 13524
rect 22379 13515 22437 13521
rect 22379 13481 22391 13515
rect 22425 13512 22437 13515
rect 24026 13512 24032 13524
rect 22425 13484 24032 13512
rect 22425 13481 22437 13484
rect 22379 13475 22437 13481
rect 24026 13472 24032 13484
rect 24084 13472 24090 13524
rect 24587 13515 24645 13521
rect 24587 13481 24599 13515
rect 24633 13512 24645 13515
rect 26145 13515 26203 13521
rect 24633 13484 25544 13512
rect 24633 13481 24645 13484
rect 24587 13475 24645 13481
rect 14844 13444 14872 13472
rect 15289 13447 15347 13453
rect 15289 13444 15301 13447
rect 14844 13416 15301 13444
rect 15289 13413 15301 13416
rect 15335 13413 15347 13447
rect 15289 13407 15347 13413
rect 15378 13404 15384 13456
rect 15436 13404 15442 13456
rect 11701 13379 11759 13385
rect 11701 13376 11713 13379
rect 11480 13348 11713 13376
rect 11480 13336 11486 13348
rect 11701 13345 11713 13348
rect 11747 13345 11759 13379
rect 11701 13339 11759 13345
rect 12161 13379 12219 13385
rect 12161 13345 12173 13379
rect 12207 13376 12219 13379
rect 12437 13379 12495 13385
rect 12207 13348 12394 13376
rect 12207 13345 12219 13348
rect 12161 13339 12219 13345
rect 6144 13280 6500 13308
rect 6144 13268 6150 13280
rect 6730 13268 6736 13320
rect 6788 13317 6794 13320
rect 6788 13308 6799 13317
rect 6788 13280 6833 13308
rect 6788 13271 6799 13280
rect 6788 13268 6794 13271
rect 7006 13268 7012 13320
rect 7064 13317 7070 13320
rect 7064 13311 7118 13317
rect 7064 13277 7072 13311
rect 7106 13277 7118 13311
rect 7064 13271 7118 13277
rect 7064 13268 7070 13271
rect 7190 13268 7196 13320
rect 7248 13268 7254 13320
rect 7466 13268 7472 13320
rect 7524 13268 7530 13320
rect 9490 13268 9496 13320
rect 9548 13308 9554 13320
rect 9548 13280 11376 13308
rect 9548 13268 9554 13280
rect 5040 13212 6040 13240
rect 5040 13200 5046 13212
rect 8386 13200 8392 13252
rect 8444 13240 8450 13252
rect 9214 13240 9220 13252
rect 8444 13212 9220 13240
rect 8444 13200 8450 13212
rect 9214 13200 9220 13212
rect 9272 13240 9278 13252
rect 11348 13249 11376 13280
rect 11333 13243 11391 13249
rect 9272 13212 11290 13240
rect 9272 13200 9278 13212
rect 3786 13172 3792 13184
rect 3528 13144 3792 13172
rect 1075 13141 1087 13144
rect 1029 13135 1087 13141
rect 3786 13132 3792 13144
rect 3844 13132 3850 13184
rect 5442 13132 5448 13184
rect 5500 13172 5506 13184
rect 5813 13175 5871 13181
rect 5813 13172 5825 13175
rect 5500 13144 5825 13172
rect 5500 13132 5506 13144
rect 5813 13141 5825 13144
rect 5859 13141 5871 13175
rect 5813 13135 5871 13141
rect 6457 13175 6515 13181
rect 6457 13141 6469 13175
rect 6503 13172 6515 13175
rect 6638 13172 6644 13184
rect 6503 13144 6644 13172
rect 6503 13141 6515 13144
rect 6457 13135 6515 13141
rect 6638 13132 6644 13144
rect 6696 13132 6702 13184
rect 7926 13132 7932 13184
rect 7984 13172 7990 13184
rect 9674 13172 9680 13184
rect 7984 13144 9680 13172
rect 7984 13132 7990 13144
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 10045 13175 10103 13181
rect 10045 13141 10057 13175
rect 10091 13172 10103 13175
rect 10226 13172 10232 13184
rect 10091 13144 10232 13172
rect 10091 13141 10103 13144
rect 10045 13135 10103 13141
rect 10226 13132 10232 13144
rect 10284 13132 10290 13184
rect 10321 13175 10379 13181
rect 10321 13141 10333 13175
rect 10367 13172 10379 13175
rect 10410 13172 10416 13184
rect 10367 13144 10416 13172
rect 10367 13141 10379 13144
rect 10321 13135 10379 13141
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 10594 13132 10600 13184
rect 10652 13132 10658 13184
rect 11262 13172 11290 13212
rect 11333 13209 11345 13243
rect 11379 13209 11391 13243
rect 12366 13240 12394 13348
rect 12437 13345 12449 13379
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 12856 13379 12914 13385
rect 12856 13345 12868 13379
rect 12902 13376 12914 13379
rect 12902 13348 13676 13376
rect 12902 13345 12914 13348
rect 12856 13339 12914 13345
rect 13648 13320 13676 13348
rect 14918 13336 14924 13388
rect 14976 13336 14982 13388
rect 15013 13379 15071 13385
rect 15013 13345 15025 13379
rect 15059 13345 15071 13379
rect 15396 13376 15424 13404
rect 15933 13379 15991 13385
rect 15933 13376 15945 13379
rect 15396 13348 15945 13376
rect 15013 13339 15071 13345
rect 15933 13345 15945 13348
rect 15979 13376 15991 13379
rect 16022 13376 16028 13388
rect 15979 13348 16028 13376
rect 15979 13345 15991 13348
rect 15933 13339 15991 13345
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13308 12587 13311
rect 12710 13308 12716 13320
rect 12575 13280 12716 13308
rect 12575 13277 12587 13280
rect 12529 13271 12587 13277
rect 12710 13268 12716 13280
rect 12768 13268 12774 13320
rect 13035 13311 13093 13317
rect 13035 13277 13047 13311
rect 13081 13308 13093 13311
rect 13170 13308 13176 13320
rect 13081 13280 13176 13308
rect 13081 13277 13093 13280
rect 13035 13271 13093 13277
rect 13170 13268 13176 13280
rect 13228 13268 13234 13320
rect 13262 13268 13268 13320
rect 13320 13268 13326 13320
rect 13630 13268 13636 13320
rect 13688 13268 13694 13320
rect 14936 13240 14964 13336
rect 11333 13203 11391 13209
rect 11440 13212 12394 13240
rect 11440 13172 11468 13212
rect 11262 13144 11468 13172
rect 11977 13175 12035 13181
rect 11977 13141 11989 13175
rect 12023 13172 12035 13175
rect 12250 13172 12256 13184
rect 12023 13144 12256 13172
rect 12023 13141 12035 13144
rect 11977 13135 12035 13141
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 12366 13172 12394 13212
rect 13924 13212 14964 13240
rect 15028 13240 15056 13339
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 21821 13379 21879 13385
rect 21821 13345 21833 13379
rect 21867 13345 21879 13379
rect 21821 13339 21879 13345
rect 21913 13379 21971 13385
rect 21913 13345 21925 13379
rect 21959 13376 21971 13379
rect 23658 13376 23664 13388
rect 21959 13348 23664 13376
rect 21959 13345 21971 13348
rect 21913 13339 21971 13345
rect 15102 13268 15108 13320
rect 15160 13308 15166 13320
rect 16117 13311 16175 13317
rect 16117 13308 16129 13311
rect 15160 13280 16129 13308
rect 15160 13268 15166 13280
rect 16117 13277 16129 13280
rect 16163 13277 16175 13311
rect 16117 13271 16175 13277
rect 16298 13268 16304 13320
rect 16356 13308 16362 13320
rect 16444 13311 16502 13317
rect 16444 13308 16456 13311
rect 16356 13280 16456 13308
rect 16356 13268 16362 13280
rect 16444 13277 16456 13280
rect 16490 13277 16502 13311
rect 16444 13271 16502 13277
rect 16574 13268 16580 13320
rect 16632 13268 16638 13320
rect 16850 13268 16856 13320
rect 16908 13268 16914 13320
rect 18325 13311 18383 13317
rect 18325 13277 18337 13311
rect 18371 13308 18383 13311
rect 18598 13308 18604 13320
rect 18371 13280 18604 13308
rect 18371 13277 18383 13280
rect 18325 13271 18383 13277
rect 18598 13268 18604 13280
rect 18656 13268 18662 13320
rect 18782 13268 18788 13320
rect 18840 13268 18846 13320
rect 19061 13311 19119 13317
rect 19061 13277 19073 13311
rect 19107 13308 19119 13311
rect 19702 13308 19708 13320
rect 19107 13280 19708 13308
rect 19107 13277 19119 13280
rect 19061 13271 19119 13277
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 20162 13268 20168 13320
rect 20220 13308 20226 13320
rect 21836 13308 21864 13339
rect 23658 13336 23664 13348
rect 23716 13336 23722 13388
rect 24029 13379 24087 13385
rect 24029 13345 24041 13379
rect 24075 13376 24087 13379
rect 25516 13376 25544 13484
rect 26145 13481 26157 13515
rect 26191 13512 26203 13515
rect 26878 13512 26884 13524
rect 26191 13484 26884 13512
rect 26191 13481 26203 13484
rect 26145 13475 26203 13481
rect 26878 13472 26884 13484
rect 26936 13472 26942 13524
rect 27614 13472 27620 13524
rect 27672 13512 27678 13524
rect 28261 13515 28319 13521
rect 28261 13512 28273 13515
rect 27672 13484 28273 13512
rect 27672 13472 27678 13484
rect 28261 13481 28273 13484
rect 28307 13481 28319 13515
rect 28261 13475 28319 13481
rect 29270 13472 29276 13524
rect 29328 13512 29334 13524
rect 30009 13515 30067 13521
rect 30009 13512 30021 13515
rect 29328 13484 30021 13512
rect 29328 13472 29334 13484
rect 30009 13481 30021 13484
rect 30055 13481 30067 13515
rect 30009 13475 30067 13481
rect 30282 13472 30288 13524
rect 30340 13512 30346 13524
rect 30377 13515 30435 13521
rect 30377 13512 30389 13515
rect 30340 13484 30389 13512
rect 30340 13472 30346 13484
rect 30377 13481 30389 13484
rect 30423 13481 30435 13515
rect 30377 13475 30435 13481
rect 30466 13404 30472 13456
rect 30524 13404 30530 13456
rect 26786 13385 26792 13388
rect 26748 13379 26792 13385
rect 26748 13376 26760 13379
rect 24075 13348 24394 13376
rect 25516 13348 26760 13376
rect 24075 13345 24087 13348
rect 24029 13339 24087 13345
rect 24366 13326 24394 13348
rect 26748 13345 26760 13348
rect 26748 13339 26792 13345
rect 26786 13336 26792 13339
rect 26844 13336 26850 13388
rect 28350 13336 28356 13388
rect 28408 13376 28414 13388
rect 28629 13379 28687 13385
rect 28629 13376 28641 13379
rect 28408 13348 28641 13376
rect 28408 13336 28414 13348
rect 28629 13345 28641 13348
rect 28675 13345 28687 13379
rect 28629 13339 28687 13345
rect 28905 13379 28963 13385
rect 28905 13345 28917 13379
rect 28951 13376 28963 13379
rect 30006 13376 30012 13388
rect 28951 13348 30012 13376
rect 28951 13345 28963 13348
rect 28905 13339 28963 13345
rect 30006 13336 30012 13348
rect 30064 13336 30070 13388
rect 30484 13376 30512 13404
rect 30561 13379 30619 13385
rect 30561 13376 30573 13379
rect 30484 13348 30573 13376
rect 30561 13345 30573 13348
rect 30607 13345 30619 13379
rect 30561 13339 30619 13345
rect 24584 13329 24642 13335
rect 24584 13326 24596 13329
rect 22094 13308 22100 13320
rect 20220 13280 22100 13308
rect 20220 13268 20226 13280
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 22462 13317 22468 13320
rect 22419 13311 22468 13317
rect 22419 13277 22431 13311
rect 22465 13277 22468 13311
rect 22419 13271 22468 13277
rect 22462 13268 22468 13271
rect 22520 13268 22526 13320
rect 22646 13268 22652 13320
rect 22704 13268 22710 13320
rect 24118 13268 24124 13320
rect 24176 13268 24182 13320
rect 24366 13298 24596 13326
rect 24584 13295 24596 13298
rect 24630 13295 24642 13329
rect 24584 13289 24642 13295
rect 24857 13311 24915 13317
rect 24857 13277 24869 13311
rect 24903 13308 24915 13311
rect 25038 13308 25044 13320
rect 24903 13280 25044 13308
rect 24903 13277 24915 13280
rect 24857 13271 24915 13277
rect 25038 13268 25044 13280
rect 25096 13268 25102 13320
rect 26421 13311 26479 13317
rect 26421 13277 26433 13311
rect 26467 13308 26479 13311
rect 26602 13308 26608 13320
rect 26467 13280 26608 13308
rect 26467 13277 26479 13280
rect 26421 13271 26479 13277
rect 26602 13268 26608 13280
rect 26660 13268 26666 13320
rect 26878 13268 26884 13320
rect 26936 13268 26942 13320
rect 27157 13311 27215 13317
rect 27157 13277 27169 13311
rect 27203 13308 27215 13311
rect 27338 13308 27344 13320
rect 27203 13280 27344 13308
rect 27203 13277 27215 13280
rect 27157 13271 27215 13277
rect 27338 13268 27344 13280
rect 27396 13268 27402 13320
rect 15028 13212 16160 13240
rect 13924 13172 13952 13212
rect 12366 13144 13952 13172
rect 14366 13132 14372 13184
rect 14424 13132 14430 13184
rect 14458 13132 14464 13184
rect 14516 13172 14522 13184
rect 15028 13172 15056 13212
rect 14516 13144 15056 13172
rect 14516 13132 14522 13144
rect 15746 13132 15752 13184
rect 15804 13132 15810 13184
rect 16132 13172 16160 13212
rect 18690 13172 18696 13184
rect 16132 13144 18696 13172
rect 18690 13132 18696 13144
rect 18748 13132 18754 13184
rect 20346 13132 20352 13184
rect 20404 13132 20410 13184
rect 21637 13175 21695 13181
rect 21637 13141 21649 13175
rect 21683 13172 21695 13175
rect 24118 13172 24124 13184
rect 21683 13144 24124 13172
rect 21683 13141 21695 13144
rect 21637 13135 21695 13141
rect 24118 13132 24124 13144
rect 24176 13132 24182 13184
rect 24302 13132 24308 13184
rect 24360 13172 24366 13184
rect 29546 13172 29552 13184
rect 24360 13144 29552 13172
rect 24360 13132 24366 13144
rect 29546 13132 29552 13144
rect 29604 13132 29610 13184
rect 30282 13132 30288 13184
rect 30340 13172 30346 13184
rect 31202 13172 31208 13184
rect 30340 13144 31208 13172
rect 30340 13132 30346 13144
rect 31202 13132 31208 13144
rect 31260 13132 31266 13184
rect 552 13082 30912 13104
rect 552 13030 4193 13082
rect 4245 13030 4257 13082
rect 4309 13030 4321 13082
rect 4373 13030 4385 13082
rect 4437 13030 4449 13082
rect 4501 13030 11783 13082
rect 11835 13030 11847 13082
rect 11899 13030 11911 13082
rect 11963 13030 11975 13082
rect 12027 13030 12039 13082
rect 12091 13030 19373 13082
rect 19425 13030 19437 13082
rect 19489 13030 19501 13082
rect 19553 13030 19565 13082
rect 19617 13030 19629 13082
rect 19681 13030 26963 13082
rect 27015 13030 27027 13082
rect 27079 13030 27091 13082
rect 27143 13030 27155 13082
rect 27207 13030 27219 13082
rect 27271 13030 30912 13082
rect 552 13008 30912 13030
rect 3142 12928 3148 12980
rect 3200 12968 3206 12980
rect 3513 12971 3571 12977
rect 3513 12968 3525 12971
rect 3200 12940 3525 12968
rect 3200 12928 3206 12940
rect 3513 12937 3525 12940
rect 3559 12937 3571 12971
rect 3513 12931 3571 12937
rect 3602 12928 3608 12980
rect 3660 12968 3666 12980
rect 5718 12968 5724 12980
rect 3660 12940 5724 12968
rect 3660 12928 3666 12940
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 7190 12968 7196 12980
rect 5951 12940 7196 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 7466 12928 7472 12980
rect 7524 12968 7530 12980
rect 8757 12971 8815 12977
rect 8757 12968 8769 12971
rect 7524 12940 8769 12968
rect 7524 12928 7530 12940
rect 8757 12937 8769 12940
rect 8803 12937 8815 12971
rect 8757 12931 8815 12937
rect 9306 12928 9312 12980
rect 9364 12968 9370 12980
rect 9364 12940 9628 12968
rect 9364 12928 9370 12940
rect 937 12835 995 12841
rect 937 12801 949 12835
rect 983 12832 995 12835
rect 1302 12832 1308 12844
rect 983 12804 1308 12832
rect 983 12801 995 12804
rect 937 12795 995 12801
rect 1302 12792 1308 12804
rect 1360 12792 1366 12844
rect 1443 12835 1501 12841
rect 1443 12801 1455 12835
rect 1489 12832 1501 12835
rect 2130 12832 2136 12844
rect 1489 12804 2136 12832
rect 1489 12801 1501 12804
rect 1443 12795 1501 12801
rect 2130 12792 2136 12804
rect 2188 12792 2194 12844
rect 3053 12835 3111 12841
rect 3053 12801 3065 12835
rect 3099 12832 3111 12835
rect 4344 12835 4402 12841
rect 4344 12832 4356 12835
rect 3099 12804 4356 12832
rect 3099 12801 3111 12804
rect 3053 12795 3111 12801
rect 4344 12801 4356 12804
rect 4390 12801 4402 12835
rect 4344 12795 4402 12801
rect 4614 12792 4620 12844
rect 4672 12792 4678 12844
rect 5736 12832 5764 12928
rect 7834 12860 7840 12912
rect 7892 12900 7898 12912
rect 9033 12903 9091 12909
rect 9033 12900 9045 12903
rect 7892 12872 9045 12900
rect 7892 12860 7898 12872
rect 9033 12869 9045 12872
rect 9079 12869 9091 12903
rect 9033 12863 9091 12869
rect 9490 12860 9496 12912
rect 9548 12860 9554 12912
rect 6638 12839 6644 12844
rect 6595 12833 6644 12839
rect 5736 12830 6040 12832
rect 6104 12830 6500 12832
rect 5736 12804 6500 12830
rect 6012 12802 6132 12804
rect 1673 12767 1731 12773
rect 1673 12733 1685 12767
rect 1719 12764 1731 12767
rect 3234 12764 3240 12776
rect 1719 12736 3240 12764
rect 1719 12733 1731 12736
rect 1673 12727 1731 12733
rect 3234 12724 3240 12736
rect 3292 12724 3298 12776
rect 3421 12767 3479 12773
rect 3421 12733 3433 12767
rect 3467 12733 3479 12767
rect 3421 12727 3479 12733
rect 3436 12696 3464 12727
rect 3602 12724 3608 12776
rect 3660 12764 3666 12776
rect 3697 12767 3755 12773
rect 3697 12764 3709 12767
rect 3660 12736 3709 12764
rect 3660 12724 3666 12736
rect 3697 12733 3709 12736
rect 3743 12733 3755 12767
rect 3697 12727 3755 12733
rect 3786 12724 3792 12776
rect 3844 12764 3850 12776
rect 3881 12767 3939 12773
rect 3881 12764 3893 12767
rect 3844 12736 3893 12764
rect 3844 12724 3850 12736
rect 3881 12733 3893 12736
rect 3927 12733 3939 12767
rect 5350 12764 5356 12776
rect 3881 12727 3939 12733
rect 3994 12736 5356 12764
rect 3994 12696 4022 12736
rect 5350 12724 5356 12736
rect 5408 12724 5414 12776
rect 6089 12767 6147 12773
rect 6089 12764 6101 12767
rect 6012 12736 6101 12764
rect 3436 12668 4022 12696
rect 6012 12640 6040 12736
rect 6089 12733 6101 12736
rect 6135 12733 6147 12767
rect 6472 12764 6500 12804
rect 6595 12799 6607 12833
rect 6641 12799 6644 12833
rect 6595 12793 6644 12799
rect 6638 12792 6644 12793
rect 6696 12792 6702 12844
rect 6730 12792 6736 12844
rect 6788 12832 6794 12844
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6788 12804 6837 12832
rect 6788 12792 6794 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 8312 12804 9260 12832
rect 8312 12764 8340 12804
rect 6472 12736 8340 12764
rect 8389 12767 8447 12773
rect 6089 12727 6147 12733
rect 8389 12733 8401 12767
rect 8435 12764 8447 12767
rect 8846 12764 8852 12776
rect 8435 12736 8852 12764
rect 8435 12733 8447 12736
rect 8389 12727 8447 12733
rect 8846 12724 8852 12736
rect 8904 12724 8910 12776
rect 9232 12773 9260 12804
rect 9508 12773 9536 12860
rect 9600 12832 9628 12940
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 12529 12971 12587 12977
rect 11480 12940 12488 12968
rect 11480 12928 11486 12940
rect 11330 12860 11336 12912
rect 11388 12900 11394 12912
rect 12460 12900 12488 12940
rect 12529 12937 12541 12971
rect 12575 12968 12587 12971
rect 12802 12968 12808 12980
rect 12575 12940 12808 12968
rect 12575 12937 12587 12940
rect 12529 12931 12587 12937
rect 12802 12928 12808 12940
rect 12860 12928 12866 12980
rect 16206 12928 16212 12980
rect 16264 12968 16270 12980
rect 16850 12968 16856 12980
rect 16264 12940 16856 12968
rect 16264 12928 16270 12940
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 17954 12928 17960 12980
rect 18012 12968 18018 12980
rect 18233 12971 18291 12977
rect 18233 12968 18245 12971
rect 18012 12940 18245 12968
rect 18012 12928 18018 12940
rect 18233 12937 18245 12940
rect 18279 12937 18291 12971
rect 18966 12968 18972 12980
rect 18233 12931 18291 12937
rect 18708 12940 18972 12968
rect 13446 12900 13452 12912
rect 11388 12872 12112 12900
rect 12460 12872 13452 12900
rect 11388 12860 11394 12872
rect 9600 12826 9720 12832
rect 9600 12804 9680 12826
rect 8941 12767 8999 12773
rect 8941 12733 8953 12767
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 9217 12767 9275 12773
rect 9217 12733 9229 12767
rect 9263 12733 9275 12767
rect 9217 12727 9275 12733
rect 9493 12767 9551 12773
rect 9493 12733 9505 12767
rect 9539 12733 9551 12767
rect 9493 12727 9551 12733
rect 8205 12699 8263 12705
rect 8205 12665 8217 12699
rect 8251 12696 8263 12699
rect 8251 12668 8892 12696
rect 8251 12665 8263 12668
rect 8205 12659 8263 12665
rect 8864 12640 8892 12668
rect 1403 12631 1461 12637
rect 1403 12597 1415 12631
rect 1449 12628 1461 12631
rect 1670 12628 1676 12640
rect 1449 12600 1676 12628
rect 1449 12597 1461 12600
rect 1403 12591 1461 12597
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 3234 12588 3240 12640
rect 3292 12588 3298 12640
rect 3970 12588 3976 12640
rect 4028 12628 4034 12640
rect 4347 12631 4405 12637
rect 4347 12628 4359 12631
rect 4028 12600 4359 12628
rect 4028 12588 4034 12600
rect 4347 12597 4359 12600
rect 4393 12597 4405 12631
rect 4347 12591 4405 12597
rect 5994 12588 6000 12640
rect 6052 12588 6058 12640
rect 6454 12588 6460 12640
rect 6512 12628 6518 12640
rect 6555 12631 6613 12637
rect 6555 12628 6567 12631
rect 6512 12600 6567 12628
rect 6512 12588 6518 12600
rect 6555 12597 6567 12600
rect 6601 12628 6613 12631
rect 7098 12628 7104 12640
rect 6601 12600 7104 12628
rect 6601 12597 6613 12600
rect 6555 12591 6613 12597
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 7466 12588 7472 12640
rect 7524 12628 7530 12640
rect 8573 12631 8631 12637
rect 8573 12628 8585 12631
rect 7524 12600 8585 12628
rect 7524 12588 7530 12600
rect 8573 12597 8585 12600
rect 8619 12597 8631 12631
rect 8573 12591 8631 12597
rect 8846 12588 8852 12640
rect 8904 12588 8910 12640
rect 8956 12628 8984 12727
rect 9232 12696 9260 12727
rect 9582 12724 9588 12776
rect 9640 12724 9646 12776
rect 9674 12774 9680 12804
rect 9732 12774 9738 12826
rect 9766 12792 9772 12844
rect 9824 12832 9830 12844
rect 10048 12835 10106 12841
rect 10048 12832 10060 12835
rect 9824 12804 10060 12832
rect 9824 12792 9830 12804
rect 10048 12801 10060 12804
rect 10094 12801 10106 12835
rect 10048 12795 10106 12801
rect 10321 12835 10379 12841
rect 10321 12801 10333 12835
rect 10367 12830 10379 12835
rect 10502 12830 10508 12844
rect 10367 12802 10508 12830
rect 10367 12801 10379 12802
rect 10321 12795 10379 12801
rect 10502 12792 10508 12802
rect 10560 12792 10566 12844
rect 11146 12832 11152 12844
rect 10704 12804 11152 12832
rect 9912 12767 9970 12773
rect 9912 12733 9924 12767
rect 9958 12764 9970 12767
rect 10704 12764 10732 12804
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 11514 12792 11520 12844
rect 11572 12832 11578 12844
rect 12084 12841 12112 12872
rect 13446 12860 13452 12872
rect 13504 12860 13510 12912
rect 12069 12835 12127 12841
rect 11572 12804 11836 12832
rect 11572 12792 11578 12804
rect 9958 12736 10732 12764
rect 9958 12733 9970 12736
rect 9912 12727 9970 12733
rect 10778 12724 10784 12776
rect 10836 12764 10842 12776
rect 10836 12736 11008 12764
rect 10836 12724 10842 12736
rect 10980 12696 11008 12736
rect 11330 12724 11336 12776
rect 11388 12764 11394 12776
rect 11388 12736 11655 12764
rect 11388 12724 11394 12736
rect 11627 12696 11655 12736
rect 11698 12724 11704 12776
rect 11756 12724 11762 12776
rect 11808 12773 11836 12804
rect 12069 12801 12081 12835
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 12618 12792 12624 12844
rect 12676 12832 12682 12844
rect 12676 12804 13216 12832
rect 12676 12792 12682 12804
rect 13188 12776 13216 12804
rect 13906 12792 13912 12844
rect 13964 12832 13970 12844
rect 14004 12835 14062 12841
rect 14004 12832 14016 12835
rect 13964 12804 14016 12832
rect 13964 12792 13970 12804
rect 14004 12801 14016 12804
rect 14050 12801 14062 12835
rect 14004 12795 14062 12801
rect 15194 12792 15200 12844
rect 15252 12832 15258 12844
rect 16212 12835 16270 12841
rect 16212 12832 16224 12835
rect 15252 12804 16224 12832
rect 15252 12792 15258 12804
rect 16212 12801 16224 12804
rect 16258 12801 16270 12835
rect 16212 12795 16270 12801
rect 16390 12792 16396 12844
rect 16448 12792 16454 12844
rect 16485 12835 16543 12841
rect 16485 12801 16497 12835
rect 16531 12832 16543 12835
rect 16666 12832 16672 12844
rect 16531 12804 16672 12832
rect 16531 12801 16543 12804
rect 16485 12795 16543 12801
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 16776 12804 18460 12832
rect 11793 12767 11851 12773
rect 11793 12733 11805 12767
rect 11839 12764 11851 12767
rect 12158 12764 12164 12776
rect 11839 12736 12164 12764
rect 11839 12733 11851 12736
rect 11793 12727 11851 12733
rect 12158 12724 12164 12736
rect 12216 12764 12222 12776
rect 12345 12767 12403 12773
rect 12345 12764 12357 12767
rect 12216 12736 12357 12764
rect 12216 12724 12222 12736
rect 12345 12733 12357 12736
rect 12391 12733 12403 12767
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12345 12727 12403 12733
rect 12544 12736 12817 12764
rect 12544 12708 12572 12736
rect 12805 12733 12817 12736
rect 12851 12733 12863 12767
rect 12805 12727 12863 12733
rect 12986 12724 12992 12776
rect 13044 12764 13050 12776
rect 13081 12767 13139 12773
rect 13081 12764 13093 12767
rect 13044 12736 13093 12764
rect 13044 12724 13050 12736
rect 13081 12733 13093 12736
rect 13127 12733 13139 12767
rect 13081 12727 13139 12733
rect 13170 12724 13176 12776
rect 13228 12724 13234 12776
rect 13354 12724 13360 12776
rect 13412 12724 13418 12776
rect 13538 12724 13544 12776
rect 13596 12724 13602 12776
rect 14277 12767 14335 12773
rect 14277 12764 14289 12767
rect 13648 12736 14289 12764
rect 12526 12696 12532 12708
rect 9232 12668 9444 12696
rect 10980 12668 11468 12696
rect 11627 12668 12532 12696
rect 9214 12628 9220 12640
rect 8956 12600 9220 12628
rect 9214 12588 9220 12600
rect 9272 12588 9278 12640
rect 9306 12588 9312 12640
rect 9364 12588 9370 12640
rect 9416 12628 9444 12668
rect 11330 12628 11336 12640
rect 9416 12600 11336 12628
rect 11330 12588 11336 12600
rect 11388 12588 11394 12640
rect 11440 12628 11468 12668
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 13648 12696 13676 12736
rect 14277 12733 14289 12736
rect 14323 12733 14335 12767
rect 14277 12727 14335 12733
rect 14642 12724 14648 12776
rect 14700 12764 14706 12776
rect 15102 12764 15108 12776
rect 14700 12736 15108 12764
rect 14700 12724 14706 12736
rect 15102 12724 15108 12736
rect 15160 12764 15166 12776
rect 15749 12767 15807 12773
rect 15749 12764 15761 12767
rect 15160 12736 15761 12764
rect 15160 12724 15166 12736
rect 15749 12733 15761 12736
rect 15795 12733 15807 12767
rect 16076 12767 16134 12773
rect 16076 12764 16088 12767
rect 15749 12727 15807 12733
rect 15856 12736 16088 12764
rect 12636 12668 13676 12696
rect 12636 12637 12664 12668
rect 15194 12656 15200 12708
rect 15252 12696 15258 12708
rect 15856 12696 15884 12736
rect 16076 12733 16088 12736
rect 16122 12764 16134 12767
rect 16408 12764 16436 12792
rect 16776 12776 16804 12804
rect 16122 12736 16436 12764
rect 16122 12733 16134 12736
rect 16076 12727 16134 12733
rect 16758 12724 16764 12776
rect 16816 12724 16822 12776
rect 18138 12724 18144 12776
rect 18196 12724 18202 12776
rect 18432 12773 18460 12804
rect 18598 12792 18604 12844
rect 18656 12792 18662 12844
rect 18708 12832 18736 12940
rect 18966 12928 18972 12940
rect 19024 12928 19030 12980
rect 20346 12928 20352 12980
rect 20404 12928 20410 12980
rect 22646 12928 22652 12980
rect 22704 12968 22710 12980
rect 23109 12971 23167 12977
rect 23109 12968 23121 12971
rect 22704 12940 23121 12968
rect 22704 12928 22710 12940
rect 23109 12937 23121 12940
rect 23155 12937 23167 12971
rect 23109 12931 23167 12937
rect 23566 12928 23572 12980
rect 23624 12968 23630 12980
rect 23842 12968 23848 12980
rect 23624 12940 23848 12968
rect 23624 12928 23630 12940
rect 23842 12928 23848 12940
rect 23900 12928 23906 12980
rect 24486 12928 24492 12980
rect 24544 12968 24550 12980
rect 25685 12971 25743 12977
rect 25685 12968 25697 12971
rect 24544 12940 25697 12968
rect 24544 12928 24550 12940
rect 25685 12937 25697 12940
rect 25731 12937 25743 12971
rect 25685 12931 25743 12937
rect 28721 12971 28779 12977
rect 28721 12937 28733 12971
rect 28767 12968 28779 12971
rect 28902 12968 28908 12980
rect 28767 12940 28908 12968
rect 28767 12937 28779 12940
rect 28721 12931 28779 12937
rect 28902 12928 28908 12940
rect 28960 12928 28966 12980
rect 29086 12928 29092 12980
rect 29144 12968 29150 12980
rect 29365 12971 29423 12977
rect 29365 12968 29377 12971
rect 29144 12940 29377 12968
rect 29144 12928 29150 12940
rect 29365 12937 29377 12940
rect 29411 12937 29423 12971
rect 29365 12931 29423 12937
rect 29454 12928 29460 12980
rect 29512 12928 29518 12980
rect 29638 12928 29644 12980
rect 29696 12928 29702 12980
rect 29822 12928 29828 12980
rect 29880 12968 29886 12980
rect 29917 12971 29975 12977
rect 29917 12968 29929 12971
rect 29880 12940 29929 12968
rect 29880 12928 29886 12940
rect 29917 12937 29929 12940
rect 29963 12937 29975 12971
rect 29917 12931 29975 12937
rect 19156 12835 19214 12841
rect 19156 12832 19168 12835
rect 18708 12804 19168 12832
rect 19156 12801 19168 12804
rect 19202 12801 19214 12835
rect 20364 12832 20392 12928
rect 29472 12900 29500 12928
rect 30193 12903 30251 12909
rect 30193 12900 30205 12903
rect 29472 12872 30205 12900
rect 30193 12869 30205 12872
rect 30239 12869 30251 12903
rect 30193 12863 30251 12869
rect 21364 12835 21422 12841
rect 21364 12832 21376 12835
rect 20364 12804 21376 12832
rect 19156 12795 19214 12801
rect 21364 12801 21376 12804
rect 21410 12801 21422 12835
rect 21364 12795 21422 12801
rect 22922 12792 22928 12844
rect 22980 12832 22986 12844
rect 24308 12835 24366 12841
rect 24308 12832 24320 12835
rect 22980 12804 24320 12832
rect 22980 12792 22986 12804
rect 24308 12801 24320 12804
rect 24354 12801 24366 12835
rect 24308 12795 24366 12801
rect 24946 12792 24952 12844
rect 25004 12832 25010 12844
rect 26602 12832 26608 12844
rect 25004 12804 26608 12832
rect 25004 12792 25010 12804
rect 26602 12792 26608 12804
rect 26660 12792 26666 12844
rect 31202 12832 31208 12844
rect 27172 12817 31208 12832
rect 18417 12767 18475 12773
rect 18417 12733 18429 12767
rect 18463 12733 18475 12767
rect 18616 12764 18644 12792
rect 27172 12786 27205 12817
rect 27193 12783 27205 12786
rect 27239 12804 31208 12817
rect 27239 12783 27251 12804
rect 31202 12792 31208 12804
rect 31260 12792 31266 12844
rect 27193 12777 27251 12783
rect 19058 12773 19064 12776
rect 18693 12767 18751 12773
rect 18693 12764 18705 12767
rect 18616 12736 18705 12764
rect 18417 12727 18475 12733
rect 18693 12733 18705 12736
rect 18739 12733 18751 12767
rect 18693 12727 18751 12733
rect 19020 12767 19064 12773
rect 19020 12733 19032 12767
rect 19020 12727 19064 12733
rect 15252 12668 15884 12696
rect 15252 12656 15258 12668
rect 11977 12631 12035 12637
rect 11977 12628 11989 12631
rect 11440 12600 11989 12628
rect 11977 12597 11989 12600
rect 12023 12597 12035 12631
rect 11977 12591 12035 12597
rect 12621 12631 12679 12637
rect 12621 12597 12633 12631
rect 12667 12597 12679 12631
rect 12621 12591 12679 12597
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13078 12628 13084 12640
rect 12943 12600 13084 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 13170 12588 13176 12640
rect 13228 12588 13234 12640
rect 13630 12588 13636 12640
rect 13688 12628 13694 12640
rect 14007 12631 14065 12637
rect 14007 12628 14019 12631
rect 13688 12600 14019 12628
rect 13688 12588 13694 12600
rect 14007 12597 14019 12600
rect 14053 12597 14065 12631
rect 14007 12591 14065 12597
rect 15102 12588 15108 12640
rect 15160 12628 15166 12640
rect 15381 12631 15439 12637
rect 15381 12628 15393 12631
rect 15160 12600 15393 12628
rect 15160 12588 15166 12600
rect 15381 12597 15393 12600
rect 15427 12597 15439 12631
rect 15381 12591 15439 12597
rect 17586 12588 17592 12640
rect 17644 12588 17650 12640
rect 17954 12588 17960 12640
rect 18012 12588 18018 12640
rect 18432 12628 18460 12727
rect 19058 12724 19064 12727
rect 19116 12724 19122 12776
rect 19426 12724 19432 12776
rect 19484 12724 19490 12776
rect 19518 12724 19524 12776
rect 19576 12764 19582 12776
rect 20714 12764 20720 12776
rect 19576 12736 20720 12764
rect 19576 12724 19582 12736
rect 20714 12724 20720 12736
rect 20772 12724 20778 12776
rect 20901 12767 20959 12773
rect 20901 12733 20913 12767
rect 20947 12764 20959 12767
rect 21266 12764 21272 12776
rect 20947 12736 21272 12764
rect 20947 12733 20959 12736
rect 20901 12727 20959 12733
rect 21266 12724 21272 12736
rect 21324 12724 21330 12776
rect 21634 12724 21640 12776
rect 21692 12724 21698 12776
rect 23014 12724 23020 12776
rect 23072 12764 23078 12776
rect 23293 12767 23351 12773
rect 23293 12764 23305 12767
rect 23072 12736 23305 12764
rect 23072 12724 23078 12736
rect 23293 12733 23305 12736
rect 23339 12764 23351 12767
rect 23474 12764 23480 12776
rect 23339 12736 23480 12764
rect 23339 12733 23351 12736
rect 23293 12727 23351 12733
rect 23474 12724 23480 12736
rect 23532 12724 23538 12776
rect 23569 12767 23627 12773
rect 23569 12733 23581 12767
rect 23615 12733 23627 12767
rect 23569 12727 23627 12733
rect 20806 12656 20812 12708
rect 20864 12656 20870 12708
rect 23584 12696 23612 12727
rect 23658 12724 23664 12776
rect 23716 12764 23722 12776
rect 23845 12767 23903 12773
rect 23845 12764 23857 12767
rect 23716 12736 23857 12764
rect 23716 12724 23722 12736
rect 23845 12733 23857 12736
rect 23891 12733 23903 12767
rect 24581 12767 24639 12773
rect 24581 12764 24593 12767
rect 23845 12727 23903 12733
rect 23971 12736 24593 12764
rect 23750 12696 23756 12708
rect 23584 12668 23756 12696
rect 23750 12656 23756 12668
rect 23808 12656 23814 12708
rect 20990 12628 20996 12640
rect 18432 12600 20996 12628
rect 20990 12588 20996 12600
rect 21048 12588 21054 12640
rect 21367 12631 21425 12637
rect 21367 12597 21379 12631
rect 21413 12628 21425 12631
rect 21726 12628 21732 12640
rect 21413 12600 21732 12628
rect 21413 12597 21425 12600
rect 21367 12591 21425 12597
rect 21726 12588 21732 12600
rect 21784 12588 21790 12640
rect 22738 12588 22744 12640
rect 22796 12588 22802 12640
rect 23385 12631 23443 12637
rect 23385 12597 23397 12631
rect 23431 12628 23443 12631
rect 23971 12628 23999 12736
rect 24581 12733 24593 12736
rect 24627 12733 24639 12767
rect 24581 12727 24639 12733
rect 24854 12724 24860 12776
rect 24912 12764 24918 12776
rect 26053 12767 26111 12773
rect 26053 12764 26065 12767
rect 24912 12736 26065 12764
rect 24912 12724 24918 12736
rect 26053 12733 26065 12736
rect 26099 12733 26111 12767
rect 26053 12727 26111 12733
rect 26510 12724 26516 12776
rect 26568 12764 26574 12776
rect 26697 12767 26755 12773
rect 26697 12764 26709 12767
rect 26568 12736 26709 12764
rect 26568 12724 26574 12736
rect 26697 12733 26709 12736
rect 26743 12733 26755 12767
rect 26697 12727 26755 12733
rect 27433 12767 27491 12773
rect 27433 12733 27445 12767
rect 27479 12764 27491 12767
rect 28442 12764 28448 12776
rect 27479 12736 28448 12764
rect 27479 12733 27491 12736
rect 27433 12727 27491 12733
rect 28442 12724 28448 12736
rect 28500 12724 28506 12776
rect 29178 12724 29184 12776
rect 29236 12764 29242 12776
rect 29549 12767 29607 12773
rect 29549 12764 29561 12767
rect 29236 12736 29561 12764
rect 29236 12724 29242 12736
rect 29549 12733 29561 12736
rect 29595 12764 29607 12767
rect 29825 12767 29883 12773
rect 29595 12736 29776 12764
rect 29595 12733 29607 12736
rect 29549 12727 29607 12733
rect 26329 12699 26387 12705
rect 26329 12665 26341 12699
rect 26375 12665 26387 12699
rect 26329 12659 26387 12665
rect 29089 12699 29147 12705
rect 29089 12665 29101 12699
rect 29135 12696 29147 12699
rect 29270 12696 29276 12708
rect 29135 12668 29276 12696
rect 29135 12665 29147 12668
rect 29089 12659 29147 12665
rect 23431 12600 23999 12628
rect 23431 12597 23443 12600
rect 23385 12591 23443 12597
rect 24118 12588 24124 12640
rect 24176 12628 24182 12640
rect 24311 12631 24369 12637
rect 24311 12628 24323 12631
rect 24176 12600 24323 12628
rect 24176 12588 24182 12600
rect 24311 12597 24323 12600
rect 24357 12628 24369 12631
rect 24670 12628 24676 12640
rect 24357 12600 24676 12628
rect 24357 12597 24369 12600
rect 24311 12591 24369 12597
rect 24670 12588 24676 12600
rect 24728 12628 24734 12640
rect 26344 12628 26372 12659
rect 29270 12656 29276 12668
rect 29328 12656 29334 12708
rect 26786 12628 26792 12640
rect 24728 12600 26792 12628
rect 24728 12588 24734 12600
rect 26786 12588 26792 12600
rect 26844 12628 26850 12640
rect 27163 12631 27221 12637
rect 27163 12628 27175 12631
rect 26844 12600 27175 12628
rect 26844 12588 26850 12600
rect 27163 12597 27175 12600
rect 27209 12628 27221 12631
rect 27798 12628 27804 12640
rect 27209 12600 27804 12628
rect 27209 12597 27221 12600
rect 27163 12591 27221 12597
rect 27798 12588 27804 12600
rect 27856 12588 27862 12640
rect 28994 12588 29000 12640
rect 29052 12628 29058 12640
rect 29181 12631 29239 12637
rect 29181 12628 29193 12631
rect 29052 12600 29193 12628
rect 29052 12588 29058 12600
rect 29181 12597 29193 12600
rect 29227 12597 29239 12631
rect 29748 12628 29776 12736
rect 29825 12733 29837 12767
rect 29871 12764 29883 12767
rect 29914 12764 29920 12776
rect 29871 12736 29920 12764
rect 29871 12733 29883 12736
rect 29825 12727 29883 12733
rect 29914 12724 29920 12736
rect 29972 12724 29978 12776
rect 30006 12724 30012 12776
rect 30064 12764 30070 12776
rect 30101 12767 30159 12773
rect 30101 12764 30113 12767
rect 30064 12736 30113 12764
rect 30064 12724 30070 12736
rect 30101 12733 30113 12736
rect 30147 12733 30159 12767
rect 30101 12727 30159 12733
rect 30377 12767 30435 12773
rect 30377 12733 30389 12767
rect 30423 12764 30435 12767
rect 30558 12764 30564 12776
rect 30423 12736 30564 12764
rect 30423 12733 30435 12736
rect 30377 12727 30435 12733
rect 30116 12696 30144 12727
rect 30558 12724 30564 12736
rect 30616 12764 30622 12776
rect 30616 12736 30788 12764
rect 30616 12724 30622 12736
rect 30650 12696 30656 12708
rect 30116 12668 30656 12696
rect 30650 12656 30656 12668
rect 30708 12656 30714 12708
rect 30760 12628 30788 12736
rect 29748 12600 30788 12628
rect 29181 12591 29239 12597
rect 552 12538 31072 12560
rect 552 12486 7988 12538
rect 8040 12486 8052 12538
rect 8104 12486 8116 12538
rect 8168 12486 8180 12538
rect 8232 12486 8244 12538
rect 8296 12486 15578 12538
rect 15630 12486 15642 12538
rect 15694 12486 15706 12538
rect 15758 12486 15770 12538
rect 15822 12486 15834 12538
rect 15886 12486 23168 12538
rect 23220 12486 23232 12538
rect 23284 12486 23296 12538
rect 23348 12486 23360 12538
rect 23412 12486 23424 12538
rect 23476 12486 30758 12538
rect 30810 12486 30822 12538
rect 30874 12486 30886 12538
rect 30938 12486 30950 12538
rect 31002 12486 31014 12538
rect 31066 12486 31072 12538
rect 552 12464 31072 12486
rect 1026 12384 1032 12436
rect 1084 12424 1090 12436
rect 2130 12424 2136 12436
rect 1084 12396 2136 12424
rect 1084 12384 1090 12396
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 5810 12384 5816 12436
rect 5868 12384 5874 12436
rect 6181 12427 6239 12433
rect 6181 12393 6193 12427
rect 6227 12393 6239 12427
rect 6181 12387 6239 12393
rect 6196 12356 6224 12387
rect 6270 12384 6276 12436
rect 6328 12424 6334 12436
rect 6822 12424 6828 12436
rect 6328 12396 6828 12424
rect 6328 12384 6334 12396
rect 6822 12384 6828 12396
rect 6880 12384 6886 12436
rect 6923 12427 6981 12433
rect 6923 12393 6935 12427
rect 6969 12424 6981 12427
rect 7098 12424 7104 12436
rect 6969 12396 7104 12424
rect 6969 12393 6981 12396
rect 6923 12387 6981 12393
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 8481 12427 8539 12433
rect 8481 12393 8493 12427
rect 8527 12424 8539 12427
rect 9766 12424 9772 12436
rect 8527 12396 9772 12424
rect 8527 12393 8539 12396
rect 8481 12387 8539 12393
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 11238 12384 11244 12436
rect 11296 12384 11302 12436
rect 11698 12384 11704 12436
rect 11756 12424 11762 12436
rect 11756 12396 12670 12424
rect 11756 12384 11762 12396
rect 6196 12328 6598 12356
rect 1210 12248 1216 12300
rect 1268 12248 1274 12300
rect 1670 12297 1676 12300
rect 1632 12291 1676 12297
rect 1632 12257 1644 12291
rect 1632 12251 1676 12257
rect 1670 12248 1676 12251
rect 1728 12248 1734 12300
rect 3421 12291 3479 12297
rect 3421 12257 3433 12291
rect 3467 12288 3479 12291
rect 4249 12291 4307 12297
rect 3467 12260 4019 12288
rect 3467 12257 3479 12260
rect 3421 12251 3479 12257
rect 1302 12180 1308 12232
rect 1360 12180 1366 12232
rect 1762 12220 1768 12232
rect 1726 12192 1768 12220
rect 1762 12180 1768 12192
rect 1820 12180 1826 12232
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12220 2099 12223
rect 2130 12220 2136 12232
rect 2087 12192 2136 12220
rect 2087 12189 2099 12192
rect 2041 12183 2099 12189
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 3510 12180 3516 12232
rect 3568 12180 3574 12232
rect 3878 12229 3884 12232
rect 3840 12223 3884 12229
rect 3840 12189 3852 12223
rect 3840 12183 3884 12189
rect 3878 12180 3884 12183
rect 3936 12180 3942 12232
rect 3991 12231 4019 12260
rect 4249 12257 4261 12291
rect 4295 12288 4307 12291
rect 4706 12288 4712 12300
rect 4295 12260 4712 12288
rect 4295 12257 4307 12260
rect 4249 12251 4307 12257
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 5997 12291 6055 12297
rect 5997 12288 6009 12291
rect 5592 12260 6009 12288
rect 5592 12248 5598 12260
rect 5997 12257 6009 12260
rect 6043 12288 6055 12291
rect 6365 12291 6423 12297
rect 6365 12288 6377 12291
rect 6043 12260 6377 12288
rect 6043 12257 6055 12260
rect 5997 12251 6055 12257
rect 6365 12257 6377 12260
rect 6411 12257 6423 12291
rect 6570 12288 6598 12328
rect 8570 12316 8576 12368
rect 8628 12356 8634 12368
rect 8628 12328 8800 12356
rect 8628 12316 8634 12328
rect 7193 12291 7251 12297
rect 7193 12288 7205 12291
rect 6570 12260 7205 12288
rect 6365 12251 6423 12257
rect 7193 12257 7205 12260
rect 7239 12257 7251 12291
rect 8772 12288 8800 12328
rect 11072 12328 11928 12356
rect 8772 12260 9171 12288
rect 7193 12251 7251 12257
rect 3976 12225 4034 12231
rect 3976 12191 3988 12225
rect 4022 12191 4034 12225
rect 3976 12185 4034 12191
rect 6457 12223 6515 12229
rect 6457 12189 6469 12223
rect 6503 12189 6515 12223
rect 6457 12183 6515 12189
rect 5994 12112 6000 12164
rect 6052 12152 6058 12164
rect 6472 12152 6500 12183
rect 6822 12180 6828 12232
rect 6880 12220 6886 12232
rect 6920 12223 6978 12229
rect 6920 12220 6932 12223
rect 6880 12192 6932 12220
rect 6880 12180 6886 12192
rect 6920 12189 6932 12192
rect 6966 12189 6978 12223
rect 6920 12183 6978 12189
rect 8665 12223 8723 12229
rect 8665 12189 8677 12223
rect 8711 12189 8723 12223
rect 8665 12183 8723 12189
rect 6052 12124 6500 12152
rect 6052 12112 6058 12124
rect 1029 12087 1087 12093
rect 1029 12053 1041 12087
rect 1075 12084 1087 12087
rect 2130 12084 2136 12096
rect 1075 12056 2136 12084
rect 1075 12053 1087 12056
rect 1029 12047 1087 12053
rect 2130 12044 2136 12056
rect 2188 12044 2194 12096
rect 5537 12087 5595 12093
rect 5537 12053 5549 12087
rect 5583 12084 5595 12087
rect 6730 12084 6736 12096
rect 5583 12056 6736 12084
rect 5583 12053 5595 12056
rect 5537 12047 5595 12053
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 7006 12044 7012 12096
rect 7064 12084 7070 12096
rect 8478 12084 8484 12096
rect 7064 12056 8484 12084
rect 7064 12044 7070 12056
rect 8478 12044 8484 12056
rect 8536 12044 8542 12096
rect 8680 12084 8708 12183
rect 8846 12180 8852 12232
rect 8904 12220 8910 12232
rect 9143 12231 9171 12260
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 9401 12291 9459 12297
rect 9401 12288 9413 12291
rect 9364 12260 9413 12288
rect 9364 12248 9370 12260
rect 9401 12257 9413 12260
rect 9447 12257 9459 12291
rect 11072 12292 11100 12328
rect 11149 12292 11207 12297
rect 11072 12291 11207 12292
rect 11072 12264 11161 12291
rect 9401 12251 9459 12257
rect 11149 12257 11161 12264
rect 11195 12257 11207 12291
rect 11149 12251 11207 12257
rect 11514 12248 11520 12300
rect 11572 12248 11578 12300
rect 11793 12291 11851 12297
rect 11793 12257 11805 12291
rect 11839 12257 11851 12291
rect 11900 12288 11928 12328
rect 12434 12288 12440 12300
rect 11900 12260 12440 12288
rect 11793 12251 11851 12257
rect 8992 12223 9050 12229
rect 8992 12220 9004 12223
rect 8904 12192 9004 12220
rect 8904 12180 8910 12192
rect 8992 12189 9004 12192
rect 9038 12189 9050 12223
rect 8992 12183 9050 12189
rect 9128 12225 9186 12231
rect 9128 12191 9140 12225
rect 9174 12191 9186 12225
rect 9128 12185 9186 12191
rect 10778 12180 10784 12232
rect 10836 12220 10842 12232
rect 11808 12220 11836 12251
rect 12434 12248 12440 12260
rect 12492 12248 12498 12300
rect 12642 12288 12670 12396
rect 12802 12384 12808 12436
rect 12860 12424 12866 12436
rect 12995 12427 13053 12433
rect 12995 12424 13007 12427
rect 12860 12396 13007 12424
rect 12860 12384 12866 12396
rect 12995 12393 13007 12396
rect 13041 12424 13053 12427
rect 13630 12424 13636 12436
rect 13041 12396 13636 12424
rect 13041 12393 13053 12396
rect 12995 12387 13053 12393
rect 13630 12384 13636 12396
rect 13688 12424 13694 12436
rect 13688 12396 13952 12424
rect 13688 12384 13694 12396
rect 13924 12356 13952 12396
rect 14274 12384 14280 12436
rect 14332 12424 14338 12436
rect 15289 12427 15347 12433
rect 15289 12424 15301 12427
rect 14332 12396 15301 12424
rect 14332 12384 14338 12396
rect 15289 12393 15301 12396
rect 15335 12393 15347 12427
rect 15289 12387 15347 12393
rect 16114 12384 16120 12436
rect 16172 12384 16178 12436
rect 17218 12384 17224 12436
rect 17276 12424 17282 12436
rect 17411 12427 17469 12433
rect 17411 12424 17423 12427
rect 17276 12396 17423 12424
rect 17276 12384 17282 12396
rect 17411 12393 17423 12396
rect 17457 12393 17469 12427
rect 17411 12387 17469 12393
rect 18782 12384 18788 12436
rect 18840 12384 18846 12436
rect 19444 12396 19656 12424
rect 15013 12359 15071 12365
rect 15013 12356 15025 12359
rect 13924 12328 15025 12356
rect 15013 12325 15025 12328
rect 15059 12325 15071 12359
rect 15013 12319 15071 12325
rect 18874 12316 18880 12368
rect 18932 12356 18938 12368
rect 19444 12356 19472 12396
rect 18932 12328 19472 12356
rect 19628 12356 19656 12396
rect 19702 12384 19708 12436
rect 19760 12384 19766 12436
rect 20349 12427 20407 12433
rect 20349 12393 20361 12427
rect 20395 12393 20407 12427
rect 20349 12387 20407 12393
rect 20901 12427 20959 12433
rect 20901 12393 20913 12427
rect 20947 12424 20959 12427
rect 21634 12424 21640 12436
rect 20947 12396 21640 12424
rect 20947 12393 20959 12396
rect 20901 12387 20959 12393
rect 20364 12356 20392 12387
rect 21634 12384 21640 12396
rect 21692 12384 21698 12436
rect 21726 12384 21732 12436
rect 21784 12433 21790 12436
rect 21784 12424 21793 12433
rect 21910 12424 21916 12436
rect 21784 12396 21916 12424
rect 21784 12387 21793 12396
rect 21784 12384 21790 12387
rect 21910 12384 21916 12396
rect 21968 12384 21974 12436
rect 22462 12384 22468 12436
rect 22520 12424 22526 12436
rect 23109 12427 23167 12433
rect 23109 12424 23121 12427
rect 22520 12396 23121 12424
rect 22520 12384 22526 12396
rect 23109 12393 23121 12396
rect 23155 12393 23167 12427
rect 23109 12387 23167 12393
rect 23943 12427 24001 12433
rect 23943 12393 23955 12427
rect 23989 12424 24001 12427
rect 24118 12424 24124 12436
rect 23989 12396 24124 12424
rect 23989 12393 24001 12396
rect 23943 12387 24001 12393
rect 24118 12384 24124 12396
rect 24176 12384 24182 12436
rect 24578 12384 24584 12436
rect 24636 12424 24642 12436
rect 25317 12427 25375 12433
rect 25317 12424 25329 12427
rect 24636 12396 25329 12424
rect 24636 12384 24642 12396
rect 25317 12393 25329 12396
rect 25363 12393 25375 12427
rect 25317 12387 25375 12393
rect 26786 12384 26792 12436
rect 26844 12424 26850 12436
rect 26887 12427 26945 12433
rect 26887 12424 26899 12427
rect 26844 12396 26899 12424
rect 26844 12384 26850 12396
rect 26887 12393 26899 12396
rect 26933 12393 26945 12427
rect 26887 12387 26945 12393
rect 28258 12384 28264 12436
rect 28316 12384 28322 12436
rect 30190 12384 30196 12436
rect 30248 12424 30254 12436
rect 30561 12427 30619 12433
rect 30561 12424 30573 12427
rect 30248 12396 30573 12424
rect 30248 12384 30254 12396
rect 30561 12393 30573 12396
rect 30607 12393 30619 12427
rect 30561 12387 30619 12393
rect 19628 12328 20300 12356
rect 20364 12328 21220 12356
rect 18932 12316 18938 12328
rect 12642 12260 12940 12288
rect 12912 12238 12940 12260
rect 13170 12248 13176 12300
rect 13228 12288 13234 12300
rect 13265 12291 13323 12297
rect 13265 12288 13277 12291
rect 13228 12260 13277 12288
rect 13228 12248 13234 12260
rect 13265 12257 13277 12260
rect 13311 12257 13323 12291
rect 13265 12251 13323 12257
rect 13998 12248 14004 12300
rect 14056 12288 14062 12300
rect 14737 12291 14795 12297
rect 14737 12288 14749 12291
rect 14056 12260 14749 12288
rect 14056 12248 14062 12260
rect 14737 12257 14749 12260
rect 14783 12257 14795 12291
rect 15473 12291 15531 12297
rect 15473 12288 15485 12291
rect 14737 12251 14795 12257
rect 14844 12260 15485 12288
rect 12992 12241 13050 12247
rect 12992 12238 13004 12241
rect 10836 12192 11836 12220
rect 12529 12223 12587 12229
rect 10836 12180 10842 12192
rect 12529 12189 12541 12223
rect 12575 12220 12587 12223
rect 12710 12220 12716 12232
rect 12575 12192 12716 12220
rect 12575 12189 12587 12192
rect 12529 12183 12587 12189
rect 12710 12180 12716 12192
rect 12768 12180 12774 12232
rect 12912 12210 13004 12238
rect 12992 12207 13004 12210
rect 13038 12207 13050 12241
rect 12992 12201 13050 12207
rect 13446 12180 13452 12232
rect 13504 12220 13510 12232
rect 13504 12192 14234 12220
rect 13504 12180 13510 12192
rect 10318 12112 10324 12164
rect 10376 12152 10382 12164
rect 11977 12155 12035 12161
rect 11977 12152 11989 12155
rect 10376 12124 11989 12152
rect 10376 12112 10382 12124
rect 11977 12121 11989 12124
rect 12023 12121 12035 12155
rect 14206 12152 14234 12192
rect 14274 12180 14280 12232
rect 14332 12220 14338 12232
rect 14844 12220 14872 12260
rect 15473 12257 15485 12260
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12257 15807 12291
rect 15749 12251 15807 12257
rect 16301 12291 16359 12297
rect 16301 12257 16313 12291
rect 16347 12288 16359 12291
rect 16853 12291 16911 12297
rect 16853 12288 16865 12291
rect 16347 12260 16865 12288
rect 16347 12257 16359 12260
rect 16301 12251 16359 12257
rect 16853 12257 16865 12260
rect 16899 12288 16911 12291
rect 17681 12291 17739 12297
rect 16899 12260 17632 12288
rect 16899 12257 16911 12260
rect 16853 12251 16911 12257
rect 14332 12192 14872 12220
rect 14332 12180 14338 12192
rect 15764 12152 15792 12251
rect 16945 12223 17003 12229
rect 16945 12220 16957 12223
rect 14206 12124 15792 12152
rect 16776 12192 16957 12220
rect 11977 12115 12035 12121
rect 16776 12096 16804 12192
rect 16945 12189 16957 12192
rect 16991 12189 17003 12223
rect 16945 12183 17003 12189
rect 17408 12225 17466 12231
rect 17408 12191 17420 12225
rect 17454 12220 17466 12225
rect 17494 12220 17500 12232
rect 17454 12192 17500 12220
rect 17454 12191 17466 12192
rect 17408 12185 17466 12191
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 17604 12220 17632 12260
rect 17681 12257 17693 12291
rect 17727 12288 17739 12291
rect 17954 12288 17960 12300
rect 17727 12260 17960 12288
rect 17727 12257 17739 12260
rect 17681 12251 17739 12257
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 18046 12248 18052 12300
rect 18104 12288 18110 12300
rect 19337 12291 19395 12297
rect 19337 12288 19349 12291
rect 18104 12260 19349 12288
rect 18104 12248 18110 12260
rect 19337 12257 19349 12260
rect 19383 12288 19395 12291
rect 19518 12288 19524 12324
rect 19383 12272 19524 12288
rect 19576 12272 19582 12324
rect 19613 12291 19671 12297
rect 19383 12260 19564 12272
rect 19383 12257 19395 12260
rect 19337 12251 19395 12257
rect 19613 12257 19625 12291
rect 19659 12288 19671 12291
rect 19794 12288 19800 12300
rect 19659 12260 19800 12288
rect 19659 12257 19671 12260
rect 19613 12251 19671 12257
rect 19628 12222 19656 12251
rect 19794 12248 19800 12260
rect 19852 12248 19858 12300
rect 19889 12291 19947 12297
rect 19889 12257 19901 12291
rect 19935 12288 19947 12291
rect 20162 12288 20168 12300
rect 19935 12260 20168 12288
rect 19935 12257 19947 12260
rect 19889 12251 19947 12257
rect 20162 12248 20168 12260
rect 20220 12248 20226 12300
rect 20272 12288 20300 12328
rect 20533 12291 20591 12297
rect 20533 12288 20545 12291
rect 20272 12260 20545 12288
rect 20533 12257 20545 12260
rect 20579 12257 20591 12291
rect 20533 12251 20591 12257
rect 20622 12248 20628 12300
rect 20680 12288 20686 12300
rect 20809 12291 20867 12297
rect 20809 12288 20821 12291
rect 20680 12260 20821 12288
rect 20680 12248 20686 12260
rect 20809 12257 20821 12260
rect 20855 12257 20867 12291
rect 20809 12251 20867 12257
rect 21082 12248 21088 12300
rect 21140 12248 21146 12300
rect 19260 12220 19380 12222
rect 19444 12220 19656 12222
rect 17604 12194 19656 12220
rect 21192 12220 21220 12328
rect 22738 12316 22744 12368
rect 22796 12316 22802 12368
rect 26145 12359 26203 12365
rect 26145 12325 26157 12359
rect 26191 12356 26203 12359
rect 26418 12356 26424 12368
rect 26191 12328 26424 12356
rect 26191 12325 26203 12328
rect 26145 12319 26203 12325
rect 26418 12316 26424 12328
rect 26476 12316 26482 12368
rect 29914 12316 29920 12368
rect 29972 12356 29978 12368
rect 29972 12328 30420 12356
rect 29972 12316 29978 12328
rect 21266 12248 21272 12300
rect 21324 12248 21330 12300
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 21422 12260 22017 12288
rect 21422 12220 21450 12260
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 22756 12288 22784 12316
rect 22756 12260 23796 12288
rect 22005 12251 22063 12257
rect 17604 12192 19288 12194
rect 19352 12192 19472 12194
rect 21192 12192 21450 12220
rect 21726 12180 21732 12232
rect 21784 12180 21790 12232
rect 23477 12223 23535 12229
rect 23477 12189 23489 12223
rect 23523 12220 23535 12223
rect 23658 12220 23664 12232
rect 23523 12192 23664 12220
rect 23523 12189 23535 12192
rect 23477 12183 23535 12189
rect 19242 12112 19248 12164
rect 19300 12152 19306 12164
rect 20530 12152 20536 12164
rect 19300 12124 20536 12152
rect 19300 12112 19306 12124
rect 20530 12112 20536 12124
rect 20588 12112 20594 12164
rect 20625 12155 20683 12161
rect 20625 12121 20637 12155
rect 20671 12152 20683 12155
rect 20671 12124 21312 12152
rect 20671 12121 20683 12124
rect 20625 12115 20683 12121
rect 9306 12084 9312 12096
rect 8680 12056 9312 12084
rect 9306 12044 9312 12056
rect 9364 12084 9370 12096
rect 9582 12084 9588 12096
rect 9364 12056 9588 12084
rect 9364 12044 9370 12056
rect 9582 12044 9588 12056
rect 9640 12044 9646 12096
rect 10686 12044 10692 12096
rect 10744 12044 10750 12096
rect 10962 12044 10968 12096
rect 11020 12044 11026 12096
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 11701 12087 11759 12093
rect 11701 12084 11713 12087
rect 11112 12056 11713 12084
rect 11112 12044 11118 12056
rect 11701 12053 11713 12056
rect 11747 12053 11759 12087
rect 11701 12047 11759 12053
rect 12253 12087 12311 12093
rect 12253 12053 12265 12087
rect 12299 12084 12311 12087
rect 13262 12084 13268 12096
rect 12299 12056 13268 12084
rect 12299 12053 12311 12056
rect 12253 12047 12311 12053
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 14550 12044 14556 12096
rect 14608 12044 14614 12096
rect 15562 12044 15568 12096
rect 15620 12044 15626 12096
rect 16666 12044 16672 12096
rect 16724 12044 16730 12096
rect 16758 12044 16764 12096
rect 16816 12044 16822 12096
rect 17494 12044 17500 12096
rect 17552 12084 17558 12096
rect 18414 12084 18420 12096
rect 17552 12056 18420 12084
rect 17552 12044 17558 12056
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 19058 12044 19064 12096
rect 19116 12084 19122 12096
rect 19153 12087 19211 12093
rect 19153 12084 19165 12087
rect 19116 12056 19165 12084
rect 19116 12044 19122 12056
rect 19153 12053 19165 12056
rect 19199 12053 19211 12087
rect 19153 12047 19211 12053
rect 19426 12044 19432 12096
rect 19484 12044 19490 12096
rect 21284 12084 21312 12124
rect 21450 12084 21456 12096
rect 21284 12056 21456 12084
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 22370 12044 22376 12096
rect 22428 12084 22434 12096
rect 23290 12084 23296 12096
rect 22428 12056 23296 12084
rect 22428 12044 22434 12056
rect 23290 12044 23296 12056
rect 23348 12044 23354 12096
rect 23492 12084 23520 12183
rect 23658 12180 23664 12192
rect 23716 12180 23722 12232
rect 23768 12220 23796 12260
rect 24210 12248 24216 12300
rect 24268 12248 24274 12300
rect 25777 12291 25835 12297
rect 25777 12288 25789 12291
rect 25424 12260 25789 12288
rect 23940 12223 23998 12229
rect 23940 12220 23952 12223
rect 23768 12192 23952 12220
rect 23940 12189 23952 12192
rect 23986 12189 23998 12223
rect 23940 12183 23998 12189
rect 24210 12084 24216 12096
rect 23492 12056 24216 12084
rect 24210 12044 24216 12056
rect 24268 12084 24274 12096
rect 25424 12084 25452 12260
rect 25777 12257 25789 12260
rect 25823 12288 25835 12291
rect 26510 12288 26516 12300
rect 25823 12260 26516 12288
rect 25823 12257 25835 12260
rect 25777 12251 25835 12257
rect 26436 12229 26464 12260
rect 26510 12248 26516 12260
rect 26568 12288 26574 12300
rect 28074 12288 28080 12300
rect 26568 12260 28080 12288
rect 26568 12248 26574 12260
rect 28074 12248 28080 12260
rect 28132 12248 28138 12300
rect 28902 12248 28908 12300
rect 28960 12248 28966 12300
rect 30392 12297 30420 12328
rect 30377 12291 30435 12297
rect 30377 12257 30389 12291
rect 30423 12257 30435 12291
rect 30377 12251 30435 12257
rect 26421 12223 26479 12229
rect 26421 12189 26433 12223
rect 26467 12189 26479 12223
rect 26421 12183 26479 12189
rect 26878 12180 26884 12232
rect 26936 12220 26942 12232
rect 27157 12223 27215 12229
rect 26936 12192 26981 12220
rect 26936 12180 26942 12192
rect 27157 12189 27169 12223
rect 27203 12220 27215 12223
rect 27798 12220 27804 12232
rect 27203 12192 27804 12220
rect 27203 12189 27215 12192
rect 27157 12183 27215 12189
rect 27798 12180 27804 12192
rect 27856 12180 27862 12232
rect 28626 12180 28632 12232
rect 28684 12180 28690 12232
rect 24268 12056 25452 12084
rect 24268 12044 24274 12056
rect 25498 12044 25504 12096
rect 25556 12084 25562 12096
rect 30009 12087 30067 12093
rect 30009 12084 30021 12087
rect 25556 12056 30021 12084
rect 25556 12044 25562 12056
rect 30009 12053 30021 12056
rect 30055 12053 30067 12087
rect 30009 12047 30067 12053
rect 552 11994 30912 12016
rect 552 11942 4193 11994
rect 4245 11942 4257 11994
rect 4309 11942 4321 11994
rect 4373 11942 4385 11994
rect 4437 11942 4449 11994
rect 4501 11942 11783 11994
rect 11835 11942 11847 11994
rect 11899 11942 11911 11994
rect 11963 11942 11975 11994
rect 12027 11942 12039 11994
rect 12091 11942 19373 11994
rect 19425 11942 19437 11994
rect 19489 11942 19501 11994
rect 19553 11942 19565 11994
rect 19617 11942 19629 11994
rect 19681 11942 26963 11994
rect 27015 11942 27027 11994
rect 27079 11942 27091 11994
rect 27143 11942 27155 11994
rect 27207 11942 27219 11994
rect 27271 11942 30912 11994
rect 552 11920 30912 11942
rect 2774 11840 2780 11892
rect 2832 11840 2838 11892
rect 5813 11883 5871 11889
rect 3160 11852 5212 11880
rect 1443 11747 1501 11753
rect 1443 11713 1455 11747
rect 1489 11744 1501 11747
rect 3160 11744 3188 11852
rect 3237 11815 3295 11821
rect 3237 11781 3249 11815
rect 3283 11812 3295 11815
rect 3694 11812 3700 11824
rect 3283 11784 3700 11812
rect 3283 11781 3295 11784
rect 3237 11775 3295 11781
rect 3694 11772 3700 11784
rect 3752 11772 3758 11824
rect 5184 11812 5212 11852
rect 5813 11849 5825 11883
rect 5859 11880 5871 11883
rect 7282 11880 7288 11892
rect 5859 11852 7288 11880
rect 5859 11849 5871 11852
rect 5813 11843 5871 11849
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 10134 11880 10140 11892
rect 7944 11852 10140 11880
rect 5184 11784 5856 11812
rect 3510 11744 3516 11756
rect 1489 11716 3188 11744
rect 3344 11716 3516 11744
rect 1489 11713 1501 11716
rect 1443 11707 1501 11713
rect 934 11636 940 11688
rect 992 11676 998 11688
rect 1210 11676 1216 11688
rect 992 11648 1216 11676
rect 992 11636 998 11648
rect 1210 11636 1216 11648
rect 1268 11636 1274 11688
rect 1670 11636 1676 11688
rect 1728 11636 1734 11688
rect 1394 11500 1400 11552
rect 1452 11549 1458 11552
rect 1452 11540 1461 11549
rect 1452 11512 1497 11540
rect 1452 11503 1461 11512
rect 1452 11500 1458 11503
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 2958 11540 2964 11552
rect 1636 11512 2964 11540
rect 1636 11500 1642 11512
rect 2958 11500 2964 11512
rect 3016 11540 3022 11552
rect 3344 11540 3372 11716
rect 3510 11704 3516 11716
rect 3568 11744 3574 11756
rect 3789 11747 3847 11753
rect 3789 11744 3801 11747
rect 3568 11716 3801 11744
rect 3568 11704 3574 11716
rect 3789 11713 3801 11716
rect 3835 11713 3847 11747
rect 3789 11707 3847 11713
rect 4246 11704 4252 11756
rect 4304 11744 4310 11756
rect 4525 11747 4583 11753
rect 4304 11716 4349 11744
rect 4304 11704 4310 11716
rect 4525 11713 4537 11747
rect 4571 11744 4583 11747
rect 5442 11744 5448 11756
rect 4571 11716 5448 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11645 3479 11679
rect 3421 11639 3479 11645
rect 3697 11679 3755 11685
rect 3697 11645 3709 11679
rect 3743 11676 3755 11679
rect 4154 11676 4160 11688
rect 3743 11648 4160 11676
rect 3743 11645 3755 11648
rect 3697 11639 3755 11645
rect 3436 11552 3464 11639
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 5166 11636 5172 11688
rect 5224 11636 5230 11688
rect 3016 11512 3372 11540
rect 3016 11500 3022 11512
rect 3418 11500 3424 11552
rect 3476 11500 3482 11552
rect 3510 11500 3516 11552
rect 3568 11500 3574 11552
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 4255 11543 4313 11549
rect 4255 11540 4267 11543
rect 4120 11512 4267 11540
rect 4120 11500 4126 11512
rect 4255 11509 4267 11512
rect 4301 11509 4313 11543
rect 4255 11503 4313 11509
rect 4522 11500 4528 11552
rect 4580 11540 4586 11552
rect 5184 11540 5212 11636
rect 5828 11608 5856 11784
rect 5902 11704 5908 11756
rect 5960 11744 5966 11756
rect 6552 11747 6610 11753
rect 6552 11744 6564 11747
rect 5960 11716 6564 11744
rect 5960 11704 5966 11716
rect 6552 11713 6564 11716
rect 6598 11713 6610 11747
rect 6552 11707 6610 11713
rect 6825 11747 6883 11753
rect 6825 11713 6837 11747
rect 6871 11744 6883 11747
rect 7834 11744 7840 11756
rect 6871 11716 7840 11744
rect 6871 11713 6883 11716
rect 6825 11707 6883 11713
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 5994 11636 6000 11688
rect 6052 11676 6058 11688
rect 6089 11679 6147 11685
rect 6089 11676 6101 11679
rect 6052 11648 6101 11676
rect 6052 11636 6058 11648
rect 6089 11645 6101 11648
rect 6135 11645 6147 11679
rect 7944 11676 7972 11852
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 10686 11840 10692 11892
rect 10744 11880 10750 11892
rect 10744 11852 12670 11880
rect 10744 11840 10750 11852
rect 11606 11772 11612 11824
rect 11664 11812 11670 11824
rect 12069 11815 12127 11821
rect 12069 11812 12081 11815
rect 11664 11784 12081 11812
rect 11664 11772 11670 11784
rect 12069 11781 12081 11784
rect 12115 11781 12127 11815
rect 12069 11775 12127 11781
rect 12158 11772 12164 11824
rect 12216 11772 12222 11824
rect 12526 11812 12532 11824
rect 12366 11784 12532 11812
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11744 8723 11747
rect 9030 11744 9036 11756
rect 8711 11716 9036 11744
rect 8711 11713 8723 11716
rect 8665 11707 8723 11713
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 9548 11716 9812 11744
rect 9548 11704 9554 11716
rect 8573 11679 8631 11685
rect 8573 11676 8585 11679
rect 6089 11639 6147 11645
rect 6196 11648 7972 11676
rect 8036 11648 8585 11676
rect 6196 11608 6224 11648
rect 5828 11580 6224 11608
rect 7834 11568 7840 11620
rect 7892 11608 7898 11620
rect 8036 11608 8064 11648
rect 8573 11645 8585 11648
rect 8619 11645 8631 11679
rect 9585 11679 9643 11685
rect 9585 11676 9597 11679
rect 8573 11639 8631 11645
rect 9416 11648 9597 11676
rect 7892 11580 8064 11608
rect 8205 11611 8263 11617
rect 7892 11568 7898 11580
rect 8205 11577 8217 11611
rect 8251 11608 8263 11611
rect 8478 11608 8484 11620
rect 8251 11580 8484 11608
rect 8251 11577 8263 11580
rect 8205 11571 8263 11577
rect 8478 11568 8484 11580
rect 8536 11568 8542 11620
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 9125 11611 9183 11617
rect 9125 11608 9137 11611
rect 8996 11580 9137 11608
rect 8996 11568 9002 11580
rect 9125 11577 9137 11580
rect 9171 11577 9183 11611
rect 9125 11571 9183 11577
rect 4580 11512 5212 11540
rect 4580 11500 4586 11512
rect 6454 11500 6460 11552
rect 6512 11540 6518 11552
rect 6555 11543 6613 11549
rect 6555 11540 6567 11543
rect 6512 11512 6567 11540
rect 6512 11500 6518 11512
rect 6555 11509 6567 11512
rect 6601 11509 6613 11543
rect 6555 11503 6613 11509
rect 6914 11500 6920 11552
rect 6972 11540 6978 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 6972 11512 8401 11540
rect 6972 11500 6978 11512
rect 8389 11509 8401 11512
rect 8435 11509 8447 11543
rect 8389 11503 8447 11509
rect 9306 11500 9312 11552
rect 9364 11540 9370 11552
rect 9416 11549 9444 11648
rect 9585 11645 9597 11648
rect 9631 11645 9643 11679
rect 9784 11676 9812 11716
rect 9858 11704 9864 11756
rect 9916 11744 9922 11756
rect 10048 11747 10106 11753
rect 10048 11744 10060 11747
rect 9916 11716 10060 11744
rect 9916 11704 9922 11716
rect 10048 11713 10060 11716
rect 10094 11713 10106 11747
rect 10048 11707 10106 11713
rect 10226 11704 10232 11756
rect 10284 11744 10290 11756
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 10284 11716 10333 11744
rect 10284 11704 10290 11716
rect 10321 11713 10333 11716
rect 10367 11713 10379 11747
rect 11793 11747 11851 11753
rect 11793 11744 11805 11747
rect 10321 11707 10379 11713
rect 10428 11716 11805 11744
rect 10428 11676 10456 11716
rect 11793 11713 11805 11716
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 9784 11648 10456 11676
rect 9585 11639 9643 11645
rect 11146 11636 11152 11688
rect 11204 11636 11210 11688
rect 12176 11676 12204 11772
rect 12253 11679 12311 11685
rect 12253 11676 12265 11679
rect 12176 11648 12265 11676
rect 12253 11645 12265 11648
rect 12299 11645 12311 11679
rect 12366 11676 12394 11784
rect 12526 11772 12532 11784
rect 12584 11772 12590 11824
rect 12642 11812 12670 11852
rect 12710 11840 12716 11892
rect 12768 11880 12774 11892
rect 13262 11880 13268 11892
rect 12768 11852 13268 11880
rect 12768 11840 12774 11852
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 13872 11852 15884 11880
rect 13872 11840 13878 11852
rect 12642 11784 12756 11812
rect 12728 11744 12756 11784
rect 12986 11772 12992 11824
rect 13044 11812 13050 11824
rect 13357 11815 13415 11821
rect 13357 11812 13369 11815
rect 13044 11784 13369 11812
rect 13044 11772 13050 11784
rect 13357 11781 13369 11784
rect 13403 11812 13415 11815
rect 13446 11812 13452 11824
rect 13403 11784 13452 11812
rect 13403 11781 13415 11784
rect 13357 11775 13415 11781
rect 13446 11772 13452 11784
rect 13504 11772 13510 11824
rect 15856 11812 15884 11852
rect 15930 11840 15936 11892
rect 15988 11840 15994 11892
rect 17954 11880 17960 11892
rect 16040 11852 17960 11880
rect 16040 11812 16068 11852
rect 17954 11840 17960 11852
rect 18012 11840 18018 11892
rect 19794 11880 19800 11892
rect 18064 11852 19800 11880
rect 15856 11784 16068 11812
rect 16117 11815 16175 11821
rect 12728 11735 14047 11744
rect 12728 11729 14062 11735
rect 12728 11716 14016 11729
rect 14004 11695 14016 11716
rect 14050 11695 14062 11729
rect 14004 11689 14062 11695
rect 12529 11679 12587 11685
rect 12366 11672 12488 11676
rect 12529 11672 12541 11679
rect 12366 11648 12541 11672
rect 12253 11639 12311 11645
rect 12460 11645 12541 11648
rect 12575 11645 12587 11679
rect 12460 11644 12587 11645
rect 12529 11639 12587 11644
rect 12989 11679 13047 11685
rect 12989 11645 13001 11679
rect 13035 11645 13047 11679
rect 12989 11639 13047 11645
rect 9401 11543 9459 11549
rect 9401 11540 9413 11543
rect 9364 11512 9413 11540
rect 9364 11500 9370 11512
rect 9401 11509 9413 11512
rect 9447 11509 9459 11543
rect 9401 11503 9459 11509
rect 9950 11500 9956 11552
rect 10008 11540 10014 11552
rect 10051 11543 10109 11549
rect 10051 11540 10063 11543
rect 10008 11512 10063 11540
rect 10008 11500 10014 11512
rect 10051 11509 10063 11512
rect 10097 11540 10109 11543
rect 11164 11540 11192 11636
rect 11698 11568 11704 11620
rect 11756 11608 11762 11620
rect 13004 11608 13032 11639
rect 13170 11636 13176 11688
rect 13228 11636 13234 11688
rect 13262 11636 13268 11688
rect 13320 11676 13326 11688
rect 13538 11676 13544 11688
rect 13320 11648 13544 11676
rect 13320 11636 13326 11648
rect 13538 11636 13544 11648
rect 13596 11636 13602 11688
rect 14090 11636 14096 11688
rect 14148 11676 14154 11688
rect 14277 11679 14335 11685
rect 14277 11676 14289 11679
rect 14148 11648 14289 11676
rect 14148 11636 14154 11648
rect 14277 11645 14289 11648
rect 14323 11645 14335 11679
rect 15856 11676 15884 11784
rect 16117 11781 16129 11815
rect 16163 11781 16175 11815
rect 16117 11775 16175 11781
rect 16132 11744 16160 11775
rect 16899 11747 16957 11753
rect 16132 11716 16626 11744
rect 16301 11679 16359 11685
rect 16301 11676 16313 11679
rect 15856 11648 16313 11676
rect 14277 11639 14335 11645
rect 16301 11645 16313 11648
rect 16347 11645 16359 11679
rect 16301 11639 16359 11645
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11645 16451 11679
rect 16598 11676 16626 11716
rect 16899 11713 16911 11747
rect 16945 11744 16957 11747
rect 18064 11744 18092 11852
rect 19794 11840 19800 11852
rect 19852 11840 19858 11892
rect 20717 11883 20775 11889
rect 20717 11849 20729 11883
rect 20763 11880 20775 11883
rect 21726 11880 21732 11892
rect 20763 11852 21732 11880
rect 20763 11849 20775 11852
rect 20717 11843 20775 11849
rect 21726 11840 21732 11852
rect 21784 11840 21790 11892
rect 22922 11840 22928 11892
rect 22980 11840 22986 11892
rect 23290 11840 23296 11892
rect 23348 11880 23354 11892
rect 23934 11880 23940 11892
rect 23348 11852 23940 11880
rect 23348 11840 23354 11852
rect 23934 11840 23940 11852
rect 23992 11840 23998 11892
rect 26237 11883 26295 11889
rect 26237 11849 26249 11883
rect 26283 11880 26295 11883
rect 26786 11880 26792 11892
rect 26283 11852 26792 11880
rect 26283 11849 26295 11852
rect 26237 11843 26295 11849
rect 26786 11840 26792 11852
rect 26844 11840 26850 11892
rect 26878 11840 26884 11892
rect 26936 11880 26942 11892
rect 28261 11883 28319 11889
rect 28261 11880 28273 11883
rect 26936 11852 28273 11880
rect 26936 11840 26942 11852
rect 28261 11849 28273 11852
rect 28307 11849 28319 11883
rect 28261 11843 28319 11849
rect 28442 11840 28448 11892
rect 28500 11840 28506 11892
rect 28629 11883 28687 11889
rect 28629 11849 28641 11883
rect 28675 11880 28687 11883
rect 28810 11880 28816 11892
rect 28675 11852 28816 11880
rect 28675 11849 28687 11852
rect 28629 11843 28687 11849
rect 28810 11840 28816 11852
rect 28868 11840 28874 11892
rect 30282 11840 30288 11892
rect 30340 11840 30346 11892
rect 23201 11815 23259 11821
rect 23201 11781 23213 11815
rect 23247 11812 23259 11815
rect 28460 11812 28488 11840
rect 29365 11815 29423 11821
rect 29365 11812 29377 11815
rect 23247 11784 23999 11812
rect 28460 11784 29377 11812
rect 23247 11781 23259 11784
rect 23201 11775 23259 11781
rect 16945 11716 18092 11744
rect 18509 11747 18567 11753
rect 16945 11713 16957 11716
rect 16899 11707 16957 11713
rect 18509 11713 18521 11747
rect 18555 11744 18567 11747
rect 19156 11747 19214 11753
rect 19156 11744 19168 11747
rect 18555 11716 19168 11744
rect 18555 11713 18567 11716
rect 18509 11707 18567 11713
rect 19156 11713 19168 11716
rect 19202 11713 19214 11747
rect 19156 11707 19214 11713
rect 20806 11704 20812 11756
rect 20864 11744 20870 11756
rect 21364 11747 21422 11753
rect 21364 11744 21376 11747
rect 20864 11716 21376 11744
rect 20864 11704 20870 11716
rect 21364 11713 21376 11716
rect 21410 11713 21422 11747
rect 21364 11707 21422 11713
rect 21450 11704 21456 11756
rect 21508 11744 21514 11756
rect 21637 11747 21695 11753
rect 21637 11744 21649 11747
rect 21508 11716 21649 11744
rect 21508 11704 21514 11716
rect 21637 11713 21649 11716
rect 21683 11713 21695 11747
rect 23971 11744 23999 11784
rect 29365 11781 29377 11784
rect 29411 11781 29423 11815
rect 29365 11775 29423 11781
rect 30374 11772 30380 11824
rect 30432 11772 30438 11824
rect 24394 11744 24400 11756
rect 23971 11716 24400 11744
rect 21637 11707 21695 11713
rect 24394 11704 24400 11716
rect 24452 11704 24458 11756
rect 24719 11747 24777 11753
rect 24719 11713 24731 11747
rect 24765 11744 24777 11747
rect 24765 11716 25360 11744
rect 24765 11713 24777 11716
rect 24719 11707 24777 11713
rect 25332 11688 25360 11716
rect 25958 11704 25964 11756
rect 26016 11744 26022 11756
rect 26884 11747 26942 11753
rect 26884 11744 26896 11747
rect 26016 11716 26896 11744
rect 26016 11704 26022 11716
rect 26884 11713 26896 11716
rect 26930 11713 26942 11747
rect 28902 11744 28908 11756
rect 26884 11707 26942 11713
rect 28828 11716 28908 11744
rect 17129 11679 17187 11685
rect 17129 11676 17141 11679
rect 16598 11648 17141 11676
rect 16393 11639 16451 11645
rect 17129 11645 17141 11648
rect 17175 11645 17187 11679
rect 17129 11639 17187 11645
rect 11756 11580 13032 11608
rect 11756 11568 11762 11580
rect 10097 11512 11192 11540
rect 11609 11543 11667 11549
rect 10097 11509 10109 11512
rect 10051 11503 10109 11509
rect 11609 11509 11621 11543
rect 11655 11540 11667 11543
rect 12158 11540 12164 11552
rect 11655 11512 12164 11540
rect 11655 11509 11667 11512
rect 11609 11503 11667 11509
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 12342 11500 12348 11552
rect 12400 11500 12406 11552
rect 12805 11543 12863 11549
rect 12805 11509 12817 11543
rect 12851 11540 12863 11543
rect 13170 11540 13176 11552
rect 12851 11512 13176 11540
rect 12851 11509 12863 11512
rect 12805 11503 12863 11509
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 13262 11500 13268 11552
rect 13320 11540 13326 11552
rect 14007 11543 14065 11549
rect 14007 11540 14019 11543
rect 13320 11512 14019 11540
rect 13320 11500 13326 11512
rect 14007 11509 14019 11512
rect 14053 11509 14065 11543
rect 14007 11503 14065 11509
rect 14918 11500 14924 11552
rect 14976 11540 14982 11552
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 14976 11512 15393 11540
rect 14976 11500 14982 11512
rect 15381 11509 15393 11512
rect 15427 11509 15439 11543
rect 16408 11540 16436 11639
rect 18690 11636 18696 11688
rect 18748 11636 18754 11688
rect 19058 11636 19064 11688
rect 19116 11676 19122 11688
rect 19429 11679 19487 11685
rect 19429 11676 19441 11679
rect 19116 11648 19441 11676
rect 19116 11636 19122 11648
rect 19429 11645 19441 11648
rect 19475 11645 19487 11679
rect 19429 11639 19487 11645
rect 20901 11679 20959 11685
rect 20901 11645 20913 11679
rect 20947 11676 20959 11679
rect 21266 11676 21272 11688
rect 20947 11648 21272 11676
rect 20947 11645 20959 11648
rect 20901 11639 20959 11645
rect 21266 11636 21272 11648
rect 21324 11676 21330 11688
rect 22922 11676 22928 11688
rect 21324 11648 22928 11676
rect 21324 11636 21330 11648
rect 22922 11636 22928 11648
rect 22980 11636 22986 11688
rect 23290 11636 23296 11688
rect 23348 11676 23354 11688
rect 23385 11679 23443 11685
rect 23385 11676 23397 11679
rect 23348 11648 23397 11676
rect 23348 11636 23354 11648
rect 23385 11645 23397 11648
rect 23431 11645 23443 11679
rect 23385 11639 23443 11645
rect 23661 11679 23719 11685
rect 23661 11645 23673 11679
rect 23707 11645 23719 11679
rect 23661 11639 23719 11645
rect 23676 11608 23704 11639
rect 23842 11636 23848 11688
rect 23900 11636 23906 11688
rect 23934 11636 23940 11688
rect 23992 11676 23998 11688
rect 23992 11648 24164 11676
rect 23992 11636 23998 11648
rect 24136 11608 24164 11648
rect 24210 11636 24216 11688
rect 24268 11636 24274 11688
rect 24949 11679 25007 11685
rect 24949 11676 24961 11679
rect 24320 11648 24961 11676
rect 24320 11608 24348 11648
rect 24949 11645 24961 11648
rect 24995 11645 25007 11679
rect 24949 11639 25007 11645
rect 25314 11636 25320 11688
rect 25372 11636 25378 11688
rect 26418 11636 26424 11688
rect 26476 11636 26482 11688
rect 27154 11636 27160 11688
rect 27212 11636 27218 11688
rect 28828 11685 28856 11716
rect 28902 11704 28908 11716
rect 28960 11744 28966 11756
rect 29178 11744 29184 11756
rect 28960 11716 29184 11744
rect 28960 11704 28966 11716
rect 29178 11704 29184 11716
rect 29236 11704 29242 11756
rect 29270 11704 29276 11756
rect 29328 11744 29334 11756
rect 30466 11744 30472 11756
rect 29328 11716 30472 11744
rect 29328 11704 29334 11716
rect 30466 11704 30472 11716
rect 30524 11704 30530 11756
rect 31110 11744 31116 11756
rect 30576 11716 31116 11744
rect 30576 11688 30604 11716
rect 31110 11704 31116 11716
rect 31168 11704 31174 11756
rect 28813 11679 28871 11685
rect 28813 11645 28825 11679
rect 28859 11645 28871 11679
rect 28813 11639 28871 11645
rect 29086 11636 29092 11688
rect 29144 11636 29150 11688
rect 29454 11636 29460 11688
rect 29512 11676 29518 11688
rect 29549 11679 29607 11685
rect 29549 11676 29561 11679
rect 29512 11648 29561 11676
rect 29512 11636 29518 11648
rect 29549 11645 29561 11648
rect 29595 11645 29607 11679
rect 29549 11639 29607 11645
rect 29822 11636 29828 11688
rect 29880 11636 29886 11688
rect 29914 11636 29920 11688
rect 29972 11676 29978 11688
rect 30101 11679 30159 11685
rect 30101 11676 30113 11679
rect 29972 11648 30113 11676
rect 29972 11636 29978 11648
rect 30101 11645 30113 11648
rect 30147 11645 30159 11679
rect 30101 11639 30159 11645
rect 30558 11636 30564 11688
rect 30616 11636 30622 11688
rect 29840 11608 29868 11636
rect 22572 11580 24072 11608
rect 24136 11580 24348 11608
rect 28828 11580 29868 11608
rect 22572 11552 22600 11580
rect 16758 11540 16764 11552
rect 16408 11512 16764 11540
rect 15381 11503 15439 11509
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 16859 11543 16917 11549
rect 16859 11509 16871 11543
rect 16905 11540 16917 11543
rect 17218 11540 17224 11552
rect 16905 11512 17224 11540
rect 16905 11509 16917 11512
rect 16859 11503 16917 11509
rect 17218 11500 17224 11512
rect 17276 11500 17282 11552
rect 19150 11500 19156 11552
rect 19208 11549 19214 11552
rect 19208 11540 19217 11549
rect 21367 11543 21425 11549
rect 19208 11512 19253 11540
rect 19208 11503 19217 11512
rect 21367 11509 21379 11543
rect 21413 11540 21425 11543
rect 21910 11540 21916 11552
rect 21413 11512 21916 11540
rect 21413 11509 21425 11512
rect 21367 11503 21425 11509
rect 19208 11500 19214 11503
rect 21910 11500 21916 11512
rect 21968 11540 21974 11552
rect 22370 11540 22376 11552
rect 21968 11512 22376 11540
rect 21968 11500 21974 11512
rect 22370 11500 22376 11512
rect 22428 11500 22434 11552
rect 22554 11500 22560 11552
rect 22612 11500 22618 11552
rect 23477 11543 23535 11549
rect 23477 11509 23489 11543
rect 23523 11540 23535 11543
rect 23934 11540 23940 11552
rect 23523 11512 23940 11540
rect 23523 11509 23535 11512
rect 23477 11503 23535 11509
rect 23934 11500 23940 11512
rect 23992 11500 23998 11552
rect 24044 11549 24072 11580
rect 28828 11552 28856 11580
rect 24029 11543 24087 11549
rect 24029 11509 24041 11543
rect 24075 11509 24087 11543
rect 24029 11503 24087 11509
rect 24670 11500 24676 11552
rect 24728 11549 24734 11552
rect 24728 11540 24737 11549
rect 24728 11512 24773 11540
rect 24728 11503 24737 11512
rect 24728 11500 24734 11503
rect 26694 11500 26700 11552
rect 26752 11540 26758 11552
rect 26887 11543 26945 11549
rect 26887 11540 26899 11543
rect 26752 11512 26899 11540
rect 26752 11500 26758 11512
rect 26887 11509 26899 11512
rect 26933 11509 26945 11543
rect 26887 11503 26945 11509
rect 28810 11500 28816 11552
rect 28868 11500 28874 11552
rect 29086 11500 29092 11552
rect 29144 11540 29150 11552
rect 29181 11543 29239 11549
rect 29181 11540 29193 11543
rect 29144 11512 29193 11540
rect 29144 11500 29150 11512
rect 29181 11509 29193 11512
rect 29227 11540 29239 11543
rect 29454 11540 29460 11552
rect 29227 11512 29460 11540
rect 29227 11509 29239 11512
rect 29181 11503 29239 11509
rect 29454 11500 29460 11512
rect 29512 11500 29518 11552
rect 29638 11500 29644 11552
rect 29696 11500 29702 11552
rect 552 11450 31072 11472
rect 552 11398 7988 11450
rect 8040 11398 8052 11450
rect 8104 11398 8116 11450
rect 8168 11398 8180 11450
rect 8232 11398 8244 11450
rect 8296 11398 15578 11450
rect 15630 11398 15642 11450
rect 15694 11398 15706 11450
rect 15758 11398 15770 11450
rect 15822 11398 15834 11450
rect 15886 11398 23168 11450
rect 23220 11398 23232 11450
rect 23284 11398 23296 11450
rect 23348 11398 23360 11450
rect 23412 11398 23424 11450
rect 23476 11398 30758 11450
rect 30810 11398 30822 11450
rect 30874 11398 30886 11450
rect 30938 11398 30950 11450
rect 31002 11398 31014 11450
rect 31066 11398 31072 11450
rect 552 11376 31072 11398
rect 1302 11296 1308 11348
rect 1360 11296 1366 11348
rect 1762 11296 1768 11348
rect 1820 11336 1826 11348
rect 1955 11339 2013 11345
rect 1955 11336 1967 11339
rect 1820 11308 1967 11336
rect 1820 11296 1826 11308
rect 1955 11305 1967 11308
rect 2001 11336 2013 11339
rect 8386 11336 8392 11348
rect 2001 11308 5396 11336
rect 2001 11305 2013 11308
rect 1955 11299 2013 11305
rect 1029 11203 1087 11209
rect 1029 11169 1041 11203
rect 1075 11169 1087 11203
rect 1320 11200 1348 11296
rect 3605 11271 3663 11277
rect 3605 11237 3617 11271
rect 3651 11268 3663 11271
rect 3973 11271 4031 11277
rect 3651 11240 3924 11268
rect 3651 11237 3663 11240
rect 3605 11231 3663 11237
rect 1489 11203 1547 11209
rect 1489 11200 1501 11203
rect 1320 11172 1501 11200
rect 1029 11163 1087 11169
rect 1489 11169 1501 11172
rect 1535 11169 1547 11203
rect 1489 11163 1547 11169
rect 1044 11132 1072 11163
rect 1578 11160 1584 11212
rect 1636 11160 1642 11212
rect 2130 11160 2136 11212
rect 2188 11200 2194 11212
rect 2225 11203 2283 11209
rect 2225 11200 2237 11203
rect 2188 11172 2237 11200
rect 2188 11160 2194 11172
rect 2225 11169 2237 11172
rect 2271 11169 2283 11203
rect 2225 11163 2283 11169
rect 3697 11203 3755 11209
rect 3697 11169 3709 11203
rect 3743 11169 3755 11203
rect 3896 11200 3924 11240
rect 3973 11237 3985 11271
rect 4019 11268 4031 11271
rect 4062 11268 4068 11280
rect 4019 11240 4068 11268
rect 4019 11237 4031 11240
rect 3973 11231 4031 11237
rect 4062 11228 4068 11240
rect 4120 11228 4126 11280
rect 5368 11277 5396 11308
rect 5736 11308 8392 11336
rect 5353 11271 5411 11277
rect 4448 11240 5304 11268
rect 4246 11200 4252 11212
rect 3896 11172 4252 11200
rect 3697 11163 3755 11169
rect 1596 11132 1624 11160
rect 1985 11153 2043 11159
rect 1985 11150 1997 11153
rect 1964 11144 1997 11150
rect 1044 11104 1624 11132
rect 1946 11092 1952 11144
rect 2031 11119 2043 11153
rect 2004 11113 2043 11119
rect 2004 11092 2010 11113
rect 3718 10996 3746 11163
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 4448 11209 4476 11240
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 4617 11203 4675 11209
rect 4617 11169 4629 11203
rect 4663 11200 4675 11203
rect 5077 11203 5135 11209
rect 4663 11172 5028 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 3970 11092 3976 11144
rect 4028 11132 4034 11144
rect 4893 11135 4951 11141
rect 4893 11132 4905 11135
rect 4028 11104 4905 11132
rect 4028 11092 4034 11104
rect 4893 11101 4905 11104
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 4249 11067 4307 11073
rect 4249 11033 4261 11067
rect 4295 11064 4307 11067
rect 4614 11064 4620 11076
rect 4295 11036 4620 11064
rect 4295 11033 4307 11036
rect 4249 11027 4307 11033
rect 4614 11024 4620 11036
rect 4672 11024 4678 11076
rect 5000 11064 5028 11172
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 5166 11200 5172 11212
rect 5123 11172 5172 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 5276 11200 5304 11240
rect 5353 11237 5365 11271
rect 5399 11237 5411 11271
rect 5353 11231 5411 11237
rect 5736 11200 5764 11308
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 8478 11296 8484 11348
rect 8536 11296 8542 11348
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 11422 11336 11428 11348
rect 8628 11308 11428 11336
rect 8628 11296 8634 11308
rect 11422 11296 11428 11308
rect 11480 11296 11486 11348
rect 11514 11296 11520 11348
rect 11572 11296 11578 11348
rect 12802 11336 12808 11348
rect 11808 11308 12808 11336
rect 5276 11172 5764 11200
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 6362 11200 6368 11212
rect 5813 11163 5871 11169
rect 6155 11172 6368 11200
rect 5534 11092 5540 11144
rect 5592 11132 5598 11144
rect 5828 11132 5856 11163
rect 5994 11132 6000 11144
rect 5592 11104 6000 11132
rect 5592 11092 5598 11104
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 6155 11141 6183 11172
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 6822 11160 6828 11212
rect 6880 11160 6886 11212
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 8205 11203 8263 11209
rect 8205 11200 8217 11203
rect 7524 11172 8217 11200
rect 7524 11160 7530 11172
rect 8205 11169 8217 11172
rect 8251 11169 8263 11203
rect 8496 11200 8524 11296
rect 11808 11268 11836 11308
rect 12802 11296 12808 11308
rect 12860 11336 12866 11348
rect 12995 11339 13053 11345
rect 12995 11336 13007 11339
rect 12860 11308 13007 11336
rect 12860 11296 12866 11308
rect 12995 11305 13007 11308
rect 13041 11336 13053 11339
rect 13262 11336 13268 11348
rect 13041 11308 13268 11336
rect 13041 11305 13053 11308
rect 12995 11299 13053 11305
rect 13262 11296 13268 11308
rect 13320 11296 13326 11348
rect 14182 11296 14188 11348
rect 14240 11336 14246 11348
rect 15102 11336 15108 11348
rect 14240 11308 15108 11336
rect 14240 11296 14246 11308
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 16390 11296 16396 11348
rect 16448 11296 16454 11348
rect 16666 11296 16672 11348
rect 16724 11296 16730 11348
rect 18877 11339 18935 11345
rect 16868 11308 18276 11336
rect 10704 11240 11836 11268
rect 11885 11271 11943 11277
rect 9401 11203 9459 11209
rect 8496 11172 9171 11200
rect 8205 11163 8263 11169
rect 6140 11135 6198 11141
rect 6140 11101 6152 11135
rect 6186 11101 6198 11135
rect 6140 11095 6198 11101
rect 6270 11092 6276 11144
rect 6328 11092 6334 11144
rect 6454 11092 6460 11144
rect 6512 11132 6518 11144
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 6512 11104 6561 11132
rect 6512 11092 6518 11104
rect 6549 11101 6561 11104
rect 6595 11101 6607 11135
rect 6840 11132 6868 11160
rect 6840 11104 7512 11132
rect 6549 11095 6607 11101
rect 5552 11064 5580 11092
rect 5000 11036 5580 11064
rect 7484 11064 7512 11104
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 7708 11104 7941 11132
rect 7708 11092 7714 11104
rect 7929 11101 7941 11104
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 7834 11064 7840 11076
rect 7484 11036 7840 11064
rect 7834 11024 7840 11036
rect 7892 11064 7898 11076
rect 8220 11064 8248 11163
rect 8294 11092 8300 11144
rect 8352 11132 8358 11144
rect 8665 11135 8723 11141
rect 8665 11132 8677 11135
rect 8352 11104 8677 11132
rect 8352 11092 8358 11104
rect 8665 11101 8677 11104
rect 8711 11101 8723 11135
rect 8665 11095 8723 11101
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 9030 11141 9036 11144
rect 8992 11135 9036 11141
rect 8992 11132 9004 11135
rect 8904 11104 9004 11132
rect 8904 11092 8910 11104
rect 8992 11101 9004 11104
rect 8992 11095 9036 11101
rect 9030 11092 9036 11095
rect 9088 11092 9094 11144
rect 9143 11143 9171 11172
rect 9401 11169 9413 11203
rect 9447 11200 9459 11203
rect 10594 11200 10600 11212
rect 9447 11172 10600 11200
rect 9447 11169 9459 11172
rect 9401 11163 9459 11169
rect 10594 11160 10600 11172
rect 10652 11160 10658 11212
rect 9128 11137 9186 11143
rect 9128 11103 9140 11137
rect 9174 11103 9186 11137
rect 9128 11097 9186 11103
rect 9490 11092 9496 11144
rect 9548 11132 9554 11144
rect 10704 11132 10732 11240
rect 11885 11237 11897 11271
rect 11931 11268 11943 11271
rect 12066 11268 12072 11280
rect 11931 11240 12072 11268
rect 11931 11237 11943 11240
rect 11885 11231 11943 11237
rect 12066 11228 12072 11240
rect 12124 11228 12130 11280
rect 15841 11271 15899 11277
rect 15841 11268 15853 11271
rect 15120 11240 15853 11268
rect 11054 11160 11060 11212
rect 11112 11160 11118 11212
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11200 11207 11203
rect 11425 11203 11483 11209
rect 11195 11172 11376 11200
rect 11195 11169 11207 11172
rect 11149 11163 11207 11169
rect 9548 11104 10732 11132
rect 10781 11135 10839 11141
rect 9548 11092 9554 11104
rect 10781 11101 10793 11135
rect 10827 11132 10839 11135
rect 11072 11132 11100 11160
rect 10827 11104 11100 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 11348 11076 11376 11172
rect 11425 11169 11437 11203
rect 11471 11169 11483 11203
rect 11425 11163 11483 11169
rect 7892 11036 8156 11064
rect 8220 11036 8708 11064
rect 7892 11024 7898 11036
rect 5166 10996 5172 11008
rect 3718 10968 5172 10996
rect 5166 10956 5172 10968
rect 5224 10996 5230 11008
rect 6546 10996 6552 11008
rect 5224 10968 6552 10996
rect 5224 10956 5230 10968
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 8128 10996 8156 11036
rect 8389 10999 8447 11005
rect 8389 10996 8401 10999
rect 8128 10968 8401 10996
rect 8389 10965 8401 10968
rect 8435 10965 8447 10999
rect 8680 10996 8708 11036
rect 11238 11024 11244 11076
rect 11296 11024 11302 11076
rect 11330 11024 11336 11076
rect 11388 11024 11394 11076
rect 11440 11064 11468 11163
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 11701 11203 11759 11209
rect 11701 11200 11713 11203
rect 11572 11172 11713 11200
rect 11572 11160 11578 11172
rect 11701 11169 11713 11172
rect 11747 11169 11759 11203
rect 12253 11203 12311 11209
rect 12253 11200 12265 11203
rect 11701 11163 11759 11169
rect 11992 11172 12265 11200
rect 11716 11132 11744 11163
rect 11992 11132 12020 11172
rect 12253 11169 12265 11172
rect 12299 11169 12311 11203
rect 12253 11163 12311 11169
rect 12460 11172 12848 11200
rect 11716 11104 12020 11132
rect 12158 11092 12164 11144
rect 12216 11132 12222 11144
rect 12460 11132 12488 11172
rect 12216 11104 12488 11132
rect 12529 11135 12587 11141
rect 12216 11092 12222 11104
rect 12529 11101 12541 11135
rect 12575 11132 12587 11135
rect 12710 11132 12716 11144
rect 12575 11104 12716 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 12820 11132 12848 11172
rect 13078 11160 13084 11212
rect 13136 11200 13142 11212
rect 13265 11203 13323 11209
rect 13265 11200 13277 11203
rect 13136 11172 13277 11200
rect 13136 11160 13142 11172
rect 13265 11169 13277 11172
rect 13311 11169 13323 11203
rect 13265 11163 13323 11169
rect 13354 11160 13360 11212
rect 13412 11200 13418 11212
rect 14921 11203 14979 11209
rect 14921 11200 14933 11203
rect 13412 11172 14933 11200
rect 13412 11160 13418 11172
rect 14921 11169 14933 11172
rect 14967 11169 14979 11203
rect 14921 11163 14979 11169
rect 12992 11135 13050 11141
rect 12992 11132 13004 11135
rect 12820 11104 13004 11132
rect 12992 11101 13004 11104
rect 13038 11101 13050 11135
rect 12992 11095 13050 11101
rect 13170 11092 13176 11144
rect 13228 11132 13234 11144
rect 14734 11132 14740 11144
rect 13228 11104 14740 11132
rect 13228 11092 13234 11104
rect 14734 11092 14740 11104
rect 14792 11132 14798 11144
rect 15120 11132 15148 11240
rect 15841 11237 15853 11240
rect 15887 11268 15899 11271
rect 16298 11268 16304 11280
rect 15887 11240 16304 11268
rect 15887 11237 15899 11240
rect 15841 11231 15899 11237
rect 16298 11228 16304 11240
rect 16356 11228 16362 11280
rect 15194 11160 15200 11212
rect 15252 11200 15258 11212
rect 16408 11200 16436 11296
rect 15252 11172 16436 11200
rect 16684 11200 16712 11296
rect 16868 11280 16896 11308
rect 16850 11228 16856 11280
rect 16908 11228 16914 11280
rect 17589 11203 17647 11209
rect 17589 11200 17601 11203
rect 16684 11172 17601 11200
rect 15252 11160 15258 11172
rect 17589 11169 17601 11172
rect 17635 11169 17647 11203
rect 18248 11200 18276 11308
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 18966 11336 18972 11348
rect 18923 11308 18972 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 20346 11296 20352 11348
rect 20404 11336 20410 11348
rect 22002 11336 22008 11348
rect 20404 11308 22008 11336
rect 20404 11296 20410 11308
rect 22002 11296 22008 11308
rect 22060 11296 22066 11348
rect 22370 11296 22376 11348
rect 22428 11336 22434 11348
rect 23943 11339 24001 11345
rect 23943 11336 23955 11339
rect 22428 11308 23955 11336
rect 22428 11296 22434 11308
rect 23943 11305 23955 11308
rect 23989 11336 24001 11339
rect 23989 11308 25268 11336
rect 23989 11305 24001 11308
rect 23943 11299 24001 11305
rect 19150 11228 19156 11280
rect 19208 11268 19214 11280
rect 19337 11271 19395 11277
rect 19337 11268 19349 11271
rect 19208 11240 19349 11268
rect 19208 11228 19214 11240
rect 19337 11237 19349 11240
rect 19383 11268 19395 11271
rect 21358 11268 21364 11280
rect 19383 11240 21364 11268
rect 19383 11237 19395 11240
rect 19337 11231 19395 11237
rect 21358 11228 21364 11240
rect 21416 11228 21422 11280
rect 23014 11228 23020 11280
rect 23072 11268 23078 11280
rect 25240 11268 25268 11308
rect 25314 11296 25320 11348
rect 25372 11296 25378 11348
rect 26418 11296 26424 11348
rect 26476 11336 26482 11348
rect 26476 11308 27108 11336
rect 26476 11296 26482 11308
rect 26694 11268 26700 11280
rect 23072 11240 23612 11268
rect 25240 11240 26700 11268
rect 23072 11228 23078 11240
rect 19061 11203 19119 11209
rect 19061 11200 19073 11203
rect 18248 11172 19073 11200
rect 17589 11163 17647 11169
rect 19061 11169 19073 11172
rect 19107 11169 19119 11203
rect 22646 11200 22652 11212
rect 19061 11163 19119 11169
rect 21928 11172 22652 11200
rect 21765 11153 21823 11159
rect 21765 11150 21777 11153
rect 14792 11104 15148 11132
rect 14792 11092 14798 11104
rect 16758 11092 16764 11144
rect 16816 11132 16822 11144
rect 17218 11141 17224 11144
rect 16853 11135 16911 11141
rect 16853 11132 16865 11135
rect 16816 11104 16865 11132
rect 16816 11092 16822 11104
rect 16853 11101 16865 11104
rect 16899 11101 16911 11135
rect 16853 11095 16911 11101
rect 17180 11135 17224 11141
rect 17180 11101 17192 11135
rect 17180 11095 17224 11101
rect 11514 11064 11520 11076
rect 11440 11036 11520 11064
rect 11514 11024 11520 11036
rect 11572 11024 11578 11076
rect 11790 11024 11796 11076
rect 11848 11064 11854 11076
rect 12069 11067 12127 11073
rect 12069 11064 12081 11067
rect 11848 11036 12081 11064
rect 11848 11024 11854 11036
rect 12069 11033 12081 11036
rect 12115 11064 12127 11067
rect 12250 11064 12256 11076
rect 12115 11036 12256 11064
rect 12115 11033 12127 11036
rect 12069 11027 12127 11033
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 12434 11024 12440 11076
rect 12492 11024 12498 11076
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 15013 11067 15071 11073
rect 15013 11064 15025 11067
rect 14884 11036 15025 11064
rect 14884 11024 14890 11036
rect 15013 11033 15025 11036
rect 15059 11033 15071 11067
rect 15013 11027 15071 11033
rect 9858 10996 9864 11008
rect 8680 10968 9864 10996
rect 8389 10959 8447 10965
rect 9858 10956 9864 10968
rect 9916 10956 9922 11008
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 10965 10999 11023 11005
rect 10965 10996 10977 10999
rect 10652 10968 10977 10996
rect 10652 10956 10658 10968
rect 10965 10965 10977 10968
rect 11011 10965 11023 10999
rect 10965 10959 11023 10965
rect 11698 10956 11704 11008
rect 11756 10996 11762 11008
rect 12526 10996 12532 11008
rect 11756 10968 12532 10996
rect 11756 10956 11762 10968
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 13722 10956 13728 11008
rect 13780 10996 13786 11008
rect 14369 10999 14427 11005
rect 14369 10996 14381 10999
rect 13780 10968 14381 10996
rect 13780 10956 13786 10968
rect 14369 10965 14381 10968
rect 14415 10965 14427 10999
rect 14369 10959 14427 10965
rect 14734 10956 14740 11008
rect 14792 10956 14798 11008
rect 15470 10956 15476 11008
rect 15528 10956 15534 11008
rect 16868 10996 16896 11095
rect 17218 11092 17224 11095
rect 17276 11092 17282 11144
rect 17359 11135 17417 11141
rect 17359 11101 17371 11135
rect 17405 11132 17417 11135
rect 17405 11104 19012 11132
rect 17405 11101 17417 11104
rect 17359 11095 17417 11101
rect 18984 11064 19012 11104
rect 20806 11092 20812 11144
rect 20864 11092 20870 11144
rect 21082 11092 21088 11144
rect 21140 11132 21146 11144
rect 21269 11135 21327 11141
rect 21269 11132 21281 11135
rect 21140 11104 21281 11132
rect 21140 11092 21146 11104
rect 21269 11101 21281 11104
rect 21315 11101 21327 11135
rect 21269 11095 21327 11101
rect 21542 11092 21548 11144
rect 21600 11141 21606 11144
rect 21600 11135 21654 11141
rect 21600 11101 21608 11135
rect 21642 11101 21654 11135
rect 21763 11119 21777 11150
rect 21811 11132 21823 11153
rect 21928 11132 21956 11172
rect 22646 11160 22652 11172
rect 22704 11160 22710 11212
rect 23584 11200 23612 11240
rect 26694 11228 26700 11240
rect 26752 11228 26758 11280
rect 27080 11277 27108 11308
rect 27154 11296 27160 11348
rect 27212 11336 27218 11348
rect 27525 11339 27583 11345
rect 27525 11336 27537 11339
rect 27212 11308 27537 11336
rect 27212 11296 27218 11308
rect 27525 11305 27537 11308
rect 27571 11305 27583 11339
rect 27525 11299 27583 11305
rect 27706 11296 27712 11348
rect 27764 11296 27770 11348
rect 27798 11296 27804 11348
rect 27856 11296 27862 11348
rect 27890 11296 27896 11348
rect 27948 11336 27954 11348
rect 29917 11339 29975 11345
rect 29917 11336 29929 11339
rect 27948 11308 29929 11336
rect 27948 11296 27954 11308
rect 29917 11305 29929 11308
rect 29963 11305 29975 11339
rect 29917 11299 29975 11305
rect 30466 11296 30472 11348
rect 30524 11296 30530 11348
rect 27065 11271 27123 11277
rect 27065 11237 27077 11271
rect 27111 11237 27123 11271
rect 27724 11268 27752 11296
rect 27724 11240 28120 11268
rect 27065 11231 27123 11237
rect 24213 11203 24271 11209
rect 24213 11200 24225 11203
rect 23584 11172 24225 11200
rect 24213 11169 24225 11172
rect 24259 11169 24271 11203
rect 24213 11163 24271 11169
rect 25590 11160 25596 11212
rect 25648 11200 25654 11212
rect 25777 11203 25835 11209
rect 25777 11200 25789 11203
rect 25648 11172 25789 11200
rect 25648 11160 25654 11172
rect 25777 11169 25789 11172
rect 25823 11200 25835 11203
rect 26142 11200 26148 11212
rect 25823 11172 26148 11200
rect 25823 11169 25835 11172
rect 25777 11163 25835 11169
rect 26142 11160 26148 11172
rect 26200 11160 26206 11212
rect 26326 11160 26332 11212
rect 26384 11200 26390 11212
rect 26421 11203 26479 11209
rect 26421 11200 26433 11203
rect 26384 11172 26433 11200
rect 26384 11160 26390 11172
rect 26421 11169 26433 11172
rect 26467 11169 26479 11203
rect 26421 11163 26479 11169
rect 27709 11203 27767 11209
rect 27709 11169 27721 11203
rect 27755 11200 27767 11203
rect 27985 11203 28043 11209
rect 27985 11200 27997 11203
rect 27755 11172 27997 11200
rect 27755 11169 27767 11172
rect 27709 11163 27767 11169
rect 27985 11169 27997 11172
rect 28031 11169 28043 11203
rect 28092 11200 28120 11240
rect 29638 11228 29644 11280
rect 29696 11228 29702 11280
rect 28404 11203 28462 11209
rect 28404 11200 28416 11203
rect 28092 11172 28416 11200
rect 27985 11163 28043 11169
rect 28404 11169 28416 11172
rect 28450 11169 28462 11203
rect 28404 11163 28462 11169
rect 28813 11203 28871 11209
rect 28813 11169 28825 11203
rect 28859 11200 28871 11203
rect 29656 11200 29684 11228
rect 28859 11172 29684 11200
rect 28859 11169 28871 11172
rect 28813 11163 28871 11169
rect 21811 11119 21956 11132
rect 21763 11104 21956 11119
rect 21600 11095 21654 11101
rect 21600 11092 21606 11095
rect 22002 11092 22008 11144
rect 22060 11092 22066 11144
rect 22922 11092 22928 11144
rect 22980 11132 22986 11144
rect 23477 11135 23535 11141
rect 23477 11132 23489 11135
rect 22980 11104 23489 11132
rect 22980 11092 22986 11104
rect 23477 11101 23489 11104
rect 23523 11132 23535 11135
rect 23842 11132 23848 11144
rect 23523 11104 23848 11132
rect 23523 11101 23535 11104
rect 23477 11095 23535 11101
rect 23842 11092 23848 11104
rect 23900 11092 23906 11144
rect 23934 11092 23940 11144
rect 23992 11092 23998 11144
rect 24026 11092 24032 11144
rect 24084 11132 24090 11144
rect 27724 11132 27752 11163
rect 24084 11104 27752 11132
rect 24084 11092 24090 11104
rect 20824 11064 20852 11092
rect 18984 11036 20852 11064
rect 23293 11067 23351 11073
rect 23293 11033 23305 11067
rect 23339 11064 23351 11067
rect 26326 11064 26332 11076
rect 23339 11036 23520 11064
rect 23339 11033 23351 11036
rect 23293 11027 23351 11033
rect 19058 10996 19064 11008
rect 16868 10968 19064 10996
rect 19058 10956 19064 10968
rect 19116 10956 19122 11008
rect 23492 10996 23520 11036
rect 25884 11036 26332 11064
rect 25884 11008 25912 11036
rect 26326 11024 26332 11036
rect 26384 11024 26390 11076
rect 23750 10996 23756 11008
rect 23492 10968 23756 10996
rect 23750 10956 23756 10968
rect 23808 10956 23814 11008
rect 25866 10956 25872 11008
rect 25924 10956 25930 11008
rect 26234 10956 26240 11008
rect 26292 10996 26298 11008
rect 27157 10999 27215 11005
rect 27157 10996 27169 10999
rect 26292 10968 27169 10996
rect 26292 10956 26298 10968
rect 27157 10965 27169 10968
rect 27203 10965 27215 10999
rect 28000 10996 28028 11163
rect 30282 11160 30288 11212
rect 30340 11160 30346 11212
rect 28074 11092 28080 11144
rect 28132 11092 28138 11144
rect 28583 11135 28641 11141
rect 28583 11101 28595 11135
rect 28629 11132 28641 11135
rect 29546 11132 29552 11144
rect 28629 11104 29552 11132
rect 28629 11101 28641 11104
rect 28583 11095 28641 11101
rect 29546 11092 29552 11104
rect 29604 11092 29610 11144
rect 29454 10996 29460 11008
rect 28000 10968 29460 10996
rect 27157 10959 27215 10965
rect 29454 10956 29460 10968
rect 29512 10996 29518 11008
rect 30650 10996 30656 11008
rect 29512 10968 30656 10996
rect 29512 10956 29518 10968
rect 30650 10956 30656 10968
rect 30708 10956 30714 11008
rect 552 10906 30912 10928
rect 552 10854 4193 10906
rect 4245 10854 4257 10906
rect 4309 10854 4321 10906
rect 4373 10854 4385 10906
rect 4437 10854 4449 10906
rect 4501 10854 11783 10906
rect 11835 10854 11847 10906
rect 11899 10854 11911 10906
rect 11963 10854 11975 10906
rect 12027 10854 12039 10906
rect 12091 10854 19373 10906
rect 19425 10854 19437 10906
rect 19489 10854 19501 10906
rect 19553 10854 19565 10906
rect 19617 10854 19629 10906
rect 19681 10854 26963 10906
rect 27015 10854 27027 10906
rect 27079 10854 27091 10906
rect 27143 10854 27155 10906
rect 27207 10854 27219 10906
rect 27271 10854 30912 10906
rect 552 10832 30912 10854
rect 15470 10792 15476 10804
rect 2746 10764 15476 10792
rect 937 10659 995 10665
rect 937 10625 949 10659
rect 983 10656 995 10659
rect 1302 10656 1308 10668
rect 983 10628 1308 10656
rect 983 10625 995 10628
rect 937 10619 995 10625
rect 1302 10616 1308 10628
rect 1360 10616 1366 10668
rect 1443 10659 1501 10665
rect 1443 10625 1455 10659
rect 1489 10656 1501 10659
rect 2746 10656 2774 10764
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 21358 10752 21364 10804
rect 21416 10792 21422 10804
rect 21416 10764 22876 10792
rect 21416 10752 21422 10764
rect 11609 10727 11667 10733
rect 11609 10693 11621 10727
rect 11655 10724 11667 10727
rect 11698 10724 11704 10736
rect 11655 10696 11704 10724
rect 11655 10693 11667 10696
rect 11609 10687 11667 10693
rect 11698 10684 11704 10696
rect 11756 10684 11762 10736
rect 11974 10684 11980 10736
rect 12032 10724 12038 10736
rect 12710 10724 12716 10736
rect 12032 10696 12716 10724
rect 12032 10684 12038 10696
rect 12710 10684 12716 10696
rect 12768 10684 12774 10736
rect 13814 10684 13820 10736
rect 13872 10684 13878 10736
rect 3700 10659 3758 10665
rect 3700 10656 3712 10659
rect 1489 10628 2774 10656
rect 3160 10628 3712 10656
rect 1489 10625 1501 10628
rect 1443 10619 1501 10625
rect 3160 10600 3188 10628
rect 3700 10625 3712 10628
rect 3746 10625 3758 10659
rect 3700 10619 3758 10625
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 6000 10659 6058 10665
rect 6000 10656 6012 10659
rect 5408 10628 6012 10656
rect 5408 10616 5414 10628
rect 6000 10625 6012 10628
rect 6046 10625 6058 10659
rect 6362 10656 6368 10668
rect 6000 10619 6058 10625
rect 6104 10628 6368 10656
rect 6104 10600 6132 10628
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 7653 10659 7711 10665
rect 7653 10625 7665 10659
rect 7699 10656 7711 10659
rect 7834 10656 7840 10668
rect 7699 10628 7840 10656
rect 7699 10625 7711 10628
rect 7653 10619 7711 10625
rect 7834 10616 7840 10628
rect 7892 10616 7898 10668
rect 8757 10659 8815 10665
rect 8757 10656 8769 10659
rect 8266 10628 8769 10656
rect 658 10548 664 10600
rect 716 10588 722 10600
rect 1673 10591 1731 10597
rect 1673 10588 1685 10591
rect 716 10560 1685 10588
rect 716 10548 722 10560
rect 1673 10557 1685 10560
rect 1719 10557 1731 10591
rect 1673 10551 1731 10557
rect 3142 10548 3148 10600
rect 3200 10548 3206 10600
rect 3237 10591 3295 10597
rect 3237 10557 3249 10591
rect 3283 10588 3295 10591
rect 3602 10588 3608 10600
rect 3283 10560 3608 10588
rect 3283 10557 3295 10560
rect 3237 10551 3295 10557
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 3973 10591 4031 10597
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 5258 10588 5264 10600
rect 4019 10560 5264 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 5258 10548 5264 10560
rect 5316 10548 5322 10600
rect 5534 10548 5540 10600
rect 5592 10588 5598 10600
rect 5864 10591 5922 10597
rect 5592 10560 5672 10588
rect 5592 10548 5598 10560
rect 3050 10480 3056 10532
rect 3108 10480 3114 10532
rect 5350 10480 5356 10532
rect 5408 10480 5414 10532
rect 1403 10455 1461 10461
rect 1403 10421 1415 10455
rect 1449 10452 1461 10455
rect 1762 10452 1768 10464
rect 1449 10424 1768 10452
rect 1449 10421 1461 10424
rect 1403 10415 1461 10421
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 3326 10412 3332 10464
rect 3384 10452 3390 10464
rect 3703 10455 3761 10461
rect 3703 10452 3715 10455
rect 3384 10424 3715 10452
rect 3384 10412 3390 10424
rect 3703 10421 3715 10424
rect 3749 10452 3761 10455
rect 3970 10452 3976 10464
rect 3749 10424 3976 10452
rect 3749 10421 3761 10424
rect 3703 10415 3761 10421
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 5644 10452 5672 10560
rect 5864 10557 5876 10591
rect 5910 10588 5922 10591
rect 6086 10588 6092 10600
rect 5910 10560 6092 10588
rect 5910 10557 5922 10560
rect 5864 10551 5922 10557
rect 6086 10548 6092 10560
rect 6144 10548 6150 10600
rect 6178 10548 6184 10600
rect 6236 10588 6242 10600
rect 6273 10591 6331 10597
rect 6273 10588 6285 10591
rect 6236 10560 6285 10588
rect 6236 10548 6242 10560
rect 6273 10557 6285 10560
rect 6319 10557 6331 10591
rect 8266 10588 8294 10628
rect 8757 10625 8769 10628
rect 8803 10656 8815 10659
rect 8846 10656 8852 10668
rect 8803 10628 8852 10656
rect 8803 10625 8815 10628
rect 8757 10619 8815 10625
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 9950 10665 9956 10668
rect 9912 10659 9956 10665
rect 9912 10625 9924 10659
rect 9912 10619 9956 10625
rect 9950 10616 9956 10619
rect 10008 10616 10014 10668
rect 10042 10616 10048 10668
rect 10100 10616 10106 10668
rect 10321 10659 10379 10665
rect 10321 10625 10333 10659
rect 10367 10656 10379 10659
rect 10962 10656 10968 10668
rect 10367 10628 10968 10656
rect 10367 10625 10379 10628
rect 10321 10619 10379 10625
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 14274 10665 14280 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 11572 10628 13093 10656
rect 11572 10616 11578 10628
rect 13081 10625 13093 10628
rect 13127 10656 13139 10659
rect 14236 10659 14280 10665
rect 14236 10656 14248 10659
rect 13127 10628 14248 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 14236 10625 14248 10628
rect 14236 10619 14280 10625
rect 14274 10616 14280 10619
rect 14332 10616 14338 10668
rect 14415 10659 14473 10665
rect 14415 10625 14427 10659
rect 14461 10656 14473 10659
rect 14550 10656 14556 10668
rect 14461 10628 14556 10656
rect 14461 10625 14473 10628
rect 14415 10619 14473 10625
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 14645 10659 14703 10665
rect 14645 10625 14657 10659
rect 14691 10656 14703 10659
rect 14734 10656 14740 10668
rect 14691 10628 14740 10656
rect 14691 10625 14703 10628
rect 14645 10619 14703 10625
rect 14734 10616 14740 10628
rect 14792 10616 14798 10668
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 16856 10659 16914 10665
rect 16856 10656 16868 10659
rect 16632 10628 16868 10656
rect 16632 10616 16638 10628
rect 16856 10625 16868 10628
rect 16902 10625 16914 10659
rect 16856 10619 16914 10625
rect 20671 10659 20729 10665
rect 20671 10625 20683 10659
rect 20717 10656 20729 10659
rect 20717 10628 21404 10656
rect 20717 10625 20729 10628
rect 20671 10619 20729 10625
rect 21376 10600 21404 10628
rect 6273 10551 6331 10557
rect 7116 10560 8294 10588
rect 8481 10591 8539 10597
rect 7116 10532 7144 10560
rect 8481 10557 8493 10591
rect 8527 10588 8539 10591
rect 8662 10588 8668 10600
rect 8527 10560 8668 10588
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 9030 10548 9036 10600
rect 9088 10548 9094 10600
rect 9306 10588 9312 10600
rect 9140 10560 9312 10588
rect 7098 10480 7104 10532
rect 7156 10480 7162 10532
rect 7558 10480 7564 10532
rect 7616 10520 7622 10532
rect 7837 10523 7895 10529
rect 7837 10520 7849 10523
rect 7616 10492 7849 10520
rect 7616 10480 7622 10492
rect 7837 10489 7849 10492
rect 7883 10520 7895 10523
rect 8294 10520 8300 10532
rect 7883 10492 8300 10520
rect 7883 10489 7895 10492
rect 7837 10483 7895 10489
rect 8294 10480 8300 10492
rect 8352 10520 8358 10532
rect 9140 10520 9168 10560
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 9611 10591 9669 10597
rect 9611 10588 9623 10591
rect 9600 10557 9623 10588
rect 9657 10557 9669 10591
rect 9600 10551 9669 10557
rect 8352 10492 9490 10520
rect 8352 10480 8358 10492
rect 7929 10455 7987 10461
rect 7929 10452 7941 10455
rect 5644 10424 7941 10452
rect 7929 10421 7941 10424
rect 7975 10421 7987 10455
rect 7929 10415 7987 10421
rect 9214 10412 9220 10464
rect 9272 10412 9278 10464
rect 9462 10452 9490 10492
rect 9600 10452 9628 10551
rect 10686 10548 10692 10600
rect 10744 10588 10750 10600
rect 12897 10591 12955 10597
rect 12897 10588 12909 10591
rect 10744 10560 12909 10588
rect 10744 10548 10750 10560
rect 12897 10557 12909 10560
rect 12943 10588 12955 10591
rect 12943 10560 13860 10588
rect 12943 10557 12955 10560
rect 12897 10551 12955 10557
rect 11146 10480 11152 10532
rect 11204 10520 11210 10532
rect 11885 10523 11943 10529
rect 11885 10520 11897 10523
rect 11204 10492 11897 10520
rect 11204 10480 11210 10492
rect 11885 10489 11897 10492
rect 11931 10489 11943 10523
rect 11885 10483 11943 10489
rect 12437 10523 12495 10529
rect 12437 10489 12449 10523
rect 12483 10489 12495 10523
rect 12437 10483 12495 10489
rect 9462 10424 9628 10452
rect 9858 10412 9864 10464
rect 9916 10452 9922 10464
rect 11974 10452 11980 10464
rect 9916 10424 11980 10452
rect 9916 10412 9922 10424
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 12342 10412 12348 10464
rect 12400 10452 12406 10464
rect 12452 10452 12480 10483
rect 12802 10480 12808 10532
rect 12860 10480 12866 10532
rect 13078 10480 13084 10532
rect 13136 10520 13142 10532
rect 13633 10523 13691 10529
rect 13633 10520 13645 10523
rect 13136 10492 13645 10520
rect 13136 10480 13142 10492
rect 13633 10489 13645 10492
rect 13679 10489 13691 10523
rect 13832 10520 13860 10560
rect 13906 10548 13912 10600
rect 13964 10548 13970 10600
rect 16390 10548 16396 10600
rect 16448 10548 16454 10600
rect 16720 10591 16778 10597
rect 16720 10557 16732 10591
rect 16766 10588 16778 10591
rect 16942 10588 16948 10600
rect 16766 10560 16948 10588
rect 16766 10557 16778 10560
rect 16720 10551 16778 10557
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 17126 10548 17132 10600
rect 17184 10548 17190 10600
rect 18690 10548 18696 10600
rect 18748 10588 18754 10600
rect 18785 10591 18843 10597
rect 18785 10588 18797 10591
rect 18748 10560 18797 10588
rect 18748 10548 18754 10560
rect 18785 10557 18797 10560
rect 18831 10557 18843 10591
rect 18785 10551 18843 10557
rect 19058 10548 19064 10600
rect 19116 10588 19122 10600
rect 19153 10591 19211 10597
rect 19153 10588 19165 10591
rect 19116 10560 19165 10588
rect 19116 10548 19122 10560
rect 19153 10557 19165 10560
rect 19199 10588 19211 10591
rect 20165 10591 20223 10597
rect 20165 10588 20177 10591
rect 19199 10560 20177 10588
rect 19199 10557 19211 10560
rect 19153 10551 19211 10557
rect 20165 10557 20177 10560
rect 20211 10588 20223 10591
rect 20530 10588 20536 10600
rect 20211 10560 20536 10588
rect 20211 10557 20223 10560
rect 20165 10551 20223 10557
rect 20530 10548 20536 10560
rect 20588 10548 20594 10600
rect 20901 10591 20959 10597
rect 20901 10557 20913 10591
rect 20947 10588 20959 10591
rect 21174 10588 21180 10600
rect 20947 10560 21180 10588
rect 20947 10557 20959 10560
rect 20901 10551 20959 10557
rect 21174 10548 21180 10560
rect 21232 10548 21238 10600
rect 21358 10548 21364 10600
rect 21416 10548 21422 10600
rect 22554 10588 22560 10600
rect 22296 10560 22560 10588
rect 22296 10532 22324 10560
rect 22554 10548 22560 10560
rect 22612 10548 22618 10600
rect 13998 10520 14004 10532
rect 13832 10492 14004 10520
rect 13633 10483 13691 10489
rect 13998 10480 14004 10492
rect 14056 10480 14062 10532
rect 18506 10480 18512 10532
rect 18564 10480 18570 10532
rect 22278 10480 22284 10532
rect 22336 10480 22342 10532
rect 12400 10424 12480 10452
rect 12400 10412 12406 10424
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 14642 10452 14648 10464
rect 13596 10424 14648 10452
rect 13596 10412 13602 10424
rect 14642 10412 14648 10424
rect 14700 10412 14706 10464
rect 15286 10412 15292 10464
rect 15344 10452 15350 10464
rect 15749 10455 15807 10461
rect 15749 10452 15761 10455
rect 15344 10424 15761 10452
rect 15344 10412 15350 10424
rect 15749 10421 15761 10424
rect 15795 10421 15807 10455
rect 15749 10415 15807 10421
rect 17218 10412 17224 10464
rect 17276 10452 17282 10464
rect 20631 10455 20689 10461
rect 20631 10452 20643 10455
rect 17276 10424 20643 10452
rect 17276 10412 17282 10424
rect 20631 10421 20643 10424
rect 20677 10452 20689 10455
rect 21542 10452 21548 10464
rect 20677 10424 21548 10452
rect 20677 10421 20689 10424
rect 20631 10415 20689 10421
rect 21542 10412 21548 10424
rect 21600 10412 21606 10464
rect 21910 10412 21916 10464
rect 21968 10452 21974 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21968 10424 22017 10452
rect 21968 10412 21974 10424
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 22005 10415 22063 10421
rect 22370 10412 22376 10464
rect 22428 10412 22434 10464
rect 22848 10452 22876 10764
rect 23014 10752 23020 10804
rect 23072 10752 23078 10804
rect 25869 10795 25927 10801
rect 23676 10764 25268 10792
rect 23201 10591 23259 10597
rect 23201 10557 23213 10591
rect 23247 10557 23259 10591
rect 23676 10588 23704 10764
rect 23750 10616 23756 10668
rect 23808 10656 23814 10668
rect 24308 10659 24366 10665
rect 24308 10656 24320 10659
rect 23808 10628 24320 10656
rect 23808 10616 23814 10628
rect 24308 10625 24320 10628
rect 24354 10625 24366 10659
rect 24308 10619 24366 10625
rect 24394 10616 24400 10668
rect 24452 10656 24458 10668
rect 24581 10659 24639 10665
rect 24581 10656 24593 10659
rect 24452 10628 24593 10656
rect 24452 10616 24458 10628
rect 24581 10625 24593 10628
rect 24627 10625 24639 10659
rect 24581 10619 24639 10625
rect 23845 10591 23903 10597
rect 23845 10588 23857 10591
rect 23676 10560 23857 10588
rect 23201 10551 23259 10557
rect 23216 10520 23244 10551
rect 23768 10532 23796 10560
rect 23845 10557 23857 10560
rect 23891 10557 23903 10591
rect 25240 10588 25268 10764
rect 25869 10761 25881 10795
rect 25915 10792 25927 10795
rect 25958 10792 25964 10804
rect 25915 10764 25964 10792
rect 25915 10761 25927 10764
rect 25869 10755 25927 10761
rect 25958 10752 25964 10764
rect 26016 10752 26022 10804
rect 26142 10752 26148 10804
rect 26200 10792 26206 10804
rect 28166 10792 28172 10804
rect 26200 10764 28172 10792
rect 26200 10752 26206 10764
rect 28166 10752 28172 10764
rect 28224 10792 28230 10804
rect 29638 10792 29644 10804
rect 28224 10764 29644 10792
rect 28224 10752 28230 10764
rect 29638 10752 29644 10764
rect 29696 10752 29702 10804
rect 29730 10752 29736 10804
rect 29788 10792 29794 10804
rect 29788 10764 30052 10792
rect 29788 10752 29794 10764
rect 28442 10684 28448 10736
rect 28500 10684 28506 10736
rect 29178 10684 29184 10736
rect 29236 10724 29242 10736
rect 29236 10696 29960 10724
rect 29236 10684 29242 10696
rect 25314 10616 25320 10668
rect 25372 10656 25378 10668
rect 26510 10656 26516 10668
rect 25372 10628 26516 10656
rect 25372 10616 25378 10628
rect 26510 10616 26516 10628
rect 26568 10665 26574 10668
rect 26568 10659 26622 10665
rect 26568 10625 26576 10659
rect 26610 10625 26622 10659
rect 26568 10619 26622 10625
rect 26700 10657 26758 10663
rect 26700 10623 26712 10657
rect 26746 10623 26758 10657
rect 26568 10616 26574 10619
rect 26700 10617 26758 10623
rect 26234 10588 26240 10600
rect 25240 10560 26240 10588
rect 23845 10551 23903 10557
rect 26234 10548 26240 10560
rect 26292 10548 26298 10600
rect 26344 10584 26648 10588
rect 26715 10584 26743 10617
rect 26344 10560 26743 10584
rect 23658 10520 23664 10532
rect 23216 10492 23664 10520
rect 23658 10480 23664 10492
rect 23716 10480 23722 10532
rect 23750 10480 23756 10532
rect 23808 10480 23814 10532
rect 26344 10520 26372 10560
rect 26620 10556 26743 10560
rect 26973 10591 27031 10597
rect 26973 10557 26985 10591
rect 27019 10588 27031 10591
rect 27982 10588 27988 10600
rect 27019 10560 27988 10588
rect 27019 10557 27031 10560
rect 26973 10551 27031 10557
rect 27982 10548 27988 10560
rect 28040 10548 28046 10600
rect 28629 10591 28687 10597
rect 28629 10588 28641 10591
rect 28092 10560 28641 10588
rect 26160 10492 26372 10520
rect 26160 10464 26188 10492
rect 27798 10480 27804 10532
rect 27856 10520 27862 10532
rect 28092 10520 28120 10560
rect 28629 10557 28641 10560
rect 28675 10588 28687 10591
rect 28810 10588 28816 10600
rect 28675 10560 28816 10588
rect 28675 10557 28687 10560
rect 28629 10551 28687 10557
rect 28810 10548 28816 10560
rect 28868 10548 28874 10600
rect 28997 10591 29055 10597
rect 28997 10557 29009 10591
rect 29043 10588 29055 10591
rect 29086 10588 29092 10600
rect 29043 10560 29092 10588
rect 29043 10557 29055 10560
rect 28997 10551 29055 10557
rect 29086 10548 29092 10560
rect 29144 10548 29150 10600
rect 29932 10597 29960 10696
rect 30024 10656 30052 10764
rect 30098 10752 30104 10804
rect 30156 10792 30162 10804
rect 30377 10795 30435 10801
rect 30377 10792 30389 10795
rect 30156 10764 30389 10792
rect 30156 10752 30162 10764
rect 30377 10761 30389 10764
rect 30423 10761 30435 10795
rect 30377 10755 30435 10761
rect 30098 10656 30104 10668
rect 30024 10628 30104 10656
rect 30098 10616 30104 10628
rect 30156 10656 30162 10668
rect 30156 10628 30604 10656
rect 30156 10616 30162 10628
rect 30576 10597 30604 10628
rect 29365 10591 29423 10597
rect 29365 10557 29377 10591
rect 29411 10557 29423 10591
rect 29365 10551 29423 10557
rect 29917 10591 29975 10597
rect 29917 10557 29929 10591
rect 29963 10557 29975 10591
rect 30193 10591 30251 10597
rect 30193 10588 30205 10591
rect 29917 10551 29975 10557
rect 30024 10560 30205 10588
rect 27856 10492 28120 10520
rect 27856 10480 27862 10492
rect 28350 10480 28356 10532
rect 28408 10480 28414 10532
rect 29270 10520 29276 10532
rect 28460 10492 29276 10520
rect 24311 10455 24369 10461
rect 24311 10452 24323 10455
rect 22848 10424 24323 10452
rect 24311 10421 24323 10424
rect 24357 10452 24369 10455
rect 25314 10452 25320 10464
rect 24357 10424 25320 10452
rect 24357 10421 24369 10424
rect 24311 10415 24369 10421
rect 25314 10412 25320 10424
rect 25372 10412 25378 10464
rect 26142 10412 26148 10464
rect 26200 10412 26206 10464
rect 26326 10412 26332 10464
rect 26384 10452 26390 10464
rect 28460 10452 28488 10492
rect 29270 10480 29276 10492
rect 29328 10520 29334 10532
rect 29380 10520 29408 10551
rect 30024 10520 30052 10560
rect 30193 10557 30205 10560
rect 30239 10557 30251 10591
rect 30193 10551 30251 10557
rect 30561 10591 30619 10597
rect 30561 10557 30573 10591
rect 30607 10557 30619 10591
rect 30561 10551 30619 10557
rect 29328 10492 29408 10520
rect 29564 10492 30052 10520
rect 29328 10480 29334 10492
rect 26384 10424 28488 10452
rect 26384 10412 26390 10424
rect 28534 10412 28540 10464
rect 28592 10452 28598 10464
rect 29564 10461 29592 10492
rect 29549 10455 29607 10461
rect 29549 10452 29561 10455
rect 28592 10424 29561 10452
rect 28592 10412 28598 10424
rect 29549 10421 29561 10424
rect 29595 10421 29607 10455
rect 29549 10415 29607 10421
rect 29733 10455 29791 10461
rect 29733 10421 29745 10455
rect 29779 10452 29791 10455
rect 29822 10452 29828 10464
rect 29779 10424 29828 10452
rect 29779 10421 29791 10424
rect 29733 10415 29791 10421
rect 29822 10412 29828 10424
rect 29880 10412 29886 10464
rect 29914 10412 29920 10464
rect 29972 10452 29978 10464
rect 30009 10455 30067 10461
rect 30009 10452 30021 10455
rect 29972 10424 30021 10452
rect 29972 10412 29978 10424
rect 30009 10421 30021 10424
rect 30055 10421 30067 10455
rect 30009 10415 30067 10421
rect 552 10362 31072 10384
rect 552 10310 7988 10362
rect 8040 10310 8052 10362
rect 8104 10310 8116 10362
rect 8168 10310 8180 10362
rect 8232 10310 8244 10362
rect 8296 10310 15578 10362
rect 15630 10310 15642 10362
rect 15694 10310 15706 10362
rect 15758 10310 15770 10362
rect 15822 10310 15834 10362
rect 15886 10310 23168 10362
rect 23220 10310 23232 10362
rect 23284 10310 23296 10362
rect 23348 10310 23360 10362
rect 23412 10310 23424 10362
rect 23476 10310 30758 10362
rect 30810 10310 30822 10362
rect 30874 10310 30886 10362
rect 30938 10310 30950 10362
rect 31002 10310 31014 10362
rect 31066 10310 31072 10362
rect 552 10288 31072 10310
rect 1302 10248 1308 10260
rect 1044 10220 1308 10248
rect 934 10072 940 10124
rect 992 10112 998 10124
rect 1044 10121 1072 10220
rect 1302 10208 1308 10220
rect 1360 10208 1366 10260
rect 1495 10251 1553 10257
rect 1495 10217 1507 10251
rect 1541 10248 1553 10251
rect 1762 10248 1768 10260
rect 1541 10220 1768 10248
rect 1541 10217 1553 10220
rect 1495 10211 1553 10217
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 3050 10208 3056 10260
rect 3108 10208 3114 10260
rect 3703 10251 3761 10257
rect 3703 10217 3715 10251
rect 3749 10248 3761 10251
rect 4062 10248 4068 10260
rect 3749 10220 4068 10248
rect 3749 10217 3761 10220
rect 3703 10211 3761 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4890 10208 4896 10260
rect 4948 10248 4954 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 4948 10220 5457 10248
rect 4948 10208 4954 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 9030 10248 9036 10260
rect 5445 10211 5503 10217
rect 5644 10220 9036 10248
rect 1029 10115 1087 10121
rect 1029 10112 1041 10115
rect 992 10084 1041 10112
rect 992 10072 998 10084
rect 1029 10081 1041 10084
rect 1075 10081 1087 10115
rect 1029 10075 1087 10081
rect 2958 10072 2964 10124
rect 3016 10072 3022 10124
rect 3068 10112 3096 10208
rect 3068 10084 3372 10112
rect 1525 10065 1583 10071
rect 1525 10062 1537 10065
rect 1504 10056 1537 10062
rect 1486 10004 1492 10056
rect 1571 10031 1583 10065
rect 1544 10025 1583 10031
rect 1765 10047 1823 10053
rect 1544 10004 1550 10025
rect 1765 10013 1777 10047
rect 1811 10044 1823 10047
rect 1854 10044 1860 10056
rect 1811 10016 1860 10044
rect 1811 10013 1823 10016
rect 1765 10007 1823 10013
rect 1854 10004 1860 10016
rect 1912 10004 1918 10056
rect 2976 10044 3004 10072
rect 3234 10044 3240 10056
rect 2976 10016 3240 10044
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 3344 10044 3372 10084
rect 3786 10072 3792 10124
rect 3844 10112 3850 10124
rect 5644 10121 5672 10220
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9131 10251 9189 10257
rect 9131 10217 9143 10251
rect 9177 10248 9189 10251
rect 9306 10248 9312 10260
rect 9177 10220 9312 10248
rect 9177 10217 9189 10220
rect 9131 10211 9189 10217
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 13538 10248 13544 10260
rect 9732 10220 13544 10248
rect 9732 10208 9738 10220
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 14274 10208 14280 10260
rect 14332 10257 14338 10260
rect 14332 10248 14341 10257
rect 14332 10220 14377 10248
rect 14332 10211 14341 10220
rect 14332 10208 14338 10211
rect 17862 10208 17868 10260
rect 17920 10257 17926 10260
rect 17920 10248 17929 10257
rect 17920 10220 17965 10248
rect 17920 10211 17929 10220
rect 17920 10208 17926 10211
rect 18414 10208 18420 10260
rect 18472 10248 18478 10260
rect 19245 10251 19303 10257
rect 19245 10248 19257 10251
rect 18472 10220 19257 10248
rect 18472 10208 18478 10220
rect 19245 10217 19257 10220
rect 19291 10217 19303 10251
rect 19245 10211 19303 10217
rect 20346 10208 20352 10260
rect 20404 10208 20410 10260
rect 22278 10248 22284 10260
rect 20916 10220 22284 10248
rect 6546 10180 6552 10192
rect 6012 10152 6552 10180
rect 3973 10115 4031 10121
rect 3973 10112 3985 10115
rect 3844 10084 3985 10112
rect 3844 10072 3850 10084
rect 3973 10081 3985 10084
rect 4019 10081 4031 10115
rect 3973 10075 4031 10081
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10081 5687 10115
rect 5629 10075 5687 10081
rect 5915 10115 5973 10121
rect 5915 10081 5927 10115
rect 5961 10112 5973 10115
rect 6012 10112 6040 10152
rect 6546 10140 6552 10152
rect 6604 10140 6610 10192
rect 13446 10140 13452 10192
rect 13504 10140 13510 10192
rect 16209 10183 16267 10189
rect 16209 10149 16221 10183
rect 16255 10180 16267 10183
rect 20438 10180 20444 10192
rect 16255 10152 16988 10180
rect 16255 10149 16267 10152
rect 16209 10143 16267 10149
rect 5961 10084 6040 10112
rect 5961 10081 5973 10084
rect 5915 10075 5973 10081
rect 3700 10047 3758 10053
rect 3700 10044 3712 10047
rect 3344 10016 3712 10044
rect 3700 10013 3712 10016
rect 3746 10013 3758 10047
rect 3700 10007 3758 10013
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 5644 10044 5672 10075
rect 6086 10072 6092 10124
rect 6144 10112 6150 10124
rect 6181 10115 6239 10121
rect 6181 10112 6193 10115
rect 6144 10084 6193 10112
rect 6144 10072 6150 10084
rect 6181 10081 6193 10084
rect 6227 10081 6239 10115
rect 7650 10112 7656 10124
rect 6181 10075 6239 10081
rect 6288 10084 6684 10112
rect 4672 10016 5672 10044
rect 4672 10004 4678 10016
rect 2590 9936 2596 9988
rect 2648 9976 2654 9988
rect 6288 9976 6316 10084
rect 6656 10056 6684 10084
rect 7116 10084 7656 10112
rect 6362 10004 6368 10056
rect 6420 10044 6426 10056
rect 6457 10047 6515 10053
rect 6457 10044 6469 10047
rect 6420 10016 6469 10044
rect 6420 10004 6426 10016
rect 6457 10013 6469 10016
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 2648 9948 3280 9976
rect 2648 9936 2654 9948
rect 3050 9868 3056 9920
rect 3108 9868 3114 9920
rect 3252 9908 3280 9948
rect 4632 9948 6316 9976
rect 4632 9908 4660 9948
rect 3252 9880 4660 9908
rect 5261 9911 5319 9917
rect 5261 9877 5273 9911
rect 5307 9908 5319 9911
rect 5902 9908 5908 9920
rect 5307 9880 5908 9908
rect 5307 9877 5319 9880
rect 5261 9871 5319 9877
rect 5902 9868 5908 9880
rect 5960 9868 5966 9920
rect 6472 9908 6500 10007
rect 6638 10004 6644 10056
rect 6696 10004 6702 10056
rect 6822 10053 6828 10056
rect 6784 10047 6828 10053
rect 6784 10013 6796 10047
rect 6784 10007 6828 10013
rect 6822 10004 6828 10007
rect 6880 10004 6886 10056
rect 6963 10047 7021 10053
rect 6963 10013 6975 10047
rect 7009 10044 7021 10047
rect 7116 10044 7144 10084
rect 7650 10072 7656 10084
rect 7708 10072 7714 10124
rect 8573 10115 8631 10121
rect 8573 10081 8585 10115
rect 8619 10112 8631 10115
rect 9401 10115 9459 10121
rect 8619 10096 9112 10112
rect 8619 10084 9171 10096
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 9084 10071 9171 10084
rect 9401 10081 9413 10115
rect 9447 10112 9459 10115
rect 10594 10112 10600 10124
rect 9447 10084 10600 10112
rect 9447 10081 9459 10084
rect 9401 10075 9459 10081
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 13078 10112 13084 10124
rect 10796 10084 13084 10112
rect 9084 10068 9186 10071
rect 9128 10065 9186 10068
rect 7009 10016 7144 10044
rect 7193 10047 7251 10053
rect 7009 10013 7021 10016
rect 6963 10007 7021 10013
rect 7193 10013 7205 10047
rect 7239 10044 7251 10047
rect 8386 10044 8392 10056
rect 7239 10016 8392 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 8662 10004 8668 10056
rect 8720 10044 8726 10056
rect 8938 10044 8944 10056
rect 8720 10016 8944 10044
rect 8720 10004 8726 10016
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9128 10031 9140 10065
rect 9174 10031 9186 10065
rect 10796 10056 10824 10084
rect 13078 10072 13084 10084
rect 13136 10072 13142 10124
rect 13464 10112 13492 10140
rect 13725 10115 13783 10121
rect 13725 10112 13737 10115
rect 13464 10084 13737 10112
rect 13725 10081 13737 10084
rect 13771 10081 13783 10115
rect 13725 10075 13783 10081
rect 13817 10115 13875 10121
rect 13817 10081 13829 10115
rect 13863 10112 13875 10115
rect 13906 10112 13912 10124
rect 13863 10084 13912 10112
rect 13863 10081 13875 10084
rect 13817 10075 13875 10081
rect 13906 10072 13912 10084
rect 13964 10072 13970 10124
rect 16850 10072 16856 10124
rect 16908 10072 16914 10124
rect 9128 10025 9186 10031
rect 9582 10004 9588 10056
rect 9640 10044 9646 10056
rect 10778 10044 10784 10056
rect 9640 10016 10784 10044
rect 9640 10004 9646 10016
rect 10778 10004 10784 10016
rect 10836 10004 10842 10056
rect 11146 10004 11152 10056
rect 11204 10004 11210 10056
rect 11514 10053 11520 10056
rect 11476 10047 11520 10053
rect 11476 10013 11488 10047
rect 11476 10007 11520 10013
rect 11514 10004 11520 10007
rect 11572 10004 11578 10056
rect 11606 10004 11612 10056
rect 11664 10004 11670 10056
rect 11698 10004 11704 10056
rect 11756 10044 11762 10056
rect 11885 10047 11943 10053
rect 11885 10044 11897 10047
rect 11756 10016 11897 10044
rect 11756 10004 11762 10016
rect 11885 10013 11897 10016
rect 11931 10013 11943 10047
rect 14280 10047 14338 10053
rect 14280 10044 14292 10047
rect 11885 10007 11943 10013
rect 13740 10016 14292 10044
rect 13740 9988 13768 10016
rect 14280 10013 14292 10016
rect 14326 10013 14338 10047
rect 14280 10007 14338 10013
rect 14550 10004 14556 10056
rect 14608 10004 14614 10056
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10044 15991 10047
rect 16666 10044 16672 10056
rect 15979 10016 16672 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 13722 9936 13728 9988
rect 13780 9936 13786 9988
rect 7650 9908 7656 9920
rect 6472 9880 7656 9908
rect 7650 9868 7656 9880
rect 7708 9868 7714 9920
rect 9030 9868 9036 9920
rect 9088 9908 9094 9920
rect 9582 9908 9588 9920
rect 9088 9880 9588 9908
rect 9088 9868 9094 9880
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 10689 9911 10747 9917
rect 10689 9877 10701 9911
rect 10735 9908 10747 9911
rect 11054 9908 11060 9920
rect 10735 9880 11060 9908
rect 10735 9877 10747 9880
rect 10689 9871 10747 9877
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 12342 9868 12348 9920
rect 12400 9908 12406 9920
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12400 9880 13001 9908
rect 12400 9868 12406 9880
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 12989 9871 13047 9877
rect 13541 9911 13599 9917
rect 13541 9877 13553 9911
rect 13587 9908 13599 9911
rect 14550 9908 14556 9920
rect 13587 9880 14556 9908
rect 13587 9877 13599 9880
rect 13541 9871 13599 9877
rect 14550 9868 14556 9880
rect 14608 9868 14614 9920
rect 16482 9868 16488 9920
rect 16540 9868 16546 9920
rect 16960 9908 16988 10152
rect 18800 10152 20444 10180
rect 18800 10124 18828 10152
rect 20438 10140 20444 10152
rect 20496 10140 20502 10192
rect 17126 10072 17132 10124
rect 17184 10112 17190 10124
rect 18141 10115 18199 10121
rect 18141 10112 18153 10115
rect 17184 10084 18153 10112
rect 17184 10072 17190 10084
rect 18141 10081 18153 10084
rect 18187 10081 18199 10115
rect 18141 10075 18199 10081
rect 18782 10072 18788 10124
rect 18840 10072 18846 10124
rect 19797 10115 19855 10121
rect 19797 10081 19809 10115
rect 19843 10112 19855 10115
rect 19886 10112 19892 10124
rect 19843 10084 19892 10112
rect 19843 10081 19855 10084
rect 19797 10075 19855 10081
rect 19886 10072 19892 10084
rect 19944 10072 19950 10124
rect 20533 10115 20591 10121
rect 20533 10081 20545 10115
rect 20579 10081 20591 10115
rect 20533 10075 20591 10081
rect 17037 10047 17095 10053
rect 17037 10013 17049 10047
rect 17083 10044 17095 10047
rect 17218 10044 17224 10056
rect 17083 10016 17224 10044
rect 17083 10013 17095 10016
rect 17037 10007 17095 10013
rect 17218 10004 17224 10016
rect 17276 10004 17282 10056
rect 17402 10004 17408 10056
rect 17460 10004 17466 10056
rect 17911 10047 17969 10053
rect 17911 10013 17923 10047
rect 17957 10044 17969 10047
rect 19242 10044 19248 10056
rect 17957 10016 19248 10044
rect 17957 10013 17969 10016
rect 17911 10007 17969 10013
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 20548 10044 20576 10075
rect 20622 10072 20628 10124
rect 20680 10112 20686 10124
rect 20809 10115 20867 10121
rect 20809 10112 20821 10115
rect 20680 10084 20821 10112
rect 20680 10072 20686 10084
rect 20809 10081 20821 10084
rect 20855 10112 20867 10115
rect 20916 10112 20944 10220
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 23293 10251 23351 10257
rect 23293 10217 23305 10251
rect 23339 10248 23351 10251
rect 23934 10248 23940 10260
rect 23339 10220 23940 10248
rect 23339 10217 23351 10220
rect 23293 10211 23351 10217
rect 23934 10208 23940 10220
rect 23992 10208 23998 10260
rect 24210 10208 24216 10260
rect 24268 10248 24274 10260
rect 24268 10220 26096 10248
rect 24268 10208 24274 10220
rect 26068 10180 26096 10220
rect 26142 10208 26148 10260
rect 26200 10208 26206 10260
rect 26510 10208 26516 10260
rect 26568 10248 26574 10260
rect 26887 10251 26945 10257
rect 26887 10248 26899 10251
rect 26568 10220 26899 10248
rect 26568 10208 26574 10220
rect 26887 10217 26899 10220
rect 26933 10217 26945 10251
rect 26887 10211 26945 10217
rect 26326 10180 26332 10192
rect 26068 10152 26332 10180
rect 26326 10140 26332 10152
rect 26384 10140 26390 10192
rect 20855 10084 20944 10112
rect 20855 10081 20867 10084
rect 20809 10075 20867 10081
rect 20990 10072 20996 10124
rect 21048 10112 21054 10124
rect 21085 10115 21143 10121
rect 21085 10112 21097 10115
rect 21048 10084 21097 10112
rect 21048 10072 21054 10084
rect 21085 10081 21097 10084
rect 21131 10081 21143 10115
rect 21085 10075 21143 10081
rect 21266 10072 21272 10124
rect 21324 10072 21330 10124
rect 21596 10115 21654 10121
rect 21596 10112 21608 10115
rect 21468 10084 21608 10112
rect 21008 10044 21036 10072
rect 21468 10056 21496 10084
rect 21596 10081 21608 10084
rect 21642 10081 21654 10115
rect 21596 10075 21654 10081
rect 21910 10072 21916 10124
rect 21968 10072 21974 10124
rect 22005 10115 22063 10121
rect 22005 10081 22017 10115
rect 22051 10112 22063 10115
rect 22370 10112 22376 10124
rect 22051 10084 22376 10112
rect 22051 10081 22063 10084
rect 22005 10075 22063 10081
rect 22370 10072 22376 10084
rect 22428 10072 22434 10124
rect 24448 10115 24506 10121
rect 24448 10112 24460 10115
rect 24044 10084 24460 10112
rect 20548 10016 21036 10044
rect 21174 10004 21180 10056
rect 21232 10004 21238 10056
rect 21450 10004 21456 10056
rect 21508 10004 21514 10056
rect 21775 10047 21833 10053
rect 21775 10013 21787 10047
rect 21821 10044 21833 10047
rect 21928 10044 21956 10072
rect 21821 10016 21956 10044
rect 21821 10013 21833 10016
rect 21775 10007 21833 10013
rect 20625 9979 20683 9985
rect 20625 9945 20637 9979
rect 20671 9976 20683 9979
rect 21192 9976 21220 10004
rect 20671 9948 21220 9976
rect 20671 9945 20683 9948
rect 20625 9939 20683 9945
rect 19150 9908 19156 9920
rect 16960 9880 19156 9908
rect 19150 9868 19156 9880
rect 19208 9868 19214 9920
rect 19613 9911 19671 9917
rect 19613 9877 19625 9911
rect 19659 9908 19671 9911
rect 19702 9908 19708 9920
rect 19659 9880 19708 9908
rect 19659 9877 19671 9880
rect 19613 9871 19671 9877
rect 19702 9868 19708 9880
rect 19760 9868 19766 9920
rect 20898 9868 20904 9920
rect 20956 9868 20962 9920
rect 21542 9868 21548 9920
rect 21600 9908 21606 9920
rect 24044 9908 24072 10084
rect 24448 10081 24460 10084
rect 24494 10081 24506 10115
rect 24448 10075 24506 10081
rect 24780 10084 25084 10112
rect 24118 10004 24124 10056
rect 24176 10004 24182 10056
rect 24627 10047 24685 10053
rect 24627 10013 24639 10047
rect 24673 10044 24685 10047
rect 24780 10044 24808 10084
rect 25056 10056 25084 10084
rect 25774 10072 25780 10124
rect 25832 10112 25838 10124
rect 25832 10084 27752 10112
rect 25832 10072 25838 10084
rect 24673 10016 24808 10044
rect 24673 10013 24685 10016
rect 24627 10007 24685 10013
rect 24854 10004 24860 10056
rect 24912 10004 24918 10056
rect 25038 10004 25044 10056
rect 25096 10004 25102 10056
rect 26050 10004 26056 10056
rect 26108 10004 26114 10056
rect 26234 10004 26240 10056
rect 26292 10044 26298 10056
rect 26421 10047 26479 10053
rect 26421 10044 26433 10047
rect 26292 10016 26433 10044
rect 26292 10004 26298 10016
rect 26421 10013 26433 10016
rect 26467 10013 26479 10047
rect 26421 10007 26479 10013
rect 26878 10004 26884 10056
rect 26936 10004 26942 10056
rect 27157 10047 27215 10053
rect 27157 10013 27169 10047
rect 27203 10044 27215 10047
rect 27614 10044 27620 10056
rect 27203 10016 27620 10044
rect 27203 10013 27215 10016
rect 27157 10007 27215 10013
rect 27614 10004 27620 10016
rect 27672 10004 27678 10056
rect 27724 10044 27752 10084
rect 28626 10072 28632 10124
rect 28684 10072 28690 10124
rect 28905 10115 28963 10121
rect 28905 10081 28917 10115
rect 28951 10081 28963 10115
rect 28905 10075 28963 10081
rect 28920 10044 28948 10075
rect 29638 10072 29644 10124
rect 29696 10112 29702 10124
rect 30377 10115 30435 10121
rect 30377 10112 30389 10115
rect 29696 10084 30389 10112
rect 29696 10072 29702 10084
rect 30377 10081 30389 10084
rect 30423 10081 30435 10115
rect 30377 10075 30435 10081
rect 27724 10016 28948 10044
rect 24946 9908 24952 9920
rect 21600 9880 24952 9908
rect 21600 9868 21606 9880
rect 24946 9868 24952 9880
rect 25004 9868 25010 9920
rect 26068 9908 26096 10004
rect 30469 9979 30527 9985
rect 30469 9976 30481 9979
rect 28092 9948 28396 9976
rect 28092 9908 28120 9948
rect 26068 9880 28120 9908
rect 28166 9868 28172 9920
rect 28224 9908 28230 9920
rect 28261 9911 28319 9917
rect 28261 9908 28273 9911
rect 28224 9880 28273 9908
rect 28224 9868 28230 9880
rect 28261 9877 28273 9880
rect 28307 9877 28319 9911
rect 28368 9908 28396 9948
rect 29564 9948 30481 9976
rect 29564 9908 29592 9948
rect 30469 9945 30481 9948
rect 30515 9945 30527 9979
rect 30469 9939 30527 9945
rect 28368 9880 29592 9908
rect 28261 9871 28319 9877
rect 30006 9868 30012 9920
rect 30064 9868 30070 9920
rect 552 9818 30912 9840
rect 552 9766 4193 9818
rect 4245 9766 4257 9818
rect 4309 9766 4321 9818
rect 4373 9766 4385 9818
rect 4437 9766 4449 9818
rect 4501 9766 11783 9818
rect 11835 9766 11847 9818
rect 11899 9766 11911 9818
rect 11963 9766 11975 9818
rect 12027 9766 12039 9818
rect 12091 9766 19373 9818
rect 19425 9766 19437 9818
rect 19489 9766 19501 9818
rect 19553 9766 19565 9818
rect 19617 9766 19629 9818
rect 19681 9766 26963 9818
rect 27015 9766 27027 9818
rect 27079 9766 27091 9818
rect 27143 9766 27155 9818
rect 27207 9766 27219 9818
rect 27271 9766 30912 9818
rect 552 9744 30912 9766
rect 5813 9707 5871 9713
rect 3344 9676 4752 9704
rect 3344 9636 3372 9676
rect 2746 9608 3372 9636
rect 4724 9636 4752 9676
rect 5813 9673 5825 9707
rect 5859 9673 5871 9707
rect 6638 9704 6644 9716
rect 5813 9667 5871 9673
rect 6104 9676 6644 9704
rect 5166 9636 5172 9648
rect 4724 9608 5172 9636
rect 934 9528 940 9580
rect 992 9528 998 9580
rect 1443 9571 1501 9577
rect 1443 9537 1455 9571
rect 1489 9568 1501 9571
rect 2746 9568 2774 9608
rect 5166 9596 5172 9608
rect 5224 9596 5230 9648
rect 5828 9636 5856 9667
rect 6104 9636 6132 9676
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 6822 9664 6828 9716
rect 6880 9704 6886 9716
rect 7006 9704 7012 9716
rect 6880 9676 7012 9704
rect 6880 9664 6886 9676
rect 7006 9664 7012 9676
rect 7064 9664 7070 9716
rect 8938 9664 8944 9716
rect 8996 9704 9002 9716
rect 10686 9704 10692 9716
rect 8996 9676 10692 9704
rect 8996 9664 9002 9676
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 11606 9704 11612 9716
rect 11072 9676 11612 9704
rect 5276 9608 5856 9636
rect 6012 9608 6132 9636
rect 10965 9639 11023 9645
rect 1489 9540 2774 9568
rect 1489 9537 1501 9540
rect 1443 9531 1501 9537
rect 3050 9528 3056 9580
rect 3108 9568 3114 9580
rect 3792 9571 3850 9577
rect 3792 9568 3804 9571
rect 3108 9540 3804 9568
rect 3108 9528 3114 9540
rect 3792 9537 3804 9540
rect 3838 9537 3850 9571
rect 3792 9531 3850 9537
rect 3970 9528 3976 9580
rect 4028 9568 4034 9580
rect 4028 9540 4200 9568
rect 4028 9528 4034 9540
rect 1670 9460 1676 9512
rect 1728 9460 1734 9512
rect 3234 9460 3240 9512
rect 3292 9500 3298 9512
rect 3329 9503 3387 9509
rect 3329 9500 3341 9503
rect 3292 9472 3341 9500
rect 3292 9460 3298 9472
rect 3329 9469 3341 9472
rect 3375 9469 3387 9503
rect 3329 9463 3387 9469
rect 3602 9460 3608 9512
rect 3660 9500 3666 9512
rect 4065 9503 4123 9509
rect 4065 9500 4077 9503
rect 3660 9472 4077 9500
rect 3660 9460 3666 9472
rect 4065 9469 4077 9472
rect 4111 9469 4123 9503
rect 4172 9500 4200 9540
rect 4982 9528 4988 9580
rect 5040 9568 5046 9580
rect 5276 9568 5304 9608
rect 5040 9540 5304 9568
rect 5445 9571 5503 9577
rect 5040 9528 5046 9540
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 5810 9568 5816 9580
rect 5491 9540 5816 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 5810 9528 5816 9540
rect 5868 9528 5874 9580
rect 6012 9509 6040 9608
rect 10965 9605 10977 9639
rect 11011 9636 11023 9639
rect 11072 9636 11100 9676
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 17126 9704 17132 9716
rect 16408 9676 17132 9704
rect 11011 9608 11100 9636
rect 13541 9639 13599 9645
rect 11011 9605 11023 9608
rect 10965 9599 11023 9605
rect 13541 9605 13553 9639
rect 13587 9605 13599 9639
rect 13541 9599 13599 9605
rect 16117 9639 16175 9645
rect 16117 9605 16129 9639
rect 16163 9636 16175 9639
rect 16408 9636 16436 9676
rect 17126 9664 17132 9676
rect 17184 9664 17190 9716
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 21082 9704 21088 9716
rect 20772 9676 21088 9704
rect 20772 9664 20778 9676
rect 21082 9664 21088 9676
rect 21140 9664 21146 9716
rect 21358 9664 21364 9716
rect 21416 9704 21422 9716
rect 22741 9707 22799 9713
rect 22741 9704 22753 9707
rect 21416 9676 22753 9704
rect 21416 9664 21422 9676
rect 22741 9673 22753 9676
rect 22787 9673 22799 9707
rect 22741 9667 22799 9673
rect 24854 9664 24860 9716
rect 24912 9704 24918 9716
rect 26605 9707 26663 9713
rect 24912 9676 26280 9704
rect 24912 9664 24918 9676
rect 24486 9636 24492 9648
rect 16163 9608 16436 9636
rect 23676 9608 24492 9636
rect 16163 9605 16175 9608
rect 16117 9599 16175 9605
rect 6089 9571 6147 9577
rect 6089 9537 6101 9571
rect 6135 9568 6147 9571
rect 6362 9568 6368 9580
rect 6135 9540 6368 9568
rect 6135 9537 6147 9540
rect 6089 9531 6147 9537
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 6595 9571 6653 9577
rect 6595 9537 6607 9571
rect 6641 9568 6653 9571
rect 6641 9540 6960 9568
rect 6641 9537 6653 9540
rect 6595 9531 6653 9537
rect 6932 9512 6960 9540
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 9306 9577 9312 9580
rect 8941 9571 8999 9577
rect 8941 9568 8953 9571
rect 8720 9540 8953 9568
rect 8720 9528 8726 9540
rect 8941 9537 8953 9540
rect 8987 9537 8999 9571
rect 8941 9531 8999 9537
rect 9268 9571 9312 9577
rect 9268 9537 9280 9571
rect 9268 9531 9312 9537
rect 5721 9503 5779 9509
rect 4172 9472 5672 9500
rect 4065 9463 4123 9469
rect 5350 9432 5356 9444
rect 4724 9404 5356 9432
rect 1403 9367 1461 9373
rect 1403 9333 1415 9367
rect 1449 9364 1461 9367
rect 1762 9364 1768 9376
rect 1449 9336 1768 9364
rect 1449 9333 1461 9336
rect 1403 9327 1461 9333
rect 1762 9324 1768 9336
rect 1820 9324 1826 9376
rect 2961 9367 3019 9373
rect 2961 9333 2973 9367
rect 3007 9364 3019 9367
rect 3602 9364 3608 9376
rect 3007 9336 3608 9364
rect 3007 9333 3019 9336
rect 2961 9327 3019 9333
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 3795 9367 3853 9373
rect 3795 9333 3807 9367
rect 3841 9364 3853 9367
rect 4062 9364 4068 9376
rect 3841 9336 4068 9364
rect 3841 9333 3853 9336
rect 3795 9327 3853 9333
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4338 9324 4344 9376
rect 4396 9364 4402 9376
rect 4724 9364 4752 9404
rect 5350 9392 5356 9404
rect 5408 9392 5414 9444
rect 4396 9336 4752 9364
rect 4396 9324 4402 9336
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 4856 9336 5549 9364
rect 4856 9324 4862 9336
rect 5537 9333 5549 9336
rect 5583 9333 5595 9367
rect 5644 9364 5672 9472
rect 5721 9469 5733 9503
rect 5767 9469 5779 9503
rect 5721 9463 5779 9469
rect 5997 9503 6055 9509
rect 5997 9469 6009 9503
rect 6043 9469 6055 9503
rect 5997 9463 6055 9469
rect 5736 9432 5764 9463
rect 6822 9460 6828 9512
rect 6880 9460 6886 9512
rect 6914 9460 6920 9512
rect 6972 9460 6978 9512
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 8478 9500 8484 9512
rect 8435 9472 8484 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 8956 9500 8984 9531
rect 9306 9528 9312 9531
rect 9364 9528 9370 9580
rect 9490 9577 9496 9580
rect 9447 9571 9496 9577
rect 9447 9537 9459 9571
rect 9493 9537 9496 9571
rect 9447 9531 9496 9537
rect 9490 9528 9496 9531
rect 9548 9528 9554 9580
rect 9608 9540 9812 9568
rect 9608 9500 9636 9540
rect 9784 9512 9812 9540
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 11612 9571 11670 9577
rect 11612 9568 11624 9571
rect 11112 9540 11624 9568
rect 11112 9528 11118 9540
rect 11612 9537 11624 9540
rect 11658 9537 11670 9571
rect 13556 9568 13584 9599
rect 14366 9577 14372 9580
rect 14323 9571 14372 9577
rect 13556 9540 14050 9568
rect 11612 9531 11670 9537
rect 8956 9472 9636 9500
rect 9674 9460 9680 9512
rect 9732 9460 9738 9512
rect 9766 9460 9772 9512
rect 9824 9460 9830 9512
rect 11146 9460 11152 9512
rect 11204 9460 11210 9512
rect 11514 9509 11520 9512
rect 11476 9503 11520 9509
rect 11476 9469 11488 9503
rect 11476 9463 11520 9469
rect 11514 9460 11520 9463
rect 11572 9460 11578 9512
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9500 11943 9503
rect 12158 9500 12164 9512
rect 11931 9472 12164 9500
rect 11931 9469 11943 9472
rect 11885 9463 11943 9469
rect 12158 9460 12164 9472
rect 12216 9460 12222 9512
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9469 13783 9503
rect 13725 9463 13783 9469
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9500 13875 9503
rect 13906 9500 13912 9512
rect 13863 9472 13912 9500
rect 13863 9469 13875 9472
rect 13817 9463 13875 9469
rect 6178 9432 6184 9444
rect 5736 9404 6184 9432
rect 6178 9392 6184 9404
rect 6236 9392 6242 9444
rect 7558 9392 7564 9444
rect 7616 9432 7622 9444
rect 8205 9435 8263 9441
rect 7616 9404 7880 9432
rect 7616 9392 7622 9404
rect 6362 9364 6368 9376
rect 5644 9336 6368 9364
rect 5537 9327 5595 9333
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 6555 9367 6613 9373
rect 6555 9333 6567 9367
rect 6601 9364 6613 9367
rect 7098 9364 7104 9376
rect 6601 9336 7104 9364
rect 6601 9333 6613 9336
rect 6555 9327 6613 9333
rect 7098 9324 7104 9336
rect 7156 9364 7162 9376
rect 7742 9364 7748 9376
rect 7156 9336 7748 9364
rect 7156 9324 7162 9336
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 7852 9364 7880 9404
rect 8205 9401 8217 9435
rect 8251 9432 8263 9435
rect 9030 9432 9036 9444
rect 8251 9404 9036 9432
rect 8251 9401 8263 9404
rect 8205 9395 8263 9401
rect 9030 9392 9036 9404
rect 9088 9392 9094 9444
rect 13740 9432 13768 9463
rect 13906 9460 13912 9472
rect 13964 9460 13970 9512
rect 14022 9500 14050 9540
rect 14323 9537 14335 9571
rect 14369 9537 14372 9571
rect 14323 9531 14372 9537
rect 14366 9528 14372 9531
rect 14424 9528 14430 9580
rect 16390 9568 16396 9580
rect 16040 9540 16396 9568
rect 16040 9512 16068 9540
rect 16390 9528 16396 9540
rect 16448 9528 16454 9580
rect 16574 9528 16580 9580
rect 16632 9568 16638 9580
rect 16856 9571 16914 9577
rect 16856 9568 16868 9571
rect 16632 9540 16868 9568
rect 16632 9528 16638 9540
rect 16856 9537 16868 9540
rect 16902 9537 16914 9571
rect 17770 9568 17776 9580
rect 16856 9531 16914 9537
rect 17144 9540 17776 9568
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 14022 9472 14565 9500
rect 14553 9469 14565 9472
rect 14599 9469 14611 9503
rect 14553 9463 14611 9469
rect 16022 9460 16028 9512
rect 16080 9460 16086 9512
rect 16301 9503 16359 9509
rect 16301 9469 16313 9503
rect 16347 9469 16359 9503
rect 16301 9463 16359 9469
rect 16720 9503 16778 9509
rect 16720 9469 16732 9503
rect 16766 9500 16778 9503
rect 16942 9500 16948 9512
rect 16766 9472 16948 9500
rect 16766 9469 16778 9472
rect 16720 9463 16778 9469
rect 16316 9432 16344 9463
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17144 9509 17172 9540
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 19199 9571 19257 9577
rect 19199 9537 19211 9571
rect 19245 9568 19257 9571
rect 20714 9568 20720 9580
rect 19245 9540 20720 9568
rect 19245 9537 19257 9540
rect 19199 9531 19257 9537
rect 20714 9528 20720 9540
rect 20772 9528 20778 9580
rect 20806 9528 20812 9580
rect 20864 9528 20870 9580
rect 21407 9571 21465 9577
rect 21407 9537 21419 9571
rect 21453 9568 21465 9571
rect 22738 9568 22744 9580
rect 21453 9540 22744 9568
rect 21453 9537 21465 9540
rect 21407 9531 21465 9537
rect 22738 9528 22744 9540
rect 22796 9528 22802 9580
rect 17129 9503 17187 9509
rect 17129 9469 17141 9503
rect 17175 9469 17187 9503
rect 17129 9463 17187 9469
rect 17402 9460 17408 9512
rect 17460 9500 17466 9512
rect 18693 9503 18751 9509
rect 18693 9500 18705 9503
rect 17460 9472 18705 9500
rect 17460 9460 17466 9472
rect 18693 9469 18705 9472
rect 18739 9500 18751 9503
rect 19334 9500 19340 9512
rect 18739 9472 19340 9500
rect 18739 9469 18751 9472
rect 18693 9463 18751 9469
rect 19334 9460 19340 9472
rect 19392 9460 19398 9512
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9500 19487 9503
rect 19702 9500 19708 9512
rect 19475 9472 19708 9500
rect 19475 9469 19487 9472
rect 19429 9463 19487 9469
rect 19702 9460 19708 9472
rect 19760 9460 19766 9512
rect 20901 9503 20959 9509
rect 20901 9469 20913 9503
rect 20947 9469 20959 9503
rect 20901 9463 20959 9469
rect 12912 9404 13768 9432
rect 8573 9367 8631 9373
rect 8573 9364 8585 9367
rect 7852 9336 8585 9364
rect 8573 9333 8585 9336
rect 8619 9333 8631 9367
rect 8573 9327 8631 9333
rect 8662 9324 8668 9376
rect 8720 9364 8726 9376
rect 12912 9364 12940 9404
rect 13740 9376 13768 9404
rect 15212 9404 16344 9432
rect 8720 9336 12940 9364
rect 8720 9324 8726 9336
rect 12986 9324 12992 9376
rect 13044 9324 13050 9376
rect 13722 9324 13728 9376
rect 13780 9324 13786 9376
rect 14274 9324 14280 9376
rect 14332 9373 14338 9376
rect 14332 9364 14341 9373
rect 14332 9336 14377 9364
rect 14332 9327 14341 9336
rect 14332 9324 14338 9327
rect 14642 9324 14648 9376
rect 14700 9364 14706 9376
rect 15212 9364 15240 9404
rect 14700 9336 15240 9364
rect 14700 9324 14706 9336
rect 15378 9324 15384 9376
rect 15436 9364 15442 9376
rect 15657 9367 15715 9373
rect 15657 9364 15669 9367
rect 15436 9336 15669 9364
rect 15436 9324 15442 9336
rect 15657 9333 15669 9336
rect 15703 9333 15715 9367
rect 16316 9364 16344 9404
rect 17862 9392 17868 9444
rect 17920 9432 17926 9444
rect 18509 9435 18567 9441
rect 17920 9404 18368 9432
rect 17920 9392 17926 9404
rect 17954 9364 17960 9376
rect 16316 9336 17960 9364
rect 15657 9327 15715 9333
rect 17954 9324 17960 9336
rect 18012 9364 18018 9376
rect 18138 9364 18144 9376
rect 18012 9336 18144 9364
rect 18012 9324 18018 9336
rect 18138 9324 18144 9336
rect 18196 9324 18202 9376
rect 18340 9364 18368 9404
rect 18509 9401 18521 9435
rect 18555 9432 18567 9435
rect 18782 9432 18788 9444
rect 18555 9404 18788 9432
rect 18555 9401 18567 9404
rect 18509 9395 18567 9401
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 20806 9392 20812 9444
rect 20864 9432 20870 9444
rect 20916 9432 20944 9463
rect 21634 9460 21640 9512
rect 21692 9460 21698 9512
rect 21910 9460 21916 9512
rect 21968 9500 21974 9512
rect 23676 9509 23704 9608
rect 24486 9596 24492 9608
rect 24544 9596 24550 9648
rect 26252 9636 26280 9676
rect 26605 9673 26617 9707
rect 26651 9704 26663 9707
rect 26878 9704 26884 9716
rect 26651 9676 26884 9704
rect 26651 9673 26663 9676
rect 26605 9667 26663 9673
rect 26878 9664 26884 9676
rect 26936 9664 26942 9716
rect 27614 9664 27620 9716
rect 27672 9664 27678 9716
rect 27982 9664 27988 9716
rect 28040 9664 28046 9716
rect 27433 9639 27491 9645
rect 27433 9636 27445 9639
rect 26252 9608 27445 9636
rect 27433 9605 27445 9608
rect 27479 9605 27491 9639
rect 27632 9636 27660 9664
rect 27709 9639 27767 9645
rect 27709 9636 27721 9639
rect 27632 9608 27721 9636
rect 27433 9599 27491 9605
rect 27709 9605 27721 9608
rect 27755 9605 27767 9639
rect 27709 9599 27767 9605
rect 24581 9571 24639 9577
rect 24581 9568 24593 9571
rect 24136 9540 24593 9568
rect 24136 9512 24164 9540
rect 24581 9537 24593 9540
rect 24627 9537 24639 9571
rect 24581 9531 24639 9537
rect 25087 9571 25145 9577
rect 25087 9537 25099 9571
rect 25133 9568 25145 9571
rect 27246 9568 27252 9580
rect 25133 9540 25268 9568
rect 25133 9537 25145 9540
rect 25087 9531 25145 9537
rect 25240 9512 25268 9540
rect 25976 9540 27252 9568
rect 25976 9512 26004 9540
rect 27246 9528 27252 9540
rect 27304 9528 27310 9580
rect 29178 9568 29184 9580
rect 27632 9540 29184 9568
rect 23661 9503 23719 9509
rect 21968 9472 23612 9500
rect 21968 9460 21974 9472
rect 20864 9404 20944 9432
rect 23584 9432 23612 9472
rect 23661 9469 23673 9503
rect 23707 9469 23719 9503
rect 23661 9463 23719 9469
rect 24029 9503 24087 9509
rect 24029 9469 24041 9503
rect 24075 9469 24087 9503
rect 24029 9463 24087 9469
rect 24044 9432 24072 9463
rect 24118 9460 24124 9512
rect 24176 9460 24182 9512
rect 24302 9460 24308 9512
rect 24360 9500 24366 9512
rect 24946 9509 24952 9512
rect 24908 9503 24952 9509
rect 24360 9472 24716 9500
rect 24360 9460 24366 9472
rect 24578 9432 24584 9444
rect 23584 9404 24584 9432
rect 20864 9392 20870 9404
rect 24578 9392 24584 9404
rect 24636 9392 24642 9444
rect 19159 9367 19217 9373
rect 19159 9364 19171 9367
rect 18340 9336 19171 9364
rect 19159 9333 19171 9336
rect 19205 9364 19217 9367
rect 21367 9367 21425 9373
rect 21367 9364 21379 9367
rect 19205 9336 21379 9364
rect 19205 9333 19217 9336
rect 19159 9327 19217 9333
rect 21367 9333 21379 9336
rect 21413 9364 21425 9367
rect 22002 9364 22008 9376
rect 21413 9336 22008 9364
rect 21413 9333 21425 9336
rect 21367 9327 21425 9333
rect 22002 9324 22008 9336
rect 22060 9324 22066 9376
rect 23477 9367 23535 9373
rect 23477 9333 23489 9367
rect 23523 9364 23535 9367
rect 23566 9364 23572 9376
rect 23523 9336 23572 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 23566 9324 23572 9336
rect 23624 9324 23630 9376
rect 23845 9367 23903 9373
rect 23845 9333 23857 9367
rect 23891 9364 23903 9367
rect 23934 9364 23940 9376
rect 23891 9336 23940 9364
rect 23891 9333 23903 9336
rect 23845 9327 23903 9333
rect 23934 9324 23940 9336
rect 23992 9324 23998 9376
rect 24121 9367 24179 9373
rect 24121 9333 24133 9367
rect 24167 9364 24179 9367
rect 24394 9364 24400 9376
rect 24167 9336 24400 9364
rect 24167 9333 24179 9336
rect 24121 9327 24179 9333
rect 24394 9324 24400 9336
rect 24452 9324 24458 9376
rect 24688 9364 24716 9472
rect 24908 9469 24920 9503
rect 24908 9463 24952 9469
rect 24946 9460 24952 9463
rect 25004 9460 25010 9512
rect 25222 9460 25228 9512
rect 25280 9460 25286 9512
rect 25317 9503 25375 9509
rect 25317 9469 25329 9503
rect 25363 9500 25375 9503
rect 25682 9500 25688 9512
rect 25363 9472 25688 9500
rect 25363 9469 25375 9472
rect 25317 9463 25375 9469
rect 25682 9460 25688 9472
rect 25740 9460 25746 9512
rect 25958 9460 25964 9512
rect 26016 9460 26022 9512
rect 26326 9460 26332 9512
rect 26384 9500 26390 9512
rect 27632 9509 27660 9540
rect 28184 9509 28212 9540
rect 29178 9528 29184 9540
rect 29236 9528 29242 9580
rect 27617 9503 27675 9509
rect 27617 9500 27629 9503
rect 26384 9472 27629 9500
rect 26384 9460 26390 9472
rect 27617 9469 27629 9472
rect 27663 9469 27675 9503
rect 27617 9463 27675 9469
rect 27893 9503 27951 9509
rect 27893 9469 27905 9503
rect 27939 9469 27951 9503
rect 27893 9463 27951 9469
rect 28169 9503 28227 9509
rect 28169 9469 28181 9503
rect 28215 9469 28227 9503
rect 28169 9463 28227 9469
rect 28445 9503 28503 9509
rect 28445 9469 28457 9503
rect 28491 9500 28503 9503
rect 28534 9500 28540 9512
rect 28491 9472 28540 9500
rect 28491 9469 28503 9472
rect 28445 9463 28503 9469
rect 26344 9364 26372 9460
rect 26786 9392 26792 9444
rect 26844 9432 26850 9444
rect 26973 9435 27031 9441
rect 26973 9432 26985 9435
rect 26844 9404 26985 9432
rect 26844 9392 26850 9404
rect 26973 9401 26985 9404
rect 27019 9432 27031 9435
rect 27798 9432 27804 9444
rect 27019 9404 27804 9432
rect 27019 9401 27031 9404
rect 26973 9395 27031 9401
rect 27798 9392 27804 9404
rect 27856 9392 27862 9444
rect 24688 9336 26372 9364
rect 27246 9324 27252 9376
rect 27304 9364 27310 9376
rect 27908 9364 27936 9463
rect 28460 9432 28488 9463
rect 28534 9460 28540 9472
rect 28592 9460 28598 9512
rect 28000 9404 28488 9432
rect 28000 9376 28028 9404
rect 27304 9336 27936 9364
rect 27304 9324 27310 9336
rect 27982 9324 27988 9376
rect 28040 9324 28046 9376
rect 28074 9324 28080 9376
rect 28132 9364 28138 9376
rect 28261 9367 28319 9373
rect 28261 9364 28273 9367
rect 28132 9336 28273 9364
rect 28132 9324 28138 9336
rect 28261 9333 28273 9336
rect 28307 9333 28319 9367
rect 28261 9327 28319 9333
rect 552 9274 31072 9296
rect 552 9222 7988 9274
rect 8040 9222 8052 9274
rect 8104 9222 8116 9274
rect 8168 9222 8180 9274
rect 8232 9222 8244 9274
rect 8296 9222 15578 9274
rect 15630 9222 15642 9274
rect 15694 9222 15706 9274
rect 15758 9222 15770 9274
rect 15822 9222 15834 9274
rect 15886 9222 23168 9274
rect 23220 9222 23232 9274
rect 23284 9222 23296 9274
rect 23348 9222 23360 9274
rect 23412 9222 23424 9274
rect 23476 9222 30758 9274
rect 30810 9222 30822 9274
rect 30874 9222 30886 9274
rect 30938 9222 30950 9274
rect 31002 9222 31014 9274
rect 31066 9222 31072 9274
rect 552 9200 31072 9222
rect 1302 9120 1308 9172
rect 1360 9160 1366 9172
rect 2222 9160 2228 9172
rect 1360 9132 2228 9160
rect 1360 9120 1366 9132
rect 2222 9120 2228 9132
rect 2280 9120 2286 9172
rect 3703 9163 3761 9169
rect 3703 9129 3715 9163
rect 3749 9160 3761 9163
rect 4062 9160 4068 9172
rect 3749 9132 4068 9160
rect 3749 9129 3761 9132
rect 3703 9123 3761 9129
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 5261 9163 5319 9169
rect 5261 9129 5273 9163
rect 5307 9160 5319 9163
rect 6270 9160 6276 9172
rect 5307 9132 6276 9160
rect 5307 9129 5319 9132
rect 5261 9123 5319 9129
rect 6270 9120 6276 9132
rect 6328 9120 6334 9172
rect 6362 9120 6368 9172
rect 6420 9160 6426 9172
rect 7098 9160 7104 9172
rect 6420 9132 7104 9160
rect 6420 9120 6426 9132
rect 7098 9120 7104 9132
rect 7156 9120 7162 9172
rect 7190 9120 7196 9172
rect 7248 9120 7254 9172
rect 7377 9163 7435 9169
rect 7377 9129 7389 9163
rect 7423 9129 7435 9163
rect 7377 9123 7435 9129
rect 3142 9052 3148 9104
rect 3200 9052 3206 9104
rect 7208 9092 7236 9120
rect 4632 9064 7236 9092
rect 7392 9092 7420 9123
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 8119 9163 8177 9169
rect 8119 9160 8131 9163
rect 7800 9132 8131 9160
rect 7800 9120 7806 9132
rect 8119 9129 8131 9132
rect 8165 9129 8177 9163
rect 8119 9123 8177 9129
rect 9490 9120 9496 9172
rect 9548 9120 9554 9172
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 10045 9163 10103 9169
rect 10045 9160 10057 9163
rect 9732 9132 10057 9160
rect 9732 9120 9738 9132
rect 10045 9129 10057 9132
rect 10091 9129 10103 9163
rect 10045 9123 10103 9129
rect 10597 9163 10655 9169
rect 10597 9129 10609 9163
rect 10643 9129 10655 9163
rect 10597 9123 10655 9129
rect 10612 9092 10640 9123
rect 11514 9120 11520 9172
rect 11572 9160 11578 9172
rect 11615 9163 11673 9169
rect 11615 9160 11627 9163
rect 11572 9132 11627 9160
rect 11572 9120 11578 9132
rect 11615 9129 11627 9132
rect 11661 9129 11673 9163
rect 11615 9123 11673 9129
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 16482 9160 16488 9172
rect 13780 9132 16488 9160
rect 13780 9120 13786 9132
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 17862 9160 17868 9172
rect 17920 9169 17926 9172
rect 17144 9132 17868 9160
rect 7392 9064 7788 9092
rect 10612 9064 11284 9092
rect 1394 9033 1400 9036
rect 1356 9027 1400 9033
rect 1356 8993 1368 9027
rect 1356 8987 1400 8993
rect 1394 8984 1400 8987
rect 1452 8984 1458 9036
rect 1762 8984 1768 9036
rect 1820 8984 1826 9036
rect 3786 8984 3792 9036
rect 3844 9024 3850 9036
rect 3973 9027 4031 9033
rect 3973 9024 3985 9027
rect 3844 8996 3985 9024
rect 3844 8984 3850 8996
rect 3973 8993 3985 8996
rect 4019 8993 4031 9027
rect 4632 9024 4660 9064
rect 3973 8987 4031 8993
rect 4080 8996 4660 9024
rect 1029 8959 1087 8965
rect 1029 8925 1041 8959
rect 1075 8956 1087 8959
rect 1210 8956 1216 8968
rect 1075 8928 1216 8956
rect 1075 8925 1087 8928
rect 1029 8919 1087 8925
rect 1210 8916 1216 8928
rect 1268 8916 1274 8968
rect 1535 8959 1593 8965
rect 1535 8925 1547 8959
rect 1581 8956 1593 8959
rect 1581 8928 2774 8956
rect 1581 8925 1593 8928
rect 1535 8919 1593 8925
rect 2746 8820 2774 8928
rect 3234 8916 3240 8968
rect 3292 8916 3298 8968
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 3700 8961 3758 8967
rect 3700 8956 3712 8961
rect 3660 8928 3712 8956
rect 3660 8916 3666 8928
rect 3700 8927 3712 8928
rect 3746 8927 3758 8961
rect 3700 8921 3758 8927
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 4080 8956 4108 8996
rect 5626 8984 5632 9036
rect 5684 8984 5690 9036
rect 5810 8984 5816 9036
rect 5868 8984 5874 9036
rect 6457 9027 6515 9033
rect 6457 9024 6469 9027
rect 6380 8996 6469 9024
rect 6380 8968 6408 8996
rect 6457 8993 6469 8996
rect 6503 8993 6515 9027
rect 6457 8987 6515 8993
rect 6638 8984 6644 9036
rect 6696 9024 6702 9036
rect 6917 9027 6975 9033
rect 6917 9024 6929 9027
rect 6696 8996 6929 9024
rect 6696 8984 6702 8996
rect 6917 8993 6929 8996
rect 6963 9024 6975 9027
rect 7006 9024 7012 9036
rect 6963 8996 7012 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 9024 7251 9027
rect 7282 9024 7288 9036
rect 7239 8996 7288 9024
rect 7239 8993 7251 8996
rect 7193 8987 7251 8993
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 7558 8984 7564 9036
rect 7616 8984 7622 9036
rect 7650 8984 7656 9036
rect 7708 8984 7714 9036
rect 7760 9024 7788 9064
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 7760 8996 8401 9024
rect 8389 8993 8401 8996
rect 8435 8993 8447 9027
rect 8389 8987 8447 8993
rect 9306 8984 9312 9036
rect 9364 9024 9370 9036
rect 10229 9027 10287 9033
rect 9364 8996 9812 9024
rect 9364 8984 9370 8996
rect 3936 8928 4108 8956
rect 3936 8916 3942 8928
rect 4430 8916 4436 8968
rect 4488 8956 4494 8968
rect 4488 8928 5112 8956
rect 4488 8916 4494 8928
rect 5084 8888 5112 8928
rect 5534 8916 5540 8968
rect 5592 8956 5598 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5592 8928 6009 8956
rect 5592 8916 5598 8928
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6362 8916 6368 8968
rect 6420 8956 6426 8968
rect 7466 8956 7472 8968
rect 6420 8928 7472 8956
rect 6420 8916 6426 8928
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 6641 8891 6699 8897
rect 6641 8888 6653 8891
rect 5084 8860 6653 8888
rect 6641 8857 6653 8860
rect 6687 8857 6699 8891
rect 6641 8851 6699 8857
rect 6730 8848 6736 8900
rect 6788 8848 6794 8900
rect 7576 8888 7604 8984
rect 9784 8968 9812 8996
rect 10229 8993 10241 9027
rect 10275 9024 10287 9027
rect 10505 9027 10563 9033
rect 10505 9024 10517 9027
rect 10275 8996 10517 9024
rect 10275 8993 10287 8996
rect 10229 8987 10287 8993
rect 10505 8993 10517 8996
rect 10551 9024 10563 9027
rect 10594 9024 10600 9036
rect 10551 8996 10600 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 10781 9027 10839 9033
rect 10781 9024 10793 9027
rect 10744 8996 10793 9024
rect 10744 8984 10750 8996
rect 10781 8993 10793 8996
rect 10827 8993 10839 9027
rect 10781 8987 10839 8993
rect 11146 8984 11152 9036
rect 11204 8984 11210 9036
rect 11256 9024 11284 9064
rect 12802 9052 12808 9104
rect 12860 9092 12866 9104
rect 17144 9101 17172 9132
rect 17862 9120 17868 9132
rect 17920 9160 17929 9169
rect 17920 9132 17965 9160
rect 17920 9123 17929 9132
rect 17920 9120 17926 9123
rect 19334 9120 19340 9172
rect 19392 9120 19398 9172
rect 20165 9163 20223 9169
rect 20165 9129 20177 9163
rect 20211 9160 20223 9163
rect 21634 9160 21640 9172
rect 20211 9132 21640 9160
rect 20211 9129 20223 9132
rect 20165 9123 20223 9129
rect 21634 9120 21640 9132
rect 21692 9120 21698 9172
rect 21735 9163 21793 9169
rect 21735 9129 21747 9163
rect 21781 9160 21793 9163
rect 22002 9160 22008 9172
rect 21781 9132 22008 9160
rect 21781 9129 21793 9132
rect 21735 9123 21793 9129
rect 22002 9120 22008 9132
rect 22060 9120 22066 9172
rect 22646 9120 22652 9172
rect 22704 9160 22710 9172
rect 23109 9163 23167 9169
rect 23109 9160 23121 9163
rect 22704 9132 23121 9160
rect 22704 9120 22710 9132
rect 23109 9129 23121 9132
rect 23155 9129 23167 9163
rect 23109 9123 23167 9129
rect 23566 9120 23572 9172
rect 23624 9120 23630 9172
rect 23750 9120 23756 9172
rect 23808 9160 23814 9172
rect 23943 9163 24001 9169
rect 23943 9160 23955 9163
rect 23808 9132 23955 9160
rect 23808 9120 23814 9132
rect 23943 9129 23955 9132
rect 23989 9129 24001 9163
rect 23943 9123 24001 9129
rect 24118 9120 24124 9172
rect 24176 9160 24182 9172
rect 24176 9132 25176 9160
rect 24176 9120 24182 9132
rect 17129 9095 17187 9101
rect 12860 9064 13676 9092
rect 12860 9052 12866 9064
rect 13648 9033 13676 9064
rect 17129 9061 17141 9095
rect 17175 9061 17187 9095
rect 17129 9055 17187 9061
rect 11885 9027 11943 9033
rect 11885 9024 11897 9027
rect 11256 8996 11897 9024
rect 11885 8993 11897 8996
rect 11931 8993 11943 9027
rect 11885 8987 11943 8993
rect 13633 9027 13691 9033
rect 13633 8993 13645 9027
rect 13679 8993 13691 9027
rect 13633 8987 13691 8993
rect 14052 9027 14110 9033
rect 14052 8993 14064 9027
rect 14098 9024 14110 9027
rect 14366 9024 14372 9036
rect 14098 8996 14372 9024
rect 14098 8993 14110 8996
rect 14052 8987 14110 8993
rect 14366 8984 14372 8996
rect 14424 8984 14430 9036
rect 14461 9027 14519 9033
rect 14461 8993 14473 9027
rect 14507 9024 14519 9027
rect 14826 9024 14832 9036
rect 14507 8996 14832 9024
rect 14507 8993 14519 8996
rect 14461 8987 14519 8993
rect 14826 8984 14832 8996
rect 14884 8984 14890 9036
rect 14918 8984 14924 9036
rect 14976 8984 14982 9036
rect 16850 8984 16856 9036
rect 16908 9024 16914 9036
rect 17310 9024 17316 9036
rect 16908 8996 17316 9024
rect 16908 8984 16914 8996
rect 17310 8984 17316 8996
rect 17368 8984 17374 9036
rect 17402 8984 17408 9036
rect 17460 8984 17466 9036
rect 19352 9024 19380 9120
rect 19521 9095 19579 9101
rect 19521 9061 19533 9095
rect 19567 9092 19579 9095
rect 19794 9092 19800 9104
rect 19567 9064 19800 9092
rect 19567 9061 19579 9064
rect 19521 9055 19579 9061
rect 19794 9052 19800 9064
rect 19852 9052 19858 9104
rect 20622 9052 20628 9104
rect 20680 9052 20686 9104
rect 20717 9095 20775 9101
rect 20717 9061 20729 9095
rect 20763 9092 20775 9095
rect 21082 9092 21088 9104
rect 20763 9064 21088 9092
rect 20763 9061 20775 9064
rect 20717 9055 20775 9061
rect 21082 9052 21088 9064
rect 21140 9052 21146 9104
rect 19705 9027 19763 9033
rect 19705 9024 19717 9027
rect 18064 8996 18276 9024
rect 19352 8996 19717 9024
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 8168 8928 8213 8956
rect 8168 8916 8174 8928
rect 9030 8916 9036 8968
rect 9088 8956 9094 8968
rect 9088 8928 9674 8956
rect 9088 8916 9094 8928
rect 7650 8888 7656 8900
rect 6840 8860 7236 8888
rect 7576 8860 7656 8888
rect 3878 8820 3884 8832
rect 2746 8792 3884 8820
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 5445 8823 5503 8829
rect 5445 8789 5457 8823
rect 5491 8820 5503 8823
rect 6178 8820 6184 8832
rect 5491 8792 6184 8820
rect 5491 8789 5503 8792
rect 5445 8783 5503 8789
rect 6178 8780 6184 8792
rect 6236 8780 6242 8832
rect 6270 8780 6276 8832
rect 6328 8820 6334 8832
rect 6840 8820 6868 8860
rect 6328 8792 6868 8820
rect 7009 8823 7067 8829
rect 6328 8780 6334 8792
rect 7009 8789 7021 8823
rect 7055 8820 7067 8823
rect 7098 8820 7104 8832
rect 7055 8792 7104 8820
rect 7055 8789 7067 8792
rect 7009 8783 7067 8789
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 7208 8820 7236 8860
rect 7650 8848 7656 8860
rect 7708 8848 7714 8900
rect 9646 8888 9674 8928
rect 9766 8916 9772 8968
rect 9824 8916 9830 8968
rect 11164 8956 11192 8984
rect 11514 8956 11520 8968
rect 11164 8928 11520 8956
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 11612 8961 11670 8967
rect 11612 8927 11624 8961
rect 11658 8956 11670 8961
rect 11698 8956 11704 8968
rect 11658 8928 11704 8956
rect 11658 8927 11670 8928
rect 11612 8921 11670 8927
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 13906 8956 13912 8968
rect 13780 8928 13912 8956
rect 13780 8916 13786 8928
rect 13906 8916 13912 8928
rect 13964 8916 13970 8968
rect 14231 8959 14289 8965
rect 14231 8925 14243 8959
rect 14277 8956 14289 8959
rect 14936 8956 14964 8984
rect 14277 8928 14964 8956
rect 17911 8959 17969 8965
rect 14277 8925 14289 8928
rect 14231 8919 14289 8925
rect 17911 8925 17923 8959
rect 17957 8956 17969 8959
rect 18064 8956 18092 8996
rect 17957 8928 18092 8956
rect 17957 8925 17969 8928
rect 17911 8919 17969 8925
rect 18138 8916 18144 8968
rect 18196 8916 18202 8968
rect 18248 8956 18276 8996
rect 19705 8993 19717 8996
rect 19751 9024 19763 9027
rect 20349 9027 20407 9033
rect 19751 8996 20300 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 20162 8956 20168 8968
rect 18248 8928 20168 8956
rect 20162 8916 20168 8928
rect 20220 8916 20226 8968
rect 20272 8956 20300 8996
rect 20349 8993 20361 9027
rect 20395 9024 20407 9027
rect 20438 9024 20444 9036
rect 20395 8996 20444 9024
rect 20395 8993 20407 8996
rect 20349 8987 20407 8993
rect 20438 8984 20444 8996
rect 20496 9024 20502 9036
rect 20640 9024 20668 9052
rect 20496 8996 20668 9024
rect 20496 8984 20502 8996
rect 20898 8984 20904 9036
rect 20956 9024 20962 9036
rect 22005 9027 22063 9033
rect 22005 9024 22017 9027
rect 20956 8996 22017 9024
rect 20956 8984 20962 8996
rect 22005 8993 22017 8996
rect 22051 8993 22063 9027
rect 23584 9024 23612 9120
rect 25148 9092 25176 9132
rect 25222 9120 25228 9172
rect 25280 9160 25286 9172
rect 25317 9163 25375 9169
rect 25317 9160 25329 9163
rect 25280 9132 25329 9160
rect 25280 9120 25286 9132
rect 25317 9129 25329 9132
rect 25363 9129 25375 9163
rect 25317 9123 25375 9129
rect 25682 9120 25688 9172
rect 25740 9120 25746 9172
rect 25961 9163 26019 9169
rect 25961 9129 25973 9163
rect 26007 9160 26019 9163
rect 28994 9160 29000 9172
rect 26007 9132 26556 9160
rect 26007 9129 26019 9132
rect 25961 9123 26019 9129
rect 25148 9064 26464 9092
rect 24213 9027 24271 9033
rect 24213 9024 24225 9027
rect 23584 8996 24225 9024
rect 22005 8987 22063 8993
rect 24213 8993 24225 8996
rect 24259 8993 24271 9027
rect 24213 8987 24271 8993
rect 24486 8984 24492 9036
rect 24544 9024 24550 9036
rect 25869 9027 25927 9033
rect 25869 9024 25881 9027
rect 24544 8996 25881 9024
rect 24544 8984 24550 8996
rect 25869 8993 25881 8996
rect 25915 9024 25927 9027
rect 25915 8996 26004 9024
rect 25915 8993 25927 8996
rect 25869 8987 25927 8993
rect 25976 8968 26004 8996
rect 26050 8984 26056 9036
rect 26108 9024 26114 9036
rect 26436 9033 26464 9064
rect 26145 9027 26203 9033
rect 26145 9024 26157 9027
rect 26108 8996 26157 9024
rect 26108 8984 26114 8996
rect 26145 8993 26157 8996
rect 26191 8993 26203 9027
rect 26145 8987 26203 8993
rect 26421 9027 26479 9033
rect 26421 8993 26433 9027
rect 26467 8993 26479 9027
rect 26528 9024 26556 9132
rect 28736 9132 29000 9160
rect 28736 9033 28764 9132
rect 28994 9120 29000 9132
rect 29052 9120 29058 9172
rect 29362 9120 29368 9172
rect 29420 9160 29426 9172
rect 30101 9163 30159 9169
rect 30101 9160 30113 9163
rect 29420 9132 30113 9160
rect 29420 9120 29426 9132
rect 30101 9129 30113 9132
rect 30147 9129 30159 9163
rect 30101 9123 30159 9129
rect 27157 9027 27215 9033
rect 27157 9024 27169 9027
rect 26528 8996 27169 9024
rect 26421 8987 26479 8993
rect 27157 8993 27169 8996
rect 27203 8993 27215 9027
rect 27157 8987 27215 8993
rect 28721 9027 28779 9033
rect 28721 8993 28733 9027
rect 28767 8993 28779 9027
rect 28721 8987 28779 8993
rect 28997 9027 29055 9033
rect 28997 8993 29009 9027
rect 29043 9024 29055 9027
rect 30006 9024 30012 9036
rect 29043 8996 30012 9024
rect 29043 8993 29055 8996
rect 28997 8987 29055 8993
rect 30006 8984 30012 8996
rect 30064 8984 30070 9036
rect 20806 8956 20812 8968
rect 20272 8928 20812 8956
rect 20806 8916 20812 8928
rect 20864 8956 20870 8968
rect 20993 8959 21051 8965
rect 20993 8956 21005 8959
rect 20864 8928 21005 8956
rect 20864 8916 20870 8928
rect 20993 8925 21005 8928
rect 21039 8956 21051 8959
rect 21269 8959 21327 8965
rect 21269 8956 21281 8959
rect 21039 8928 21281 8956
rect 21039 8925 21051 8928
rect 20993 8919 21051 8925
rect 21269 8925 21281 8928
rect 21315 8925 21327 8959
rect 21269 8919 21327 8925
rect 21775 8959 21833 8965
rect 21775 8925 21787 8959
rect 21821 8956 21833 8959
rect 22646 8956 22652 8968
rect 21821 8928 22652 8956
rect 21821 8925 21833 8928
rect 21775 8919 21833 8925
rect 11146 8888 11152 8900
rect 9646 8860 11152 8888
rect 11146 8848 11152 8860
rect 11204 8848 11210 8900
rect 19058 8848 19064 8900
rect 19116 8888 19122 8900
rect 19889 8891 19947 8897
rect 19889 8888 19901 8891
rect 19116 8860 19901 8888
rect 19116 8848 19122 8860
rect 19889 8857 19901 8860
rect 19935 8888 19947 8891
rect 21174 8888 21180 8900
rect 19935 8860 21180 8888
rect 19935 8857 19947 8860
rect 19889 8851 19947 8857
rect 21174 8848 21180 8860
rect 21232 8848 21238 8900
rect 8846 8820 8852 8832
rect 7208 8792 8852 8820
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 9490 8780 9496 8832
rect 9548 8820 9554 8832
rect 9858 8820 9864 8832
rect 9548 8792 9864 8820
rect 9548 8780 9554 8792
rect 9858 8780 9864 8792
rect 9916 8780 9922 8832
rect 10321 8823 10379 8829
rect 10321 8789 10333 8823
rect 10367 8820 10379 8823
rect 11606 8820 11612 8832
rect 10367 8792 11612 8820
rect 10367 8789 10379 8792
rect 10321 8783 10379 8789
rect 11606 8780 11612 8792
rect 11664 8780 11670 8832
rect 12710 8780 12716 8832
rect 12768 8820 12774 8832
rect 12989 8823 13047 8829
rect 12989 8820 13001 8823
rect 12768 8792 13001 8820
rect 12768 8780 12774 8792
rect 12989 8789 13001 8792
rect 13035 8789 13047 8823
rect 12989 8783 13047 8789
rect 13449 8823 13507 8829
rect 13449 8789 13461 8823
rect 13495 8820 13507 8823
rect 14274 8820 14280 8832
rect 13495 8792 14280 8820
rect 13495 8789 13507 8792
rect 13449 8783 13507 8789
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 15102 8780 15108 8832
rect 15160 8820 15166 8832
rect 15565 8823 15623 8829
rect 15565 8820 15577 8823
rect 15160 8792 15577 8820
rect 15160 8780 15166 8792
rect 15565 8789 15577 8792
rect 15611 8789 15623 8823
rect 15565 8783 15623 8789
rect 16298 8780 16304 8832
rect 16356 8780 16362 8832
rect 16758 8780 16764 8832
rect 16816 8780 16822 8832
rect 18782 8780 18788 8832
rect 18840 8820 18846 8832
rect 19702 8820 19708 8832
rect 18840 8792 19708 8820
rect 18840 8780 18846 8792
rect 19702 8780 19708 8792
rect 19760 8780 19766 8832
rect 21284 8820 21312 8919
rect 22646 8916 22652 8928
rect 22704 8916 22710 8968
rect 23477 8959 23535 8965
rect 23477 8925 23489 8959
rect 23523 8925 23535 8959
rect 23477 8919 23535 8925
rect 23983 8959 24041 8965
rect 23983 8925 23995 8959
rect 24029 8956 24041 8959
rect 25314 8956 25320 8968
rect 24029 8928 25320 8956
rect 24029 8925 24041 8928
rect 23983 8919 24041 8925
rect 23492 8832 23520 8919
rect 25314 8916 25320 8928
rect 25372 8916 25378 8968
rect 25958 8916 25964 8968
rect 26016 8916 26022 8968
rect 26748 8959 26806 8965
rect 26748 8956 26760 8959
rect 26436 8928 26760 8956
rect 24946 8848 24952 8900
rect 25004 8888 25010 8900
rect 26436 8888 26464 8928
rect 26748 8925 26760 8928
rect 26794 8925 26806 8959
rect 26748 8919 26806 8925
rect 26878 8916 26884 8968
rect 26936 8916 26942 8968
rect 25004 8860 26464 8888
rect 25004 8848 25010 8860
rect 23474 8820 23480 8832
rect 21284 8792 23480 8820
rect 23474 8780 23480 8792
rect 23532 8780 23538 8832
rect 24578 8780 24584 8832
rect 24636 8820 24642 8832
rect 26050 8820 26056 8832
rect 24636 8792 26056 8820
rect 24636 8780 24642 8792
rect 26050 8780 26056 8792
rect 26108 8820 26114 8832
rect 26786 8820 26792 8832
rect 26108 8792 26792 8820
rect 26108 8780 26114 8792
rect 26786 8780 26792 8792
rect 26844 8820 26850 8832
rect 27982 8820 27988 8832
rect 26844 8792 27988 8820
rect 26844 8780 26850 8792
rect 27982 8780 27988 8792
rect 28040 8780 28046 8832
rect 28258 8780 28264 8832
rect 28316 8780 28322 8832
rect 552 8730 30912 8752
rect 552 8678 4193 8730
rect 4245 8678 4257 8730
rect 4309 8678 4321 8730
rect 4373 8678 4385 8730
rect 4437 8678 4449 8730
rect 4501 8678 11783 8730
rect 11835 8678 11847 8730
rect 11899 8678 11911 8730
rect 11963 8678 11975 8730
rect 12027 8678 12039 8730
rect 12091 8678 19373 8730
rect 19425 8678 19437 8730
rect 19489 8678 19501 8730
rect 19553 8678 19565 8730
rect 19617 8678 19629 8730
rect 19681 8678 26963 8730
rect 27015 8678 27027 8730
rect 27079 8678 27091 8730
rect 27143 8678 27155 8730
rect 27207 8678 27219 8730
rect 27271 8678 30912 8730
rect 552 8656 30912 8678
rect 1210 8576 1216 8628
rect 1268 8616 1274 8628
rect 2866 8616 2872 8628
rect 1268 8588 2872 8616
rect 1268 8576 1274 8588
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 3786 8616 3792 8628
rect 3252 8588 3792 8616
rect 2406 8508 2412 8560
rect 2464 8548 2470 8560
rect 3252 8548 3280 8588
rect 3786 8576 3792 8588
rect 3844 8576 3850 8628
rect 3878 8576 3884 8628
rect 3936 8616 3942 8628
rect 5077 8619 5135 8625
rect 5077 8616 5089 8619
rect 3936 8588 5089 8616
rect 3936 8576 3942 8588
rect 5077 8585 5089 8588
rect 5123 8585 5135 8619
rect 5077 8579 5135 8585
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 7377 8619 7435 8625
rect 7377 8616 7389 8619
rect 6972 8588 7389 8616
rect 6972 8576 6978 8588
rect 7377 8585 7389 8588
rect 7423 8585 7435 8619
rect 7377 8579 7435 8585
rect 8386 8576 8392 8628
rect 8444 8576 8450 8628
rect 11422 8616 11428 8628
rect 9324 8588 11428 8616
rect 2464 8520 3280 8548
rect 2464 8508 2470 8520
rect 1443 8483 1501 8489
rect 1443 8449 1455 8483
rect 1489 8480 1501 8483
rect 3252 8480 3280 8520
rect 7742 8508 7748 8560
rect 7800 8548 7806 8560
rect 8665 8551 8723 8557
rect 8665 8548 8677 8551
rect 7800 8520 8677 8548
rect 7800 8508 7806 8520
rect 8665 8517 8677 8520
rect 8711 8517 8723 8551
rect 8665 8511 8723 8517
rect 8754 8508 8760 8560
rect 8812 8548 8818 8560
rect 8941 8551 8999 8557
rect 8941 8548 8953 8551
rect 8812 8520 8953 8548
rect 8812 8508 8818 8520
rect 8941 8517 8953 8520
rect 8987 8517 8999 8551
rect 9324 8548 9352 8588
rect 11422 8576 11428 8588
rect 11480 8576 11486 8628
rect 11698 8576 11704 8628
rect 11756 8576 11762 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 12158 8616 12164 8628
rect 11931 8588 12164 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 13722 8616 13728 8628
rect 12636 8588 13728 8616
rect 8941 8511 8999 8517
rect 9048 8520 9352 8548
rect 3564 8483 3622 8489
rect 3564 8480 3576 8483
rect 1489 8452 2544 8480
rect 3252 8452 3576 8480
rect 1489 8449 1501 8452
rect 1443 8443 1501 8449
rect 2516 8424 2544 8452
rect 3564 8449 3576 8452
rect 3610 8449 3622 8483
rect 4062 8480 4068 8492
rect 3715 8471 4068 8480
rect 3564 8443 3622 8449
rect 3700 8465 4068 8471
rect 3700 8431 3712 8465
rect 3746 8452 4068 8465
rect 3746 8431 3758 8452
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 5368 8452 5856 8480
rect 3700 8425 3758 8431
rect 937 8415 995 8421
rect 937 8381 949 8415
rect 983 8412 995 8415
rect 1026 8412 1032 8424
rect 983 8384 1032 8412
rect 983 8381 995 8384
rect 937 8375 995 8381
rect 1026 8372 1032 8384
rect 1084 8372 1090 8424
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 2130 8412 2136 8424
rect 1719 8384 2136 8412
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 2130 8372 2136 8384
rect 2188 8372 2194 8424
rect 2498 8372 2504 8424
rect 2556 8372 2562 8424
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 5368 8412 5396 8452
rect 4019 8384 5396 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 1403 8279 1461 8285
rect 1403 8245 1415 8279
rect 1449 8276 1461 8279
rect 1578 8276 1584 8288
rect 1449 8248 1584 8276
rect 1449 8245 1461 8248
rect 1403 8239 1461 8245
rect 1578 8236 1584 8248
rect 1636 8236 1642 8288
rect 2774 8236 2780 8288
rect 2832 8236 2838 8288
rect 3252 8276 3280 8375
rect 5442 8372 5448 8424
rect 5500 8412 5506 8424
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 5500 8384 5549 8412
rect 5500 8372 5506 8384
rect 5537 8381 5549 8384
rect 5583 8381 5595 8415
rect 5828 8412 5856 8452
rect 5902 8440 5908 8492
rect 5960 8480 5966 8492
rect 6000 8483 6058 8489
rect 6000 8480 6012 8483
rect 5960 8452 6012 8480
rect 5960 8440 5966 8452
rect 6000 8449 6012 8452
rect 6046 8449 6058 8483
rect 6000 8443 6058 8449
rect 6178 8440 6184 8492
rect 6236 8480 6242 8492
rect 6273 8483 6331 8489
rect 6273 8480 6285 8483
rect 6236 8452 6285 8480
rect 6236 8440 6242 8452
rect 6273 8449 6285 8452
rect 6319 8449 6331 8483
rect 6273 8443 6331 8449
rect 7006 8440 7012 8492
rect 7064 8480 7070 8492
rect 7282 8480 7288 8492
rect 7064 8452 7288 8480
rect 7064 8440 7070 8452
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 9048 8480 9076 8520
rect 7668 8452 9076 8480
rect 7668 8412 7696 8452
rect 9858 8440 9864 8492
rect 9916 8480 9922 8492
rect 10140 8483 10198 8489
rect 10140 8480 10152 8483
rect 9916 8452 10152 8480
rect 9916 8440 9922 8452
rect 10140 8449 10152 8452
rect 10186 8449 10198 8483
rect 10140 8443 10198 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 11238 8480 11244 8492
rect 10459 8452 11244 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11514 8440 11520 8492
rect 11572 8480 11578 8492
rect 12636 8489 12664 8588
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 16298 8576 16304 8628
rect 16356 8616 16362 8628
rect 17957 8619 18015 8625
rect 17957 8616 17969 8619
rect 16356 8588 17969 8616
rect 16356 8576 16362 8588
rect 17957 8585 17969 8588
rect 18003 8585 18015 8619
rect 17957 8579 18015 8585
rect 18138 8576 18144 8628
rect 18196 8576 18202 8628
rect 19242 8576 19248 8628
rect 19300 8616 19306 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 19300 8588 20545 8616
rect 19300 8576 19306 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 20533 8579 20591 8585
rect 21177 8619 21235 8625
rect 21177 8585 21189 8619
rect 21223 8616 21235 8619
rect 21542 8616 21548 8628
rect 21223 8588 21548 8616
rect 21223 8585 21235 8588
rect 21177 8579 21235 8585
rect 12894 8508 12900 8560
rect 12952 8548 12958 8560
rect 13081 8551 13139 8557
rect 13081 8548 13093 8551
rect 12952 8520 13093 8548
rect 12952 8508 12958 8520
rect 13081 8517 13093 8520
rect 13127 8517 13139 8551
rect 13081 8511 13139 8517
rect 13740 8489 13768 8576
rect 12621 8483 12679 8489
rect 12621 8480 12633 8483
rect 11572 8452 12633 8480
rect 11572 8440 11578 8452
rect 12621 8449 12633 8452
rect 12667 8449 12679 8483
rect 13725 8483 13783 8489
rect 12621 8443 12679 8449
rect 12728 8452 13308 8480
rect 5828 8384 7696 8412
rect 7745 8415 7803 8421
rect 5537 8375 5595 8381
rect 7745 8381 7757 8415
rect 7791 8381 7803 8415
rect 7745 8375 7803 8381
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8412 8907 8415
rect 9030 8412 9036 8424
rect 8895 8384 9036 8412
rect 8895 8381 8907 8384
rect 8849 8375 8907 8381
rect 7760 8344 7788 8375
rect 6938 8316 7788 8344
rect 8021 8347 8079 8353
rect 3786 8276 3792 8288
rect 3252 8248 3792 8276
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 3878 8236 3884 8288
rect 3936 8276 3942 8288
rect 5534 8276 5540 8288
rect 3936 8248 5540 8276
rect 3936 8236 3942 8248
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 5994 8236 6000 8288
rect 6052 8285 6058 8288
rect 6052 8239 6061 8285
rect 6052 8236 6058 8239
rect 6178 8236 6184 8288
rect 6236 8276 6242 8288
rect 6546 8276 6552 8288
rect 6236 8248 6552 8276
rect 6236 8236 6242 8248
rect 6546 8236 6552 8248
rect 6604 8276 6610 8288
rect 6938 8276 6966 8316
rect 8021 8313 8033 8347
rect 8067 8313 8079 8347
rect 8021 8307 8079 8313
rect 6604 8248 6966 8276
rect 6604 8236 6610 8248
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 7834 8276 7840 8288
rect 7064 8248 7840 8276
rect 7064 8236 7070 8248
rect 7834 8236 7840 8248
rect 7892 8236 7898 8288
rect 8036 8276 8064 8307
rect 8588 8288 8616 8375
rect 9030 8372 9036 8384
rect 9088 8372 9094 8424
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8381 9183 8415
rect 9490 8412 9496 8424
rect 9125 8375 9183 8381
rect 9232 8384 9496 8412
rect 9140 8344 9168 8375
rect 8864 8316 9168 8344
rect 8864 8288 8892 8316
rect 8386 8276 8392 8288
rect 8036 8248 8392 8276
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 8570 8236 8576 8288
rect 8628 8236 8634 8288
rect 8846 8236 8852 8288
rect 8904 8236 8910 8288
rect 9122 8236 9128 8288
rect 9180 8276 9186 8288
rect 9232 8276 9260 8384
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8381 9643 8415
rect 9674 8388 9680 8440
rect 9732 8388 9738 8440
rect 9585 8375 9643 8381
rect 9677 8381 9689 8388
rect 9723 8381 9735 8388
rect 9677 8375 9735 8381
rect 9306 8304 9312 8356
rect 9364 8344 9370 8356
rect 9590 8344 9618 8375
rect 9766 8372 9772 8424
rect 9824 8412 9830 8424
rect 10004 8415 10062 8421
rect 10004 8412 10016 8415
rect 9824 8384 10016 8412
rect 9824 8372 9830 8384
rect 10004 8381 10016 8384
rect 10050 8381 10062 8415
rect 10004 8375 10062 8381
rect 11330 8372 11336 8424
rect 11388 8412 11394 8424
rect 12069 8415 12127 8421
rect 12069 8412 12081 8415
rect 11388 8384 12081 8412
rect 11388 8372 11394 8384
rect 12069 8381 12081 8384
rect 12115 8412 12127 8415
rect 12728 8412 12756 8452
rect 13280 8421 13308 8452
rect 13725 8449 13737 8483
rect 13771 8449 13783 8483
rect 13725 8443 13783 8449
rect 14182 8440 14188 8492
rect 14240 8440 14246 8492
rect 14274 8440 14280 8492
rect 14332 8480 14338 8492
rect 14461 8483 14519 8489
rect 14461 8480 14473 8483
rect 14332 8452 14473 8480
rect 14332 8440 14338 8452
rect 14461 8449 14473 8452
rect 14507 8449 14519 8483
rect 14461 8443 14519 8449
rect 15841 8483 15899 8489
rect 15841 8449 15853 8483
rect 15887 8480 15899 8483
rect 16396 8483 16454 8489
rect 16396 8480 16408 8483
rect 15887 8452 16408 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 16396 8449 16408 8452
rect 16442 8449 16454 8483
rect 16396 8443 16454 8449
rect 19199 8483 19257 8489
rect 19199 8449 19211 8483
rect 19245 8480 19257 8483
rect 21192 8480 21220 8579
rect 21542 8576 21548 8588
rect 21600 8576 21606 8628
rect 25406 8616 25412 8628
rect 23400 8588 25412 8616
rect 21545 8483 21603 8489
rect 19245 8452 21220 8480
rect 21382 8478 21504 8480
rect 21545 8478 21557 8483
rect 21382 8452 21557 8478
rect 19245 8449 19257 8452
rect 19199 8443 19257 8449
rect 12115 8384 12756 8412
rect 12989 8415 13047 8421
rect 12115 8381 12127 8384
rect 12069 8375 12127 8381
rect 12989 8381 13001 8415
rect 13035 8381 13047 8415
rect 12989 8375 13047 8381
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8412 13323 8415
rect 13814 8412 13820 8424
rect 13311 8384 13820 8412
rect 13311 8381 13323 8384
rect 13265 8375 13323 8381
rect 12158 8344 12164 8356
rect 9364 8316 9536 8344
rect 9590 8316 9628 8344
rect 9364 8304 9370 8316
rect 9180 8248 9260 8276
rect 9180 8236 9186 8248
rect 9398 8236 9404 8288
rect 9456 8236 9462 8288
rect 9508 8276 9536 8316
rect 9600 8276 9628 8316
rect 11072 8316 12164 8344
rect 9508 8248 9628 8276
rect 9950 8236 9956 8288
rect 10008 8276 10014 8288
rect 10686 8276 10692 8288
rect 10008 8248 10692 8276
rect 10008 8236 10014 8248
rect 10686 8236 10692 8248
rect 10744 8276 10750 8288
rect 11072 8276 11100 8316
rect 12158 8304 12164 8316
rect 12216 8304 12222 8356
rect 12250 8304 12256 8356
rect 12308 8344 12314 8356
rect 12345 8347 12403 8353
rect 12345 8344 12357 8347
rect 12308 8316 12357 8344
rect 12308 8304 12314 8316
rect 12345 8313 12357 8316
rect 12391 8313 12403 8347
rect 13004 8344 13032 8375
rect 13814 8372 13820 8384
rect 13872 8372 13878 8424
rect 14052 8415 14110 8421
rect 14052 8381 14064 8415
rect 14098 8412 14110 8415
rect 14366 8412 14372 8424
rect 14098 8384 14372 8412
rect 14098 8381 14110 8384
rect 14052 8375 14110 8381
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 15930 8372 15936 8424
rect 15988 8372 15994 8424
rect 16574 8372 16580 8424
rect 16632 8412 16638 8424
rect 16669 8415 16727 8421
rect 16669 8412 16681 8415
rect 16632 8384 16681 8412
rect 16632 8372 16638 8384
rect 16669 8381 16681 8384
rect 16715 8381 16727 8415
rect 16669 8375 16727 8381
rect 18325 8415 18383 8421
rect 18325 8381 18337 8415
rect 18371 8381 18383 8415
rect 18325 8375 18383 8381
rect 12345 8307 12403 8313
rect 12452 8316 13032 8344
rect 10744 8248 11100 8276
rect 12176 8276 12204 8304
rect 12452 8276 12480 8316
rect 18340 8288 18368 8375
rect 18690 8372 18696 8424
rect 18748 8412 18754 8424
rect 19058 8412 19064 8424
rect 18748 8384 19064 8412
rect 18748 8372 18754 8384
rect 19058 8372 19064 8384
rect 19116 8372 19122 8424
rect 19426 8372 19432 8424
rect 19484 8372 19490 8424
rect 21174 8372 21180 8424
rect 21232 8412 21238 8424
rect 21382 8412 21410 8452
rect 21476 8450 21557 8452
rect 21545 8449 21557 8450
rect 21591 8449 21603 8483
rect 21545 8443 21603 8449
rect 22051 8481 22109 8487
rect 22051 8447 22063 8481
rect 22097 8462 22109 8481
rect 23400 8480 23428 8588
rect 25406 8576 25412 8588
rect 25464 8576 25470 8628
rect 25869 8619 25927 8625
rect 25869 8585 25881 8619
rect 25915 8616 25927 8619
rect 26878 8616 26884 8628
rect 25915 8588 26884 8616
rect 25915 8585 25927 8588
rect 25869 8579 25927 8585
rect 26878 8576 26884 8588
rect 26936 8576 26942 8628
rect 28258 8576 28264 8628
rect 28316 8576 28322 8628
rect 22163 8462 23428 8480
rect 22097 8452 23428 8462
rect 22097 8447 22191 8452
rect 22051 8441 22191 8447
rect 22066 8434 22191 8441
rect 23474 8440 23480 8492
rect 23532 8440 23538 8492
rect 23661 8483 23719 8489
rect 23661 8449 23673 8483
rect 23707 8480 23719 8483
rect 24308 8483 24366 8489
rect 24308 8480 24320 8483
rect 23707 8452 24320 8480
rect 23707 8449 23719 8452
rect 23661 8443 23719 8449
rect 24308 8449 24320 8452
rect 24354 8449 24366 8483
rect 24308 8443 24366 8449
rect 26234 8440 26240 8492
rect 26292 8480 26298 8492
rect 26329 8483 26387 8489
rect 26329 8480 26341 8483
rect 26292 8452 26341 8480
rect 26292 8440 26298 8452
rect 26329 8449 26341 8452
rect 26375 8449 26387 8483
rect 26329 8443 26387 8449
rect 26510 8440 26516 8492
rect 26568 8480 26574 8492
rect 26656 8483 26714 8489
rect 26656 8480 26668 8483
rect 26568 8452 26668 8480
rect 26568 8440 26574 8452
rect 26656 8449 26668 8452
rect 26702 8449 26714 8483
rect 26656 8443 26714 8449
rect 26835 8483 26893 8489
rect 26835 8449 26847 8483
rect 26881 8480 26893 8483
rect 28276 8480 28304 8576
rect 26881 8452 28304 8480
rect 26881 8449 26893 8452
rect 26835 8443 26893 8449
rect 21232 8384 21410 8412
rect 21453 8415 21511 8421
rect 21232 8372 21238 8384
rect 21453 8381 21465 8415
rect 21499 8412 21511 8415
rect 21818 8412 21824 8424
rect 21499 8384 21824 8412
rect 21499 8381 21511 8384
rect 21453 8375 21511 8381
rect 21818 8372 21824 8384
rect 21876 8372 21882 8424
rect 22278 8372 22284 8424
rect 22336 8372 22342 8424
rect 23492 8412 23520 8440
rect 23842 8412 23848 8424
rect 23492 8384 23848 8412
rect 23842 8372 23848 8384
rect 23900 8372 23906 8424
rect 23934 8372 23940 8424
rect 23992 8412 23998 8424
rect 24581 8415 24639 8421
rect 24581 8412 24593 8415
rect 23992 8384 24593 8412
rect 23992 8372 23998 8384
rect 24581 8381 24593 8384
rect 24627 8381 24639 8415
rect 24581 8375 24639 8381
rect 25958 8372 25964 8424
rect 26016 8412 26022 8424
rect 26970 8412 26976 8424
rect 26016 8384 26976 8412
rect 26016 8372 26022 8384
rect 26970 8372 26976 8384
rect 27028 8372 27034 8424
rect 27065 8415 27123 8421
rect 27065 8381 27077 8415
rect 27111 8412 27123 8415
rect 28074 8412 28080 8424
rect 27111 8384 28080 8412
rect 27111 8381 27123 8384
rect 27065 8375 27123 8381
rect 28074 8372 28080 8384
rect 28132 8372 28138 8424
rect 28721 8415 28779 8421
rect 28721 8381 28733 8415
rect 28767 8381 28779 8415
rect 28721 8375 28779 8381
rect 29089 8415 29147 8421
rect 29089 8381 29101 8415
rect 29135 8412 29147 8415
rect 29454 8412 29460 8424
rect 29135 8384 29460 8412
rect 29135 8381 29147 8384
rect 29089 8375 29147 8381
rect 23750 8304 23756 8356
rect 23808 8304 23814 8356
rect 27982 8304 27988 8356
rect 28040 8344 28046 8356
rect 28736 8344 28764 8375
rect 29454 8372 29460 8384
rect 29512 8372 29518 8424
rect 30193 8415 30251 8421
rect 30193 8381 30205 8415
rect 30239 8412 30251 8415
rect 31386 8412 31392 8424
rect 30239 8384 31392 8412
rect 30239 8381 30251 8384
rect 30193 8375 30251 8381
rect 31386 8372 31392 8384
rect 31444 8372 31450 8424
rect 28040 8316 28764 8344
rect 29641 8347 29699 8353
rect 28040 8304 28046 8316
rect 29641 8313 29653 8347
rect 29687 8344 29699 8347
rect 30006 8344 30012 8356
rect 29687 8316 30012 8344
rect 29687 8313 29699 8316
rect 29641 8307 29699 8313
rect 30006 8304 30012 8316
rect 30064 8304 30070 8356
rect 12176 8248 12480 8276
rect 10744 8236 10750 8248
rect 12802 8236 12808 8288
rect 12860 8236 12866 8288
rect 14918 8236 14924 8288
rect 14976 8276 14982 8288
rect 16390 8276 16396 8288
rect 16448 8285 16454 8288
rect 14976 8248 16396 8276
rect 14976 8236 14982 8248
rect 16390 8236 16396 8248
rect 16448 8239 16457 8285
rect 16448 8236 16454 8239
rect 18322 8236 18328 8288
rect 18380 8236 18386 8288
rect 19150 8236 19156 8288
rect 19208 8285 19214 8288
rect 19208 8276 19217 8285
rect 21269 8279 21327 8285
rect 19208 8248 19253 8276
rect 19208 8239 19217 8248
rect 21269 8245 21281 8279
rect 21315 8276 21327 8279
rect 21358 8276 21364 8288
rect 21315 8248 21364 8276
rect 21315 8245 21327 8248
rect 21269 8239 21327 8245
rect 19208 8236 19214 8239
rect 21358 8236 21364 8248
rect 21416 8236 21422 8288
rect 21450 8236 21456 8288
rect 21508 8276 21514 8288
rect 22011 8279 22069 8285
rect 22011 8276 22023 8279
rect 21508 8248 22023 8276
rect 21508 8236 21514 8248
rect 22011 8245 22023 8248
rect 22057 8276 22069 8279
rect 23566 8276 23572 8288
rect 22057 8248 23572 8276
rect 22057 8245 22069 8248
rect 22011 8239 22069 8245
rect 23566 8236 23572 8248
rect 23624 8236 23630 8288
rect 23768 8276 23796 8304
rect 24210 8276 24216 8288
rect 23768 8248 24216 8276
rect 24210 8236 24216 8248
rect 24268 8276 24274 8288
rect 24311 8279 24369 8285
rect 24311 8276 24323 8279
rect 24268 8248 24323 8276
rect 24268 8236 24274 8248
rect 24311 8245 24323 8248
rect 24357 8245 24369 8279
rect 24311 8239 24369 8245
rect 25222 8236 25228 8288
rect 25280 8276 25286 8288
rect 26602 8276 26608 8288
rect 25280 8248 26608 8276
rect 25280 8236 25286 8248
rect 26602 8236 26608 8248
rect 26660 8276 26666 8288
rect 27062 8276 27068 8288
rect 26660 8248 27068 8276
rect 26660 8236 26666 8248
rect 27062 8236 27068 8248
rect 27120 8236 27126 8288
rect 27798 8236 27804 8288
rect 27856 8276 27862 8288
rect 28169 8279 28227 8285
rect 28169 8276 28181 8279
rect 27856 8248 28181 8276
rect 27856 8236 27862 8248
rect 28169 8245 28181 8248
rect 28215 8245 28227 8279
rect 28169 8239 28227 8245
rect 28534 8236 28540 8288
rect 28592 8236 28598 8288
rect 29270 8236 29276 8288
rect 29328 8276 29334 8288
rect 29365 8279 29423 8285
rect 29365 8276 29377 8279
rect 29328 8248 29377 8276
rect 29328 8236 29334 8248
rect 29365 8245 29377 8248
rect 29411 8245 29423 8279
rect 29365 8239 29423 8245
rect 29730 8236 29736 8288
rect 29788 8236 29794 8288
rect 30098 8236 30104 8288
rect 30156 8276 30162 8288
rect 30285 8279 30343 8285
rect 30285 8276 30297 8279
rect 30156 8248 30297 8276
rect 30156 8236 30162 8248
rect 30285 8245 30297 8248
rect 30331 8245 30343 8279
rect 30285 8239 30343 8245
rect 552 8186 31072 8208
rect 552 8134 7988 8186
rect 8040 8134 8052 8186
rect 8104 8134 8116 8186
rect 8168 8134 8180 8186
rect 8232 8134 8244 8186
rect 8296 8134 15578 8186
rect 15630 8134 15642 8186
rect 15694 8134 15706 8186
rect 15758 8134 15770 8186
rect 15822 8134 15834 8186
rect 15886 8134 23168 8186
rect 23220 8134 23232 8186
rect 23284 8134 23296 8186
rect 23348 8134 23360 8186
rect 23412 8134 23424 8186
rect 23476 8134 30758 8186
rect 30810 8134 30822 8186
rect 30874 8134 30886 8186
rect 30938 8134 30950 8186
rect 31002 8134 31014 8186
rect 31066 8134 31072 8186
rect 552 8112 31072 8134
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 1679 8075 1737 8081
rect 1679 8072 1691 8075
rect 1636 8044 1691 8072
rect 1636 8032 1642 8044
rect 1679 8041 1691 8044
rect 1725 8072 1737 8075
rect 1725 8044 2774 8072
rect 1725 8041 1737 8044
rect 1679 8035 1737 8041
rect 2746 8004 2774 8044
rect 3510 8032 3516 8084
rect 3568 8072 3574 8084
rect 3568 8044 4936 8072
rect 3568 8032 3574 8044
rect 3602 8004 3608 8016
rect 2746 7976 3608 8004
rect 3602 7964 3608 7976
rect 3660 7964 3666 8016
rect 4908 8004 4936 8044
rect 5442 8032 5448 8084
rect 5500 8072 5506 8084
rect 8297 8075 8355 8081
rect 8297 8072 8309 8075
rect 5500 8044 8309 8072
rect 5500 8032 5506 8044
rect 8297 8041 8309 8044
rect 8343 8041 8355 8075
rect 8297 8035 8355 8041
rect 8386 8032 8392 8084
rect 8444 8072 8450 8084
rect 9131 8075 9189 8081
rect 9131 8072 9143 8075
rect 8444 8044 9143 8072
rect 8444 8032 8450 8044
rect 9131 8041 9143 8044
rect 9177 8072 9189 8075
rect 9490 8072 9496 8084
rect 9177 8044 9496 8072
rect 9177 8041 9189 8044
rect 9131 8035 9189 8041
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 10870 8032 10876 8084
rect 10928 8072 10934 8084
rect 11698 8072 11704 8084
rect 10928 8044 11704 8072
rect 10928 8032 10934 8044
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 12075 8075 12133 8081
rect 12075 8041 12087 8075
rect 12121 8072 12133 8075
rect 14283 8075 14341 8081
rect 14283 8072 14295 8075
rect 12121 8044 14295 8072
rect 12121 8041 12133 8044
rect 12075 8035 12133 8041
rect 14283 8041 14295 8044
rect 14329 8072 14341 8075
rect 14918 8072 14924 8084
rect 14329 8044 14924 8072
rect 14329 8041 14341 8044
rect 14283 8035 14341 8041
rect 14918 8032 14924 8044
rect 14976 8032 14982 8084
rect 15286 8032 15292 8084
rect 15344 8032 15350 8084
rect 16390 8032 16396 8084
rect 16448 8072 16454 8084
rect 16583 8075 16641 8081
rect 16583 8072 16595 8075
rect 16448 8044 16595 8072
rect 16448 8032 16454 8044
rect 16583 8041 16595 8044
rect 16629 8041 16641 8075
rect 16583 8035 16641 8041
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 19886 8072 19892 8084
rect 18196 8044 19892 8072
rect 18196 8032 18202 8044
rect 19886 8032 19892 8044
rect 19944 8032 19950 8084
rect 20162 8032 20168 8084
rect 20220 8032 20226 8084
rect 22462 8072 22468 8084
rect 21100 8044 22468 8072
rect 5905 8007 5963 8013
rect 5905 8004 5917 8007
rect 4908 7976 5917 8004
rect 5905 7973 5917 7976
rect 5951 7973 5963 8007
rect 6362 8004 6368 8016
rect 5905 7967 5963 7973
rect 6012 7976 6368 8004
rect 6012 7948 6040 7976
rect 6362 7964 6368 7976
rect 6420 7964 6426 8016
rect 10410 7964 10416 8016
rect 10468 8004 10474 8016
rect 11606 8004 11612 8016
rect 10468 7976 11612 8004
rect 10468 7964 10474 7976
rect 11606 7964 11612 7976
rect 11664 7964 11670 8016
rect 1118 7896 1124 7948
rect 1176 7896 1182 7948
rect 5442 7936 5448 7948
rect 1872 7908 5448 7936
rect 1026 7828 1032 7880
rect 1084 7868 1090 7880
rect 1213 7871 1271 7877
rect 1213 7868 1225 7871
rect 1084 7840 1225 7868
rect 1084 7828 1090 7840
rect 1213 7837 1225 7840
rect 1259 7868 1271 7871
rect 1486 7868 1492 7880
rect 1259 7840 1492 7868
rect 1259 7837 1271 7840
rect 1213 7831 1271 7837
rect 1486 7828 1492 7840
rect 1544 7828 1550 7880
rect 1719 7871 1777 7877
rect 1719 7837 1731 7871
rect 1765 7868 1777 7871
rect 1872 7868 1900 7908
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 5994 7896 6000 7948
rect 6052 7896 6058 7948
rect 6273 7939 6331 7945
rect 6273 7905 6285 7939
rect 6319 7936 6331 7939
rect 6319 7908 6500 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 1765 7840 1900 7868
rect 1765 7837 1777 7840
rect 1719 7831 1777 7837
rect 1946 7828 1952 7880
rect 2004 7828 2010 7880
rect 3510 7828 3516 7880
rect 3568 7828 3574 7880
rect 3694 7828 3700 7880
rect 3752 7868 3758 7880
rect 3878 7877 3884 7880
rect 3840 7871 3884 7877
rect 3840 7868 3852 7871
rect 3752 7840 3852 7868
rect 3752 7828 3758 7840
rect 3840 7837 3852 7840
rect 3840 7831 3884 7837
rect 3878 7828 3884 7831
rect 3936 7828 3942 7880
rect 4019 7871 4077 7877
rect 4019 7837 4031 7871
rect 4065 7868 4077 7871
rect 4154 7868 4160 7880
rect 4065 7840 4160 7868
rect 4065 7837 4077 7840
rect 4019 7831 4077 7837
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 6362 7868 6368 7880
rect 4295 7840 6368 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 6362 7828 6368 7840
rect 6420 7828 6426 7880
rect 6472 7877 6500 7908
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 7156 7908 7205 7936
rect 7156 7896 7162 7908
rect 7193 7905 7205 7908
rect 7239 7905 7251 7939
rect 7193 7899 7251 7905
rect 8665 7939 8723 7945
rect 8665 7905 8677 7939
rect 8711 7936 8723 7939
rect 9030 7936 9036 7948
rect 8711 7908 9036 7936
rect 8711 7905 8723 7908
rect 8665 7899 8723 7905
rect 9030 7896 9036 7908
rect 9088 7936 9094 7948
rect 11057 7939 11115 7945
rect 11057 7936 11069 7939
rect 9088 7908 11069 7936
rect 9088 7896 9094 7908
rect 11057 7905 11069 7908
rect 11103 7905 11115 7939
rect 11057 7899 11115 7905
rect 12345 7939 12403 7945
rect 12345 7905 12357 7939
rect 12391 7936 12403 7939
rect 12802 7936 12808 7948
rect 12391 7908 12808 7936
rect 12391 7905 12403 7908
rect 12345 7899 12403 7905
rect 12802 7896 12808 7908
rect 12860 7896 12866 7948
rect 15304 7936 15332 8032
rect 20990 7964 20996 8016
rect 21048 7964 21054 8016
rect 14476 7908 15332 7936
rect 6953 7889 7011 7895
rect 6953 7886 6965 7889
rect 6932 7880 6965 7886
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7868 6515 7871
rect 6638 7868 6644 7880
rect 6503 7840 6644 7868
rect 6503 7837 6515 7840
rect 6457 7831 6515 7837
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 6822 7877 6828 7880
rect 6784 7871 6828 7877
rect 6784 7837 6796 7871
rect 6784 7831 6828 7837
rect 6822 7828 6828 7831
rect 6880 7828 6886 7880
rect 6914 7828 6920 7880
rect 6999 7855 7011 7889
rect 6972 7849 7011 7855
rect 6972 7828 6978 7849
rect 9122 7828 9128 7880
rect 9180 7877 9186 7880
rect 9180 7871 9229 7877
rect 9180 7837 9183 7871
rect 9217 7837 9229 7871
rect 9180 7831 9229 7837
rect 9180 7828 9186 7831
rect 9398 7828 9404 7880
rect 9456 7828 9462 7880
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 11296 7840 11345 7868
rect 11296 7828 11302 7840
rect 11333 7837 11345 7840
rect 11379 7868 11391 7871
rect 11609 7871 11667 7877
rect 11609 7868 11621 7871
rect 11379 7840 11621 7868
rect 11379 7837 11391 7840
rect 11333 7831 11391 7837
rect 11609 7837 11621 7840
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 12115 7871 12173 7877
rect 12115 7837 12127 7871
rect 12161 7868 12173 7871
rect 12710 7868 12716 7880
rect 12161 7840 12716 7868
rect 12161 7837 12173 7840
rect 12115 7831 12173 7837
rect 4908 7772 6132 7800
rect 934 7692 940 7744
rect 992 7692 998 7744
rect 1486 7692 1492 7744
rect 1544 7732 1550 7744
rect 3053 7735 3111 7741
rect 3053 7732 3065 7735
rect 1544 7704 3065 7732
rect 1544 7692 1550 7704
rect 3053 7701 3065 7704
rect 3099 7701 3111 7735
rect 3053 7695 3111 7701
rect 3142 7692 3148 7744
rect 3200 7732 3206 7744
rect 4908 7732 4936 7772
rect 3200 7704 4936 7732
rect 3200 7692 3206 7704
rect 5534 7692 5540 7744
rect 5592 7692 5598 7744
rect 6104 7732 6132 7772
rect 10505 7735 10563 7741
rect 10505 7732 10517 7735
rect 6104 7704 10517 7732
rect 10505 7701 10517 7704
rect 10551 7701 10563 7735
rect 11627 7732 11655 7831
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 13814 7828 13820 7880
rect 13872 7828 13878 7880
rect 14323 7871 14381 7877
rect 14323 7837 14335 7871
rect 14369 7868 14381 7871
rect 14476 7868 14504 7908
rect 15930 7896 15936 7948
rect 15988 7936 15994 7948
rect 16117 7939 16175 7945
rect 16117 7936 16129 7939
rect 15988 7908 16129 7936
rect 15988 7896 15994 7908
rect 16117 7905 16129 7908
rect 16163 7905 16175 7939
rect 16117 7899 16175 7905
rect 18652 7939 18710 7945
rect 18652 7905 18664 7939
rect 18698 7936 18710 7939
rect 20717 7939 20775 7945
rect 18698 7908 19196 7936
rect 18698 7905 18710 7908
rect 18652 7899 18710 7905
rect 14369 7840 14504 7868
rect 14369 7837 14381 7840
rect 14323 7831 14381 7837
rect 14550 7828 14556 7880
rect 14608 7828 14614 7880
rect 14734 7828 14740 7880
rect 14792 7868 14798 7880
rect 15948 7868 15976 7896
rect 16613 7889 16671 7895
rect 16613 7886 16625 7889
rect 14792 7840 15976 7868
rect 14792 7828 14798 7840
rect 16390 7828 16396 7880
rect 16448 7868 16454 7880
rect 16611 7868 16625 7886
rect 16448 7855 16625 7868
rect 16659 7855 16671 7889
rect 19168 7880 19196 7908
rect 20717 7905 20729 7939
rect 20763 7936 20775 7939
rect 21008 7936 21036 7964
rect 21100 7945 21128 8044
rect 22462 8032 22468 8044
rect 22520 8032 22526 8084
rect 22646 8032 22652 8084
rect 22704 8072 22710 8084
rect 23109 8075 23167 8081
rect 23109 8072 23121 8075
rect 22704 8044 23121 8072
rect 22704 8032 22710 8044
rect 23109 8041 23121 8044
rect 23155 8041 23167 8075
rect 23109 8035 23167 8041
rect 23566 8032 23572 8084
rect 23624 8072 23630 8084
rect 23943 8075 24001 8081
rect 23943 8072 23955 8075
rect 23624 8044 23955 8072
rect 23624 8032 23630 8044
rect 23943 8041 23955 8044
rect 23989 8041 24001 8075
rect 23943 8035 24001 8041
rect 25314 8032 25320 8084
rect 25372 8032 25378 8084
rect 26694 8032 26700 8084
rect 26752 8072 26758 8084
rect 28074 8072 28080 8084
rect 26752 8044 28080 8072
rect 26752 8032 26758 8044
rect 28074 8032 28080 8044
rect 28132 8072 28138 8084
rect 28175 8075 28233 8081
rect 28175 8072 28187 8075
rect 28132 8044 28187 8072
rect 28132 8032 28138 8044
rect 28175 8041 28187 8044
rect 28221 8041 28233 8075
rect 28175 8035 28233 8041
rect 29546 8032 29552 8084
rect 29604 8032 29610 8084
rect 25884 7976 27568 8004
rect 25884 7945 25912 7976
rect 27540 7948 27568 7976
rect 20763 7908 21036 7936
rect 21085 7939 21143 7945
rect 20763 7905 20775 7908
rect 20717 7899 20775 7905
rect 21085 7905 21097 7939
rect 21131 7905 21143 7939
rect 22005 7939 22063 7945
rect 22005 7936 22017 7939
rect 21085 7899 21143 7905
rect 21192 7908 22017 7936
rect 16448 7849 16671 7855
rect 16448 7840 16639 7849
rect 16448 7828 16454 7840
rect 16850 7828 16856 7880
rect 16908 7828 16914 7880
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 18831 7871 18889 7877
rect 18831 7837 18843 7871
rect 18877 7868 18889 7871
rect 18966 7868 18972 7880
rect 18877 7840 18972 7868
rect 18877 7837 18889 7840
rect 18831 7831 18889 7837
rect 13832 7800 13860 7828
rect 13004 7772 13860 7800
rect 12250 7732 12256 7744
rect 11627 7704 12256 7732
rect 10505 7695 10563 7701
rect 12250 7692 12256 7704
rect 12308 7732 12314 7744
rect 13004 7732 13032 7772
rect 15654 7760 15660 7812
rect 15712 7760 15718 7812
rect 12308 7704 13032 7732
rect 12308 7692 12314 7704
rect 13446 7692 13452 7744
rect 13504 7692 13510 7744
rect 14366 7692 14372 7744
rect 14424 7732 14430 7744
rect 15010 7732 15016 7744
rect 14424 7704 15016 7732
rect 14424 7692 14430 7704
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 17954 7692 17960 7744
rect 18012 7692 18018 7744
rect 18340 7732 18368 7831
rect 18966 7828 18972 7840
rect 19024 7828 19030 7880
rect 19058 7828 19064 7880
rect 19116 7828 19122 7880
rect 19150 7828 19156 7880
rect 19208 7828 19214 7880
rect 20533 7803 20591 7809
rect 20533 7769 20545 7803
rect 20579 7800 20591 7803
rect 21192 7800 21220 7908
rect 22005 7905 22017 7908
rect 22051 7905 22063 7939
rect 24213 7939 24271 7945
rect 24213 7936 24225 7939
rect 22005 7899 22063 7905
rect 22848 7908 24225 7936
rect 22848 7880 22876 7908
rect 24213 7905 24225 7908
rect 24259 7905 24271 7939
rect 24213 7899 24271 7905
rect 25869 7939 25927 7945
rect 25869 7905 25881 7939
rect 25915 7905 25927 7939
rect 25869 7899 25927 7905
rect 26145 7939 26203 7945
rect 26145 7905 26157 7939
rect 26191 7936 26203 7939
rect 26326 7936 26332 7948
rect 26191 7908 26332 7936
rect 26191 7905 26203 7908
rect 26145 7899 26203 7905
rect 26326 7896 26332 7908
rect 26384 7896 26390 7948
rect 26418 7896 26424 7948
rect 26476 7896 26482 7948
rect 26697 7939 26755 7945
rect 26697 7905 26709 7939
rect 26743 7936 26755 7939
rect 26786 7936 26792 7948
rect 26743 7908 26792 7936
rect 26743 7905 26755 7908
rect 26697 7899 26755 7905
rect 26786 7896 26792 7908
rect 26844 7896 26850 7948
rect 26878 7896 26884 7948
rect 26936 7936 26942 7948
rect 26973 7939 27031 7945
rect 26973 7936 26985 7939
rect 26936 7908 26985 7936
rect 26936 7896 26942 7908
rect 26973 7905 26985 7908
rect 27019 7905 27031 7939
rect 26973 7899 27031 7905
rect 27062 7896 27068 7948
rect 27120 7936 27126 7948
rect 27249 7939 27307 7945
rect 27249 7936 27261 7939
rect 27120 7908 27261 7936
rect 27120 7896 27126 7908
rect 27249 7905 27261 7908
rect 27295 7905 27307 7939
rect 27249 7899 27307 7905
rect 27522 7896 27528 7948
rect 27580 7896 27586 7948
rect 27617 7939 27675 7945
rect 27617 7905 27629 7939
rect 27663 7936 27675 7939
rect 27982 7936 27988 7948
rect 27663 7908 27988 7936
rect 27663 7905 27675 7908
rect 27617 7899 27675 7905
rect 27982 7896 27988 7908
rect 28040 7896 28046 7948
rect 28442 7896 28448 7948
rect 28500 7896 28506 7948
rect 29638 7896 29644 7948
rect 29696 7936 29702 7948
rect 30098 7936 30104 7948
rect 29696 7908 30104 7936
rect 29696 7896 29702 7908
rect 30098 7896 30104 7908
rect 30156 7896 30162 7948
rect 21266 7828 21272 7880
rect 21324 7828 21330 7880
rect 21450 7828 21456 7880
rect 21508 7868 21514 7880
rect 21596 7871 21654 7877
rect 21596 7868 21608 7871
rect 21508 7840 21608 7868
rect 21508 7828 21514 7840
rect 21596 7837 21608 7840
rect 21642 7837 21654 7871
rect 21596 7831 21654 7837
rect 21775 7871 21833 7877
rect 21775 7837 21787 7871
rect 21821 7868 21833 7871
rect 22646 7868 22652 7880
rect 21821 7840 22652 7868
rect 21821 7837 21833 7840
rect 21775 7831 21833 7837
rect 22646 7828 22652 7840
rect 22704 7828 22710 7880
rect 22830 7828 22836 7880
rect 22888 7828 22894 7880
rect 23198 7828 23204 7880
rect 23256 7868 23262 7880
rect 23477 7871 23535 7877
rect 23477 7868 23489 7871
rect 23256 7840 23489 7868
rect 23256 7828 23262 7840
rect 23477 7837 23489 7840
rect 23523 7837 23535 7871
rect 23477 7831 23535 7837
rect 23983 7871 24041 7877
rect 23983 7837 23995 7871
rect 24029 7868 24041 7871
rect 26050 7868 26056 7880
rect 24029 7840 26056 7868
rect 24029 7837 24041 7840
rect 23983 7831 24041 7837
rect 26050 7828 26056 7840
rect 26108 7828 26114 7880
rect 26436 7868 26464 7896
rect 27706 7868 27712 7880
rect 26436 7840 27712 7868
rect 27706 7828 27712 7840
rect 27764 7828 27770 7880
rect 28166 7828 28172 7880
rect 28224 7879 28230 7880
rect 28224 7873 28246 7879
rect 28234 7839 28246 7873
rect 28224 7833 28246 7839
rect 28224 7828 28230 7833
rect 20579 7772 21220 7800
rect 26513 7803 26571 7809
rect 20579 7769 20591 7772
rect 20533 7763 20591 7769
rect 26513 7769 26525 7803
rect 26559 7800 26571 7803
rect 26559 7772 27752 7800
rect 26559 7769 26571 7772
rect 26513 7763 26571 7769
rect 18690 7732 18696 7744
rect 18340 7704 18696 7732
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 18874 7692 18880 7744
rect 18932 7732 18938 7744
rect 19426 7732 19432 7744
rect 18932 7704 19432 7732
rect 18932 7692 18938 7704
rect 19426 7692 19432 7704
rect 19484 7692 19490 7744
rect 20901 7735 20959 7741
rect 20901 7701 20913 7735
rect 20947 7732 20959 7735
rect 22830 7732 22836 7744
rect 20947 7704 22836 7732
rect 20947 7701 20959 7704
rect 20901 7695 20959 7701
rect 22830 7692 22836 7704
rect 22888 7692 22894 7744
rect 25682 7692 25688 7744
rect 25740 7692 25746 7744
rect 25958 7692 25964 7744
rect 26016 7692 26022 7744
rect 26786 7692 26792 7744
rect 26844 7692 26850 7744
rect 27724 7732 27752 7772
rect 28258 7732 28264 7744
rect 27724 7704 28264 7732
rect 28258 7692 28264 7704
rect 28316 7692 28322 7744
rect 28810 7692 28816 7744
rect 28868 7732 28874 7744
rect 29917 7735 29975 7741
rect 29917 7732 29929 7735
rect 28868 7704 29929 7732
rect 28868 7692 28874 7704
rect 29917 7701 29929 7704
rect 29963 7701 29975 7735
rect 29917 7695 29975 7701
rect 552 7642 30912 7664
rect 552 7590 4193 7642
rect 4245 7590 4257 7642
rect 4309 7590 4321 7642
rect 4373 7590 4385 7642
rect 4437 7590 4449 7642
rect 4501 7590 11783 7642
rect 11835 7590 11847 7642
rect 11899 7590 11911 7642
rect 11963 7590 11975 7642
rect 12027 7590 12039 7642
rect 12091 7590 19373 7642
rect 19425 7590 19437 7642
rect 19489 7590 19501 7642
rect 19553 7590 19565 7642
rect 19617 7590 19629 7642
rect 19681 7590 26963 7642
rect 27015 7590 27027 7642
rect 27079 7590 27091 7642
rect 27143 7590 27155 7642
rect 27207 7590 27219 7642
rect 27271 7590 30912 7642
rect 552 7568 30912 7590
rect 934 7488 940 7540
rect 992 7528 998 7540
rect 2961 7531 3019 7537
rect 992 7500 2544 7528
rect 992 7488 998 7500
rect 2130 7392 2136 7404
rect 1458 7383 2136 7392
rect 1433 7377 2136 7383
rect 1433 7343 1445 7377
rect 1479 7364 2136 7377
rect 1479 7343 1491 7364
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 2516 7392 2544 7500
rect 2961 7497 2973 7531
rect 3007 7528 3019 7531
rect 3050 7528 3056 7540
rect 3007 7500 3056 7528
rect 3007 7497 3019 7500
rect 2961 7491 3019 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 3510 7528 3516 7540
rect 3344 7500 3516 7528
rect 3344 7401 3372 7500
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 3602 7488 3608 7540
rect 3660 7528 3666 7540
rect 4062 7528 4068 7540
rect 3660 7500 4068 7528
rect 3660 7488 3666 7500
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 5810 7488 5816 7540
rect 5868 7488 5874 7540
rect 6822 7528 6828 7540
rect 6104 7500 6828 7528
rect 5537 7463 5595 7469
rect 5537 7429 5549 7463
rect 5583 7460 5595 7463
rect 5994 7460 6000 7472
rect 5583 7432 6000 7460
rect 5583 7429 5595 7432
rect 5537 7423 5595 7429
rect 5994 7420 6000 7432
rect 6052 7420 6058 7472
rect 3694 7401 3700 7404
rect 3329 7395 3387 7401
rect 2516 7364 2912 7392
rect 1433 7337 1491 7343
rect 937 7327 995 7333
rect 937 7293 949 7327
rect 983 7324 995 7327
rect 1026 7324 1032 7336
rect 983 7296 1032 7324
rect 983 7293 995 7296
rect 937 7287 995 7293
rect 1026 7284 1032 7296
rect 1084 7284 1090 7336
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 2884 7324 2912 7364
rect 3329 7361 3341 7395
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 3656 7395 3700 7401
rect 3656 7361 3668 7395
rect 3656 7355 3700 7361
rect 3694 7352 3700 7355
rect 3752 7352 3758 7404
rect 3835 7395 3893 7401
rect 3835 7361 3847 7395
rect 3881 7392 3893 7395
rect 6104 7392 6132 7500
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7006 7488 7012 7540
rect 7064 7528 7070 7540
rect 9674 7528 9680 7540
rect 7064 7500 9680 7528
rect 7064 7488 7070 7500
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 13446 7528 13452 7540
rect 10980 7500 13452 7528
rect 7558 7420 7564 7472
rect 7616 7460 7622 7472
rect 7929 7463 7987 7469
rect 7929 7460 7941 7463
rect 7616 7432 7941 7460
rect 7616 7420 7622 7432
rect 7929 7429 7941 7432
rect 7975 7429 7987 7463
rect 7929 7423 7987 7429
rect 8757 7463 8815 7469
rect 8757 7429 8769 7463
rect 8803 7429 8815 7463
rect 8757 7423 8815 7429
rect 3881 7364 6132 7392
rect 3881 7361 3893 7364
rect 3835 7355 3893 7361
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6546 7392 6552 7404
rect 6328 7364 6552 7392
rect 6328 7352 6334 7364
rect 6546 7352 6552 7364
rect 6604 7392 6610 7404
rect 6825 7395 6883 7401
rect 6604 7364 6649 7392
rect 6604 7352 6610 7364
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 7742 7392 7748 7404
rect 6871 7364 7748 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 8772 7392 8800 7423
rect 9398 7401 9404 7404
rect 9360 7395 9404 7401
rect 8772 7364 9260 7392
rect 4065 7327 4123 7333
rect 4065 7324 4077 7327
rect 1719 7296 2774 7324
rect 2884 7296 4077 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 2746 7256 2774 7296
rect 4065 7293 4077 7296
rect 4111 7293 4123 7327
rect 4065 7287 4123 7293
rect 5718 7284 5724 7336
rect 5776 7284 5782 7336
rect 5902 7284 5908 7336
rect 5960 7324 5966 7336
rect 5997 7327 6055 7333
rect 5997 7324 6009 7327
rect 5960 7296 6009 7324
rect 5960 7284 5966 7296
rect 5997 7293 6009 7296
rect 6043 7293 6055 7327
rect 5997 7287 6055 7293
rect 6089 7327 6147 7333
rect 6089 7293 6101 7327
rect 6135 7324 6147 7327
rect 6638 7324 6644 7336
rect 6135 7296 6644 7324
rect 6135 7293 6147 7296
rect 6089 7287 6147 7293
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7324 8723 7327
rect 8941 7327 8999 7333
rect 8711 7296 8892 7324
rect 8711 7293 8723 7296
rect 8665 7287 8723 7293
rect 3234 7256 3240 7268
rect 2746 7228 3240 7256
rect 3234 7216 3240 7228
rect 3292 7216 3298 7268
rect 8570 7256 8576 7268
rect 7576 7228 8576 7256
rect 7576 7200 7604 7228
rect 8570 7216 8576 7228
rect 8628 7216 8634 7268
rect 1403 7191 1461 7197
rect 1403 7157 1415 7191
rect 1449 7188 1461 7191
rect 1578 7188 1584 7200
rect 1449 7160 1584 7188
rect 1449 7157 1461 7160
rect 1403 7151 1461 7157
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 2958 7148 2964 7200
rect 3016 7188 3022 7200
rect 5169 7191 5227 7197
rect 5169 7188 5181 7191
rect 3016 7160 5181 7188
rect 3016 7148 3022 7160
rect 5169 7157 5181 7160
rect 5215 7157 5227 7191
rect 5169 7151 5227 7157
rect 6546 7148 6552 7200
rect 6604 7197 6610 7200
rect 6604 7188 6613 7197
rect 6914 7188 6920 7200
rect 6604 7160 6920 7188
rect 6604 7151 6613 7160
rect 6604 7148 6610 7151
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7558 7148 7564 7200
rect 7616 7148 7622 7200
rect 8478 7148 8484 7200
rect 8536 7148 8542 7200
rect 8864 7188 8892 7296
rect 8941 7293 8953 7327
rect 8987 7293 8999 7327
rect 8941 7287 8999 7293
rect 8956 7256 8984 7287
rect 9030 7284 9036 7336
rect 9088 7284 9094 7336
rect 9232 7324 9260 7364
rect 9360 7361 9372 7395
rect 9360 7355 9404 7361
rect 9398 7352 9404 7355
rect 9456 7352 9462 7404
rect 9539 7395 9597 7401
rect 9539 7361 9551 7395
rect 9585 7392 9597 7395
rect 10980 7392 11008 7500
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 13817 7531 13875 7537
rect 13817 7497 13829 7531
rect 13863 7528 13875 7531
rect 13998 7528 14004 7540
rect 13863 7500 14004 7528
rect 13863 7497 13875 7500
rect 13817 7491 13875 7497
rect 13998 7488 14004 7500
rect 14056 7488 14062 7540
rect 14550 7488 14556 7540
rect 14608 7528 14614 7540
rect 16945 7531 17003 7537
rect 16945 7528 16957 7531
rect 14608 7500 16957 7528
rect 14608 7488 14614 7500
rect 16945 7497 16957 7500
rect 16991 7497 17003 7531
rect 18325 7531 18383 7537
rect 16945 7491 17003 7497
rect 17144 7500 18276 7528
rect 12802 7420 12808 7472
rect 12860 7460 12866 7472
rect 13078 7460 13084 7472
rect 12860 7432 13084 7460
rect 12860 7420 12866 7432
rect 13078 7420 13084 7432
rect 13136 7460 13142 7472
rect 16577 7463 16635 7469
rect 13136 7432 13676 7460
rect 13136 7420 13142 7432
rect 9585 7364 11008 7392
rect 9585 7361 9597 7364
rect 9539 7355 9597 7361
rect 11238 7352 11244 7404
rect 11296 7352 11302 7404
rect 11747 7395 11805 7401
rect 11747 7361 11759 7395
rect 11793 7392 11805 7395
rect 12342 7392 12348 7404
rect 11793 7364 12348 7392
rect 11793 7361 11805 7364
rect 11747 7355 11805 7361
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 9232 7296 9781 7324
rect 9769 7293 9781 7296
rect 9815 7293 9827 7327
rect 9769 7287 9827 7293
rect 10962 7284 10968 7336
rect 11020 7324 11026 7336
rect 11882 7324 11888 7336
rect 11020 7296 11888 7324
rect 11020 7284 11026 7296
rect 11882 7284 11888 7296
rect 11940 7284 11946 7336
rect 11977 7327 12035 7333
rect 11977 7293 11989 7327
rect 12023 7324 12035 7327
rect 12710 7324 12716 7336
rect 12023 7296 12716 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 13648 7333 13676 7432
rect 16577 7429 16589 7463
rect 16623 7460 16635 7463
rect 16666 7460 16672 7472
rect 16623 7432 16672 7460
rect 16623 7429 16635 7432
rect 16577 7423 16635 7429
rect 16666 7420 16672 7432
rect 16724 7420 16730 7472
rect 13814 7352 13820 7404
rect 13872 7392 13878 7404
rect 14734 7392 14740 7404
rect 13872 7364 14740 7392
rect 13872 7352 13878 7364
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 14918 7392 14924 7404
rect 14844 7364 14924 7392
rect 13633 7327 13691 7333
rect 13633 7293 13645 7327
rect 13679 7293 13691 7327
rect 14093 7327 14151 7333
rect 14093 7324 14105 7327
rect 13633 7287 13691 7293
rect 13832 7296 14105 7324
rect 9122 7256 9128 7268
rect 8956 7228 9128 7256
rect 9122 7216 9128 7228
rect 9180 7216 9186 7268
rect 13832 7200 13860 7296
rect 14093 7293 14105 7296
rect 14139 7293 14151 7327
rect 14093 7287 14151 7293
rect 14185 7327 14243 7333
rect 14185 7293 14197 7327
rect 14231 7293 14243 7327
rect 14185 7287 14243 7293
rect 14200 7256 14228 7287
rect 14458 7284 14464 7336
rect 14516 7324 14522 7336
rect 14844 7324 14872 7364
rect 14918 7352 14924 7364
rect 14976 7392 14982 7404
rect 15064 7395 15122 7401
rect 15064 7392 15076 7395
rect 14976 7364 15076 7392
rect 14976 7352 14982 7364
rect 15064 7361 15076 7364
rect 15110 7361 15122 7395
rect 15064 7355 15122 7361
rect 15243 7395 15301 7401
rect 15243 7361 15255 7395
rect 15289 7392 15301 7395
rect 15378 7392 15384 7404
rect 15289 7364 15384 7392
rect 15289 7361 15301 7364
rect 15243 7355 15301 7361
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 15470 7352 15476 7404
rect 15528 7352 15534 7404
rect 17144 7333 17172 7500
rect 18248 7472 18276 7500
rect 18325 7497 18337 7531
rect 18371 7528 18383 7531
rect 19058 7528 19064 7540
rect 18371 7500 19064 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 19058 7488 19064 7500
rect 19116 7488 19122 7540
rect 20640 7500 22692 7528
rect 17773 7463 17831 7469
rect 17773 7429 17785 7463
rect 17819 7429 17831 7463
rect 17773 7423 17831 7429
rect 17788 7392 17816 7423
rect 18046 7420 18052 7472
rect 18104 7420 18110 7472
rect 18230 7420 18236 7472
rect 18288 7420 18294 7472
rect 18874 7392 18880 7404
rect 17788 7364 18880 7392
rect 18874 7352 18880 7364
rect 18932 7352 18938 7404
rect 19058 7401 19064 7404
rect 19020 7395 19064 7401
rect 19020 7361 19032 7395
rect 19020 7355 19064 7361
rect 19058 7352 19064 7355
rect 19116 7352 19122 7404
rect 19199 7395 19257 7401
rect 19199 7361 19211 7395
rect 19245 7392 19257 7395
rect 20640 7392 20668 7500
rect 20714 7420 20720 7472
rect 20772 7420 20778 7472
rect 22664 7460 22692 7500
rect 22738 7488 22744 7540
rect 22796 7488 22802 7540
rect 24670 7528 24676 7540
rect 22848 7500 24676 7528
rect 22848 7460 22876 7500
rect 24670 7488 24676 7500
rect 24728 7488 24734 7540
rect 25038 7488 25044 7540
rect 25096 7528 25102 7540
rect 25685 7531 25743 7537
rect 25685 7528 25697 7531
rect 25096 7500 25697 7528
rect 25096 7488 25102 7500
rect 25685 7497 25697 7500
rect 25731 7497 25743 7531
rect 25685 7491 25743 7497
rect 26694 7488 26700 7540
rect 26752 7488 26758 7540
rect 28718 7488 28724 7540
rect 28776 7488 28782 7540
rect 22664 7432 22876 7460
rect 19245 7364 20668 7392
rect 20901 7395 20959 7401
rect 19245 7361 19257 7364
rect 19199 7355 19257 7361
rect 20901 7361 20913 7395
rect 20947 7392 20959 7395
rect 21174 7392 21180 7404
rect 20947 7364 21180 7392
rect 20947 7361 20959 7364
rect 20901 7355 20959 7361
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 21407 7395 21465 7401
rect 21407 7361 21419 7395
rect 21453 7392 21465 7395
rect 21453 7364 23980 7392
rect 21453 7361 21465 7364
rect 21407 7355 21465 7361
rect 14516 7296 14872 7324
rect 17129 7327 17187 7333
rect 14516 7284 14522 7296
rect 17129 7293 17141 7327
rect 17175 7293 17187 7327
rect 17129 7287 17187 7293
rect 17402 7284 17408 7336
rect 17460 7284 17466 7336
rect 17681 7327 17739 7333
rect 17681 7293 17693 7327
rect 17727 7293 17739 7327
rect 17681 7287 17739 7293
rect 14826 7256 14832 7268
rect 14200 7228 14832 7256
rect 14826 7216 14832 7228
rect 14884 7216 14890 7268
rect 16482 7216 16488 7268
rect 16540 7256 16546 7268
rect 17696 7256 17724 7287
rect 17862 7284 17868 7336
rect 17920 7324 17926 7336
rect 17957 7327 18015 7333
rect 17957 7324 17969 7327
rect 17920 7296 17969 7324
rect 17920 7284 17926 7296
rect 17957 7293 17969 7296
rect 18003 7293 18015 7327
rect 17957 7287 18015 7293
rect 18046 7284 18052 7336
rect 18104 7284 18110 7336
rect 18138 7284 18144 7336
rect 18196 7324 18202 7336
rect 18233 7327 18291 7333
rect 18233 7324 18245 7327
rect 18196 7296 18245 7324
rect 18196 7284 18202 7296
rect 18233 7293 18245 7296
rect 18279 7293 18291 7327
rect 18233 7287 18291 7293
rect 18322 7284 18328 7336
rect 18380 7324 18386 7336
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 18380 7296 18521 7324
rect 18380 7284 18386 7296
rect 18509 7293 18521 7296
rect 18555 7293 18567 7327
rect 18509 7287 18567 7293
rect 18690 7284 18696 7336
rect 18748 7284 18754 7336
rect 19429 7327 19487 7333
rect 19429 7324 19441 7327
rect 18800 7296 19441 7324
rect 18064 7256 18092 7284
rect 18800 7256 18828 7296
rect 19429 7293 19441 7296
rect 19475 7293 19487 7327
rect 19429 7287 19487 7293
rect 21634 7284 21640 7336
rect 21692 7284 21698 7336
rect 23842 7284 23848 7336
rect 23900 7284 23906 7336
rect 23952 7324 23980 7364
rect 24026 7352 24032 7404
rect 24084 7392 24090 7404
rect 24308 7395 24366 7401
rect 24308 7392 24320 7395
rect 24084 7364 24320 7392
rect 24084 7352 24090 7364
rect 24308 7361 24320 7364
rect 24354 7361 24366 7395
rect 24308 7355 24366 7361
rect 24394 7352 24400 7404
rect 24452 7392 24458 7404
rect 24581 7395 24639 7401
rect 24581 7392 24593 7395
rect 24452 7364 24593 7392
rect 24452 7352 24458 7364
rect 24581 7361 24593 7364
rect 24627 7361 24639 7395
rect 24581 7355 24639 7361
rect 24946 7352 24952 7404
rect 25004 7352 25010 7404
rect 26418 7352 26424 7404
rect 26476 7352 26482 7404
rect 26712 7392 26740 7488
rect 28902 7420 28908 7472
rect 28960 7460 28966 7472
rect 29273 7463 29331 7469
rect 29273 7460 29285 7463
rect 28960 7432 29285 7460
rect 28960 7420 28966 7432
rect 29273 7429 29285 7432
rect 29319 7429 29331 7463
rect 29273 7423 29331 7429
rect 27024 7395 27082 7401
rect 27024 7392 27036 7395
rect 26712 7364 27036 7392
rect 27024 7361 27036 7364
rect 27070 7361 27082 7395
rect 27024 7355 27082 7361
rect 27203 7395 27261 7401
rect 27203 7361 27215 7395
rect 27249 7392 27261 7395
rect 27798 7392 27804 7404
rect 27249 7364 27804 7392
rect 27249 7361 27261 7364
rect 27203 7355 27261 7361
rect 27798 7352 27804 7364
rect 27856 7352 27862 7404
rect 29914 7392 29920 7404
rect 28736 7364 29920 7392
rect 24964 7324 24992 7352
rect 23952 7296 24992 7324
rect 25038 7284 25044 7336
rect 25096 7324 25102 7336
rect 25866 7324 25872 7336
rect 25096 7296 25872 7324
rect 25096 7284 25102 7296
rect 25866 7284 25872 7296
rect 25924 7324 25930 7336
rect 26053 7327 26111 7333
rect 26053 7324 26065 7327
rect 25924 7296 26065 7324
rect 25924 7284 25930 7296
rect 26053 7293 26065 7296
rect 26099 7293 26111 7327
rect 26436 7324 26464 7352
rect 26697 7327 26755 7333
rect 26697 7324 26709 7327
rect 26436 7296 26709 7324
rect 26053 7287 26111 7293
rect 26697 7293 26709 7296
rect 26743 7293 26755 7327
rect 26697 7287 26755 7293
rect 27433 7327 27491 7333
rect 27433 7293 27445 7327
rect 27479 7324 27491 7327
rect 28736 7324 28764 7364
rect 29914 7352 29920 7364
rect 29972 7352 29978 7404
rect 27479 7296 28764 7324
rect 29181 7327 29239 7333
rect 27479 7293 27491 7296
rect 27433 7287 27491 7293
rect 29181 7293 29193 7327
rect 29227 7293 29239 7327
rect 29181 7287 29239 7293
rect 16540 7228 17954 7256
rect 18064 7228 18828 7256
rect 16540 7216 16546 7228
rect 10594 7188 10600 7200
rect 8864 7160 10600 7188
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 11054 7148 11060 7200
rect 11112 7148 11118 7200
rect 11707 7191 11765 7197
rect 11707 7157 11719 7191
rect 11753 7188 11765 7191
rect 12066 7188 12072 7200
rect 11753 7160 12072 7188
rect 11753 7157 11765 7160
rect 11707 7151 11765 7157
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 12618 7148 12624 7200
rect 12676 7188 12682 7200
rect 13081 7191 13139 7197
rect 13081 7188 13093 7191
rect 12676 7160 13093 7188
rect 12676 7148 12682 7160
rect 13081 7157 13093 7160
rect 13127 7157 13139 7191
rect 13081 7151 13139 7157
rect 13814 7148 13820 7200
rect 13872 7148 13878 7200
rect 13909 7191 13967 7197
rect 13909 7157 13921 7191
rect 13955 7188 13967 7191
rect 15378 7188 15384 7200
rect 13955 7160 15384 7188
rect 13955 7157 13967 7160
rect 13909 7151 13967 7157
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 17218 7148 17224 7200
rect 17276 7148 17282 7200
rect 17494 7148 17500 7200
rect 17552 7148 17558 7200
rect 17926 7188 17954 7228
rect 23198 7216 23204 7268
rect 23256 7216 23262 7268
rect 23566 7216 23572 7268
rect 23624 7216 23630 7268
rect 26326 7216 26332 7268
rect 26384 7216 26390 7268
rect 29196 7256 29224 7287
rect 29270 7284 29276 7336
rect 29328 7324 29334 7336
rect 29457 7327 29515 7333
rect 29457 7324 29469 7327
rect 29328 7296 29469 7324
rect 29328 7284 29334 7296
rect 29457 7293 29469 7296
rect 29503 7293 29515 7327
rect 29457 7287 29515 7293
rect 29730 7256 29736 7268
rect 29196 7228 29736 7256
rect 18230 7188 18236 7200
rect 17926 7160 18236 7188
rect 18230 7148 18236 7160
rect 18288 7148 18294 7200
rect 19242 7148 19248 7200
rect 19300 7188 19306 7200
rect 21358 7188 21364 7200
rect 21416 7197 21422 7200
rect 19300 7160 21364 7188
rect 19300 7148 19306 7160
rect 21358 7148 21364 7160
rect 21416 7151 21425 7197
rect 21416 7148 21422 7151
rect 21910 7148 21916 7200
rect 21968 7188 21974 7200
rect 23216 7188 23244 7216
rect 29564 7200 29592 7228
rect 29730 7216 29736 7228
rect 29788 7216 29794 7268
rect 21968 7160 23244 7188
rect 21968 7148 21974 7160
rect 24210 7148 24216 7200
rect 24268 7188 24274 7200
rect 24311 7191 24369 7197
rect 24311 7188 24323 7191
rect 24268 7160 24323 7188
rect 24268 7148 24274 7160
rect 24311 7157 24323 7160
rect 24357 7157 24369 7191
rect 24311 7151 24369 7157
rect 24670 7148 24676 7200
rect 24728 7188 24734 7200
rect 28442 7188 28448 7200
rect 24728 7160 28448 7188
rect 24728 7148 24734 7160
rect 28442 7148 28448 7160
rect 28500 7148 28506 7200
rect 28994 7148 29000 7200
rect 29052 7148 29058 7200
rect 29546 7148 29552 7200
rect 29604 7148 29610 7200
rect 552 7098 31072 7120
rect 552 7046 7988 7098
rect 8040 7046 8052 7098
rect 8104 7046 8116 7098
rect 8168 7046 8180 7098
rect 8232 7046 8244 7098
rect 8296 7046 15578 7098
rect 15630 7046 15642 7098
rect 15694 7046 15706 7098
rect 15758 7046 15770 7098
rect 15822 7046 15834 7098
rect 15886 7046 23168 7098
rect 23220 7046 23232 7098
rect 23284 7046 23296 7098
rect 23348 7046 23360 7098
rect 23412 7046 23424 7098
rect 23476 7046 30758 7098
rect 30810 7046 30822 7098
rect 30874 7046 30886 7098
rect 30938 7046 30950 7098
rect 31002 7046 31014 7098
rect 31066 7046 31072 7098
rect 552 7024 31072 7046
rect 1578 6944 1584 6996
rect 1636 6993 1642 6996
rect 1636 6984 1645 6993
rect 1636 6956 1681 6984
rect 1636 6947 1645 6956
rect 1636 6944 1642 6947
rect 2130 6944 2136 6996
rect 2188 6984 2194 6996
rect 3142 6984 3148 6996
rect 2188 6956 3148 6984
rect 2188 6944 2194 6956
rect 3142 6944 3148 6956
rect 3200 6944 3206 6996
rect 3234 6944 3240 6996
rect 3292 6984 3298 6996
rect 5442 6984 5448 6996
rect 3292 6956 5448 6984
rect 3292 6944 3298 6956
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 6089 6987 6147 6993
rect 6089 6953 6101 6987
rect 6135 6984 6147 6987
rect 6454 6984 6460 6996
rect 6135 6956 6460 6984
rect 6135 6953 6147 6956
rect 6089 6947 6147 6953
rect 6454 6944 6460 6956
rect 6512 6944 6518 6996
rect 6914 6944 6920 6996
rect 6972 6993 6978 6996
rect 6972 6984 6981 6993
rect 9131 6987 9189 6993
rect 9131 6984 9143 6987
rect 6972 6956 9143 6984
rect 6972 6947 6981 6956
rect 9131 6953 9143 6956
rect 9177 6984 9189 6987
rect 9490 6984 9496 6996
rect 9177 6956 9496 6984
rect 9177 6953 9189 6956
rect 9131 6947 9189 6953
rect 6972 6944 6978 6947
rect 9490 6944 9496 6956
rect 9548 6944 9554 6996
rect 10502 6944 10508 6996
rect 10560 6944 10566 6996
rect 10686 6944 10692 6996
rect 10744 6984 10750 6996
rect 11425 6987 11483 6993
rect 11425 6984 11437 6987
rect 10744 6956 11437 6984
rect 10744 6944 10750 6956
rect 11425 6953 11437 6956
rect 11471 6953 11483 6987
rect 11425 6947 11483 6953
rect 11698 6944 11704 6996
rect 11756 6944 11762 6996
rect 11977 6987 12035 6993
rect 11977 6953 11989 6987
rect 12023 6953 12035 6987
rect 11977 6947 12035 6953
rect 3602 6916 3608 6928
rect 3252 6888 3608 6916
rect 1029 6851 1087 6857
rect 1029 6817 1041 6851
rect 1075 6848 1087 6851
rect 2314 6848 2320 6860
rect 1075 6820 2320 6848
rect 1075 6817 1087 6820
rect 1029 6811 1087 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 3252 6857 3280 6888
rect 3602 6876 3608 6888
rect 3660 6876 3666 6928
rect 6178 6876 6184 6928
rect 6236 6876 6242 6928
rect 11606 6876 11612 6928
rect 11664 6916 11670 6928
rect 11992 6916 12020 6947
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 12627 6987 12685 6993
rect 12627 6984 12639 6987
rect 12124 6956 12639 6984
rect 12124 6944 12130 6956
rect 12627 6953 12639 6956
rect 12673 6984 12685 6987
rect 14458 6984 14464 6996
rect 12673 6956 14464 6984
rect 12673 6953 12685 6956
rect 12627 6947 12685 6953
rect 14458 6944 14464 6956
rect 14516 6944 14522 6996
rect 14829 6987 14887 6993
rect 14829 6953 14841 6987
rect 14875 6953 14887 6987
rect 14829 6947 14887 6953
rect 11664 6888 12020 6916
rect 14844 6916 14872 6947
rect 15470 6944 15476 6996
rect 15528 6984 15534 6996
rect 15657 6987 15715 6993
rect 15657 6984 15669 6987
rect 15528 6956 15669 6984
rect 15528 6944 15534 6956
rect 15657 6953 15669 6956
rect 15703 6953 15715 6987
rect 15657 6947 15715 6953
rect 16850 6944 16856 6996
rect 16908 6944 16914 6996
rect 18230 6944 18236 6996
rect 18288 6984 18294 6996
rect 21266 6984 21272 6996
rect 18288 6956 21272 6984
rect 18288 6944 18294 6956
rect 21266 6944 21272 6956
rect 21324 6944 21330 6996
rect 21450 6944 21456 6996
rect 21508 6984 21514 6996
rect 22287 6987 22345 6993
rect 22287 6984 22299 6987
rect 21508 6956 22299 6984
rect 21508 6944 21514 6956
rect 22287 6953 22299 6956
rect 22333 6953 22345 6987
rect 22287 6947 22345 6953
rect 24587 6987 24645 6993
rect 24587 6953 24599 6987
rect 24633 6984 24645 6987
rect 24854 6984 24860 6996
rect 24633 6956 24860 6984
rect 24633 6953 24645 6956
rect 24587 6947 24645 6953
rect 24854 6944 24860 6956
rect 24912 6944 24918 6996
rect 24946 6944 24952 6996
rect 25004 6984 25010 6996
rect 25961 6987 26019 6993
rect 25961 6984 25973 6987
rect 25004 6956 25973 6984
rect 25004 6944 25010 6956
rect 25961 6953 25973 6956
rect 26007 6953 26019 6987
rect 25961 6947 26019 6953
rect 28074 6944 28080 6996
rect 28132 6984 28138 6996
rect 28175 6987 28233 6993
rect 28175 6984 28187 6987
rect 28132 6956 28187 6984
rect 28132 6944 28138 6956
rect 28175 6953 28187 6956
rect 28221 6953 28233 6987
rect 28175 6947 28233 6953
rect 16868 6916 16896 6944
rect 14844 6888 16896 6916
rect 23937 6919 23995 6925
rect 11664 6876 11670 6888
rect 23937 6885 23949 6919
rect 23983 6916 23995 6919
rect 24026 6916 24032 6928
rect 23983 6888 24032 6916
rect 23983 6885 23995 6888
rect 23937 6879 23995 6885
rect 24026 6876 24032 6888
rect 24084 6876 24090 6928
rect 3237 6851 3295 6857
rect 3237 6817 3249 6851
rect 3283 6817 3295 6851
rect 3237 6811 3295 6817
rect 3510 6808 3516 6860
rect 3568 6808 3574 6860
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6848 4307 6851
rect 4982 6848 4988 6860
rect 4295 6820 4988 6848
rect 4295 6817 4307 6820
rect 4249 6811 4307 6817
rect 4982 6808 4988 6820
rect 5040 6808 5046 6860
rect 5997 6851 6055 6857
rect 5997 6817 6009 6851
rect 6043 6848 6055 6851
rect 6086 6848 6092 6860
rect 6043 6820 6092 6848
rect 6043 6817 6055 6820
rect 5997 6811 6055 6817
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 6196 6848 6224 6876
rect 6273 6851 6331 6857
rect 6273 6848 6285 6851
rect 6196 6820 6285 6848
rect 6273 6817 6285 6820
rect 6319 6817 6331 6851
rect 7193 6851 7251 6857
rect 6273 6811 6331 6817
rect 6840 6820 7144 6848
rect 1121 6783 1179 6789
rect 1121 6780 1133 6783
rect 1044 6752 1133 6780
rect 1044 6724 1072 6752
rect 1121 6749 1133 6752
rect 1167 6749 1179 6783
rect 1121 6743 1179 6749
rect 1627 6785 1685 6791
rect 1627 6751 1639 6785
rect 1673 6780 1685 6785
rect 1762 6780 1768 6792
rect 1673 6752 1768 6780
rect 1673 6751 1685 6752
rect 1627 6745 1685 6751
rect 1762 6740 1768 6752
rect 1820 6740 1826 6792
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6780 1915 6783
rect 1903 6752 2774 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 1026 6672 1032 6724
rect 1084 6672 1090 6724
rect 845 6647 903 6653
rect 845 6613 857 6647
rect 891 6644 903 6647
rect 2038 6644 2044 6656
rect 891 6616 2044 6644
rect 891 6613 903 6616
rect 845 6607 903 6613
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 2746 6644 2774 6752
rect 3694 6740 3700 6792
rect 3752 6780 3758 6792
rect 3840 6783 3898 6789
rect 3840 6780 3852 6783
rect 3752 6752 3852 6780
rect 3752 6740 3758 6752
rect 3840 6749 3852 6752
rect 3886 6749 3898 6783
rect 3840 6743 3898 6749
rect 4019 6783 4077 6789
rect 4019 6749 4031 6783
rect 4065 6780 4077 6783
rect 4065 6752 6132 6780
rect 4065 6749 4077 6752
rect 4019 6743 4077 6749
rect 5810 6672 5816 6724
rect 5868 6672 5874 6724
rect 4890 6644 4896 6656
rect 2746 6616 4896 6644
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 5350 6604 5356 6656
rect 5408 6604 5414 6656
rect 6104 6644 6132 6752
rect 6454 6740 6460 6792
rect 6512 6780 6518 6792
rect 6638 6780 6644 6792
rect 6512 6752 6644 6780
rect 6512 6740 6518 6752
rect 6638 6740 6644 6752
rect 6696 6780 6702 6792
rect 6840 6780 6868 6820
rect 6696 6752 6868 6780
rect 6696 6740 6702 6752
rect 6914 6740 6920 6792
rect 6972 6740 6978 6792
rect 7116 6780 7144 6820
rect 7193 6817 7205 6851
rect 7239 6848 7251 6851
rect 8754 6848 8760 6860
rect 7239 6820 8760 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 8754 6808 8760 6820
rect 8812 6808 8818 6860
rect 9030 6808 9036 6860
rect 9088 6808 9094 6860
rect 10962 6848 10968 6860
rect 9324 6820 10968 6848
rect 8665 6783 8723 6789
rect 8665 6780 8677 6783
rect 7116 6752 8677 6780
rect 8665 6749 8677 6752
rect 8711 6780 8723 6783
rect 9048 6780 9076 6808
rect 8711 6752 9076 6780
rect 9171 6783 9229 6789
rect 8711 6749 8723 6752
rect 8665 6743 8723 6749
rect 9171 6749 9183 6783
rect 9217 6780 9229 6783
rect 9324 6780 9352 6820
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 11146 6808 11152 6860
rect 11204 6808 11210 6860
rect 11241 6851 11299 6857
rect 11241 6817 11253 6851
rect 11287 6848 11299 6851
rect 11330 6848 11336 6860
rect 11287 6820 11336 6848
rect 11287 6817 11299 6820
rect 11241 6811 11299 6817
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 11517 6851 11575 6857
rect 11517 6848 11529 6851
rect 11491 6817 11529 6848
rect 11563 6848 11575 6851
rect 11563 6820 11658 6848
rect 11563 6817 11575 6820
rect 11491 6811 11575 6817
rect 11491 6798 11519 6811
rect 9217 6752 9352 6780
rect 9401 6783 9459 6789
rect 9217 6749 9229 6752
rect 9171 6743 9229 6749
rect 9401 6749 9413 6783
rect 9447 6780 9459 6783
rect 9447 6752 10364 6780
rect 9447 6749 9459 6752
rect 9401 6743 9459 6749
rect 8478 6672 8484 6724
rect 8536 6672 8542 6724
rect 10336 6712 10364 6752
rect 11432 6770 11519 6798
rect 11630 6780 11658 6820
rect 11698 6808 11704 6860
rect 11756 6848 11762 6860
rect 11793 6851 11851 6857
rect 11793 6848 11805 6851
rect 11756 6820 11805 6848
rect 11756 6808 11762 6820
rect 11793 6817 11805 6820
rect 11839 6817 11851 6851
rect 11793 6811 11851 6817
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 12250 6848 12256 6860
rect 12207 6820 12256 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 12250 6808 12256 6820
rect 12308 6808 12314 6860
rect 12802 6848 12808 6860
rect 12360 6820 12808 6848
rect 12360 6780 12388 6820
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 12894 6808 12900 6860
rect 12952 6808 12958 6860
rect 12986 6808 12992 6860
rect 13044 6808 13050 6860
rect 13630 6808 13636 6860
rect 13688 6808 13694 6860
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 14737 6851 14795 6857
rect 14737 6848 14749 6851
rect 14700 6820 14749 6848
rect 14700 6808 14706 6820
rect 14737 6817 14749 6820
rect 14783 6817 14795 6851
rect 14737 6811 14795 6817
rect 15013 6851 15071 6857
rect 15013 6817 15025 6851
rect 15059 6817 15071 6851
rect 15013 6811 15071 6817
rect 10965 6715 11023 6721
rect 10965 6712 10977 6715
rect 10336 6684 10977 6712
rect 10965 6681 10977 6684
rect 11011 6681 11023 6715
rect 11432 6712 11460 6770
rect 11630 6752 12388 6780
rect 12667 6783 12725 6789
rect 12667 6749 12679 6783
rect 12713 6780 12725 6783
rect 13004 6780 13032 6808
rect 12713 6752 13032 6780
rect 13648 6780 13676 6808
rect 15028 6780 15056 6811
rect 15194 6808 15200 6860
rect 15252 6808 15258 6860
rect 15841 6851 15899 6857
rect 15841 6817 15853 6851
rect 15887 6817 15899 6851
rect 15841 6811 15899 6817
rect 13648 6752 15056 6780
rect 15856 6780 15884 6811
rect 16482 6808 16488 6860
rect 16540 6808 16546 6860
rect 17954 6848 17960 6860
rect 16592 6820 17960 6848
rect 16298 6780 16304 6792
rect 15856 6752 16304 6780
rect 12713 6749 12725 6752
rect 12667 6743 12725 6749
rect 16298 6740 16304 6752
rect 16356 6780 16362 6792
rect 16592 6780 16620 6820
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 19334 6857 19340 6860
rect 19296 6851 19340 6857
rect 19296 6848 19308 6851
rect 18064 6820 19308 6848
rect 16356 6752 16620 6780
rect 16761 6783 16819 6789
rect 16356 6740 16362 6752
rect 16761 6749 16773 6783
rect 16807 6749 16819 6783
rect 16761 6743 16819 6749
rect 10965 6675 11023 6681
rect 11348 6684 11460 6712
rect 7926 6644 7932 6656
rect 6104 6616 7932 6644
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 8294 6604 8300 6656
rect 8352 6604 8358 6656
rect 8496 6644 8524 6672
rect 9306 6644 9312 6656
rect 8496 6616 9312 6644
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 11348 6644 11376 6684
rect 13814 6672 13820 6724
rect 13872 6712 13878 6724
rect 14553 6715 14611 6721
rect 13872 6684 14136 6712
rect 13872 6672 13878 6684
rect 9456 6616 11376 6644
rect 9456 6604 9462 6616
rect 11882 6604 11888 6656
rect 11940 6644 11946 6656
rect 14001 6647 14059 6653
rect 14001 6644 14013 6647
rect 11940 6616 14013 6644
rect 11940 6604 11946 6616
rect 14001 6613 14013 6616
rect 14047 6613 14059 6647
rect 14108 6644 14136 6684
rect 14553 6681 14565 6715
rect 14599 6712 14611 6715
rect 16666 6712 16672 6724
rect 14599 6684 16672 6712
rect 14599 6681 14611 6684
rect 14553 6675 14611 6681
rect 16666 6672 16672 6684
rect 16724 6672 16730 6724
rect 15470 6644 15476 6656
rect 14108 6616 15476 6644
rect 14001 6607 14059 6613
rect 15470 6604 15476 6616
rect 15528 6604 15534 6656
rect 16301 6647 16359 6653
rect 16301 6613 16313 6647
rect 16347 6644 16359 6647
rect 16390 6644 16396 6656
rect 16347 6616 16396 6644
rect 16347 6613 16359 6616
rect 16301 6607 16359 6613
rect 16390 6604 16396 6616
rect 16448 6604 16454 6656
rect 16574 6604 16580 6656
rect 16632 6644 16638 6656
rect 16776 6644 16804 6743
rect 16942 6740 16948 6792
rect 17000 6780 17006 6792
rect 17088 6783 17146 6789
rect 17088 6780 17100 6783
rect 17000 6752 17100 6780
rect 17000 6740 17006 6752
rect 17088 6749 17100 6752
rect 17134 6749 17146 6783
rect 17088 6743 17146 6749
rect 17218 6740 17224 6792
rect 17276 6780 17282 6792
rect 17276 6752 17321 6780
rect 17276 6740 17282 6752
rect 17494 6740 17500 6792
rect 17552 6740 17558 6792
rect 17678 6740 17684 6792
rect 17736 6780 17742 6792
rect 18064 6780 18092 6820
rect 19296 6817 19308 6820
rect 19296 6811 19340 6817
rect 19334 6808 19340 6811
rect 19392 6808 19398 6860
rect 20530 6848 20536 6860
rect 19628 6820 20536 6848
rect 18966 6780 18972 6792
rect 17736 6752 18092 6780
rect 18248 6752 18972 6780
rect 17736 6740 17742 6752
rect 18248 6644 18276 6752
rect 18966 6740 18972 6752
rect 19024 6740 19030 6792
rect 19475 6783 19533 6789
rect 19475 6749 19487 6783
rect 19521 6780 19533 6783
rect 19628 6780 19656 6820
rect 20530 6808 20536 6820
rect 20588 6808 20594 6860
rect 21174 6808 21180 6860
rect 21232 6848 21238 6860
rect 21821 6851 21879 6857
rect 21821 6848 21833 6851
rect 21232 6820 21833 6848
rect 21232 6808 21238 6820
rect 21821 6817 21833 6820
rect 21867 6848 21879 6851
rect 21910 6848 21916 6860
rect 21867 6820 21916 6848
rect 21867 6817 21879 6820
rect 21821 6811 21879 6817
rect 21910 6808 21916 6820
rect 21968 6808 21974 6860
rect 24857 6851 24915 6857
rect 22480 6820 23244 6848
rect 19521 6752 19656 6780
rect 19705 6783 19763 6789
rect 19521 6749 19533 6752
rect 19475 6743 19533 6749
rect 19705 6749 19717 6783
rect 19751 6780 19763 6783
rect 20622 6780 20628 6792
rect 19751 6752 20628 6780
rect 19751 6749 19763 6752
rect 19705 6743 19763 6749
rect 20622 6740 20628 6752
rect 20680 6740 20686 6792
rect 21542 6740 21548 6792
rect 21600 6740 21606 6792
rect 22327 6783 22385 6789
rect 22327 6749 22339 6783
rect 22373 6780 22385 6783
rect 22480 6780 22508 6820
rect 23216 6792 23244 6820
rect 23500 6820 24538 6848
rect 22373 6752 22508 6780
rect 22373 6749 22385 6752
rect 22327 6743 22385 6749
rect 22554 6740 22560 6792
rect 22612 6740 22618 6792
rect 23198 6740 23204 6792
rect 23256 6740 23262 6792
rect 16632 6616 18276 6644
rect 16632 6604 16638 6616
rect 18782 6604 18788 6656
rect 18840 6604 18846 6656
rect 19334 6604 19340 6656
rect 19392 6644 19398 6656
rect 20070 6644 20076 6656
rect 19392 6616 20076 6644
rect 19392 6604 19398 6616
rect 20070 6604 20076 6616
rect 20128 6604 20134 6656
rect 20993 6647 21051 6653
rect 20993 6613 21005 6647
rect 21039 6644 21051 6647
rect 23500 6644 23528 6820
rect 23566 6740 23572 6792
rect 23624 6780 23630 6792
rect 24121 6783 24179 6789
rect 24121 6780 24133 6783
rect 23624 6752 24133 6780
rect 23624 6740 23630 6752
rect 24121 6749 24133 6752
rect 24167 6749 24179 6783
rect 24510 6780 24538 6820
rect 24857 6817 24869 6851
rect 24903 6848 24915 6851
rect 25682 6848 25688 6860
rect 24903 6820 25688 6848
rect 24903 6817 24915 6820
rect 24857 6811 24915 6817
rect 25682 6808 25688 6820
rect 25740 6808 25746 6860
rect 26418 6808 26424 6860
rect 26476 6848 26482 6860
rect 27249 6851 27307 6857
rect 27249 6848 27261 6851
rect 26476 6820 27261 6848
rect 26476 6808 26482 6820
rect 27249 6817 27261 6820
rect 27295 6817 27307 6851
rect 27249 6811 27307 6817
rect 27706 6808 27712 6860
rect 27764 6808 27770 6860
rect 28350 6808 28356 6860
rect 28408 6808 28414 6860
rect 28445 6851 28503 6857
rect 28445 6817 28457 6851
rect 28491 6848 28503 6851
rect 29822 6848 29828 6860
rect 28491 6820 29828 6848
rect 28491 6817 28503 6820
rect 28445 6811 28503 6817
rect 29822 6808 29828 6820
rect 29880 6808 29886 6860
rect 24584 6783 24642 6789
rect 24584 6780 24596 6783
rect 24510 6752 24596 6780
rect 24121 6743 24179 6749
rect 24584 6749 24596 6752
rect 24630 6749 24642 6783
rect 24584 6743 24642 6749
rect 21039 6616 23528 6644
rect 24136 6644 24164 6743
rect 26234 6740 26240 6792
rect 26292 6780 26298 6792
rect 26694 6780 26700 6792
rect 26292 6752 26700 6780
rect 26292 6740 26298 6752
rect 26694 6740 26700 6752
rect 26752 6740 26758 6792
rect 28215 6783 28273 6789
rect 28215 6749 28227 6783
rect 28261 6780 28273 6783
rect 28368 6780 28396 6808
rect 28261 6752 28396 6780
rect 28261 6749 28273 6752
rect 28215 6743 28273 6749
rect 25866 6672 25872 6724
rect 25924 6712 25930 6724
rect 25924 6684 27752 6712
rect 25924 6672 25930 6684
rect 24486 6644 24492 6656
rect 24136 6616 24492 6644
rect 21039 6613 21051 6616
rect 20993 6607 21051 6613
rect 24486 6604 24492 6616
rect 24544 6644 24550 6656
rect 26418 6644 26424 6656
rect 24544 6616 26424 6644
rect 24544 6604 24550 6616
rect 26418 6604 26424 6616
rect 26476 6604 26482 6656
rect 26510 6604 26516 6656
rect 26568 6644 26574 6656
rect 26878 6644 26884 6656
rect 26568 6616 26884 6644
rect 26568 6604 26574 6616
rect 26878 6604 26884 6616
rect 26936 6604 26942 6656
rect 27338 6604 27344 6656
rect 27396 6604 27402 6656
rect 27724 6644 27752 6684
rect 29086 6644 29092 6656
rect 27724 6616 29092 6644
rect 29086 6604 29092 6616
rect 29144 6604 29150 6656
rect 29733 6647 29791 6653
rect 29733 6613 29745 6647
rect 29779 6644 29791 6647
rect 31202 6644 31208 6656
rect 29779 6616 31208 6644
rect 29779 6613 29791 6616
rect 29733 6607 29791 6613
rect 31202 6604 31208 6616
rect 31260 6604 31266 6656
rect 552 6554 30912 6576
rect 552 6502 4193 6554
rect 4245 6502 4257 6554
rect 4309 6502 4321 6554
rect 4373 6502 4385 6554
rect 4437 6502 4449 6554
rect 4501 6502 11783 6554
rect 11835 6502 11847 6554
rect 11899 6502 11911 6554
rect 11963 6502 11975 6554
rect 12027 6502 12039 6554
rect 12091 6502 19373 6554
rect 19425 6502 19437 6554
rect 19489 6502 19501 6554
rect 19553 6502 19565 6554
rect 19617 6502 19629 6554
rect 19681 6502 26963 6554
rect 27015 6502 27027 6554
rect 27079 6502 27091 6554
rect 27143 6502 27155 6554
rect 27207 6502 27219 6554
rect 27271 6502 30912 6554
rect 552 6480 30912 6502
rect 5350 6440 5356 6452
rect 3344 6412 5356 6440
rect 1443 6307 1501 6313
rect 1443 6273 1455 6307
rect 1489 6304 1501 6307
rect 3344 6304 3372 6412
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 5442 6400 5448 6452
rect 5500 6440 5506 6452
rect 5813 6443 5871 6449
rect 5813 6440 5825 6443
rect 5500 6412 5825 6440
rect 5500 6400 5506 6412
rect 5813 6409 5825 6412
rect 5859 6409 5871 6443
rect 8294 6440 8300 6452
rect 5813 6403 5871 6409
rect 6104 6412 8300 6440
rect 4890 6332 4896 6384
rect 4948 6372 4954 6384
rect 5537 6375 5595 6381
rect 5537 6372 5549 6375
rect 4948 6344 5549 6372
rect 4948 6332 4954 6344
rect 5537 6341 5549 6344
rect 5583 6341 5595 6375
rect 5537 6335 5595 6341
rect 1489 6276 3372 6304
rect 1489 6273 1501 6276
rect 1443 6267 1501 6273
rect 3510 6264 3516 6316
rect 3568 6264 3574 6316
rect 3694 6313 3700 6316
rect 3656 6307 3700 6313
rect 3656 6273 3668 6307
rect 3656 6267 3700 6273
rect 3694 6264 3700 6267
rect 3752 6264 3758 6316
rect 3835 6307 3893 6313
rect 3835 6273 3847 6307
rect 3881 6304 3893 6307
rect 6104 6304 6132 6412
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 8849 6443 8907 6449
rect 8849 6440 8861 6443
rect 8404 6412 8861 6440
rect 7926 6332 7932 6384
rect 7984 6332 7990 6384
rect 8404 6372 8432 6412
rect 8849 6409 8861 6412
rect 8895 6409 8907 6443
rect 8849 6403 8907 6409
rect 9122 6400 9128 6452
rect 9180 6400 9186 6452
rect 9214 6400 9220 6452
rect 9272 6440 9278 6452
rect 9401 6443 9459 6449
rect 9401 6440 9413 6443
rect 9272 6412 9413 6440
rect 9272 6400 9278 6412
rect 9401 6409 9413 6412
rect 9447 6409 9459 6443
rect 9401 6403 9459 6409
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 11333 6443 11391 6449
rect 11333 6440 11345 6443
rect 9732 6412 11345 6440
rect 9732 6400 9738 6412
rect 11333 6409 11345 6412
rect 11379 6409 11391 6443
rect 11333 6403 11391 6409
rect 11422 6400 11428 6452
rect 11480 6440 11486 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11480 6412 11805 6440
rect 11480 6400 11486 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 13173 6443 13231 6449
rect 13173 6409 13185 6443
rect 13219 6440 13231 6443
rect 14458 6440 14464 6452
rect 13219 6412 14464 6440
rect 13219 6409 13231 6412
rect 13173 6403 13231 6409
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 16482 6400 16488 6452
rect 16540 6400 16546 6452
rect 16666 6400 16672 6452
rect 16724 6400 16730 6452
rect 16850 6400 16856 6452
rect 16908 6440 16914 6452
rect 17678 6440 17684 6452
rect 16908 6412 17684 6440
rect 16908 6400 16914 6412
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 19886 6440 19892 6452
rect 18012 6412 19892 6440
rect 18012 6400 18018 6412
rect 19886 6400 19892 6412
rect 19944 6400 19950 6452
rect 21634 6440 21640 6452
rect 19996 6412 21640 6440
rect 8662 6372 8668 6384
rect 8036 6344 8432 6372
rect 8588 6344 8668 6372
rect 3881 6276 6132 6304
rect 3881 6273 3893 6276
rect 3835 6267 3893 6273
rect 6454 6264 6460 6316
rect 6512 6264 6518 6316
rect 6595 6307 6653 6313
rect 6595 6273 6607 6307
rect 6641 6273 6653 6307
rect 6595 6267 6653 6273
rect 937 6239 995 6245
rect 937 6205 949 6239
rect 983 6236 995 6239
rect 1578 6236 1584 6248
rect 983 6208 1584 6236
rect 983 6205 995 6208
rect 937 6199 995 6205
rect 1044 6100 1072 6208
rect 1578 6196 1584 6208
rect 1636 6196 1642 6248
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 2130 6236 2136 6248
rect 1719 6208 2136 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 2130 6196 2136 6208
rect 2188 6196 2194 6248
rect 3329 6239 3387 6245
rect 3329 6205 3341 6239
rect 3375 6236 3387 6239
rect 3528 6236 3556 6264
rect 3375 6208 3556 6236
rect 4065 6239 4123 6245
rect 3375 6205 3387 6208
rect 3329 6199 3387 6205
rect 4065 6205 4077 6239
rect 4111 6236 4123 6239
rect 4798 6236 4804 6248
rect 4111 6208 4804 6236
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 5721 6239 5779 6245
rect 5721 6236 5733 6239
rect 5644 6208 5733 6236
rect 5644 6180 5672 6208
rect 5721 6205 5733 6208
rect 5767 6205 5779 6239
rect 5721 6199 5779 6205
rect 5902 6196 5908 6248
rect 5960 6236 5966 6248
rect 5997 6239 6055 6245
rect 5997 6236 6009 6239
rect 5960 6208 6009 6236
rect 5960 6196 5966 6208
rect 5997 6205 6009 6208
rect 6043 6205 6055 6239
rect 5997 6199 6055 6205
rect 6089 6239 6147 6245
rect 6089 6205 6101 6239
rect 6135 6236 6147 6239
rect 6472 6236 6500 6264
rect 6135 6208 6500 6236
rect 6610 6236 6638 6267
rect 6730 6264 6736 6316
rect 6788 6304 6794 6316
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6788 6276 6837 6304
rect 6788 6264 6794 6276
rect 6825 6273 6837 6276
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 7466 6264 7472 6316
rect 7524 6304 7530 6316
rect 8036 6304 8064 6344
rect 7524 6276 8064 6304
rect 7524 6264 7530 6276
rect 6914 6236 6920 6248
rect 6610 6208 6920 6236
rect 6135 6205 6147 6208
rect 6089 6199 6147 6205
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 7650 6196 7656 6248
rect 7708 6196 7714 6248
rect 8588 6245 8616 6344
rect 8662 6332 8668 6344
rect 8720 6372 8726 6384
rect 8720 6344 9260 6372
rect 8720 6332 8726 6344
rect 9030 6264 9036 6316
rect 9088 6264 9094 6316
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6205 8723 6239
rect 8665 6199 8723 6205
rect 8941 6239 8999 6245
rect 8941 6205 8953 6239
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 5626 6128 5632 6180
rect 5684 6128 5690 6180
rect 7668 6168 7696 6196
rect 8478 6168 8484 6180
rect 7668 6140 8484 6168
rect 8478 6128 8484 6140
rect 8536 6168 8542 6180
rect 8680 6168 8708 6199
rect 8536 6140 8708 6168
rect 8536 6128 8542 6140
rect 1302 6100 1308 6112
rect 1044 6072 1308 6100
rect 1302 6060 1308 6072
rect 1360 6060 1366 6112
rect 1403 6103 1461 6109
rect 1403 6069 1415 6103
rect 1449 6100 1461 6103
rect 1578 6100 1584 6112
rect 1449 6072 1584 6100
rect 1449 6069 1461 6072
rect 1403 6063 1461 6069
rect 1578 6060 1584 6072
rect 1636 6100 1642 6112
rect 1762 6100 1768 6112
rect 1636 6072 1768 6100
rect 1636 6060 1642 6072
rect 1762 6060 1768 6072
rect 1820 6100 1826 6112
rect 2406 6100 2412 6112
rect 1820 6072 2412 6100
rect 1820 6060 1826 6072
rect 2406 6060 2412 6072
rect 2464 6060 2470 6112
rect 2961 6103 3019 6109
rect 2961 6069 2973 6103
rect 3007 6100 3019 6103
rect 4522 6100 4528 6112
rect 3007 6072 4528 6100
rect 3007 6069 3019 6072
rect 2961 6063 3019 6069
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 5166 6060 5172 6112
rect 5224 6060 5230 6112
rect 6546 6060 6552 6112
rect 6604 6109 6610 6112
rect 6604 6100 6613 6109
rect 6604 6072 6649 6100
rect 6604 6063 6613 6072
rect 6604 6060 6610 6063
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 8389 6103 8447 6109
rect 8389 6100 8401 6103
rect 6788 6072 8401 6100
rect 6788 6060 6794 6072
rect 8389 6069 8401 6072
rect 8435 6069 8447 6103
rect 8956 6100 8984 6199
rect 9048 6168 9076 6264
rect 9232 6245 9260 6344
rect 11054 6332 11060 6384
rect 11112 6372 11118 6384
rect 12897 6375 12955 6381
rect 11112 6344 12848 6372
rect 11112 6332 11118 6344
rect 9306 6264 9312 6316
rect 9364 6304 9370 6316
rect 9999 6307 10057 6313
rect 9364 6276 9628 6304
rect 9364 6264 9370 6276
rect 9217 6239 9275 6245
rect 9217 6205 9229 6239
rect 9263 6205 9275 6239
rect 9217 6199 9275 6205
rect 9493 6239 9551 6245
rect 9493 6205 9505 6239
rect 9539 6205 9551 6239
rect 9600 6236 9628 6276
rect 9999 6273 10011 6307
rect 10045 6304 10057 6307
rect 12618 6304 12624 6316
rect 10045 6276 12624 6304
rect 10045 6273 10057 6276
rect 9999 6267 10057 6273
rect 12618 6264 12624 6276
rect 12676 6264 12682 6316
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 9600 6208 10241 6236
rect 9493 6199 9551 6205
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 11977 6215 12035 6221
rect 9508 6168 9536 6199
rect 11977 6181 11989 6215
rect 12023 6181 12035 6215
rect 12250 6196 12256 6248
rect 12308 6196 12314 6248
rect 12526 6196 12532 6248
rect 12584 6196 12590 6248
rect 12820 6245 12848 6344
rect 12897 6341 12909 6375
rect 12943 6372 12955 6375
rect 14366 6372 14372 6384
rect 12943 6344 14372 6372
rect 12943 6341 12955 6344
rect 12897 6335 12955 6341
rect 14366 6332 14372 6344
rect 14424 6332 14430 6384
rect 13814 6304 13820 6316
rect 13096 6276 13820 6304
rect 13096 6245 13124 6276
rect 13814 6264 13820 6276
rect 13872 6264 13878 6316
rect 14274 6264 14280 6316
rect 14332 6304 14338 6316
rect 14461 6307 14519 6313
rect 14461 6304 14473 6307
rect 14332 6276 14473 6304
rect 14332 6264 14338 6276
rect 14461 6273 14473 6276
rect 14507 6273 14519 6307
rect 14461 6267 14519 6273
rect 15102 6264 15108 6316
rect 15160 6304 15166 6316
rect 15160 6276 15205 6304
rect 15160 6264 15166 6276
rect 15378 6264 15384 6316
rect 15436 6264 15442 6316
rect 16390 6264 16396 6316
rect 16448 6264 16454 6316
rect 16500 6304 16528 6400
rect 18233 6375 18291 6381
rect 18233 6341 18245 6375
rect 18279 6372 18291 6375
rect 19702 6372 19708 6384
rect 18279 6344 19708 6372
rect 18279 6341 18291 6344
rect 18233 6335 18291 6341
rect 19702 6332 19708 6344
rect 19760 6332 19766 6384
rect 16500 6276 17540 6304
rect 12805 6239 12863 6245
rect 12805 6205 12817 6239
rect 12851 6236 12863 6239
rect 13081 6239 13139 6245
rect 13081 6236 13093 6239
rect 12851 6208 13093 6236
rect 12851 6205 12863 6208
rect 12805 6199 12863 6205
rect 13081 6205 13093 6208
rect 13127 6205 13139 6239
rect 13081 6199 13139 6205
rect 13357 6239 13415 6245
rect 13357 6205 13369 6239
rect 13403 6236 13415 6239
rect 13725 6239 13783 6245
rect 13725 6236 13737 6239
rect 13403 6208 13737 6236
rect 13403 6205 13415 6208
rect 13357 6199 13415 6205
rect 13725 6205 13737 6208
rect 13771 6205 13783 6239
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13725 6199 13783 6205
rect 13832 6208 14013 6236
rect 11977 6175 12035 6181
rect 9048 6140 9536 6168
rect 9398 6100 9404 6112
rect 8956 6072 9404 6100
rect 8389 6063 8447 6069
rect 9398 6060 9404 6072
rect 9456 6060 9462 6112
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 9959 6103 10017 6109
rect 9959 6100 9971 6103
rect 9548 6072 9971 6100
rect 9548 6060 9554 6072
rect 9959 6069 9971 6072
rect 10005 6069 10017 6103
rect 9959 6063 10017 6069
rect 10134 6060 10140 6112
rect 10192 6100 10198 6112
rect 11698 6100 11704 6112
rect 10192 6072 11704 6100
rect 10192 6060 10198 6072
rect 11698 6060 11704 6072
rect 11756 6100 11762 6112
rect 11992 6100 12020 6175
rect 12544 6168 12572 6196
rect 13372 6168 13400 6199
rect 12544 6140 13400 6168
rect 13630 6128 13636 6180
rect 13688 6168 13694 6180
rect 13832 6168 13860 6208
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 14645 6239 14703 6245
rect 14645 6205 14657 6239
rect 14691 6236 14703 6239
rect 14734 6236 14740 6248
rect 14691 6208 14740 6236
rect 14691 6205 14703 6208
rect 14645 6199 14703 6205
rect 14734 6196 14740 6208
rect 14792 6196 14798 6248
rect 13688 6140 13860 6168
rect 13688 6128 13694 6140
rect 13906 6128 13912 6180
rect 13964 6168 13970 6180
rect 14185 6171 14243 6177
rect 14185 6168 14197 6171
rect 13964 6140 14197 6168
rect 13964 6128 13970 6140
rect 14185 6137 14197 6140
rect 14231 6137 14243 6171
rect 16408 6168 16436 6264
rect 16853 6239 16911 6245
rect 16853 6205 16865 6239
rect 16899 6236 16911 6239
rect 17310 6236 17316 6248
rect 16899 6208 17316 6236
rect 16899 6205 16911 6208
rect 16853 6199 16911 6205
rect 17310 6196 17316 6208
rect 17368 6196 17374 6248
rect 16942 6168 16948 6180
rect 16408 6140 16948 6168
rect 14185 6131 14243 6137
rect 16942 6128 16948 6140
rect 17000 6128 17006 6180
rect 17126 6128 17132 6180
rect 17184 6128 17190 6180
rect 17512 6168 17540 6276
rect 17604 6302 18092 6304
rect 18156 6302 18920 6304
rect 17604 6276 18920 6302
rect 17604 6245 17632 6276
rect 18064 6274 18184 6276
rect 17589 6239 17647 6245
rect 17589 6205 17601 6239
rect 17635 6205 17647 6239
rect 17589 6199 17647 6205
rect 17865 6239 17923 6245
rect 17865 6205 17877 6239
rect 17911 6236 17923 6239
rect 17954 6236 17960 6248
rect 17911 6208 17960 6236
rect 17911 6205 17923 6208
rect 17865 6199 17923 6205
rect 17954 6196 17960 6208
rect 18012 6236 18018 6248
rect 18892 6245 18920 6276
rect 19334 6264 19340 6316
rect 19392 6264 19398 6316
rect 19996 6304 20024 6412
rect 21634 6400 21640 6412
rect 21692 6400 21698 6452
rect 22281 6443 22339 6449
rect 22281 6409 22293 6443
rect 22327 6440 22339 6443
rect 22554 6440 22560 6452
rect 22327 6412 22560 6440
rect 22327 6409 22339 6412
rect 22281 6403 22339 6409
rect 22554 6400 22560 6412
rect 22612 6400 22618 6452
rect 23198 6400 23204 6452
rect 23256 6440 23262 6452
rect 26329 6443 26387 6449
rect 26329 6440 26341 6443
rect 23256 6412 26341 6440
rect 23256 6400 23262 6412
rect 26329 6409 26341 6412
rect 26375 6409 26387 6443
rect 28537 6443 28595 6449
rect 28537 6440 28549 6443
rect 26329 6403 26387 6409
rect 26436 6412 28549 6440
rect 22830 6332 22836 6384
rect 22888 6372 22894 6384
rect 24302 6372 24308 6384
rect 22888 6344 24308 6372
rect 22888 6332 22894 6344
rect 24302 6332 24308 6344
rect 24360 6332 24366 6384
rect 24394 6332 24400 6384
rect 24452 6332 24458 6384
rect 26050 6332 26056 6384
rect 26108 6372 26114 6384
rect 26436 6372 26464 6412
rect 28537 6409 28549 6412
rect 28583 6409 28595 6443
rect 28537 6403 28595 6409
rect 26108 6344 26464 6372
rect 26108 6332 26114 6344
rect 20254 6304 20260 6316
rect 19812 6276 20024 6304
rect 20088 6276 20260 6304
rect 18141 6239 18199 6245
rect 18141 6236 18153 6239
rect 18012 6208 18153 6236
rect 18012 6196 18018 6208
rect 18141 6205 18153 6208
rect 18187 6205 18199 6239
rect 18141 6199 18199 6205
rect 18417 6239 18475 6245
rect 18417 6205 18429 6239
rect 18463 6205 18475 6239
rect 18417 6199 18475 6205
rect 18877 6239 18935 6245
rect 18877 6205 18889 6239
rect 18923 6236 18935 6239
rect 19058 6236 19064 6248
rect 18923 6208 19064 6236
rect 18923 6205 18935 6208
rect 18877 6199 18935 6205
rect 18432 6168 18460 6199
rect 19058 6196 19064 6208
rect 19116 6196 19122 6248
rect 19153 6239 19211 6245
rect 19153 6205 19165 6239
rect 19199 6236 19211 6239
rect 19242 6236 19248 6248
rect 19199 6208 19248 6236
rect 19199 6205 19211 6208
rect 19153 6199 19211 6205
rect 19242 6196 19248 6208
rect 19300 6196 19306 6248
rect 19518 6168 19524 6180
rect 17512 6140 19524 6168
rect 19518 6128 19524 6140
rect 19576 6128 19582 6180
rect 11756 6072 12020 6100
rect 12069 6103 12127 6109
rect 11756 6060 11762 6072
rect 12069 6069 12081 6103
rect 12115 6100 12127 6103
rect 12158 6100 12164 6112
rect 12115 6072 12164 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 12342 6060 12348 6112
rect 12400 6060 12406 6112
rect 12618 6060 12624 6112
rect 12676 6060 12682 6112
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 13541 6103 13599 6109
rect 13541 6100 13553 6103
rect 12768 6072 13553 6100
rect 12768 6060 12774 6072
rect 13541 6069 13553 6072
rect 13587 6069 13599 6103
rect 13541 6063 13599 6069
rect 13817 6103 13875 6109
rect 13817 6069 13829 6103
rect 13863 6100 13875 6103
rect 14550 6100 14556 6112
rect 13863 6072 14556 6100
rect 13863 6069 13875 6072
rect 13817 6063 13875 6069
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 14918 6060 14924 6112
rect 14976 6100 14982 6112
rect 15111 6103 15169 6109
rect 15111 6100 15123 6103
rect 14976 6072 15123 6100
rect 14976 6060 14982 6072
rect 15111 6069 15123 6072
rect 15157 6069 15169 6103
rect 15111 6063 15169 6069
rect 17402 6060 17408 6112
rect 17460 6060 17466 6112
rect 17678 6060 17684 6112
rect 17736 6060 17742 6112
rect 17954 6060 17960 6112
rect 18012 6060 18018 6112
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 18874 6100 18880 6112
rect 18739 6072 18880 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 18874 6060 18880 6072
rect 18932 6060 18938 6112
rect 19705 6103 19763 6109
rect 19705 6069 19717 6103
rect 19751 6100 19763 6103
rect 19812 6100 19840 6276
rect 19886 6196 19892 6248
rect 19944 6196 19950 6248
rect 19978 6196 19984 6248
rect 20036 6196 20042 6248
rect 19904 6168 19932 6196
rect 20088 6168 20116 6276
rect 20254 6264 20260 6276
rect 20312 6264 20318 6316
rect 20444 6307 20502 6313
rect 20444 6304 20456 6307
rect 20364 6276 20456 6304
rect 20364 6248 20392 6276
rect 20444 6273 20456 6276
rect 20490 6273 20502 6307
rect 20444 6267 20502 6273
rect 22097 6307 22155 6313
rect 22097 6273 22109 6307
rect 22143 6304 22155 6307
rect 24026 6304 24032 6316
rect 22143 6276 24032 6304
rect 22143 6273 22155 6276
rect 22097 6267 22155 6273
rect 24026 6264 24032 6276
rect 24084 6264 24090 6316
rect 20346 6196 20352 6248
rect 20404 6196 20410 6248
rect 20714 6196 20720 6248
rect 20772 6196 20778 6248
rect 22465 6239 22523 6245
rect 22465 6205 22477 6239
rect 22511 6236 22523 6239
rect 22741 6239 22799 6245
rect 22741 6236 22753 6239
rect 22511 6208 22753 6236
rect 22511 6205 22523 6208
rect 22465 6199 22523 6205
rect 22741 6205 22753 6208
rect 22787 6236 22799 6239
rect 22830 6236 22836 6248
rect 22787 6208 22836 6236
rect 22787 6205 22799 6208
rect 22741 6199 22799 6205
rect 22830 6196 22836 6208
rect 22888 6196 22894 6248
rect 23017 6239 23075 6245
rect 23017 6212 23029 6239
rect 22940 6205 23029 6212
rect 23063 6205 23075 6239
rect 22940 6199 23075 6205
rect 24121 6239 24179 6245
rect 24121 6205 24133 6239
rect 24167 6236 24179 6239
rect 24320 6236 24348 6332
rect 24412 6245 24440 6332
rect 24486 6264 24492 6316
rect 24544 6264 24550 6316
rect 25038 6311 25044 6316
rect 24995 6305 25044 6311
rect 24995 6271 25007 6305
rect 25041 6271 25044 6305
rect 24995 6265 25044 6271
rect 25038 6264 25044 6265
rect 25096 6264 25102 6316
rect 25225 6307 25283 6313
rect 25225 6273 25237 6307
rect 25271 6304 25283 6307
rect 25958 6304 25964 6316
rect 25271 6276 25964 6304
rect 25271 6273 25283 6276
rect 25225 6267 25283 6273
rect 25958 6264 25964 6276
rect 26016 6264 26022 6316
rect 26234 6264 26240 6316
rect 26292 6304 26298 6316
rect 27160 6307 27218 6313
rect 27160 6304 27172 6307
rect 26292 6276 27172 6304
rect 26292 6264 26298 6276
rect 27160 6273 27172 6276
rect 27206 6273 27218 6307
rect 27160 6267 27218 6273
rect 27246 6264 27252 6316
rect 27304 6304 27310 6316
rect 27522 6304 27528 6316
rect 27304 6276 27528 6304
rect 27304 6264 27310 6276
rect 27522 6264 27528 6276
rect 27580 6304 27586 6316
rect 27580 6276 29224 6304
rect 27580 6264 27586 6276
rect 24167 6208 24348 6236
rect 24397 6239 24455 6245
rect 24167 6205 24179 6208
rect 24121 6199 24179 6205
rect 24397 6205 24409 6239
rect 24443 6236 24455 6239
rect 25590 6236 25596 6248
rect 24443 6208 25596 6236
rect 24443 6205 24455 6208
rect 24397 6199 24455 6205
rect 22940 6184 23060 6199
rect 25590 6196 25596 6208
rect 25648 6196 25654 6248
rect 26418 6196 26424 6248
rect 26476 6236 26482 6248
rect 26697 6239 26755 6245
rect 26697 6236 26709 6239
rect 26476 6208 26709 6236
rect 26476 6196 26482 6208
rect 26697 6205 26709 6208
rect 26743 6205 26755 6239
rect 26697 6199 26755 6205
rect 26786 6196 26792 6248
rect 26844 6236 26850 6248
rect 29196 6245 29224 6276
rect 27433 6239 27491 6245
rect 27433 6236 27445 6239
rect 26844 6208 27445 6236
rect 26844 6196 26850 6208
rect 27433 6205 27445 6208
rect 27479 6205 27491 6239
rect 27433 6199 27491 6205
rect 29181 6239 29239 6245
rect 29181 6205 29193 6239
rect 29227 6236 29239 6239
rect 30558 6236 30564 6248
rect 29227 6208 30564 6236
rect 29227 6205 29239 6208
rect 29181 6199 29239 6205
rect 30558 6196 30564 6208
rect 30616 6196 30622 6248
rect 22940 6168 22968 6184
rect 19904 6140 20116 6168
rect 22066 6140 22968 6168
rect 23952 6140 24624 6168
rect 19751 6072 19840 6100
rect 20447 6103 20505 6109
rect 19751 6069 19763 6072
rect 19705 6063 19763 6069
rect 20447 6069 20459 6103
rect 20493 6100 20505 6103
rect 20990 6100 20996 6112
rect 20493 6072 20996 6100
rect 20493 6069 20505 6072
rect 20447 6063 20505 6069
rect 20990 6060 20996 6072
rect 21048 6060 21054 6112
rect 21450 6060 21456 6112
rect 21508 6100 21514 6112
rect 22066 6100 22094 6140
rect 22756 6112 22784 6140
rect 21508 6072 22094 6100
rect 21508 6060 21514 6072
rect 22554 6060 22560 6112
rect 22612 6060 22618 6112
rect 22738 6060 22744 6112
rect 22796 6060 22802 6112
rect 22833 6103 22891 6109
rect 22833 6069 22845 6103
rect 22879 6100 22891 6103
rect 23750 6100 23756 6112
rect 22879 6072 23756 6100
rect 22879 6069 22891 6072
rect 22833 6063 22891 6069
rect 23750 6060 23756 6072
rect 23808 6060 23814 6112
rect 23952 6109 23980 6140
rect 23937 6103 23995 6109
rect 23937 6069 23949 6103
rect 23983 6069 23995 6103
rect 23937 6063 23995 6069
rect 24213 6103 24271 6109
rect 24213 6069 24225 6103
rect 24259 6100 24271 6103
rect 24486 6100 24492 6112
rect 24259 6072 24492 6100
rect 24259 6069 24271 6072
rect 24213 6063 24271 6069
rect 24486 6060 24492 6072
rect 24544 6060 24550 6112
rect 24596 6100 24624 6140
rect 24762 6100 24768 6112
rect 24596 6072 24768 6100
rect 24762 6060 24768 6072
rect 24820 6060 24826 6112
rect 24854 6060 24860 6112
rect 24912 6100 24918 6112
rect 24955 6103 25013 6109
rect 24955 6100 24967 6103
rect 24912 6072 24967 6100
rect 24912 6060 24918 6072
rect 24955 6069 24967 6072
rect 25001 6100 25013 6103
rect 26326 6100 26332 6112
rect 25001 6072 26332 6100
rect 25001 6069 25013 6072
rect 24955 6063 25013 6069
rect 26326 6060 26332 6072
rect 26384 6100 26390 6112
rect 27163 6103 27221 6109
rect 27163 6100 27175 6103
rect 26384 6072 27175 6100
rect 26384 6060 26390 6072
rect 27163 6069 27175 6072
rect 27209 6100 27221 6103
rect 27890 6100 27896 6112
rect 27209 6072 27896 6100
rect 27209 6069 27221 6072
rect 27163 6063 27221 6069
rect 27890 6060 27896 6072
rect 27948 6060 27954 6112
rect 28626 6060 28632 6112
rect 28684 6100 28690 6112
rect 28997 6103 29055 6109
rect 28997 6100 29009 6103
rect 28684 6072 29009 6100
rect 28684 6060 28690 6072
rect 28997 6069 29009 6072
rect 29043 6069 29055 6103
rect 28997 6063 29055 6069
rect 552 6010 31072 6032
rect 552 5958 7988 6010
rect 8040 5958 8052 6010
rect 8104 5958 8116 6010
rect 8168 5958 8180 6010
rect 8232 5958 8244 6010
rect 8296 5958 15578 6010
rect 15630 5958 15642 6010
rect 15694 5958 15706 6010
rect 15758 5958 15770 6010
rect 15822 5958 15834 6010
rect 15886 5958 23168 6010
rect 23220 5958 23232 6010
rect 23284 5958 23296 6010
rect 23348 5958 23360 6010
rect 23412 5958 23424 6010
rect 23476 5958 30758 6010
rect 30810 5958 30822 6010
rect 30874 5958 30886 6010
rect 30938 5958 30950 6010
rect 31002 5958 31014 6010
rect 31066 5958 31072 6010
rect 552 5936 31072 5958
rect 845 5899 903 5905
rect 845 5865 857 5899
rect 891 5896 903 5899
rect 1854 5896 1860 5908
rect 891 5868 1860 5896
rect 891 5865 903 5868
rect 845 5859 903 5865
rect 1854 5856 1860 5868
rect 1912 5856 1918 5908
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3568 5868 4077 5896
rect 3568 5856 3574 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 4433 5899 4491 5905
rect 4433 5865 4445 5899
rect 4479 5896 4491 5899
rect 5074 5896 5080 5908
rect 4479 5868 5080 5896
rect 4479 5865 4491 5868
rect 4433 5859 4491 5865
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 5166 5856 5172 5908
rect 5224 5856 5230 5908
rect 5629 5899 5687 5905
rect 5629 5865 5641 5899
rect 5675 5896 5687 5899
rect 6270 5896 6276 5908
rect 5675 5868 6276 5896
rect 5675 5865 5687 5868
rect 5629 5859 5687 5865
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 6362 5856 6368 5908
rect 6420 5856 6426 5908
rect 6454 5856 6460 5908
rect 6512 5896 6518 5908
rect 7374 5896 7380 5908
rect 6512 5868 7380 5896
rect 6512 5856 6518 5868
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 8478 5856 8484 5908
rect 8536 5896 8542 5908
rect 10134 5896 10140 5908
rect 8536 5868 10140 5896
rect 8536 5856 8542 5868
rect 10134 5856 10140 5868
rect 10192 5856 10198 5908
rect 12434 5896 12440 5908
rect 10244 5868 12440 5896
rect 5184 5828 5212 5856
rect 6086 5828 6092 5840
rect 2746 5800 5212 5828
rect 5552 5800 6092 5828
rect 1029 5763 1087 5769
rect 1029 5729 1041 5763
rect 1075 5729 1087 5763
rect 1029 5723 1087 5729
rect 934 5652 940 5704
rect 992 5692 998 5704
rect 1044 5692 1072 5723
rect 1578 5720 1584 5772
rect 1636 5769 1642 5772
rect 1636 5763 1690 5769
rect 1636 5729 1644 5763
rect 1678 5729 1690 5763
rect 2746 5760 2774 5800
rect 5552 5772 5580 5800
rect 6086 5788 6092 5800
rect 6144 5828 6150 5840
rect 6144 5800 7696 5828
rect 6144 5788 6150 5800
rect 3878 5760 3884 5772
rect 1636 5723 1690 5729
rect 1964 5732 2774 5760
rect 3160 5732 3884 5760
rect 1636 5720 1642 5723
rect 1801 5713 1859 5719
rect 992 5664 1072 5692
rect 992 5652 998 5664
rect 1302 5652 1308 5704
rect 1360 5652 1366 5704
rect 1801 5679 1813 5713
rect 1847 5692 1859 5713
rect 1964 5692 1992 5732
rect 1847 5679 1992 5692
rect 1801 5673 1992 5679
rect 1826 5664 1992 5673
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 3160 5692 3188 5732
rect 3878 5720 3884 5732
rect 3936 5720 3942 5772
rect 3970 5720 3976 5772
rect 4028 5720 4034 5772
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4617 5763 4675 5769
rect 4617 5760 4629 5763
rect 4212 5732 4629 5760
rect 4212 5720 4218 5732
rect 4617 5729 4629 5732
rect 4663 5729 4675 5763
rect 4617 5723 4675 5729
rect 4890 5720 4896 5772
rect 4948 5720 4954 5772
rect 5534 5720 5540 5772
rect 5592 5720 5598 5772
rect 5905 5763 5963 5769
rect 5905 5729 5917 5763
rect 5951 5729 5963 5763
rect 5905 5723 5963 5729
rect 6273 5763 6331 5769
rect 6273 5729 6285 5763
rect 6319 5760 6331 5763
rect 6454 5760 6460 5772
rect 6319 5732 6460 5760
rect 6319 5729 6331 5732
rect 6273 5723 6331 5729
rect 5920 5692 5948 5723
rect 2087 5664 3188 5692
rect 3344 5664 5948 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 2866 5584 2872 5636
rect 2924 5624 2930 5636
rect 3344 5624 3372 5664
rect 2924 5596 3372 5624
rect 2924 5584 2930 5596
rect 4706 5584 4712 5636
rect 4764 5584 4770 5636
rect 6288 5624 6316 5723
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 6564 5769 6592 5800
rect 7668 5772 7696 5800
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5729 6607 5763
rect 6825 5763 6883 5769
rect 6825 5760 6837 5763
rect 6549 5723 6607 5729
rect 6748 5732 6837 5760
rect 6748 5704 6776 5732
rect 6825 5729 6837 5732
rect 6871 5729 6883 5763
rect 6825 5723 6883 5729
rect 7006 5720 7012 5772
rect 7064 5760 7070 5772
rect 7101 5763 7159 5769
rect 7101 5760 7113 5763
rect 7064 5732 7113 5760
rect 7064 5720 7070 5732
rect 7101 5729 7113 5732
rect 7147 5760 7159 5763
rect 7282 5760 7288 5772
rect 7147 5732 7288 5760
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 7377 5763 7435 5769
rect 7377 5729 7389 5763
rect 7423 5760 7435 5763
rect 7558 5760 7564 5772
rect 7423 5732 7564 5760
rect 7423 5729 7435 5732
rect 7377 5723 7435 5729
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 7650 5720 7656 5772
rect 7708 5720 7714 5772
rect 7926 5720 7932 5772
rect 7984 5760 7990 5772
rect 8846 5760 8852 5772
rect 7984 5732 8852 5760
rect 7984 5720 7990 5732
rect 8846 5720 8852 5732
rect 8904 5760 8910 5772
rect 10244 5769 10272 5868
rect 12434 5856 12440 5868
rect 12492 5896 12498 5908
rect 13630 5896 13636 5908
rect 12492 5868 13636 5896
rect 12492 5856 12498 5868
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 16022 5896 16028 5908
rect 13924 5868 16028 5896
rect 10594 5788 10600 5840
rect 10652 5788 10658 5840
rect 11054 5788 11060 5840
rect 11112 5788 11118 5840
rect 11146 5788 11152 5840
rect 11204 5788 11210 5840
rect 13924 5828 13952 5868
rect 16022 5856 16028 5868
rect 16080 5896 16086 5908
rect 16482 5896 16488 5908
rect 16080 5868 16488 5896
rect 16080 5856 16086 5868
rect 16482 5856 16488 5868
rect 16540 5856 16546 5908
rect 16574 5856 16580 5908
rect 16632 5905 16638 5908
rect 16632 5896 16641 5905
rect 17126 5896 17132 5908
rect 16632 5868 17132 5896
rect 16632 5859 16641 5868
rect 16632 5856 16638 5859
rect 17126 5856 17132 5868
rect 17184 5856 17190 5908
rect 17954 5856 17960 5908
rect 18012 5856 18018 5908
rect 19058 5856 19064 5908
rect 19116 5896 19122 5908
rect 19116 5868 20300 5896
rect 19116 5856 19122 5868
rect 13648 5800 13952 5828
rect 10229 5763 10287 5769
rect 8904 5732 10183 5760
rect 8904 5720 8910 5732
rect 6730 5652 6736 5704
rect 6788 5652 6794 5704
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7837 5695 7895 5701
rect 7837 5692 7849 5695
rect 6972 5664 7849 5692
rect 6972 5652 6978 5664
rect 7837 5661 7849 5664
rect 7883 5661 7895 5695
rect 7837 5655 7895 5661
rect 8018 5652 8024 5704
rect 8076 5692 8082 5704
rect 8386 5701 8392 5704
rect 8164 5695 8222 5701
rect 8164 5692 8176 5695
rect 8076 5664 8176 5692
rect 8076 5652 8082 5664
rect 8164 5661 8176 5664
rect 8210 5661 8222 5695
rect 8164 5655 8222 5661
rect 8343 5695 8392 5701
rect 8343 5661 8355 5695
rect 8389 5661 8392 5695
rect 8343 5655 8392 5661
rect 8386 5652 8392 5655
rect 8444 5652 8450 5704
rect 8570 5652 8576 5704
rect 8628 5652 8634 5704
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5692 10011 5695
rect 10042 5692 10048 5704
rect 9999 5664 10048 5692
rect 9999 5661 10011 5664
rect 9953 5655 10011 5661
rect 10042 5652 10048 5664
rect 10100 5652 10106 5704
rect 10155 5692 10183 5732
rect 10229 5729 10241 5763
rect 10275 5729 10287 5763
rect 10229 5723 10287 5729
rect 10505 5763 10563 5769
rect 10505 5729 10517 5763
rect 10551 5760 10563 5763
rect 10612 5760 10640 5788
rect 10551 5732 10640 5760
rect 10781 5763 10839 5769
rect 10551 5729 10563 5732
rect 10505 5723 10563 5729
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 11072 5760 11100 5788
rect 10827 5732 11100 5760
rect 11164 5760 11192 5788
rect 11241 5763 11299 5769
rect 11241 5760 11253 5763
rect 11164 5732 11253 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 11241 5729 11253 5732
rect 11287 5760 11299 5763
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 11287 5732 11345 5760
rect 11287 5729 11299 5732
rect 11241 5723 11299 5729
rect 11333 5729 11345 5732
rect 11379 5729 11391 5763
rect 11333 5723 11391 5729
rect 10796 5692 10824 5723
rect 11422 5720 11428 5772
rect 11480 5760 11486 5772
rect 12345 5763 12403 5769
rect 11480 5732 12112 5760
rect 11480 5720 11486 5732
rect 10155 5664 10824 5692
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 11609 5695 11667 5701
rect 11609 5692 11621 5695
rect 11112 5664 11621 5692
rect 11112 5652 11118 5664
rect 11609 5661 11621 5664
rect 11655 5661 11667 5695
rect 11609 5655 11667 5661
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 12084 5701 12112 5732
rect 12345 5729 12357 5763
rect 12391 5760 12403 5763
rect 12618 5760 12624 5772
rect 12391 5732 12624 5760
rect 12391 5729 12403 5732
rect 12345 5723 12403 5729
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 11936 5695 11994 5701
rect 11936 5692 11948 5695
rect 11848 5664 11948 5692
rect 11848 5652 11854 5664
rect 11936 5661 11948 5664
rect 11982 5661 11994 5695
rect 11936 5655 11994 5661
rect 12072 5695 12130 5701
rect 12072 5661 12084 5695
rect 12118 5661 12130 5695
rect 12072 5655 12130 5661
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 13648 5692 13676 5800
rect 13725 5763 13783 5769
rect 13725 5729 13737 5763
rect 13771 5760 13783 5763
rect 13771 5732 14320 5760
rect 13771 5729 13783 5732
rect 13725 5723 13783 5729
rect 12492 5664 13676 5692
rect 12492 5652 12498 5664
rect 13814 5652 13820 5704
rect 13872 5652 13878 5704
rect 14182 5701 14188 5704
rect 14144 5695 14188 5701
rect 14144 5661 14156 5695
rect 14144 5655 14188 5661
rect 14182 5652 14188 5655
rect 14240 5652 14246 5704
rect 14292 5701 14320 5732
rect 14366 5720 14372 5772
rect 14424 5760 14430 5772
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 14424 5732 14565 5760
rect 14424 5720 14430 5732
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 16853 5763 16911 5769
rect 16853 5729 16865 5763
rect 16899 5760 16911 5763
rect 16942 5760 16948 5772
rect 16899 5732 16948 5760
rect 16899 5729 16911 5732
rect 16853 5723 16911 5729
rect 16942 5720 16948 5732
rect 17000 5720 17006 5772
rect 17972 5760 18000 5856
rect 20272 5828 20300 5868
rect 20346 5856 20352 5908
rect 20404 5856 20410 5908
rect 20714 5856 20720 5908
rect 20772 5896 20778 5908
rect 21269 5899 21327 5905
rect 21269 5896 21281 5899
rect 20772 5868 21281 5896
rect 20772 5856 20778 5868
rect 21269 5865 21281 5868
rect 21315 5865 21327 5899
rect 21269 5859 21327 5865
rect 22379 5899 22437 5905
rect 22379 5865 22391 5899
rect 22425 5896 22437 5899
rect 22922 5896 22928 5908
rect 22425 5868 22928 5896
rect 22425 5865 22437 5868
rect 22379 5859 22437 5865
rect 22922 5856 22928 5868
rect 22980 5856 22986 5908
rect 23382 5856 23388 5908
rect 23440 5896 23446 5908
rect 23440 5868 27568 5896
rect 23440 5856 23446 5868
rect 20272 5800 21956 5828
rect 19061 5763 19119 5769
rect 19061 5760 19073 5763
rect 17972 5732 19073 5760
rect 19061 5729 19073 5732
rect 19107 5729 19119 5763
rect 19061 5723 19119 5729
rect 19518 5720 19524 5772
rect 19576 5760 19582 5772
rect 20717 5763 20775 5769
rect 20717 5760 20729 5763
rect 19576 5732 20729 5760
rect 19576 5720 19582 5732
rect 20717 5729 20729 5732
rect 20763 5760 20775 5763
rect 20898 5760 20904 5772
rect 20763 5732 20904 5760
rect 20763 5729 20775 5732
rect 20717 5723 20775 5729
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 21008 5769 21036 5800
rect 20993 5763 21051 5769
rect 20993 5729 21005 5763
rect 21039 5729 21051 5763
rect 20993 5723 21051 5729
rect 21450 5720 21456 5772
rect 21508 5720 21514 5772
rect 21818 5720 21824 5772
rect 21876 5720 21882 5772
rect 21928 5760 21956 5800
rect 25590 5788 25596 5840
rect 25648 5828 25654 5840
rect 25648 5800 26648 5828
rect 25648 5788 25654 5800
rect 21928 5732 22508 5760
rect 14280 5695 14338 5701
rect 14280 5661 14292 5695
rect 14326 5661 14338 5695
rect 14280 5655 14338 5661
rect 16022 5652 16028 5704
rect 16080 5692 16086 5704
rect 16666 5701 16672 5704
rect 16117 5695 16175 5701
rect 16117 5692 16129 5695
rect 16080 5664 16129 5692
rect 16080 5652 16086 5664
rect 16117 5661 16129 5664
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 16623 5695 16672 5701
rect 16623 5661 16635 5695
rect 16669 5661 16672 5695
rect 16623 5655 16672 5661
rect 16666 5652 16672 5655
rect 16724 5652 16730 5704
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5692 18383 5695
rect 18506 5692 18512 5704
rect 18371 5664 18512 5692
rect 18371 5661 18383 5664
rect 18325 5655 18383 5661
rect 18506 5652 18512 5664
rect 18564 5652 18570 5704
rect 18690 5701 18696 5704
rect 18652 5695 18696 5701
rect 18652 5661 18664 5695
rect 18652 5655 18696 5661
rect 18690 5652 18696 5655
rect 18748 5652 18754 5704
rect 18782 5652 18788 5704
rect 18840 5652 18846 5704
rect 20438 5652 20444 5704
rect 20496 5692 20502 5704
rect 21468 5692 21496 5720
rect 20496 5664 21496 5692
rect 20496 5652 20502 5664
rect 21910 5652 21916 5704
rect 21968 5652 21974 5704
rect 22370 5652 22376 5704
rect 22428 5652 22434 5704
rect 22480 5692 22508 5732
rect 22554 5720 22560 5772
rect 22612 5760 22618 5772
rect 22649 5763 22707 5769
rect 22649 5760 22661 5763
rect 22612 5732 22661 5760
rect 22612 5720 22618 5732
rect 22649 5729 22661 5732
rect 22695 5729 22707 5763
rect 24121 5763 24179 5769
rect 24121 5760 24133 5763
rect 22649 5723 22707 5729
rect 23971 5732 24133 5760
rect 23566 5692 23572 5704
rect 22480 5664 23572 5692
rect 23566 5652 23572 5664
rect 23624 5652 23630 5704
rect 4816 5596 6316 5624
rect 3326 5516 3332 5568
rect 3384 5516 3390 5568
rect 3789 5559 3847 5565
rect 3789 5525 3801 5559
rect 3835 5556 3847 5559
rect 3878 5556 3884 5568
rect 3835 5528 3884 5556
rect 3835 5525 3847 5528
rect 3789 5519 3847 5525
rect 3878 5516 3884 5528
rect 3936 5516 3942 5568
rect 3970 5516 3976 5568
rect 4028 5556 4034 5568
rect 4816 5556 4844 5596
rect 6454 5584 6460 5636
rect 6512 5624 6518 5636
rect 7469 5627 7527 5633
rect 7469 5624 7481 5627
rect 6512 5596 7481 5624
rect 6512 5584 6518 5596
rect 7469 5593 7481 5596
rect 7515 5593 7527 5627
rect 7469 5587 7527 5593
rect 9398 5584 9404 5636
rect 9456 5624 9462 5636
rect 10597 5627 10655 5633
rect 10597 5624 10609 5627
rect 9456 5596 10609 5624
rect 9456 5584 9462 5596
rect 10597 5593 10609 5596
rect 10643 5593 10655 5627
rect 10597 5587 10655 5593
rect 10962 5584 10968 5636
rect 11020 5624 11026 5636
rect 11238 5624 11244 5636
rect 11020 5596 11244 5624
rect 11020 5584 11026 5596
rect 11238 5584 11244 5596
rect 11296 5584 11302 5636
rect 11514 5584 11520 5636
rect 11572 5584 11578 5636
rect 20533 5627 20591 5633
rect 20533 5593 20545 5627
rect 20579 5624 20591 5627
rect 21450 5624 21456 5636
rect 20579 5596 21456 5624
rect 20579 5593 20591 5596
rect 20533 5587 20591 5593
rect 21450 5584 21456 5596
rect 21508 5584 21514 5636
rect 23971 5624 23999 5732
rect 24121 5729 24133 5732
rect 24167 5729 24179 5763
rect 24121 5723 24179 5729
rect 24394 5720 24400 5772
rect 24452 5769 24458 5772
rect 24452 5763 24506 5769
rect 24452 5729 24460 5763
rect 24494 5729 24506 5763
rect 24452 5723 24506 5729
rect 24452 5720 24458 5723
rect 24762 5720 24768 5772
rect 24820 5760 24826 5772
rect 24857 5763 24915 5769
rect 24857 5760 24869 5763
rect 24820 5732 24869 5760
rect 24820 5720 24826 5732
rect 24857 5729 24869 5732
rect 24903 5729 24915 5763
rect 24857 5723 24915 5729
rect 26418 5720 26424 5772
rect 26476 5720 26482 5772
rect 26620 5769 26648 5800
rect 26718 5800 27476 5828
rect 26605 5763 26663 5769
rect 26605 5729 26617 5763
rect 26651 5760 26663 5763
rect 26718 5760 26746 5800
rect 26651 5732 26746 5760
rect 26651 5729 26663 5732
rect 26605 5723 26663 5729
rect 26786 5720 26792 5772
rect 26844 5760 26850 5772
rect 26881 5763 26939 5769
rect 26881 5760 26893 5763
rect 26844 5732 26893 5760
rect 26844 5720 26850 5732
rect 26881 5729 26893 5732
rect 26927 5729 26939 5763
rect 26881 5723 26939 5729
rect 27157 5763 27215 5769
rect 27157 5729 27169 5763
rect 27203 5760 27215 5763
rect 27246 5760 27252 5772
rect 27203 5732 27252 5760
rect 27203 5729 27215 5732
rect 27157 5723 27215 5729
rect 27246 5720 27252 5732
rect 27304 5720 27310 5772
rect 27448 5769 27476 5800
rect 27433 5763 27491 5769
rect 27433 5729 27445 5763
rect 27479 5729 27491 5763
rect 27540 5760 27568 5868
rect 27614 5856 27620 5908
rect 27672 5896 27678 5908
rect 29365 5899 29423 5905
rect 29365 5896 29377 5899
rect 27672 5868 29377 5896
rect 27672 5856 27678 5868
rect 29365 5865 29377 5868
rect 29411 5865 29423 5899
rect 29365 5859 29423 5865
rect 28261 5763 28319 5769
rect 27540 5732 28028 5760
rect 27433 5723 27491 5729
rect 24029 5695 24087 5701
rect 24029 5661 24041 5695
rect 24075 5692 24087 5695
rect 24584 5695 24642 5701
rect 24584 5692 24596 5695
rect 24075 5664 24596 5692
rect 24075 5661 24087 5664
rect 24029 5655 24087 5661
rect 24584 5661 24596 5664
rect 24630 5661 24642 5695
rect 24584 5655 24642 5661
rect 24670 5652 24676 5704
rect 24728 5692 24734 5704
rect 25866 5692 25872 5704
rect 24728 5664 25872 5692
rect 24728 5652 24734 5664
rect 25866 5652 25872 5664
rect 25924 5652 25930 5704
rect 26436 5692 26464 5720
rect 27522 5692 27528 5704
rect 26436 5664 27528 5692
rect 27522 5652 27528 5664
rect 27580 5652 27586 5704
rect 27890 5701 27896 5704
rect 27852 5695 27896 5701
rect 27852 5661 27864 5695
rect 27852 5655 27896 5661
rect 27890 5652 27896 5655
rect 27948 5652 27954 5704
rect 28000 5701 28028 5732
rect 28261 5729 28273 5763
rect 28307 5760 28319 5763
rect 28534 5760 28540 5772
rect 28307 5732 28540 5760
rect 28307 5729 28319 5732
rect 28261 5723 28319 5729
rect 28534 5720 28540 5732
rect 28592 5720 28598 5772
rect 27988 5695 28046 5701
rect 27988 5661 28000 5695
rect 28034 5661 28046 5695
rect 27988 5655 28046 5661
rect 24118 5624 24124 5636
rect 23971 5596 24124 5624
rect 24118 5584 24124 5596
rect 24176 5584 24182 5636
rect 26234 5624 26240 5636
rect 25516 5596 26240 5624
rect 4028 5528 4844 5556
rect 4028 5516 4034 5528
rect 5166 5516 5172 5568
rect 5224 5516 5230 5568
rect 6638 5516 6644 5568
rect 6696 5516 6702 5568
rect 6914 5516 6920 5568
rect 6972 5516 6978 5568
rect 7193 5559 7251 5565
rect 7193 5525 7205 5559
rect 7239 5556 7251 5559
rect 7374 5556 7380 5568
rect 7239 5528 7380 5556
rect 7239 5525 7251 5528
rect 7193 5519 7251 5525
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 7834 5516 7840 5568
rect 7892 5556 7898 5568
rect 9582 5556 9588 5568
rect 7892 5528 9588 5556
rect 7892 5516 7898 5528
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 9766 5516 9772 5568
rect 9824 5556 9830 5568
rect 10045 5559 10103 5565
rect 10045 5556 10057 5559
rect 9824 5528 10057 5556
rect 9824 5516 9830 5528
rect 10045 5525 10057 5528
rect 10091 5525 10103 5559
rect 10045 5519 10103 5525
rect 10321 5559 10379 5565
rect 10321 5525 10333 5559
rect 10367 5556 10379 5559
rect 10502 5556 10508 5568
rect 10367 5528 10508 5556
rect 10367 5525 10379 5528
rect 10321 5519 10379 5525
rect 10502 5516 10508 5528
rect 10560 5516 10566 5568
rect 11057 5559 11115 5565
rect 11057 5525 11069 5559
rect 11103 5556 11115 5559
rect 11330 5556 11336 5568
rect 11103 5528 11336 5556
rect 11103 5525 11115 5528
rect 11057 5519 11115 5525
rect 11330 5516 11336 5528
rect 11388 5516 11394 5568
rect 15841 5559 15899 5565
rect 15841 5525 15853 5559
rect 15887 5556 15899 5559
rect 16390 5556 16396 5568
rect 15887 5528 16396 5556
rect 15887 5525 15899 5528
rect 15841 5519 15899 5525
rect 16390 5516 16396 5528
rect 16448 5516 16454 5568
rect 18138 5516 18144 5568
rect 18196 5516 18202 5568
rect 18230 5516 18236 5568
rect 18288 5556 18294 5568
rect 19242 5556 19248 5568
rect 18288 5528 19248 5556
rect 18288 5516 18294 5528
rect 19242 5516 19248 5528
rect 19300 5516 19306 5568
rect 19978 5516 19984 5568
rect 20036 5556 20042 5568
rect 20714 5556 20720 5568
rect 20036 5528 20720 5556
rect 20036 5516 20042 5528
rect 20714 5516 20720 5528
rect 20772 5516 20778 5568
rect 20806 5516 20812 5568
rect 20864 5516 20870 5568
rect 21637 5559 21695 5565
rect 21637 5525 21649 5559
rect 21683 5556 21695 5559
rect 22554 5556 22560 5568
rect 21683 5528 22560 5556
rect 21683 5525 21695 5528
rect 21637 5519 21695 5525
rect 22554 5516 22560 5528
rect 22612 5516 22618 5568
rect 22738 5516 22744 5568
rect 22796 5556 22802 5568
rect 25516 5556 25544 5596
rect 26234 5584 26240 5596
rect 26292 5584 26298 5636
rect 26421 5627 26479 5633
rect 26421 5593 26433 5627
rect 26467 5624 26479 5627
rect 26786 5624 26792 5636
rect 26467 5596 26792 5624
rect 26467 5593 26479 5596
rect 26421 5587 26479 5593
rect 26786 5584 26792 5596
rect 26844 5584 26850 5636
rect 22796 5528 25544 5556
rect 22796 5516 22802 5528
rect 26142 5516 26148 5568
rect 26200 5516 26206 5568
rect 26602 5516 26608 5568
rect 26660 5556 26666 5568
rect 26697 5559 26755 5565
rect 26697 5556 26709 5559
rect 26660 5528 26709 5556
rect 26660 5516 26666 5528
rect 26697 5525 26709 5528
rect 26743 5525 26755 5559
rect 26697 5519 26755 5525
rect 26878 5516 26884 5568
rect 26936 5556 26942 5568
rect 26973 5559 27031 5565
rect 26973 5556 26985 5559
rect 26936 5528 26985 5556
rect 26936 5516 26942 5528
rect 26973 5525 26985 5528
rect 27019 5525 27031 5559
rect 26973 5519 27031 5525
rect 27249 5559 27307 5565
rect 27249 5525 27261 5559
rect 27295 5556 27307 5559
rect 28166 5556 28172 5568
rect 27295 5528 28172 5556
rect 27295 5525 27307 5528
rect 27249 5519 27307 5525
rect 28166 5516 28172 5528
rect 28224 5516 28230 5568
rect 552 5466 30912 5488
rect 552 5414 4193 5466
rect 4245 5414 4257 5466
rect 4309 5414 4321 5466
rect 4373 5414 4385 5466
rect 4437 5414 4449 5466
rect 4501 5414 11783 5466
rect 11835 5414 11847 5466
rect 11899 5414 11911 5466
rect 11963 5414 11975 5466
rect 12027 5414 12039 5466
rect 12091 5414 19373 5466
rect 19425 5414 19437 5466
rect 19489 5414 19501 5466
rect 19553 5414 19565 5466
rect 19617 5414 19629 5466
rect 19681 5414 26963 5466
rect 27015 5414 27027 5466
rect 27079 5414 27091 5466
rect 27143 5414 27155 5466
rect 27207 5414 27219 5466
rect 27271 5414 30912 5466
rect 552 5392 30912 5414
rect 934 5312 940 5364
rect 992 5352 998 5364
rect 2498 5352 2504 5364
rect 992 5324 2504 5352
rect 992 5312 998 5324
rect 2498 5312 2504 5324
rect 2556 5352 2562 5364
rect 3237 5355 3295 5361
rect 2556 5324 2820 5352
rect 2556 5312 2562 5324
rect 937 5219 995 5225
rect 937 5185 949 5219
rect 983 5216 995 5219
rect 1302 5216 1308 5228
rect 983 5188 1308 5216
rect 983 5185 995 5188
rect 937 5179 995 5185
rect 1302 5176 1308 5188
rect 1360 5176 1366 5228
rect 1443 5219 1501 5225
rect 1443 5185 1455 5219
rect 1489 5216 1501 5219
rect 2590 5216 2596 5228
rect 1489 5188 2596 5216
rect 1489 5185 1501 5188
rect 1443 5179 1501 5185
rect 2590 5176 2596 5188
rect 2648 5176 2654 5228
rect 1673 5151 1731 5157
rect 1673 5117 1685 5151
rect 1719 5148 1731 5151
rect 2314 5148 2320 5160
rect 1719 5120 2320 5148
rect 1719 5117 1731 5120
rect 1673 5111 1731 5117
rect 2314 5108 2320 5120
rect 2372 5108 2378 5160
rect 2792 5148 2820 5324
rect 3237 5321 3249 5355
rect 3283 5352 3295 5355
rect 4982 5352 4988 5364
rect 3283 5324 4988 5352
rect 3283 5321 3295 5324
rect 3237 5315 3295 5321
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 6546 5352 6552 5364
rect 6104 5324 6552 5352
rect 2866 5176 2872 5228
rect 2924 5216 2930 5228
rect 3234 5216 3240 5228
rect 2924 5188 3240 5216
rect 2924 5176 2930 5188
rect 3234 5176 3240 5188
rect 3292 5216 3298 5228
rect 6104 5225 6132 5324
rect 6546 5312 6552 5324
rect 6604 5352 6610 5364
rect 6822 5352 6828 5364
rect 6604 5324 6828 5352
rect 6604 5312 6610 5324
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 8754 5352 8760 5364
rect 7064 5324 8760 5352
rect 7064 5312 7070 5324
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 9214 5312 9220 5364
rect 9272 5352 9278 5364
rect 11146 5352 11152 5364
rect 9272 5324 11152 5352
rect 9272 5312 9278 5324
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 15657 5355 15715 5361
rect 15657 5321 15669 5355
rect 15703 5352 15715 5355
rect 16666 5352 16672 5364
rect 15703 5324 16672 5352
rect 15703 5321 15715 5324
rect 15657 5315 15715 5321
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 16942 5312 16948 5364
rect 17000 5352 17006 5364
rect 21358 5352 21364 5364
rect 17000 5324 21364 5352
rect 17000 5312 17006 5324
rect 21358 5312 21364 5324
rect 21416 5312 21422 5364
rect 21542 5312 21548 5364
rect 21600 5352 21606 5364
rect 24670 5352 24676 5364
rect 21600 5324 24676 5352
rect 21600 5312 21606 5324
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 24762 5312 24768 5364
rect 24820 5352 24826 5364
rect 26053 5355 26111 5361
rect 26053 5352 26065 5355
rect 24820 5324 26065 5352
rect 24820 5312 24826 5324
rect 26053 5321 26065 5324
rect 26099 5321 26111 5355
rect 29457 5355 29515 5361
rect 29457 5352 29469 5355
rect 26053 5315 26111 5321
rect 26160 5324 29469 5352
rect 8113 5287 8171 5293
rect 8113 5253 8125 5287
rect 8159 5284 8171 5287
rect 26160 5284 26188 5324
rect 29457 5321 29469 5324
rect 29503 5321 29515 5355
rect 29457 5315 29515 5321
rect 8159 5256 8708 5284
rect 8159 5253 8171 5256
rect 8113 5247 8171 5253
rect 3513 5219 3571 5225
rect 3513 5216 3525 5219
rect 3292 5188 3525 5216
rect 3292 5176 3298 5188
rect 3513 5185 3525 5188
rect 3559 5185 3571 5219
rect 3976 5219 4034 5225
rect 3976 5216 3988 5219
rect 3513 5179 3571 5185
rect 3855 5188 3988 5216
rect 3421 5151 3479 5157
rect 3421 5148 3433 5151
rect 2792 5120 3433 5148
rect 3421 5117 3433 5120
rect 3467 5117 3479 5151
rect 3855 5148 3883 5188
rect 3976 5185 3988 5188
rect 4022 5185 4034 5219
rect 3976 5179 4034 5185
rect 6089 5219 6147 5225
rect 6089 5185 6101 5219
rect 6135 5185 6147 5219
rect 6089 5179 6147 5185
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 6552 5219 6610 5225
rect 6552 5216 6564 5219
rect 6328 5188 6564 5216
rect 6328 5176 6334 5188
rect 6552 5185 6564 5188
rect 6598 5185 6610 5219
rect 6552 5179 6610 5185
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 7466 5216 7472 5228
rect 6788 5188 7472 5216
rect 6788 5176 6794 5188
rect 7466 5176 7472 5188
rect 7524 5216 7530 5228
rect 7926 5216 7932 5228
rect 7524 5188 7932 5216
rect 7524 5176 7530 5188
rect 7926 5176 7932 5188
rect 7984 5176 7990 5228
rect 8478 5176 8484 5228
rect 8536 5216 8542 5228
rect 8536 5188 8616 5216
rect 8536 5176 8542 5188
rect 3421 5111 3479 5117
rect 3620 5120 3883 5148
rect 4249 5151 4307 5157
rect 3053 5083 3111 5089
rect 3053 5049 3065 5083
rect 3099 5080 3111 5083
rect 3620 5080 3648 5120
rect 4249 5117 4261 5151
rect 4295 5148 4307 5151
rect 4522 5148 4528 5160
rect 4295 5120 4528 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 6825 5151 6883 5157
rect 8588 5153 8616 5188
rect 8680 5214 8708 5256
rect 25792 5256 26188 5284
rect 9496 5217 9554 5223
rect 9496 5216 9508 5217
rect 8864 5214 9508 5216
rect 8680 5188 9508 5214
rect 8680 5186 8892 5188
rect 9496 5183 9508 5188
rect 9542 5183 9554 5217
rect 9496 5177 9554 5183
rect 9766 5176 9772 5228
rect 9824 5176 9830 5228
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 11704 5219 11762 5225
rect 11704 5216 11716 5219
rect 11195 5188 11716 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11704 5185 11716 5188
rect 11750 5185 11762 5219
rect 11704 5179 11762 5185
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 12158 5216 12164 5228
rect 12023 5188 12164 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 13357 5219 13415 5225
rect 13357 5185 13369 5219
rect 13403 5216 13415 5219
rect 14096 5219 14154 5225
rect 14096 5216 14108 5219
rect 13403 5188 14108 5216
rect 13403 5185 13415 5188
rect 13357 5179 13415 5185
rect 14096 5185 14108 5188
rect 14142 5185 14154 5219
rect 14096 5179 14154 5185
rect 14182 5176 14188 5228
rect 14240 5176 14246 5228
rect 14550 5176 14556 5228
rect 14608 5176 14614 5228
rect 16114 5176 16120 5228
rect 16172 5216 16178 5228
rect 16304 5219 16362 5225
rect 16304 5216 16316 5219
rect 16172 5188 16316 5216
rect 16172 5176 16178 5188
rect 16304 5185 16316 5188
rect 16350 5185 16362 5219
rect 16304 5179 16362 5185
rect 16577 5219 16635 5225
rect 16577 5185 16589 5219
rect 16623 5216 16635 5219
rect 17402 5216 17408 5228
rect 16623 5188 17408 5216
rect 16623 5185 16635 5188
rect 16577 5179 16635 5185
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 18138 5176 18144 5228
rect 18196 5216 18202 5228
rect 19156 5219 19214 5225
rect 19156 5216 19168 5219
rect 18196 5188 19168 5216
rect 18196 5176 18202 5188
rect 19156 5185 19168 5188
rect 19202 5185 19214 5219
rect 19156 5179 19214 5185
rect 19260 5188 20668 5216
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 6871 5120 8524 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 8018 5080 8024 5092
rect 3099 5052 3648 5080
rect 7760 5052 8024 5080
rect 3099 5049 3111 5052
rect 3053 5043 3111 5049
rect 1403 5015 1461 5021
rect 1403 4981 1415 5015
rect 1449 5012 1461 5015
rect 1578 5012 1584 5024
rect 1449 4984 1584 5012
rect 1449 4981 1461 4984
rect 1403 4975 1461 4981
rect 1578 4972 1584 4984
rect 1636 5012 1642 5024
rect 1762 5012 1768 5024
rect 1636 4984 1768 5012
rect 1636 4972 1642 4984
rect 1762 4972 1768 4984
rect 1820 4972 1826 5024
rect 3970 4972 3976 5024
rect 4028 5021 4034 5024
rect 4028 5012 4037 5021
rect 5353 5015 5411 5021
rect 4028 4984 4073 5012
rect 4028 4975 4037 4984
rect 5353 4981 5365 5015
rect 5399 5012 5411 5015
rect 5442 5012 5448 5024
rect 5399 4984 5448 5012
rect 5399 4981 5411 4984
rect 5353 4975 5411 4981
rect 4028 4972 4034 4975
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 6555 5015 6613 5021
rect 6555 4981 6567 5015
rect 6601 5012 6613 5015
rect 6914 5012 6920 5024
rect 6601 4984 6920 5012
rect 6601 4981 6613 4984
rect 6555 4975 6613 4981
rect 6914 4972 6920 4984
rect 6972 5012 6978 5024
rect 7760 5012 7788 5052
rect 8018 5040 8024 5052
rect 8076 5040 8082 5092
rect 6972 4984 7788 5012
rect 6972 4972 6978 4984
rect 7834 4972 7840 5024
rect 7892 5012 7898 5024
rect 8389 5015 8447 5021
rect 8389 5012 8401 5015
rect 7892 4984 8401 5012
rect 7892 4972 7898 4984
rect 8389 4981 8401 4984
rect 8435 4981 8447 5015
rect 8496 5012 8524 5120
rect 8581 5147 8639 5153
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 8581 5113 8593 5147
rect 8627 5113 8639 5147
rect 8581 5107 8639 5113
rect 8772 5120 8861 5148
rect 8772 5092 8800 5120
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 9033 5151 9091 5157
rect 9033 5117 9045 5151
rect 9079 5117 9091 5151
rect 9033 5111 9091 5117
rect 8754 5040 8760 5092
rect 8812 5040 8818 5092
rect 9048 5080 9076 5111
rect 9582 5108 9588 5160
rect 9640 5148 9646 5160
rect 9640 5120 11008 5148
rect 9640 5108 9646 5120
rect 8864 5052 9076 5080
rect 10980 5080 11008 5120
rect 11054 5108 11060 5160
rect 11112 5148 11118 5160
rect 11241 5151 11299 5157
rect 11241 5148 11253 5151
rect 11112 5120 11253 5148
rect 11112 5108 11118 5120
rect 11241 5117 11253 5120
rect 11287 5117 11299 5151
rect 13446 5148 13452 5160
rect 11241 5111 11299 5117
rect 11348 5120 13452 5148
rect 11348 5080 11376 5120
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 13633 5151 13691 5157
rect 13633 5117 13645 5151
rect 13679 5148 13691 5151
rect 13722 5148 13728 5160
rect 13679 5120 13728 5148
rect 13679 5117 13691 5120
rect 13633 5111 13691 5117
rect 13722 5108 13728 5120
rect 13780 5108 13786 5160
rect 13960 5151 14018 5157
rect 13960 5117 13972 5151
rect 14006 5148 14018 5151
rect 14200 5148 14228 5176
rect 14006 5120 14228 5148
rect 14369 5151 14427 5157
rect 14006 5117 14018 5120
rect 13960 5111 14018 5117
rect 14369 5117 14381 5151
rect 14415 5148 14427 5151
rect 14568 5148 14596 5176
rect 14415 5120 14596 5148
rect 14415 5117 14427 5120
rect 14369 5111 14427 5117
rect 15838 5108 15844 5160
rect 15896 5108 15902 5160
rect 17310 5108 17316 5160
rect 17368 5148 17374 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 17368 5120 18061 5148
rect 17368 5108 17374 5120
rect 18049 5117 18061 5120
rect 18095 5148 18107 5151
rect 18230 5148 18236 5160
rect 18095 5120 18236 5148
rect 18095 5117 18107 5120
rect 18049 5111 18107 5117
rect 18230 5108 18236 5120
rect 18288 5108 18294 5160
rect 18506 5108 18512 5160
rect 18564 5148 18570 5160
rect 18693 5151 18751 5157
rect 18693 5148 18705 5151
rect 18564 5120 18705 5148
rect 18564 5108 18570 5120
rect 18693 5117 18705 5120
rect 18739 5117 18751 5151
rect 18693 5111 18751 5117
rect 18966 5108 18972 5160
rect 19024 5148 19030 5160
rect 19260 5148 19288 5188
rect 19024 5120 19288 5148
rect 19429 5151 19487 5157
rect 19024 5108 19030 5120
rect 19429 5117 19441 5151
rect 19475 5148 19487 5151
rect 19702 5148 19708 5160
rect 19475 5120 19708 5148
rect 19475 5117 19487 5120
rect 19429 5111 19487 5117
rect 19702 5108 19708 5120
rect 19760 5108 19766 5160
rect 10980 5052 11376 5080
rect 8864 5024 8892 5052
rect 17954 5040 17960 5092
rect 18012 5040 18018 5092
rect 18325 5083 18383 5089
rect 18325 5049 18337 5083
rect 18371 5049 18383 5083
rect 18325 5043 18383 5049
rect 8665 5015 8723 5021
rect 8665 5012 8677 5015
rect 8496 4984 8677 5012
rect 8389 4975 8447 4981
rect 8665 4981 8677 4984
rect 8711 4981 8723 5015
rect 8665 4975 8723 4981
rect 8846 4972 8852 5024
rect 8904 4972 8910 5024
rect 9030 4972 9036 5024
rect 9088 5012 9094 5024
rect 9499 5015 9557 5021
rect 9499 5012 9511 5015
rect 9088 4984 9511 5012
rect 9088 4972 9094 4984
rect 9499 4981 9511 4984
rect 9545 4981 9557 5015
rect 9499 4975 9557 4981
rect 11698 4972 11704 5024
rect 11756 5021 11762 5024
rect 11756 5012 11765 5021
rect 16307 5015 16365 5021
rect 11756 4984 11801 5012
rect 11756 4975 11765 4984
rect 16307 4981 16319 5015
rect 16353 5012 16365 5015
rect 16574 5012 16580 5024
rect 16353 4984 16580 5012
rect 16353 4981 16365 4984
rect 16307 4975 16365 4981
rect 11756 4972 11762 4975
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 18340 5012 18368 5043
rect 18690 5012 18696 5024
rect 18340 4984 18696 5012
rect 18690 4972 18696 4984
rect 18748 5012 18754 5024
rect 18966 5012 18972 5024
rect 18748 4984 18972 5012
rect 18748 4972 18754 4984
rect 18966 4972 18972 4984
rect 19024 5012 19030 5024
rect 19159 5015 19217 5021
rect 19159 5012 19171 5015
rect 19024 4984 19171 5012
rect 19024 4972 19030 4984
rect 19159 4981 19171 4984
rect 19205 4981 19217 5015
rect 20640 5012 20668 5188
rect 20714 5176 20720 5228
rect 20772 5176 20778 5228
rect 20809 5219 20867 5225
rect 20809 5185 20821 5219
rect 20855 5216 20867 5219
rect 21364 5219 21422 5225
rect 21364 5216 21376 5219
rect 20855 5188 21376 5216
rect 20855 5185 20867 5188
rect 20809 5179 20867 5185
rect 21364 5185 21376 5188
rect 21410 5185 21422 5219
rect 21364 5179 21422 5185
rect 21450 5176 21456 5228
rect 21508 5216 21514 5228
rect 21637 5219 21695 5225
rect 21637 5216 21649 5219
rect 21508 5188 21649 5216
rect 21508 5176 21514 5188
rect 21637 5185 21649 5188
rect 21683 5185 21695 5219
rect 21637 5179 21695 5185
rect 23750 5176 23756 5228
rect 23808 5216 23814 5228
rect 23808 5188 23980 5216
rect 23808 5176 23814 5188
rect 20732 5148 20760 5176
rect 20901 5151 20959 5157
rect 20901 5148 20913 5151
rect 20732 5120 20913 5148
rect 20901 5117 20913 5120
rect 20947 5117 20959 5151
rect 20901 5111 20959 5117
rect 20990 5108 20996 5160
rect 21048 5148 21054 5160
rect 21228 5151 21286 5157
rect 21228 5148 21240 5151
rect 21048 5120 21240 5148
rect 21048 5108 21054 5120
rect 21228 5117 21240 5120
rect 21274 5117 21286 5151
rect 21228 5111 21286 5117
rect 21910 5108 21916 5160
rect 21968 5148 21974 5160
rect 23845 5151 23903 5157
rect 23845 5148 23857 5151
rect 21968 5120 23857 5148
rect 21968 5108 21974 5120
rect 23845 5117 23857 5120
rect 23891 5117 23903 5151
rect 23952 5148 23980 5188
rect 24026 5176 24032 5228
rect 24084 5216 24090 5228
rect 24308 5219 24366 5225
rect 24308 5216 24320 5219
rect 24084 5188 24320 5216
rect 24084 5176 24090 5188
rect 24308 5185 24320 5188
rect 24354 5185 24366 5219
rect 24308 5179 24366 5185
rect 24670 5176 24676 5228
rect 24728 5216 24734 5228
rect 25792 5216 25820 5256
rect 28442 5244 28448 5296
rect 28500 5284 28506 5296
rect 28537 5287 28595 5293
rect 28537 5284 28549 5287
rect 28500 5256 28549 5284
rect 28500 5244 28506 5256
rect 28537 5253 28549 5256
rect 28583 5253 28595 5287
rect 28537 5247 28595 5253
rect 29178 5244 29184 5296
rect 29236 5244 29242 5296
rect 24728 5188 25820 5216
rect 24728 5176 24734 5188
rect 26326 5176 26332 5228
rect 26384 5216 26390 5228
rect 27160 5219 27218 5225
rect 27160 5216 27172 5219
rect 26384 5188 27172 5216
rect 26384 5176 26390 5188
rect 27160 5185 27172 5188
rect 27206 5185 27218 5219
rect 27160 5179 27218 5185
rect 27433 5219 27491 5225
rect 27433 5185 27445 5219
rect 27479 5216 27491 5219
rect 28994 5216 29000 5228
rect 27479 5188 29000 5216
rect 27479 5185 27491 5188
rect 27433 5179 27491 5185
rect 28994 5176 29000 5188
rect 29052 5176 29058 5228
rect 24581 5151 24639 5157
rect 24581 5148 24593 5151
rect 23952 5120 24593 5148
rect 23845 5111 23903 5117
rect 24581 5117 24593 5120
rect 24627 5117 24639 5151
rect 24581 5111 24639 5117
rect 26234 5108 26240 5160
rect 26292 5108 26298 5160
rect 26418 5108 26424 5160
rect 26476 5148 26482 5160
rect 29196 5157 29224 5244
rect 26697 5151 26755 5157
rect 26697 5148 26709 5151
rect 26476 5120 26709 5148
rect 26476 5108 26482 5120
rect 26697 5117 26709 5120
rect 26743 5117 26755 5151
rect 29181 5151 29239 5157
rect 26697 5111 26755 5117
rect 26804 5120 29132 5148
rect 23293 5083 23351 5089
rect 23293 5080 23305 5083
rect 22391 5052 23305 5080
rect 22391 5012 22419 5052
rect 23293 5049 23305 5052
rect 23339 5080 23351 5083
rect 23658 5080 23664 5092
rect 23339 5052 23664 5080
rect 23339 5049 23351 5052
rect 23293 5043 23351 5049
rect 23658 5040 23664 5052
rect 23716 5040 23722 5092
rect 23750 5040 23756 5092
rect 23808 5080 23814 5092
rect 23934 5080 23940 5092
rect 23808 5052 23940 5080
rect 23808 5040 23814 5052
rect 23934 5040 23940 5052
rect 23992 5040 23998 5092
rect 26510 5040 26516 5092
rect 26568 5080 26574 5092
rect 26804 5080 26832 5120
rect 26568 5052 26832 5080
rect 29104 5080 29132 5120
rect 29181 5117 29193 5151
rect 29227 5117 29239 5151
rect 29181 5111 29239 5117
rect 29273 5151 29331 5157
rect 29273 5117 29285 5151
rect 29319 5117 29331 5151
rect 29273 5111 29331 5117
rect 29288 5080 29316 5111
rect 29104 5052 29316 5080
rect 26568 5040 26574 5052
rect 20640 4984 22419 5012
rect 19159 4975 19217 4981
rect 22462 4972 22468 5024
rect 22520 5012 22526 5024
rect 22741 5015 22799 5021
rect 22741 5012 22753 5015
rect 22520 4984 22753 5012
rect 22520 4972 22526 4984
rect 22741 4981 22753 4984
rect 22787 4981 22799 5015
rect 22741 4975 22799 4981
rect 22922 4972 22928 5024
rect 22980 5012 22986 5024
rect 24311 5015 24369 5021
rect 24311 5012 24323 5015
rect 22980 4984 24323 5012
rect 22980 4972 22986 4984
rect 24311 4981 24323 4984
rect 24357 4981 24369 5015
rect 24311 4975 24369 4981
rect 24946 4972 24952 5024
rect 25004 5012 25010 5024
rect 25685 5015 25743 5021
rect 25685 5012 25697 5015
rect 25004 4984 25697 5012
rect 25004 4972 25010 4984
rect 25685 4981 25697 4984
rect 25731 4981 25743 5015
rect 25685 4975 25743 4981
rect 27163 5015 27221 5021
rect 27163 4981 27175 5015
rect 27209 5012 27221 5015
rect 27890 5012 27896 5024
rect 27209 4984 27896 5012
rect 27209 4981 27221 4984
rect 27163 4975 27221 4981
rect 27890 4972 27896 4984
rect 27948 4972 27954 5024
rect 28994 4972 29000 5024
rect 29052 4972 29058 5024
rect 552 4922 31072 4944
rect 552 4870 7988 4922
rect 8040 4870 8052 4922
rect 8104 4870 8116 4922
rect 8168 4870 8180 4922
rect 8232 4870 8244 4922
rect 8296 4870 15578 4922
rect 15630 4870 15642 4922
rect 15694 4870 15706 4922
rect 15758 4870 15770 4922
rect 15822 4870 15834 4922
rect 15886 4870 23168 4922
rect 23220 4870 23232 4922
rect 23284 4870 23296 4922
rect 23348 4870 23360 4922
rect 23412 4870 23424 4922
rect 23476 4870 30758 4922
rect 30810 4870 30822 4922
rect 30874 4870 30886 4922
rect 30938 4870 30950 4922
rect 31002 4870 31014 4922
rect 31066 4870 31072 4922
rect 552 4848 31072 4870
rect 842 4768 848 4820
rect 900 4808 906 4820
rect 937 4811 995 4817
rect 937 4808 949 4811
rect 900 4780 949 4808
rect 900 4768 906 4780
rect 937 4777 949 4780
rect 983 4777 995 4811
rect 2866 4808 2872 4820
rect 937 4771 995 4777
rect 1136 4780 2872 4808
rect 1136 4681 1164 4780
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 3142 4768 3148 4820
rect 3200 4768 3206 4820
rect 5537 4811 5595 4817
rect 3252 4780 4936 4808
rect 3252 4740 3280 4780
rect 3068 4712 3280 4740
rect 4908 4740 4936 4780
rect 5537 4777 5549 4811
rect 5583 4808 5595 4811
rect 6270 4808 6276 4820
rect 5583 4780 6276 4808
rect 5583 4777 5595 4780
rect 5537 4771 5595 4777
rect 6270 4768 6276 4780
rect 6328 4768 6334 4820
rect 6914 4768 6920 4820
rect 6972 4817 6978 4820
rect 6972 4808 6981 4817
rect 6972 4780 7017 4808
rect 6972 4771 6981 4780
rect 6972 4768 6978 4771
rect 7834 4768 7840 4820
rect 7892 4768 7898 4820
rect 8478 4768 8484 4820
rect 8536 4808 8542 4820
rect 9214 4808 9220 4820
rect 8536 4780 9220 4808
rect 8536 4768 8542 4780
rect 9214 4768 9220 4780
rect 9272 4768 9278 4820
rect 10689 4811 10747 4817
rect 10689 4777 10701 4811
rect 10735 4808 10747 4811
rect 11422 4808 11428 4820
rect 10735 4780 11428 4808
rect 10735 4777 10747 4780
rect 10689 4771 10747 4777
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 11698 4768 11704 4820
rect 11756 4808 11762 4820
rect 12075 4811 12133 4817
rect 12075 4808 12087 4811
rect 11756 4780 12087 4808
rect 11756 4768 11762 4780
rect 12075 4777 12087 4780
rect 12121 4777 12133 4811
rect 12075 4771 12133 4777
rect 14182 4768 14188 4820
rect 14240 4808 14246 4820
rect 14283 4811 14341 4817
rect 14283 4808 14295 4811
rect 14240 4780 14295 4808
rect 14240 4768 14246 4780
rect 14283 4777 14295 4780
rect 14329 4777 14341 4811
rect 14283 4771 14341 4777
rect 16574 4768 16580 4820
rect 16632 4817 16638 4820
rect 16632 4808 16641 4817
rect 16632 4780 16677 4808
rect 16632 4771 16641 4780
rect 16632 4768 16638 4771
rect 17954 4768 17960 4820
rect 18012 4768 18018 4820
rect 18141 4811 18199 4817
rect 18141 4777 18153 4811
rect 18187 4808 18199 4811
rect 18690 4808 18696 4820
rect 18187 4780 18696 4808
rect 18187 4777 18199 4780
rect 18141 4771 18199 4777
rect 18690 4768 18696 4780
rect 18748 4768 18754 4820
rect 18791 4811 18849 4817
rect 18791 4777 18803 4811
rect 18837 4808 18849 4811
rect 18966 4808 18972 4820
rect 18837 4780 18972 4808
rect 18837 4777 18849 4780
rect 18791 4771 18849 4777
rect 18966 4768 18972 4780
rect 19024 4768 19030 4820
rect 27065 4811 27123 4817
rect 27065 4808 27077 4811
rect 19720 4780 27077 4808
rect 4908 4712 5948 4740
rect 1121 4675 1179 4681
rect 1121 4641 1133 4675
rect 1167 4641 1179 4675
rect 1121 4635 1179 4641
rect 1302 4632 1308 4684
rect 1360 4632 1366 4684
rect 1578 4632 1584 4684
rect 1636 4681 1642 4684
rect 1636 4675 1690 4681
rect 1636 4641 1644 4675
rect 1678 4641 1690 4675
rect 2774 4672 2780 4684
rect 1636 4635 1690 4641
rect 1964 4644 2780 4672
rect 1636 4632 1642 4635
rect 1801 4625 1859 4631
rect 1801 4591 1813 4625
rect 1847 4604 1859 4625
rect 1964 4604 1992 4644
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 1847 4591 1992 4604
rect 1801 4585 1992 4591
rect 1826 4576 1992 4585
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4604 2099 4607
rect 3068 4604 3096 4712
rect 3513 4675 3571 4681
rect 3513 4641 3525 4675
rect 3559 4672 3571 4675
rect 3602 4672 3608 4684
rect 3559 4644 3608 4672
rect 3559 4641 3571 4644
rect 3513 4635 3571 4641
rect 3602 4632 3608 4644
rect 3660 4632 3666 4684
rect 4172 4644 5304 4672
rect 3840 4607 3898 4613
rect 3840 4604 3852 4607
rect 2087 4576 3096 4604
rect 3528 4576 3852 4604
rect 2087 4573 2099 4576
rect 2041 4567 2099 4573
rect 3528 4548 3556 4576
rect 3840 4573 3852 4576
rect 3886 4573 3898 4607
rect 3840 4567 3898 4573
rect 4019 4607 4077 4613
rect 4019 4573 4031 4607
rect 4065 4604 4077 4607
rect 4172 4604 4200 4644
rect 5276 4616 5304 4644
rect 5810 4632 5816 4684
rect 5868 4632 5874 4684
rect 5920 4672 5948 4712
rect 7852 4672 7880 4768
rect 15933 4743 15991 4749
rect 15933 4709 15945 4743
rect 15979 4740 15991 4743
rect 16114 4740 16120 4752
rect 15979 4712 16120 4740
rect 15979 4709 15991 4712
rect 15933 4703 15991 4709
rect 16114 4700 16120 4712
rect 16172 4700 16178 4752
rect 5920 4644 7880 4672
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4672 8631 4675
rect 8619 4644 9168 4672
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 4065 4576 4200 4604
rect 4249 4607 4307 4613
rect 4065 4573 4077 4576
rect 4019 4567 4077 4573
rect 4249 4573 4261 4607
rect 4295 4604 4307 4607
rect 4890 4604 4896 4616
rect 4295 4576 4896 4604
rect 4295 4573 4307 4576
rect 4249 4567 4307 4573
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 5258 4564 5264 4616
rect 5316 4564 5322 4616
rect 5994 4604 6000 4616
rect 5368 4576 6000 4604
rect 3510 4496 3516 4548
rect 3568 4496 3574 4548
rect 5368 4536 5396 4576
rect 5994 4564 6000 4576
rect 6052 4564 6058 4616
rect 6454 4564 6460 4616
rect 6512 4564 6518 4616
rect 6963 4607 7021 4613
rect 6963 4573 6975 4607
rect 7009 4604 7021 4607
rect 7098 4604 7104 4616
rect 7009 4576 7104 4604
rect 7009 4573 7021 4576
rect 6963 4567 7021 4573
rect 7098 4564 7104 4576
rect 7156 4564 7162 4616
rect 7190 4564 7196 4616
rect 7248 4564 7254 4616
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4604 8723 4607
rect 8846 4604 8852 4616
rect 8711 4576 8852 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 8846 4564 8852 4576
rect 8904 4564 8910 4616
rect 9030 4613 9036 4616
rect 8992 4607 9036 4613
rect 8992 4573 9004 4607
rect 8992 4567 9036 4573
rect 9030 4564 9036 4567
rect 9088 4564 9094 4616
rect 9140 4613 9168 4644
rect 9398 4632 9404 4684
rect 9456 4632 9462 4684
rect 11149 4675 11207 4681
rect 11149 4641 11161 4675
rect 11195 4672 11207 4675
rect 11195 4644 12296 4672
rect 11195 4641 11207 4644
rect 11149 4635 11207 4641
rect 12158 4613 12164 4616
rect 9128 4607 9186 4613
rect 9128 4573 9140 4607
rect 9174 4573 9186 4607
rect 11609 4607 11667 4613
rect 11609 4604 11621 4607
rect 9128 4567 9186 4573
rect 11256 4576 11621 4604
rect 5084 4508 5396 4536
rect 3528 4468 3556 4496
rect 5084 4468 5112 4508
rect 3528 4440 5112 4468
rect 5810 4428 5816 4480
rect 5868 4468 5874 4480
rect 7282 4468 7288 4480
rect 5868 4440 7288 4468
rect 5868 4428 5874 4440
rect 7282 4428 7288 4440
rect 7340 4428 7346 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11256 4477 11284 4576
rect 11609 4573 11621 4576
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 12115 4607 12164 4613
rect 12115 4573 12127 4607
rect 12161 4573 12164 4607
rect 12115 4567 12164 4573
rect 12158 4564 12164 4567
rect 12216 4564 12222 4616
rect 12268 4604 12296 4644
rect 12342 4632 12348 4684
rect 12400 4632 12406 4684
rect 13725 4675 13783 4681
rect 13725 4641 13737 4675
rect 13771 4672 13783 4675
rect 13771 4644 14320 4672
rect 13771 4641 13783 4644
rect 13725 4635 13783 4641
rect 12526 4604 12532 4616
rect 12268 4576 12532 4604
rect 12526 4564 12532 4576
rect 12584 4604 12590 4616
rect 13814 4604 13820 4616
rect 12584 4576 13820 4604
rect 12584 4564 12590 4576
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 14292 4613 14320 4644
rect 14458 4632 14464 4684
rect 14516 4672 14522 4684
rect 14553 4675 14611 4681
rect 14553 4672 14565 4675
rect 14516 4644 14565 4672
rect 14516 4632 14522 4644
rect 14553 4641 14565 4644
rect 14599 4641 14611 4675
rect 14553 4635 14611 4641
rect 16853 4675 16911 4681
rect 16853 4641 16865 4675
rect 16899 4672 16911 4675
rect 17678 4672 17684 4684
rect 16899 4644 17684 4672
rect 16899 4641 16911 4644
rect 16853 4635 16911 4641
rect 17678 4632 17684 4644
rect 17736 4632 17742 4684
rect 17972 4672 18000 4768
rect 17972 4644 18736 4672
rect 14280 4607 14338 4613
rect 14280 4573 14292 4607
rect 14326 4573 14338 4607
rect 14280 4567 14338 4573
rect 16114 4564 16120 4616
rect 16172 4564 16178 4616
rect 16390 4564 16396 4616
rect 16448 4604 16454 4616
rect 16580 4607 16638 4613
rect 16580 4604 16592 4607
rect 16448 4576 16592 4604
rect 16448 4564 16454 4576
rect 16580 4573 16592 4576
rect 16626 4573 16638 4607
rect 16580 4567 16638 4573
rect 18325 4607 18383 4613
rect 18325 4573 18337 4607
rect 18371 4604 18383 4607
rect 18506 4604 18512 4616
rect 18371 4576 18512 4604
rect 18371 4573 18383 4576
rect 18325 4567 18383 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 18708 4604 18736 4644
rect 18874 4632 18880 4684
rect 18932 4672 18938 4684
rect 19061 4675 19119 4681
rect 19061 4672 19073 4675
rect 18932 4644 19073 4672
rect 18932 4632 18938 4644
rect 19061 4641 19073 4644
rect 19107 4641 19119 4675
rect 19061 4635 19119 4641
rect 18788 4607 18846 4613
rect 18788 4604 18800 4607
rect 18708 4576 18800 4604
rect 18788 4573 18800 4576
rect 18834 4573 18846 4607
rect 18788 4567 18846 4573
rect 11241 4471 11299 4477
rect 11241 4468 11253 4471
rect 11112 4440 11253 4468
rect 11112 4428 11118 4440
rect 11241 4437 11253 4440
rect 11287 4437 11299 4471
rect 11241 4431 11299 4437
rect 13446 4428 13452 4480
rect 13504 4468 13510 4480
rect 16132 4468 16160 4564
rect 13504 4440 16160 4468
rect 13504 4428 13510 4440
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 19720 4468 19748 4780
rect 27065 4777 27077 4780
rect 27111 4777 27123 4811
rect 27065 4771 27123 4777
rect 27890 4768 27896 4820
rect 27948 4808 27954 4820
rect 27991 4811 28049 4817
rect 27991 4808 28003 4811
rect 27948 4780 28003 4808
rect 27948 4768 27954 4780
rect 27991 4777 28003 4780
rect 28037 4808 28049 4811
rect 28350 4808 28356 4820
rect 28037 4780 28356 4808
rect 28037 4777 28049 4780
rect 27991 4771 28049 4777
rect 28350 4768 28356 4780
rect 28408 4768 28414 4820
rect 20530 4700 20536 4752
rect 20588 4740 20594 4752
rect 21634 4740 21640 4752
rect 20588 4712 21640 4740
rect 20588 4700 20594 4712
rect 21634 4700 21640 4712
rect 21692 4700 21698 4752
rect 26694 4700 26700 4752
rect 26752 4740 26758 4752
rect 26752 4712 26924 4740
rect 26752 4700 26758 4712
rect 19794 4632 19800 4684
rect 19852 4672 19858 4684
rect 20717 4675 20775 4681
rect 20717 4672 20729 4675
rect 19852 4644 20729 4672
rect 19852 4632 19858 4644
rect 20717 4641 20729 4644
rect 20763 4672 20775 4675
rect 20898 4672 20904 4684
rect 20763 4644 20904 4672
rect 20763 4641 20775 4644
rect 20717 4635 20775 4641
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 20993 4675 21051 4681
rect 20993 4641 21005 4675
rect 21039 4641 21051 4675
rect 20993 4635 21051 4641
rect 21008 4604 21036 4635
rect 21266 4632 21272 4684
rect 21324 4632 21330 4684
rect 21450 4632 21456 4684
rect 21508 4672 21514 4684
rect 21821 4675 21879 4681
rect 21821 4672 21833 4675
rect 21508 4644 21833 4672
rect 21508 4632 21514 4644
rect 21821 4641 21833 4644
rect 21867 4672 21879 4675
rect 21910 4672 21916 4684
rect 21867 4644 21916 4672
rect 21867 4641 21879 4644
rect 21821 4635 21879 4641
rect 21910 4632 21916 4644
rect 21968 4632 21974 4684
rect 22462 4632 22468 4684
rect 22520 4632 22526 4684
rect 22554 4632 22560 4684
rect 22612 4632 22618 4684
rect 23937 4675 23995 4681
rect 23937 4641 23949 4675
rect 23983 4672 23995 4675
rect 23983 4644 24532 4672
rect 23983 4641 23995 4644
rect 23937 4635 23995 4641
rect 22002 4604 22008 4616
rect 19812 4576 22008 4604
rect 19812 4548 19840 4576
rect 22002 4564 22008 4576
rect 22060 4564 22066 4616
rect 22186 4613 22192 4616
rect 22148 4607 22192 4613
rect 22148 4573 22160 4607
rect 22148 4567 22192 4573
rect 22186 4564 22192 4567
rect 22244 4564 22250 4616
rect 22327 4607 22385 4613
rect 22327 4573 22339 4607
rect 22373 4604 22385 4607
rect 22480 4604 22508 4632
rect 22373 4576 22508 4604
rect 22373 4573 22385 4576
rect 22327 4567 22385 4573
rect 24026 4564 24032 4616
rect 24084 4564 24090 4616
rect 24394 4613 24400 4616
rect 24356 4607 24400 4613
rect 24356 4573 24368 4607
rect 24356 4567 24400 4573
rect 24394 4564 24400 4567
rect 24452 4564 24458 4616
rect 24504 4615 24532 4644
rect 24578 4632 24584 4684
rect 24636 4672 24642 4684
rect 24765 4675 24823 4681
rect 24765 4672 24777 4675
rect 24636 4644 24777 4672
rect 24636 4632 24642 4644
rect 24765 4641 24777 4644
rect 24811 4641 24823 4675
rect 24765 4635 24823 4641
rect 24854 4632 24860 4684
rect 24912 4672 24918 4684
rect 26896 4681 26924 4712
rect 26789 4675 26847 4681
rect 26789 4672 26801 4675
rect 24912 4644 26801 4672
rect 24912 4632 24918 4644
rect 26789 4641 26801 4644
rect 26835 4641 26847 4675
rect 26789 4635 26847 4641
rect 26881 4675 26939 4681
rect 26881 4641 26893 4675
rect 26927 4641 26939 4675
rect 26881 4635 26939 4641
rect 24492 4609 24550 4615
rect 24492 4575 24504 4609
rect 24538 4575 24550 4609
rect 24492 4569 24550 4575
rect 25406 4564 25412 4616
rect 25464 4604 25470 4616
rect 26804 4604 26832 4635
rect 27522 4632 27528 4684
rect 27580 4672 27586 4684
rect 27890 4672 27896 4684
rect 27580 4644 27896 4672
rect 27580 4632 27586 4644
rect 27890 4632 27896 4644
rect 27948 4632 27954 4684
rect 28994 4672 29000 4684
rect 28184 4644 29000 4672
rect 27430 4604 27436 4616
rect 25464 4576 26740 4604
rect 26804 4576 27436 4604
rect 25464 4564 25470 4576
rect 19794 4496 19800 4548
rect 19852 4496 19858 4548
rect 20533 4539 20591 4545
rect 20533 4505 20545 4539
rect 20579 4536 20591 4539
rect 20579 4508 21864 4536
rect 20579 4505 20591 4508
rect 20533 4499 20591 4505
rect 21836 4480 21864 4508
rect 25424 4508 26648 4536
rect 17920 4440 19748 4468
rect 17920 4428 17926 4440
rect 20346 4428 20352 4480
rect 20404 4428 20410 4480
rect 20809 4471 20867 4477
rect 20809 4437 20821 4471
rect 20855 4468 20867 4471
rect 21266 4468 21272 4480
rect 20855 4440 21272 4468
rect 20855 4437 20867 4440
rect 20809 4431 20867 4437
rect 21266 4428 21272 4440
rect 21324 4428 21330 4480
rect 21358 4428 21364 4480
rect 21416 4468 21422 4480
rect 21453 4471 21511 4477
rect 21453 4468 21465 4471
rect 21416 4440 21465 4468
rect 21416 4428 21422 4440
rect 21453 4437 21465 4440
rect 21499 4437 21511 4471
rect 21453 4431 21511 4437
rect 21818 4428 21824 4480
rect 21876 4428 21882 4480
rect 22278 4428 22284 4480
rect 22336 4468 22342 4480
rect 25424 4468 25452 4508
rect 22336 4440 25452 4468
rect 22336 4428 22342 4440
rect 26050 4428 26056 4480
rect 26108 4428 26114 4480
rect 26620 4477 26648 4508
rect 26605 4471 26663 4477
rect 26605 4437 26617 4471
rect 26651 4437 26663 4471
rect 26712 4468 26740 4576
rect 27430 4564 27436 4576
rect 27488 4604 27494 4616
rect 27798 4604 27804 4616
rect 27488 4576 27804 4604
rect 27488 4564 27494 4576
rect 27798 4564 27804 4576
rect 27856 4564 27862 4616
rect 28031 4607 28089 4613
rect 28031 4573 28043 4607
rect 28077 4604 28089 4607
rect 28184 4604 28212 4644
rect 28994 4632 29000 4644
rect 29052 4632 29058 4684
rect 28077 4576 28212 4604
rect 28077 4573 28089 4576
rect 28031 4567 28089 4573
rect 28258 4564 28264 4616
rect 28316 4564 28322 4616
rect 29365 4539 29423 4545
rect 29365 4505 29377 4539
rect 29411 4505 29423 4539
rect 29365 4499 29423 4505
rect 29380 4468 29408 4499
rect 26712 4440 29408 4468
rect 26605 4431 26663 4437
rect 552 4378 30912 4400
rect 552 4326 4193 4378
rect 4245 4326 4257 4378
rect 4309 4326 4321 4378
rect 4373 4326 4385 4378
rect 4437 4326 4449 4378
rect 4501 4326 11783 4378
rect 11835 4326 11847 4378
rect 11899 4326 11911 4378
rect 11963 4326 11975 4378
rect 12027 4326 12039 4378
rect 12091 4326 19373 4378
rect 19425 4326 19437 4378
rect 19489 4326 19501 4378
rect 19553 4326 19565 4378
rect 19617 4326 19629 4378
rect 19681 4326 26963 4378
rect 27015 4326 27027 4378
rect 27079 4326 27091 4378
rect 27143 4326 27155 4378
rect 27207 4326 27219 4378
rect 27271 4326 30912 4378
rect 552 4304 30912 4326
rect 5626 4264 5632 4276
rect 3160 4236 5632 4264
rect 937 4131 995 4137
rect 937 4097 949 4131
rect 983 4128 995 4131
rect 1302 4128 1308 4140
rect 983 4100 1308 4128
rect 983 4097 995 4100
rect 937 4091 995 4097
rect 1302 4088 1308 4100
rect 1360 4088 1366 4140
rect 1486 4137 1492 4140
rect 1443 4131 1492 4137
rect 1443 4097 1455 4131
rect 1489 4097 1492 4131
rect 1443 4091 1492 4097
rect 1486 4088 1492 4091
rect 1544 4088 1550 4140
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 2682 4128 2688 4140
rect 1719 4100 2688 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 1026 4020 1032 4072
rect 1084 4060 1090 4072
rect 3160 4060 3188 4236
rect 5626 4224 5632 4236
rect 5684 4224 5690 4276
rect 6822 4264 6828 4276
rect 5920 4236 6828 4264
rect 5350 4156 5356 4208
rect 5408 4196 5414 4208
rect 5920 4196 5948 4236
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 8754 4224 8760 4276
rect 8812 4264 8818 4276
rect 11885 4267 11943 4273
rect 8812 4236 11284 4264
rect 8812 4224 8818 4236
rect 9398 4196 9404 4208
rect 5408 4168 5948 4196
rect 8864 4168 9404 4196
rect 5408 4156 5414 4168
rect 8864 4140 8892 4168
rect 9398 4156 9404 4168
rect 9456 4156 9462 4208
rect 11256 4196 11284 4236
rect 11885 4233 11897 4267
rect 11931 4264 11943 4267
rect 12158 4264 12164 4276
rect 11931 4236 12164 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 12526 4224 12532 4276
rect 12584 4224 12590 4276
rect 14550 4264 14556 4276
rect 13832 4236 14556 4264
rect 13832 4196 13860 4236
rect 14550 4224 14556 4236
rect 14608 4224 14614 4276
rect 17494 4224 17500 4276
rect 17552 4264 17558 4276
rect 17552 4236 18460 4264
rect 17552 4224 17558 4236
rect 11256 4168 13860 4196
rect 18432 4196 18460 4236
rect 18506 4224 18512 4276
rect 18564 4264 18570 4276
rect 18969 4267 19027 4273
rect 18969 4264 18981 4267
rect 18564 4236 18981 4264
rect 18564 4224 18570 4236
rect 18969 4233 18981 4236
rect 19015 4233 19027 4267
rect 21542 4264 21548 4276
rect 18969 4227 19027 4233
rect 19904 4236 21548 4264
rect 19904 4196 19932 4236
rect 21542 4224 21548 4236
rect 21600 4224 21606 4276
rect 21634 4224 21640 4276
rect 21692 4264 21698 4276
rect 23566 4264 23572 4276
rect 21692 4236 23572 4264
rect 21692 4224 21698 4236
rect 23566 4224 23572 4236
rect 23624 4224 23630 4276
rect 24210 4264 24216 4276
rect 23998 4236 24216 4264
rect 18432 4168 19932 4196
rect 22186 4156 22192 4208
rect 22244 4196 22250 4208
rect 22244 4168 22600 4196
rect 22244 4156 22250 4168
rect 3234 4088 3240 4140
rect 3292 4088 3298 4140
rect 3326 4088 3332 4140
rect 3384 4128 3390 4140
rect 3976 4131 4034 4137
rect 3976 4128 3988 4131
rect 3384 4100 3988 4128
rect 3384 4088 3390 4100
rect 3976 4097 3988 4100
rect 4022 4097 4034 4131
rect 3976 4091 4034 4097
rect 4982 4088 4988 4140
rect 5040 4088 5046 4140
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 6368 4131 6426 4137
rect 6368 4128 6380 4131
rect 5592 4100 6380 4128
rect 5592 4088 5598 4100
rect 6368 4097 6380 4100
rect 6414 4097 6426 4131
rect 6368 4091 6426 4097
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4128 8079 4131
rect 8386 4128 8392 4140
rect 8067 4100 8392 4128
rect 8067 4097 8079 4100
rect 8021 4091 8079 4097
rect 8386 4088 8392 4100
rect 8444 4088 8450 4140
rect 8846 4088 8852 4140
rect 8904 4088 8910 4140
rect 9493 4131 9551 4137
rect 9493 4128 9505 4131
rect 9048 4100 9505 4128
rect 1084 4032 3188 4060
rect 1084 4020 1090 4032
rect 3252 3992 3280 4088
rect 3418 4020 3424 4072
rect 3476 4020 3482 4072
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4029 3571 4063
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 3513 4023 3571 4029
rect 3620 4032 4261 4060
rect 3528 3992 3556 4023
rect 3252 3964 3556 3992
rect 1403 3927 1461 3933
rect 1403 3893 1415 3927
rect 1449 3924 1461 3927
rect 1762 3924 1768 3936
rect 1449 3896 1768 3924
rect 1449 3893 1461 3896
rect 1403 3887 1461 3893
rect 1762 3884 1768 3896
rect 1820 3884 1826 3936
rect 2774 3884 2780 3936
rect 2832 3884 2838 3936
rect 3237 3927 3295 3933
rect 3237 3893 3249 3927
rect 3283 3924 3295 3927
rect 3620 3924 3648 4032
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 5000 3992 5028 4088
rect 9048 4072 9076 4100
rect 9493 4097 9505 4100
rect 9539 4128 9551 4131
rect 9539 4100 9996 4128
rect 9539 4097 9551 4100
rect 9493 4091 9551 4097
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 5905 4063 5963 4069
rect 5905 4060 5917 4063
rect 5868 4032 5917 4060
rect 5868 4020 5874 4032
rect 5905 4029 5917 4032
rect 5951 4029 5963 4063
rect 6641 4063 6699 4069
rect 6641 4060 6653 4063
rect 5905 4023 5963 4029
rect 6012 4032 6653 4060
rect 6012 3992 6040 4032
rect 6641 4029 6653 4032
rect 6687 4029 6699 4063
rect 6641 4023 6699 4029
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 8573 4063 8631 4069
rect 8573 4060 8585 4063
rect 7708 4032 8585 4060
rect 7708 4020 7714 4032
rect 8573 4029 8585 4032
rect 8619 4029 8631 4063
rect 8941 4063 8999 4069
rect 8941 4060 8953 4063
rect 8573 4023 8631 4029
rect 8680 4032 8953 4060
rect 5000 3964 6040 3992
rect 8478 3952 8484 4004
rect 8536 3992 8542 4004
rect 8680 3992 8708 4032
rect 8941 4029 8953 4032
rect 8987 4029 8999 4063
rect 8941 4023 8999 4029
rect 9030 4020 9036 4072
rect 9088 4020 9094 4072
rect 9214 4020 9220 4072
rect 9272 4020 9278 4072
rect 9306 4020 9312 4072
rect 9364 4020 9370 4072
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9861 4063 9919 4069
rect 9861 4060 9873 4063
rect 9456 4032 9873 4060
rect 9456 4020 9462 4032
rect 9861 4029 9873 4032
rect 9907 4029 9919 4063
rect 9968 4060 9996 4100
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10324 4131 10382 4137
rect 10324 4128 10336 4131
rect 10100 4100 10336 4128
rect 10100 4088 10106 4100
rect 10324 4097 10336 4100
rect 10370 4097 10382 4131
rect 10324 4091 10382 4097
rect 10502 4088 10508 4140
rect 10560 4128 10566 4140
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 10560 4100 10609 4128
rect 10560 4088 10566 4100
rect 10597 4097 10609 4100
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 13173 4131 13231 4137
rect 11296 4100 12296 4128
rect 11296 4088 11302 4100
rect 12268 4069 12296 4100
rect 13173 4097 13185 4131
rect 13219 4128 13231 4131
rect 13998 4128 14004 4140
rect 13219 4100 14004 4128
rect 13219 4097 13231 4100
rect 13173 4091 13231 4097
rect 13998 4088 14004 4100
rect 14056 4128 14062 4140
rect 14182 4137 14188 4140
rect 14144 4131 14188 4137
rect 14144 4128 14156 4131
rect 14056 4100 14156 4128
rect 14056 4088 14062 4100
rect 14144 4097 14156 4100
rect 14144 4091 14188 4097
rect 14182 4088 14188 4091
rect 14240 4088 14246 4140
rect 14280 4129 14338 4135
rect 14280 4095 14292 4129
rect 14326 4095 14338 4129
rect 14280 4089 14338 4095
rect 10188 4063 10246 4069
rect 10188 4060 10200 4063
rect 9968 4032 10200 4060
rect 9861 4023 9919 4029
rect 10188 4029 10200 4032
rect 10234 4029 10246 4063
rect 10188 4023 10246 4029
rect 12253 4063 12311 4069
rect 12253 4029 12265 4063
rect 12299 4029 12311 4063
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12253 4023 12311 4029
rect 12360 4032 12909 4060
rect 12360 3992 12388 4032
rect 12897 4029 12909 4032
rect 12943 4060 12955 4063
rect 12943 4032 13584 4060
rect 12943 4029 12955 4032
rect 12897 4023 12955 4029
rect 8536 3964 8708 3992
rect 8772 3964 9536 3992
rect 8536 3952 8542 3964
rect 3283 3896 3648 3924
rect 3283 3893 3295 3896
rect 3237 3887 3295 3893
rect 3970 3884 3976 3936
rect 4028 3933 4034 3936
rect 4028 3924 4037 3933
rect 4028 3896 4073 3924
rect 4028 3887 4037 3896
rect 4028 3884 4034 3887
rect 5534 3884 5540 3936
rect 5592 3884 5598 3936
rect 5994 3884 6000 3936
rect 6052 3924 6058 3936
rect 6371 3927 6429 3933
rect 6371 3924 6383 3927
rect 6052 3896 6383 3924
rect 6052 3884 6058 3896
rect 6371 3893 6383 3896
rect 6417 3893 6429 3927
rect 6371 3887 6429 3893
rect 8389 3927 8447 3933
rect 8389 3893 8401 3927
rect 8435 3924 8447 3927
rect 8570 3924 8576 3936
rect 8435 3896 8576 3924
rect 8435 3893 8447 3896
rect 8389 3887 8447 3893
rect 8570 3884 8576 3896
rect 8628 3884 8634 3936
rect 8772 3933 8800 3964
rect 8757 3927 8815 3933
rect 8757 3893 8769 3927
rect 8803 3893 8815 3927
rect 8757 3887 8815 3893
rect 9033 3927 9091 3933
rect 9033 3893 9045 3927
rect 9079 3924 9091 3927
rect 9306 3924 9312 3936
rect 9079 3896 9312 3924
rect 9079 3893 9091 3896
rect 9033 3887 9091 3893
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 9508 3924 9536 3964
rect 11256 3964 12388 3992
rect 12437 3995 12495 4001
rect 9674 3924 9680 3936
rect 9508 3896 9680 3924
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 9858 3884 9864 3936
rect 9916 3924 9922 3936
rect 11256 3924 11284 3964
rect 12437 3961 12449 3995
rect 12483 3992 12495 3995
rect 13446 3992 13452 4004
rect 12483 3964 13452 3992
rect 12483 3961 12495 3964
rect 12437 3955 12495 3961
rect 13446 3952 13452 3964
rect 13504 3952 13510 4004
rect 13556 3992 13584 4032
rect 13630 4020 13636 4072
rect 13688 4060 13694 4072
rect 13725 4063 13783 4069
rect 13725 4060 13737 4063
rect 13688 4032 13737 4060
rect 13688 4020 13694 4032
rect 13725 4029 13737 4032
rect 13771 4029 13783 4063
rect 13725 4023 13783 4029
rect 13814 4020 13820 4072
rect 13872 4020 13878 4072
rect 14295 4060 14323 4089
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 16942 4135 16948 4140
rect 16899 4129 16948 4135
rect 14516 4100 16804 4128
rect 14516 4088 14522 4100
rect 13924 4032 14323 4060
rect 13924 4004 13952 4032
rect 14366 4020 14372 4072
rect 14424 4060 14430 4072
rect 14553 4063 14611 4069
rect 14553 4060 14565 4063
rect 14424 4032 14565 4060
rect 14424 4020 14430 4032
rect 14553 4029 14565 4032
rect 14599 4029 14611 4063
rect 14553 4023 14611 4029
rect 14642 4020 14648 4072
rect 14700 4060 14706 4072
rect 16206 4060 16212 4072
rect 14700 4032 16212 4060
rect 14700 4020 14706 4032
rect 16206 4020 16212 4032
rect 16264 4060 16270 4072
rect 16301 4063 16359 4069
rect 16301 4060 16313 4063
rect 16264 4032 16313 4060
rect 16264 4020 16270 4032
rect 16301 4029 16313 4032
rect 16347 4029 16359 4063
rect 16301 4023 16359 4029
rect 16390 4020 16396 4072
rect 16448 4020 16454 4072
rect 16776 4060 16804 4100
rect 16899 4095 16911 4129
rect 16945 4095 16948 4129
rect 16899 4089 16948 4095
rect 16942 4088 16948 4089
rect 17000 4088 17006 4140
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 17862 4128 17868 4140
rect 17175 4100 17868 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 19306 4100 19748 4128
rect 19306 4060 19334 4100
rect 16776 4032 19334 4060
rect 19521 4063 19579 4069
rect 19521 4029 19533 4063
rect 19567 4060 19579 4063
rect 19610 4060 19616 4072
rect 19567 4032 19616 4060
rect 19567 4029 19579 4032
rect 19521 4023 19579 4029
rect 19610 4020 19616 4032
rect 19668 4020 19674 4072
rect 19720 4060 19748 4100
rect 20346 4088 20352 4140
rect 20404 4128 20410 4140
rect 20625 4131 20683 4137
rect 20404 4100 20449 4128
rect 20404 4088 20410 4100
rect 20625 4097 20637 4131
rect 20671 4128 20683 4131
rect 20806 4128 20812 4140
rect 20671 4100 20812 4128
rect 20671 4097 20683 4100
rect 20625 4091 20683 4097
rect 20806 4088 20812 4100
rect 20864 4088 20870 4140
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4128 22063 4131
rect 22370 4128 22376 4140
rect 22051 4100 22376 4128
rect 22051 4097 22063 4100
rect 22005 4091 22063 4097
rect 22370 4088 22376 4100
rect 22428 4088 22434 4140
rect 22572 4137 22600 4168
rect 22830 4156 22836 4208
rect 22888 4196 22894 4208
rect 22888 4168 23152 4196
rect 22888 4156 22894 4168
rect 22557 4131 22615 4137
rect 22557 4097 22569 4131
rect 22603 4128 22615 4131
rect 22603 4100 22968 4128
rect 22603 4097 22615 4100
rect 22557 4091 22615 4097
rect 22940 4072 22968 4100
rect 19794 4069 19800 4072
rect 19789 4060 19800 4069
rect 19720 4032 19800 4060
rect 19789 4023 19800 4032
rect 19794 4020 19800 4023
rect 19852 4020 19858 4072
rect 19889 4063 19947 4069
rect 19889 4029 19901 4063
rect 19935 4060 19947 4063
rect 19978 4060 19984 4072
rect 19935 4032 19984 4060
rect 19935 4029 19947 4032
rect 19889 4023 19947 4029
rect 13556 3964 13676 3992
rect 9916 3896 11284 3924
rect 9916 3884 9922 3896
rect 12066 3884 12072 3936
rect 12124 3884 12130 3936
rect 13538 3884 13544 3936
rect 13596 3884 13602 3936
rect 13648 3924 13676 3964
rect 13906 3952 13912 4004
rect 13964 3952 13970 4004
rect 18877 3995 18935 4001
rect 18877 3961 18889 3995
rect 18923 3992 18935 3995
rect 19904 3992 19932 4023
rect 19978 4020 19984 4032
rect 20036 4020 20042 4072
rect 22281 4063 22339 4069
rect 22281 4029 22293 4063
rect 22327 4060 22339 4063
rect 22646 4060 22652 4072
rect 22327 4032 22652 4060
rect 22327 4029 22339 4032
rect 22281 4023 22339 4029
rect 22646 4020 22652 4032
rect 22704 4020 22710 4072
rect 22922 4020 22928 4072
rect 22980 4020 22986 4072
rect 23017 4063 23075 4069
rect 23017 4029 23029 4063
rect 23063 4060 23075 4063
rect 23124 4060 23152 4168
rect 23998 4137 24026 4236
rect 24210 4224 24216 4236
rect 24268 4224 24274 4276
rect 23998 4131 24077 4137
rect 23998 4100 24031 4131
rect 24019 4097 24031 4100
rect 24065 4097 24077 4131
rect 24019 4091 24077 4097
rect 24535 4131 24593 4137
rect 24535 4097 24547 4131
rect 24581 4128 24593 4131
rect 24670 4128 24676 4140
rect 24581 4100 24676 4128
rect 24581 4097 24593 4100
rect 24535 4091 24593 4097
rect 24670 4088 24676 4100
rect 24728 4088 24734 4140
rect 24762 4088 24768 4140
rect 24820 4088 24826 4140
rect 26050 4088 26056 4140
rect 26108 4128 26114 4140
rect 26700 4131 26758 4137
rect 26700 4128 26712 4131
rect 26108 4100 26712 4128
rect 26108 4088 26114 4100
rect 26700 4097 26712 4100
rect 26746 4097 26758 4131
rect 26700 4091 26758 4097
rect 26786 4088 26792 4140
rect 26844 4128 26850 4140
rect 26973 4131 27031 4137
rect 26973 4128 26985 4131
rect 26844 4100 26985 4128
rect 26844 4088 26850 4100
rect 26973 4097 26985 4100
rect 27019 4097 27031 4131
rect 26973 4091 27031 4097
rect 23063 4032 23152 4060
rect 23293 4063 23351 4069
rect 23063 4029 23075 4032
rect 23017 4023 23075 4029
rect 23293 4029 23305 4063
rect 23339 4060 23351 4063
rect 23661 4063 23719 4069
rect 23661 4060 23673 4063
rect 23339 4032 23673 4060
rect 23339 4029 23351 4032
rect 23293 4023 23351 4029
rect 23661 4029 23673 4032
rect 23707 4060 23719 4063
rect 25222 4060 25228 4072
rect 23707 4032 25228 4060
rect 23707 4029 23719 4032
rect 23661 4023 23719 4029
rect 25222 4020 25228 4032
rect 25280 4020 25286 4072
rect 26234 4060 26240 4072
rect 25424 4032 26240 4060
rect 18923 3964 19932 3992
rect 23124 3964 24164 3992
rect 18923 3961 18935 3964
rect 18877 3955 18935 3961
rect 14274 3924 14280 3936
rect 13648 3896 14280 3924
rect 14274 3884 14280 3896
rect 14332 3884 14338 3936
rect 15841 3927 15899 3933
rect 15841 3893 15853 3927
rect 15887 3924 15899 3927
rect 16022 3924 16028 3936
rect 15887 3896 16028 3924
rect 15887 3893 15899 3896
rect 15841 3887 15899 3893
rect 16022 3884 16028 3896
rect 16080 3884 16086 3936
rect 16117 3927 16175 3933
rect 16117 3893 16129 3927
rect 16163 3924 16175 3927
rect 16666 3924 16672 3936
rect 16163 3896 16672 3924
rect 16163 3893 16175 3896
rect 16117 3887 16175 3893
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 16859 3927 16917 3933
rect 16859 3893 16871 3927
rect 16905 3924 16917 3927
rect 17034 3924 17040 3936
rect 16905 3896 17040 3924
rect 16905 3893 16917 3896
rect 16859 3887 16917 3893
rect 17034 3884 17040 3896
rect 17092 3884 17098 3936
rect 17218 3884 17224 3936
rect 17276 3924 17282 3936
rect 18233 3927 18291 3933
rect 18233 3924 18245 3927
rect 17276 3896 18245 3924
rect 17276 3884 17282 3896
rect 18233 3893 18245 3896
rect 18279 3893 18291 3927
rect 18233 3887 18291 3893
rect 19334 3884 19340 3936
rect 19392 3884 19398 3936
rect 19613 3927 19671 3933
rect 19613 3893 19625 3927
rect 19659 3924 19671 3927
rect 19702 3924 19708 3936
rect 19659 3896 19708 3924
rect 19659 3893 19671 3896
rect 19613 3887 19671 3893
rect 19702 3884 19708 3896
rect 19760 3884 19766 3936
rect 20355 3927 20413 3933
rect 20355 3893 20367 3927
rect 20401 3924 20413 3927
rect 20990 3924 20996 3936
rect 20401 3896 20996 3924
rect 20401 3893 20413 3896
rect 20355 3887 20413 3893
rect 20990 3884 20996 3896
rect 21048 3884 21054 3936
rect 22830 3884 22836 3936
rect 22888 3884 22894 3936
rect 23124 3933 23152 3964
rect 23109 3927 23167 3933
rect 23109 3893 23121 3927
rect 23155 3893 23167 3927
rect 23109 3887 23167 3893
rect 23477 3927 23535 3933
rect 23477 3893 23489 3927
rect 23523 3924 23535 3927
rect 24026 3924 24032 3936
rect 23523 3896 24032 3924
rect 23523 3893 23535 3896
rect 23477 3887 23535 3893
rect 24026 3884 24032 3896
rect 24084 3884 24090 3936
rect 24136 3924 24164 3964
rect 24394 3924 24400 3936
rect 24136 3896 24400 3924
rect 24394 3884 24400 3896
rect 24452 3884 24458 3936
rect 24486 3884 24492 3936
rect 24544 3933 24550 3936
rect 24544 3924 24553 3933
rect 24544 3896 24589 3924
rect 24544 3887 24553 3896
rect 24544 3884 24550 3887
rect 25130 3884 25136 3936
rect 25188 3924 25194 3936
rect 25424 3924 25452 4032
rect 26234 4020 26240 4032
rect 26292 4020 26298 4072
rect 25188 3896 25452 3924
rect 25188 3884 25194 3896
rect 26050 3884 26056 3936
rect 26108 3884 26114 3936
rect 26694 3884 26700 3936
rect 26752 3933 26758 3936
rect 26752 3887 26761 3933
rect 26752 3884 26758 3887
rect 28074 3884 28080 3936
rect 28132 3884 28138 3936
rect 552 3834 31072 3856
rect 552 3782 7988 3834
rect 8040 3782 8052 3834
rect 8104 3782 8116 3834
rect 8168 3782 8180 3834
rect 8232 3782 8244 3834
rect 8296 3782 15578 3834
rect 15630 3782 15642 3834
rect 15694 3782 15706 3834
rect 15758 3782 15770 3834
rect 15822 3782 15834 3834
rect 15886 3782 23168 3834
rect 23220 3782 23232 3834
rect 23284 3782 23296 3834
rect 23348 3782 23360 3834
rect 23412 3782 23424 3834
rect 23476 3782 30758 3834
rect 30810 3782 30822 3834
rect 30874 3782 30886 3834
rect 30938 3782 30950 3834
rect 31002 3782 31014 3834
rect 31066 3782 31072 3834
rect 552 3760 31072 3782
rect 750 3680 756 3732
rect 808 3720 814 3732
rect 1029 3723 1087 3729
rect 1029 3720 1041 3723
rect 808 3692 1041 3720
rect 808 3680 814 3692
rect 1029 3689 1041 3692
rect 1075 3689 1087 3723
rect 1029 3683 1087 3689
rect 1305 3723 1363 3729
rect 1305 3689 1317 3723
rect 1351 3720 1363 3723
rect 4522 3720 4528 3732
rect 1351 3692 2084 3720
rect 1351 3689 1363 3692
rect 1305 3683 1363 3689
rect 1118 3612 1124 3664
rect 1176 3652 1182 3664
rect 2056 3652 2084 3692
rect 2746 3692 4528 3720
rect 2746 3652 2774 3692
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 6546 3720 6552 3732
rect 5592 3692 6552 3720
rect 5592 3680 5598 3692
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7745 3723 7803 3729
rect 7745 3720 7757 3723
rect 7156 3692 7757 3720
rect 7156 3680 7162 3692
rect 7745 3689 7757 3692
rect 7791 3689 7803 3723
rect 7745 3683 7803 3689
rect 9214 3680 9220 3732
rect 9272 3720 9278 3732
rect 10502 3720 10508 3732
rect 9272 3692 10508 3720
rect 9272 3680 9278 3692
rect 10502 3680 10508 3692
rect 10560 3720 10566 3732
rect 10962 3720 10968 3732
rect 10560 3692 10968 3720
rect 10560 3680 10566 3692
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 12066 3680 12072 3732
rect 12124 3720 12130 3732
rect 12124 3692 13492 3720
rect 12124 3680 12130 3692
rect 1176 3624 1808 3652
rect 2056 3624 2774 3652
rect 2869 3655 2927 3661
rect 1176 3612 1182 3624
rect 1210 3544 1216 3596
rect 1268 3544 1274 3596
rect 1780 3593 1808 3624
rect 2869 3621 2881 3655
rect 2915 3652 2927 3655
rect 3234 3652 3240 3664
rect 2915 3624 3240 3652
rect 2915 3621 2927 3624
rect 2869 3615 2927 3621
rect 3234 3612 3240 3624
rect 3292 3612 3298 3664
rect 3602 3612 3608 3664
rect 3660 3612 3666 3664
rect 5994 3612 6000 3664
rect 6052 3612 6058 3664
rect 10781 3655 10839 3661
rect 10781 3621 10793 3655
rect 10827 3652 10839 3655
rect 10827 3624 11750 3652
rect 10827 3621 10839 3624
rect 10781 3615 10839 3621
rect 1489 3587 1547 3593
rect 1489 3553 1501 3587
rect 1535 3553 1547 3587
rect 1489 3547 1547 3553
rect 1765 3587 1823 3593
rect 1765 3553 1777 3587
rect 1811 3553 1823 3587
rect 1765 3547 1823 3553
rect 2501 3587 2559 3593
rect 2501 3553 2513 3587
rect 2547 3584 2559 3587
rect 3620 3584 3648 3612
rect 2547 3556 3648 3584
rect 3896 3556 4200 3584
rect 2547 3553 2559 3556
rect 2501 3547 2559 3553
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 1504 3516 1532 3547
rect 3896 3525 3924 3556
rect 992 3488 1532 3516
rect 3237 3519 3295 3525
rect 992 3476 998 3488
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3513 3519 3571 3525
rect 3513 3516 3525 3519
rect 3283 3488 3525 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 3513 3485 3525 3488
rect 3559 3485 3571 3519
rect 3513 3479 3571 3485
rect 3840 3519 3924 3525
rect 3840 3485 3852 3519
rect 3886 3488 3924 3519
rect 3886 3485 3898 3488
rect 3840 3479 3898 3485
rect 1581 3451 1639 3457
rect 1581 3417 1593 3451
rect 1627 3448 1639 3451
rect 1670 3448 1676 3460
rect 1627 3420 1676 3448
rect 1627 3417 1639 3420
rect 1581 3411 1639 3417
rect 1670 3408 1676 3420
rect 1728 3408 1734 3460
rect 3528 3380 3556 3479
rect 3970 3476 3976 3528
rect 4028 3476 4034 3528
rect 4172 3516 4200 3556
rect 4246 3544 4252 3596
rect 4304 3544 4310 3596
rect 6012 3584 6040 3612
rect 6178 3584 6184 3596
rect 6012 3556 6184 3584
rect 6178 3544 6184 3556
rect 6236 3593 6242 3596
rect 6236 3587 6290 3593
rect 6236 3553 6244 3587
rect 6278 3553 6290 3587
rect 6236 3547 6290 3553
rect 6236 3544 6242 3547
rect 6546 3544 6552 3596
rect 6604 3544 6610 3596
rect 6638 3544 6644 3596
rect 6696 3544 6702 3596
rect 7098 3544 7104 3596
rect 7156 3584 7162 3596
rect 7282 3584 7288 3596
rect 7156 3556 7288 3584
rect 7156 3544 7162 3556
rect 7282 3544 7288 3556
rect 7340 3584 7346 3596
rect 8110 3584 8116 3596
rect 7340 3556 8116 3584
rect 7340 3544 7346 3556
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 9306 3544 9312 3596
rect 9364 3584 9370 3596
rect 9401 3587 9459 3593
rect 9401 3584 9413 3587
rect 9364 3556 9413 3584
rect 9364 3544 9370 3556
rect 9401 3553 9413 3556
rect 9447 3553 9459 3587
rect 9401 3547 9459 3553
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 11057 3587 11115 3593
rect 11057 3584 11069 3587
rect 9548 3556 11069 3584
rect 9548 3544 9554 3556
rect 11057 3553 11069 3556
rect 11103 3553 11115 3587
rect 11722 3584 11750 3624
rect 13464 3584 13492 3692
rect 14182 3680 14188 3732
rect 14240 3720 14246 3732
rect 14283 3723 14341 3729
rect 14283 3720 14295 3723
rect 14240 3692 14295 3720
rect 14240 3680 14246 3692
rect 14283 3689 14295 3692
rect 14329 3689 14341 3723
rect 14283 3683 14341 3689
rect 16206 3680 16212 3732
rect 16264 3720 16270 3732
rect 16482 3720 16488 3732
rect 16264 3692 16488 3720
rect 16264 3680 16270 3692
rect 16482 3680 16488 3692
rect 16540 3680 16546 3732
rect 16574 3680 16580 3732
rect 16632 3729 16638 3732
rect 16632 3720 16641 3729
rect 18791 3723 18849 3729
rect 16632 3692 16677 3720
rect 16632 3683 16641 3692
rect 18791 3689 18803 3723
rect 18837 3720 18849 3723
rect 18966 3720 18972 3732
rect 18837 3692 18972 3720
rect 18837 3689 18849 3692
rect 18791 3683 18849 3689
rect 16632 3680 16638 3683
rect 18966 3680 18972 3692
rect 19024 3680 19030 3732
rect 20990 3680 20996 3732
rect 21048 3720 21054 3732
rect 21542 3720 21548 3732
rect 21048 3692 21548 3720
rect 21048 3680 21054 3692
rect 21542 3680 21548 3692
rect 21600 3720 21606 3732
rect 21735 3723 21793 3729
rect 21735 3720 21747 3723
rect 21600 3692 21747 3720
rect 21600 3680 21606 3692
rect 21735 3689 21747 3692
rect 21781 3689 21793 3723
rect 21735 3683 21793 3689
rect 22830 3680 22836 3732
rect 22888 3680 22894 3732
rect 22922 3680 22928 3732
rect 22980 3720 22986 3732
rect 23943 3723 24001 3729
rect 23943 3720 23955 3723
rect 22980 3692 23955 3720
rect 22980 3680 22986 3692
rect 23943 3689 23955 3692
rect 23989 3720 24001 3723
rect 24118 3720 24124 3732
rect 23989 3692 24124 3720
rect 23989 3689 24001 3692
rect 23943 3683 24001 3689
rect 24118 3680 24124 3692
rect 24176 3680 24182 3732
rect 24578 3680 24584 3732
rect 24636 3720 24642 3732
rect 26510 3720 26516 3732
rect 24636 3692 26516 3720
rect 24636 3680 24642 3692
rect 26510 3680 26516 3692
rect 26568 3720 26574 3732
rect 26568 3692 26648 3720
rect 26568 3680 26574 3692
rect 13725 3655 13783 3661
rect 13725 3621 13737 3655
rect 13771 3652 13783 3655
rect 13906 3652 13912 3664
rect 13771 3624 13912 3652
rect 13771 3621 13783 3624
rect 13725 3615 13783 3621
rect 13906 3612 13912 3624
rect 13964 3612 13970 3664
rect 20441 3655 20499 3661
rect 20441 3621 20453 3655
rect 20487 3652 20499 3655
rect 22848 3652 22876 3680
rect 20487 3624 21404 3652
rect 22848 3624 23612 3652
rect 20487 3621 20499 3624
rect 20441 3615 20499 3621
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 11722 3556 12115 3584
rect 13464 3556 14565 3584
rect 11057 3547 11115 3553
rect 4172 3488 5580 3516
rect 5442 3380 5448 3392
rect 3528 3352 5448 3380
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 5552 3380 5580 3488
rect 5626 3476 5632 3528
rect 5684 3476 5690 3528
rect 5810 3476 5816 3528
rect 5868 3516 5874 3528
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 5868 3488 5917 3516
rect 5868 3476 5874 3488
rect 5905 3485 5917 3488
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 6411 3519 6469 3525
rect 6411 3485 6423 3519
rect 6457 3516 6469 3519
rect 6564 3516 6592 3544
rect 6457 3488 6592 3516
rect 6457 3485 6469 3488
rect 6411 3479 6469 3485
rect 8386 3476 8392 3528
rect 8444 3476 8450 3528
rect 8665 3519 8723 3525
rect 8665 3485 8677 3519
rect 8711 3516 8723 3519
rect 8846 3516 8852 3528
rect 8711 3488 8852 3516
rect 8711 3485 8723 3488
rect 8665 3479 8723 3485
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 9030 3525 9036 3528
rect 8992 3519 9036 3525
rect 8992 3485 9004 3519
rect 8992 3479 9036 3485
rect 9030 3476 9036 3479
rect 9088 3476 9094 3528
rect 9171 3519 9229 3525
rect 9171 3485 9183 3519
rect 9217 3516 9229 3519
rect 9766 3516 9772 3528
rect 9217 3488 9772 3516
rect 9217 3485 9229 3488
rect 9171 3479 9229 3485
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3516 11391 3519
rect 11514 3516 11520 3528
rect 11379 3488 11520 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 11514 3476 11520 3488
rect 11572 3476 11578 3528
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 11054 3408 11060 3460
rect 11112 3448 11118 3460
rect 11624 3448 11652 3479
rect 11790 3476 11796 3528
rect 11848 3516 11854 3528
rect 12087 3527 12115 3556
rect 14553 3553 14565 3556
rect 14599 3553 14611 3587
rect 14553 3547 14611 3553
rect 15933 3587 15991 3593
rect 15933 3553 15945 3587
rect 15979 3584 15991 3587
rect 15979 3556 16623 3584
rect 15979 3553 15991 3556
rect 15933 3547 15991 3553
rect 11936 3519 11994 3525
rect 11936 3516 11948 3519
rect 11848 3488 11948 3516
rect 11848 3476 11854 3488
rect 11936 3485 11948 3488
rect 11982 3485 11994 3519
rect 11936 3479 11994 3485
rect 12072 3521 12130 3527
rect 12072 3487 12084 3521
rect 12118 3487 12130 3521
rect 12072 3481 12130 3487
rect 12342 3476 12348 3528
rect 12400 3476 12406 3528
rect 13538 3476 13544 3528
rect 13596 3476 13602 3528
rect 13814 3476 13820 3528
rect 13872 3476 13878 3528
rect 14274 3476 14280 3528
rect 14332 3476 14338 3528
rect 16114 3476 16120 3528
rect 16172 3476 16178 3528
rect 16595 3527 16623 3556
rect 16666 3544 16672 3596
rect 16724 3584 16730 3596
rect 16853 3587 16911 3593
rect 16853 3584 16865 3587
rect 16724 3556 16865 3584
rect 16724 3544 16730 3556
rect 16853 3553 16865 3556
rect 16899 3553 16911 3587
rect 16853 3547 16911 3553
rect 18233 3587 18291 3593
rect 18233 3553 18245 3587
rect 18279 3584 18291 3587
rect 19061 3587 19119 3593
rect 18279 3556 18828 3584
rect 18279 3553 18291 3556
rect 18233 3547 18291 3553
rect 16580 3521 16638 3527
rect 16580 3487 16592 3521
rect 16626 3487 16638 3521
rect 16580 3481 16638 3487
rect 18325 3519 18383 3525
rect 18325 3485 18337 3519
rect 18371 3516 18383 3519
rect 18506 3516 18512 3528
rect 18371 3488 18512 3516
rect 18371 3485 18383 3488
rect 18325 3479 18383 3485
rect 18506 3476 18512 3488
rect 18564 3476 18570 3528
rect 18800 3525 18828 3556
rect 19061 3553 19073 3587
rect 19107 3584 19119 3587
rect 19334 3584 19340 3596
rect 19107 3556 19340 3584
rect 19107 3553 19119 3556
rect 19061 3547 19119 3553
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 20533 3587 20591 3593
rect 20533 3553 20545 3587
rect 20579 3553 20591 3587
rect 20533 3547 20591 3553
rect 20809 3587 20867 3593
rect 20809 3553 20821 3587
rect 20855 3584 20867 3587
rect 20990 3584 20996 3596
rect 20855 3556 20996 3584
rect 20855 3553 20867 3556
rect 20809 3547 20867 3553
rect 18788 3519 18846 3525
rect 18788 3485 18800 3519
rect 18834 3485 18846 3519
rect 18788 3479 18846 3485
rect 19242 3476 19248 3528
rect 19300 3516 19306 3528
rect 20548 3516 20576 3547
rect 20990 3544 20996 3556
rect 21048 3544 21054 3596
rect 19300 3488 20576 3516
rect 21269 3519 21327 3525
rect 19300 3476 19306 3488
rect 21269 3485 21281 3519
rect 21315 3485 21327 3519
rect 21376 3516 21404 3624
rect 21818 3544 21824 3596
rect 21876 3584 21882 3596
rect 22005 3587 22063 3593
rect 22005 3584 22017 3587
rect 21876 3556 22017 3584
rect 21876 3544 21882 3556
rect 22005 3553 22017 3556
rect 22051 3553 22063 3587
rect 23584 3584 23612 3624
rect 24213 3587 24271 3593
rect 24213 3584 24225 3587
rect 23584 3556 24225 3584
rect 22005 3547 22063 3553
rect 24213 3553 24225 3556
rect 24259 3553 24271 3587
rect 24213 3547 24271 3553
rect 24486 3544 24492 3596
rect 24544 3544 24550 3596
rect 25498 3544 25504 3596
rect 25556 3584 25562 3596
rect 26620 3593 26648 3692
rect 26694 3680 26700 3732
rect 26752 3680 26758 3732
rect 26712 3652 26740 3680
rect 26973 3655 27031 3661
rect 26973 3652 26985 3655
rect 26712 3624 26985 3652
rect 26973 3621 26985 3624
rect 27019 3621 27031 3655
rect 26973 3615 27031 3621
rect 27614 3612 27620 3664
rect 27672 3652 27678 3664
rect 27798 3652 27804 3664
rect 27672 3624 27804 3652
rect 27672 3612 27678 3624
rect 27798 3612 27804 3624
rect 27856 3612 27862 3664
rect 25685 3587 25743 3593
rect 25685 3584 25697 3587
rect 25556 3556 25697 3584
rect 25556 3544 25562 3556
rect 25685 3553 25697 3556
rect 25731 3584 25743 3587
rect 26605 3587 26663 3593
rect 25731 3556 26556 3584
rect 25731 3553 25743 3556
rect 25685 3547 25743 3553
rect 21732 3519 21790 3525
rect 21732 3516 21744 3519
rect 21376 3488 21744 3516
rect 21269 3479 21327 3485
rect 21732 3485 21744 3488
rect 21778 3485 21790 3519
rect 21732 3479 21790 3485
rect 23477 3519 23535 3525
rect 23477 3485 23489 3519
rect 23523 3516 23535 3519
rect 23750 3516 23756 3528
rect 23523 3488 23756 3516
rect 23523 3485 23535 3488
rect 23477 3479 23535 3485
rect 11112 3420 11652 3448
rect 11112 3408 11118 3420
rect 9214 3380 9220 3392
rect 5552 3352 9220 3380
rect 9214 3340 9220 3352
rect 9272 3340 9278 3392
rect 13556 3380 13584 3476
rect 19978 3408 19984 3460
rect 20036 3448 20042 3460
rect 20898 3448 20904 3460
rect 20036 3420 20904 3448
rect 20036 3408 20042 3420
rect 20898 3408 20904 3420
rect 20956 3448 20962 3460
rect 21284 3448 21312 3479
rect 23750 3476 23756 3488
rect 23808 3476 23814 3528
rect 23842 3476 23848 3528
rect 23900 3516 23906 3528
rect 23940 3519 23998 3525
rect 23940 3516 23952 3519
rect 23900 3488 23952 3516
rect 23900 3476 23906 3488
rect 23940 3485 23952 3488
rect 23986 3485 23998 3519
rect 24504 3516 24532 3544
rect 25869 3519 25927 3525
rect 25869 3516 25881 3519
rect 24504 3488 25881 3516
rect 23940 3479 23998 3485
rect 25869 3485 25881 3488
rect 25915 3485 25927 3519
rect 26528 3516 26556 3556
rect 26605 3553 26617 3587
rect 26651 3553 26663 3587
rect 26605 3547 26663 3553
rect 26697 3587 26755 3593
rect 26697 3553 26709 3587
rect 26743 3584 26755 3587
rect 27341 3587 27399 3593
rect 27341 3584 27353 3587
rect 26743 3556 27353 3584
rect 26743 3553 26755 3556
rect 26697 3547 26755 3553
rect 27341 3553 27353 3556
rect 27387 3553 27399 3587
rect 27341 3547 27399 3553
rect 26712 3516 26740 3547
rect 27890 3544 27896 3596
rect 27948 3544 27954 3596
rect 28258 3525 28264 3528
rect 26528 3488 26740 3516
rect 28220 3519 28264 3525
rect 25869 3479 25927 3485
rect 28220 3485 28232 3519
rect 28220 3479 28264 3485
rect 28258 3476 28264 3479
rect 28316 3476 28322 3528
rect 28399 3519 28457 3525
rect 28399 3485 28411 3519
rect 28445 3516 28457 3519
rect 28534 3516 28540 3528
rect 28445 3488 28540 3516
rect 28445 3485 28457 3488
rect 28399 3479 28457 3485
rect 28534 3476 28540 3488
rect 28592 3476 28598 3528
rect 28629 3519 28687 3525
rect 28629 3485 28641 3519
rect 28675 3516 28687 3519
rect 28810 3516 28816 3528
rect 28675 3488 28816 3516
rect 28675 3485 28687 3488
rect 28629 3479 28687 3485
rect 28810 3476 28816 3488
rect 28868 3476 28874 3528
rect 20956 3420 21312 3448
rect 20956 3408 20962 3420
rect 25774 3408 25780 3460
rect 25832 3448 25838 3460
rect 29733 3451 29791 3457
rect 25832 3420 26556 3448
rect 25832 3408 25838 3420
rect 16390 3380 16396 3392
rect 13556 3352 16396 3380
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 16482 3340 16488 3392
rect 16540 3380 16546 3392
rect 19518 3380 19524 3392
rect 16540 3352 19524 3380
rect 16540 3340 16546 3352
rect 19518 3340 19524 3352
rect 19576 3340 19582 3392
rect 23290 3340 23296 3392
rect 23348 3340 23354 3392
rect 25314 3340 25320 3392
rect 25372 3340 25378 3392
rect 26418 3340 26424 3392
rect 26476 3340 26482 3392
rect 26528 3380 26556 3420
rect 29733 3417 29745 3451
rect 29779 3417 29791 3451
rect 29733 3411 29791 3417
rect 29748 3380 29776 3411
rect 26528 3352 29776 3380
rect 552 3290 30912 3312
rect 552 3238 4193 3290
rect 4245 3238 4257 3290
rect 4309 3238 4321 3290
rect 4373 3238 4385 3290
rect 4437 3238 4449 3290
rect 4501 3238 11783 3290
rect 11835 3238 11847 3290
rect 11899 3238 11911 3290
rect 11963 3238 11975 3290
rect 12027 3238 12039 3290
rect 12091 3238 19373 3290
rect 19425 3238 19437 3290
rect 19489 3238 19501 3290
rect 19553 3238 19565 3290
rect 19617 3238 19629 3290
rect 19681 3238 26963 3290
rect 27015 3238 27027 3290
rect 27079 3238 27091 3290
rect 27143 3238 27155 3290
rect 27207 3238 27219 3290
rect 27271 3238 30912 3290
rect 552 3216 30912 3238
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 5537 3179 5595 3185
rect 5537 3176 5549 3179
rect 5316 3148 5549 3176
rect 5316 3136 5322 3148
rect 5537 3145 5549 3148
rect 5583 3145 5595 3179
rect 7282 3176 7288 3188
rect 5537 3139 5595 3145
rect 5644 3148 7288 3176
rect 5442 3068 5448 3120
rect 5500 3108 5506 3120
rect 5644 3108 5672 3148
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 9858 3176 9864 3188
rect 8168 3148 9864 3176
rect 8168 3136 8174 3148
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 10962 3136 10968 3188
rect 11020 3176 11026 3188
rect 13265 3179 13323 3185
rect 11020 3148 13216 3176
rect 11020 3136 11026 3148
rect 5500 3080 5672 3108
rect 5500 3068 5506 3080
rect 8846 3068 8852 3120
rect 8904 3108 8910 3120
rect 8904 3080 9076 3108
rect 8904 3068 8910 3080
rect 937 3043 995 3049
rect 937 3009 949 3043
rect 983 3040 995 3043
rect 1302 3040 1308 3052
rect 983 3012 1308 3040
rect 983 3009 995 3012
rect 937 3003 995 3009
rect 1302 3000 1308 3012
rect 1360 3000 1366 3052
rect 2958 3040 2964 3052
rect 1458 3031 2964 3040
rect 1433 3025 2964 3031
rect 1433 2991 1445 3025
rect 1479 3012 2964 3025
rect 1479 2991 1491 3012
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3040 3111 3043
rect 4062 3040 4068 3052
rect 3099 3012 4068 3040
rect 3099 3009 3111 3012
rect 3053 3003 3111 3009
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4203 3043 4261 3049
rect 4203 3009 4215 3043
rect 4249 3040 4261 3043
rect 4614 3040 4620 3052
rect 4249 3012 4620 3040
rect 4249 3009 4261 3012
rect 4203 3003 4261 3009
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 5994 3000 6000 3052
rect 6052 3040 6058 3052
rect 6089 3043 6147 3049
rect 6089 3040 6101 3043
rect 6052 3012 6101 3040
rect 6052 3000 6058 3012
rect 6089 3009 6101 3012
rect 6135 3009 6147 3043
rect 6089 3003 6147 3009
rect 6196 3031 6595 3040
rect 6196 3025 6610 3031
rect 6196 3012 6564 3025
rect 1433 2985 1491 2991
rect 1670 2932 1676 2984
rect 1728 2932 1734 2984
rect 3234 2932 3240 2984
rect 3292 2972 3298 2984
rect 3510 2972 3516 2984
rect 3292 2944 3516 2972
rect 3292 2932 3298 2944
rect 3510 2932 3516 2944
rect 3568 2972 3574 2984
rect 3697 2975 3755 2981
rect 3697 2972 3709 2975
rect 3568 2944 3709 2972
rect 3568 2932 3574 2944
rect 3697 2941 3709 2944
rect 3743 2941 3755 2975
rect 3697 2935 3755 2941
rect 4433 2975 4491 2981
rect 4433 2941 4445 2975
rect 4479 2972 4491 2975
rect 5166 2972 5172 2984
rect 4479 2944 5172 2972
rect 4479 2941 4491 2944
rect 4433 2935 4491 2941
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 6196 2972 6224 3012
rect 6552 2991 6564 3012
rect 6598 2991 6610 3025
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 8570 3040 8576 3052
rect 7800 3012 8576 3040
rect 7800 3000 7806 3012
rect 8570 3000 8576 3012
rect 8628 3040 8634 3052
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 8628 3012 8769 3040
rect 8628 3000 8634 3012
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 6552 2985 6610 2991
rect 9048 2981 9076 3080
rect 9496 3043 9554 3049
rect 9496 3040 9508 3043
rect 9416 3012 9508 3040
rect 5552 2944 6224 2972
rect 6825 2975 6883 2981
rect 5552 2848 5580 2944
rect 6825 2941 6837 2975
rect 6871 2972 6883 2975
rect 8205 2975 8263 2981
rect 6871 2944 8156 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 1403 2839 1461 2845
rect 1403 2805 1415 2839
rect 1449 2836 1461 2839
rect 1762 2836 1768 2848
rect 1449 2808 1768 2836
rect 1449 2805 1461 2808
rect 1403 2799 1461 2805
rect 1762 2796 1768 2808
rect 1820 2796 1826 2848
rect 4154 2796 4160 2848
rect 4212 2845 4218 2848
rect 4212 2836 4221 2845
rect 4522 2836 4528 2848
rect 4212 2808 4528 2836
rect 4212 2799 4221 2808
rect 4212 2796 4218 2799
rect 4522 2796 4528 2808
rect 4580 2796 4586 2848
rect 5534 2796 5540 2848
rect 5592 2796 5598 2848
rect 5718 2796 5724 2848
rect 5776 2836 5782 2848
rect 6555 2839 6613 2845
rect 6555 2836 6567 2839
rect 5776 2808 6567 2836
rect 5776 2796 5782 2808
rect 6555 2805 6567 2808
rect 6601 2836 6613 2839
rect 6914 2836 6920 2848
rect 6601 2808 6920 2836
rect 6601 2805 6613 2808
rect 6555 2799 6613 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 8128 2836 8156 2944
rect 8205 2941 8217 2975
rect 8251 2972 8263 2975
rect 9033 2975 9091 2981
rect 8251 2944 8984 2972
rect 8251 2941 8263 2944
rect 8205 2935 8263 2941
rect 8481 2907 8539 2913
rect 8481 2873 8493 2907
rect 8527 2904 8539 2907
rect 8846 2904 8852 2916
rect 8527 2876 8852 2904
rect 8527 2873 8539 2876
rect 8481 2867 8539 2873
rect 8846 2864 8852 2876
rect 8904 2864 8910 2916
rect 8956 2904 8984 2944
rect 9033 2941 9045 2975
rect 9079 2941 9091 2975
rect 9416 2972 9444 3012
rect 9496 3009 9508 3012
rect 9542 3009 9554 3043
rect 9496 3003 9554 3009
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 9769 3043 9827 3049
rect 9769 3040 9781 3043
rect 9732 3012 9781 3040
rect 9732 3000 9738 3012
rect 9769 3009 9781 3012
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 11704 3043 11762 3049
rect 11704 3040 11716 3043
rect 11195 3012 11716 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 11704 3009 11716 3012
rect 11750 3009 11762 3043
rect 13188 3040 13216 3148
rect 13265 3145 13277 3179
rect 13311 3176 13323 3179
rect 14274 3176 14280 3188
rect 13311 3148 14280 3176
rect 13311 3145 13323 3148
rect 13265 3139 13323 3145
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 16942 3136 16948 3188
rect 17000 3176 17006 3188
rect 25958 3176 25964 3188
rect 17000 3148 25964 3176
rect 17000 3136 17006 3148
rect 25958 3136 25964 3148
rect 26016 3136 26022 3188
rect 30006 3176 30012 3188
rect 26068 3148 30012 3176
rect 22925 3111 22983 3117
rect 22925 3077 22937 3111
rect 22971 3108 22983 3111
rect 23842 3108 23848 3120
rect 22971 3080 23848 3108
rect 22971 3077 22983 3080
rect 22925 3071 22983 3077
rect 23842 3068 23848 3080
rect 23900 3068 23906 3120
rect 25498 3068 25504 3120
rect 25556 3068 25562 3120
rect 25866 3068 25872 3120
rect 25924 3108 25930 3120
rect 26068 3108 26096 3148
rect 30006 3136 30012 3148
rect 30064 3136 30070 3188
rect 25924 3080 26096 3108
rect 28629 3111 28687 3117
rect 25924 3068 25930 3080
rect 28629 3077 28641 3111
rect 28675 3077 28687 3111
rect 28629 3071 28687 3077
rect 14139 3043 14197 3049
rect 13188 3012 13768 3040
rect 11704 3003 11762 3009
rect 9033 2935 9091 2941
rect 9146 2944 9444 2972
rect 9146 2904 9174 2944
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 11112 2944 11253 2972
rect 11112 2932 11118 2944
rect 11241 2941 11253 2944
rect 11287 2941 11299 2975
rect 11241 2935 11299 2941
rect 11330 2932 11336 2984
rect 11388 2972 11394 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11388 2944 11989 2972
rect 11388 2932 11394 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 13630 2932 13636 2984
rect 13688 2932 13694 2984
rect 13740 2972 13768 3012
rect 14139 3009 14151 3043
rect 14185 3040 14197 3043
rect 15102 3040 15108 3052
rect 14185 3012 15108 3040
rect 14185 3009 14197 3012
rect 14139 3003 14197 3009
rect 15102 3000 15108 3012
rect 15160 3000 15166 3052
rect 16022 3000 16028 3052
rect 16080 3040 16086 3052
rect 16304 3043 16362 3049
rect 16304 3040 16316 3043
rect 16080 3012 16316 3040
rect 16080 3000 16086 3012
rect 16304 3009 16316 3012
rect 16350 3009 16362 3043
rect 16304 3003 16362 3009
rect 16390 3000 16396 3052
rect 16448 3040 16454 3052
rect 16577 3043 16635 3049
rect 16577 3040 16589 3043
rect 16448 3012 16589 3040
rect 16448 3000 16454 3012
rect 16577 3009 16589 3012
rect 16623 3009 16635 3043
rect 16577 3003 16635 3009
rect 17957 3043 18015 3049
rect 17957 3009 17969 3043
rect 18003 3040 18015 3043
rect 19156 3043 19214 3049
rect 19156 3040 19168 3043
rect 18003 3012 19168 3040
rect 18003 3009 18015 3012
rect 17957 3003 18015 3009
rect 19156 3009 19168 3012
rect 19202 3009 19214 3043
rect 19156 3003 19214 3009
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 21364 3043 21422 3049
rect 21364 3040 21376 3043
rect 20855 3012 21376 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 21364 3009 21376 3012
rect 21410 3009 21422 3043
rect 21364 3003 21422 3009
rect 23290 3000 23296 3052
rect 23348 3040 23354 3052
rect 24308 3043 24366 3049
rect 24308 3040 24320 3043
rect 23348 3012 24320 3040
rect 23348 3000 23354 3012
rect 24308 3009 24320 3012
rect 24354 3009 24366 3043
rect 24308 3003 24366 3009
rect 24394 3000 24400 3052
rect 24452 3040 24458 3052
rect 24581 3043 24639 3049
rect 24581 3040 24593 3043
rect 24452 3012 24593 3040
rect 24452 3000 24458 3012
rect 24581 3009 24593 3012
rect 24627 3009 24639 3043
rect 24581 3003 24639 3009
rect 14274 2972 14280 2984
rect 13740 2944 14280 2972
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 14366 2932 14372 2984
rect 14424 2932 14430 2984
rect 15841 2975 15899 2981
rect 15841 2941 15853 2975
rect 15887 2972 15899 2975
rect 16114 2972 16120 2984
rect 15887 2944 16120 2972
rect 15887 2941 15899 2944
rect 15841 2935 15899 2941
rect 16114 2932 16120 2944
rect 16172 2972 16178 2984
rect 18141 2975 18199 2981
rect 16172 2944 17264 2972
rect 16172 2932 16178 2944
rect 8956 2876 9174 2904
rect 9306 2836 9312 2848
rect 8128 2808 9312 2836
rect 9306 2796 9312 2808
rect 9364 2796 9370 2848
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 9499 2839 9557 2845
rect 9499 2836 9511 2839
rect 9456 2808 9511 2836
rect 9456 2796 9462 2808
rect 9499 2805 9511 2808
rect 9545 2805 9557 2839
rect 9499 2799 9557 2805
rect 11698 2796 11704 2848
rect 11756 2845 11762 2848
rect 11756 2836 11765 2845
rect 11756 2808 11801 2836
rect 11756 2799 11765 2808
rect 11756 2796 11762 2799
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 14099 2839 14157 2845
rect 14099 2836 14111 2839
rect 13964 2808 14111 2836
rect 13964 2796 13970 2808
rect 14099 2805 14111 2808
rect 14145 2836 14157 2839
rect 15010 2836 15016 2848
rect 14145 2808 15016 2836
rect 14145 2805 14157 2808
rect 14099 2799 14157 2805
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 15194 2796 15200 2848
rect 15252 2836 15258 2848
rect 15473 2839 15531 2845
rect 15473 2836 15485 2839
rect 15252 2808 15485 2836
rect 15252 2796 15258 2808
rect 15473 2805 15485 2808
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 16307 2839 16365 2845
rect 16307 2805 16319 2839
rect 16353 2836 16365 2839
rect 16574 2836 16580 2848
rect 16353 2808 16580 2836
rect 16353 2805 16365 2808
rect 16307 2799 16365 2805
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 17236 2836 17264 2944
rect 18141 2941 18153 2975
rect 18187 2972 18199 2975
rect 18506 2972 18512 2984
rect 18187 2944 18512 2972
rect 18187 2941 18199 2944
rect 18141 2935 18199 2941
rect 18506 2932 18512 2944
rect 18564 2972 18570 2984
rect 18693 2975 18751 2981
rect 18693 2972 18705 2975
rect 18564 2944 18705 2972
rect 18564 2932 18570 2944
rect 18693 2941 18705 2944
rect 18739 2941 18751 2975
rect 18693 2935 18751 2941
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2972 19487 2975
rect 19702 2972 19708 2984
rect 19475 2944 19708 2972
rect 19475 2941 19487 2944
rect 19429 2935 19487 2941
rect 19702 2932 19708 2944
rect 19760 2932 19766 2984
rect 20898 2932 20904 2984
rect 20956 2932 20962 2984
rect 21266 2932 21272 2984
rect 21324 2972 21330 2984
rect 21637 2975 21695 2981
rect 21637 2972 21649 2975
rect 21324 2944 21649 2972
rect 21324 2932 21330 2944
rect 21637 2941 21649 2944
rect 21683 2941 21695 2975
rect 21637 2935 21695 2941
rect 22646 2932 22652 2984
rect 22704 2972 22710 2984
rect 23569 2975 23627 2981
rect 22704 2944 23336 2972
rect 22704 2932 22710 2944
rect 23201 2907 23259 2913
rect 23201 2873 23213 2907
rect 23247 2873 23259 2907
rect 23308 2904 23336 2944
rect 23569 2941 23581 2975
rect 23615 2972 23627 2975
rect 23750 2972 23756 2984
rect 23615 2944 23756 2972
rect 23615 2941 23627 2944
rect 23569 2935 23627 2941
rect 23750 2932 23756 2944
rect 23808 2972 23814 2984
rect 23845 2975 23903 2981
rect 23845 2972 23857 2975
rect 23808 2944 23857 2972
rect 23808 2932 23814 2944
rect 23845 2941 23857 2944
rect 23891 2941 23903 2975
rect 25516 2972 25544 3068
rect 26142 3000 26148 3052
rect 26200 3040 26206 3052
rect 26700 3043 26758 3049
rect 26700 3040 26712 3043
rect 26200 3012 26712 3040
rect 26200 3000 26206 3012
rect 26700 3009 26712 3012
rect 26746 3009 26758 3043
rect 26700 3003 26758 3009
rect 27062 3000 27068 3052
rect 27120 3040 27126 3052
rect 28644 3040 28672 3071
rect 27120 3012 28672 3040
rect 27120 3000 27126 3012
rect 23845 2935 23903 2941
rect 23952 2944 25544 2972
rect 23952 2904 23980 2944
rect 26234 2932 26240 2984
rect 26292 2932 26298 2984
rect 26602 2932 26608 2984
rect 26660 2972 26666 2984
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26660 2944 26985 2972
rect 26660 2932 26666 2944
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 26973 2935 27031 2941
rect 27430 2932 27436 2984
rect 27488 2972 27494 2984
rect 28445 2975 28503 2981
rect 28445 2972 28457 2975
rect 27488 2944 28457 2972
rect 27488 2932 27494 2944
rect 28445 2941 28457 2944
rect 28491 2941 28503 2975
rect 28445 2935 28503 2941
rect 23308 2876 23980 2904
rect 23201 2867 23259 2873
rect 18233 2839 18291 2845
rect 18233 2836 18245 2839
rect 17236 2808 18245 2836
rect 18233 2805 18245 2808
rect 18279 2805 18291 2839
rect 18233 2799 18291 2805
rect 18966 2796 18972 2848
rect 19024 2836 19030 2848
rect 19159 2839 19217 2845
rect 19159 2836 19171 2839
rect 19024 2808 19171 2836
rect 19024 2796 19030 2808
rect 19159 2805 19171 2808
rect 19205 2805 19217 2839
rect 19159 2799 19217 2805
rect 21367 2839 21425 2845
rect 21367 2805 21379 2839
rect 21413 2836 21425 2839
rect 21542 2836 21548 2848
rect 21413 2808 21548 2836
rect 21413 2805 21425 2808
rect 21367 2799 21425 2805
rect 21542 2796 21548 2808
rect 21600 2796 21606 2848
rect 23216 2836 23244 2867
rect 23842 2836 23848 2848
rect 23216 2808 23848 2836
rect 23842 2796 23848 2808
rect 23900 2796 23906 2848
rect 24118 2796 24124 2848
rect 24176 2836 24182 2848
rect 24311 2839 24369 2845
rect 24311 2836 24323 2839
rect 24176 2808 24323 2836
rect 24176 2796 24182 2808
rect 24311 2805 24323 2808
rect 24357 2805 24369 2839
rect 24311 2799 24369 2805
rect 24670 2796 24676 2848
rect 24728 2836 24734 2848
rect 25685 2839 25743 2845
rect 25685 2836 25697 2839
rect 24728 2808 25697 2836
rect 24728 2796 24734 2808
rect 25685 2805 25697 2808
rect 25731 2805 25743 2839
rect 25685 2799 25743 2805
rect 26694 2796 26700 2848
rect 26752 2845 26758 2848
rect 26752 2836 26761 2845
rect 26752 2808 26797 2836
rect 26752 2799 26761 2808
rect 26752 2796 26758 2799
rect 27614 2796 27620 2848
rect 27672 2836 27678 2848
rect 28077 2839 28135 2845
rect 28077 2836 28089 2839
rect 27672 2808 28089 2836
rect 27672 2796 27678 2808
rect 28077 2805 28089 2808
rect 28123 2805 28135 2839
rect 28077 2799 28135 2805
rect 552 2746 31072 2768
rect 552 2694 7988 2746
rect 8040 2694 8052 2746
rect 8104 2694 8116 2746
rect 8168 2694 8180 2746
rect 8232 2694 8244 2746
rect 8296 2694 15578 2746
rect 15630 2694 15642 2746
rect 15694 2694 15706 2746
rect 15758 2694 15770 2746
rect 15822 2694 15834 2746
rect 15886 2694 23168 2746
rect 23220 2694 23232 2746
rect 23284 2694 23296 2746
rect 23348 2694 23360 2746
rect 23412 2694 23424 2746
rect 23476 2694 30758 2746
rect 30810 2694 30822 2746
rect 30874 2694 30886 2746
rect 30938 2694 30950 2746
rect 31002 2694 31014 2746
rect 31066 2694 31072 2746
rect 552 2672 31072 2694
rect 658 2592 664 2644
rect 716 2632 722 2644
rect 937 2635 995 2641
rect 937 2632 949 2635
rect 716 2604 949 2632
rect 716 2592 722 2604
rect 937 2601 949 2604
rect 983 2601 995 2635
rect 937 2595 995 2601
rect 1394 2592 1400 2644
rect 1452 2632 1458 2644
rect 1946 2632 1952 2644
rect 1452 2604 1952 2632
rect 1452 2592 1458 2604
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 2038 2592 2044 2644
rect 2096 2632 2102 2644
rect 5718 2632 5724 2644
rect 2096 2604 5724 2632
rect 2096 2592 2102 2604
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 6457 2635 6515 2641
rect 6457 2632 6469 2635
rect 5868 2604 6469 2632
rect 5868 2592 5874 2604
rect 6457 2601 6469 2604
rect 6503 2601 6515 2635
rect 6457 2595 6515 2601
rect 6914 2592 6920 2644
rect 6972 2592 6978 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7469 2635 7527 2641
rect 7469 2632 7481 2635
rect 7248 2604 7481 2632
rect 7248 2592 7254 2604
rect 7469 2601 7481 2604
rect 7515 2601 7527 2635
rect 8211 2635 8269 2641
rect 8211 2632 8223 2635
rect 7469 2595 7527 2601
rect 7576 2604 8223 2632
rect 3050 2524 3056 2576
rect 3108 2564 3114 2576
rect 3108 2536 5764 2564
rect 3108 2524 3114 2536
rect 1026 2456 1032 2508
rect 1084 2496 1090 2508
rect 1121 2499 1179 2505
rect 1121 2496 1133 2499
rect 1084 2468 1133 2496
rect 1084 2456 1090 2468
rect 1121 2465 1133 2468
rect 1167 2465 1179 2499
rect 1121 2459 1179 2465
rect 1632 2499 1690 2505
rect 1632 2465 1644 2499
rect 1678 2496 1690 2499
rect 1946 2496 1952 2508
rect 1678 2468 1952 2496
rect 1678 2465 1690 2468
rect 1632 2459 1690 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2041 2499 2099 2505
rect 2041 2465 2053 2499
rect 2087 2496 2099 2499
rect 3789 2499 3847 2505
rect 3789 2496 3801 2499
rect 2087 2468 3801 2496
rect 2087 2465 2099 2468
rect 2041 2459 2099 2465
rect 3789 2465 3801 2468
rect 3835 2496 3847 2499
rect 5074 2496 5080 2508
rect 3835 2468 5080 2496
rect 3835 2465 3847 2468
rect 3789 2459 3847 2465
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 5736 2496 5764 2536
rect 6086 2524 6092 2576
rect 6144 2524 6150 2576
rect 6932 2564 6960 2592
rect 7576 2564 7604 2604
rect 8211 2601 8223 2604
rect 8257 2632 8269 2635
rect 8386 2632 8392 2644
rect 8257 2604 8392 2632
rect 8257 2601 8269 2604
rect 8211 2595 8269 2601
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 9766 2592 9772 2644
rect 9824 2592 9830 2644
rect 10042 2592 10048 2644
rect 10100 2592 10106 2644
rect 10321 2635 10379 2641
rect 10321 2601 10333 2635
rect 10367 2601 10379 2635
rect 10321 2595 10379 2601
rect 6932 2536 7604 2564
rect 10336 2564 10364 2595
rect 10594 2592 10600 2644
rect 10652 2592 10658 2644
rect 10870 2592 10876 2644
rect 10928 2632 10934 2644
rect 10928 2604 11652 2632
rect 10928 2592 10934 2604
rect 11514 2564 11520 2576
rect 10336 2536 11520 2564
rect 11514 2524 11520 2536
rect 11572 2524 11578 2576
rect 5994 2496 6000 2508
rect 5736 2468 6000 2496
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6104 2496 6132 2524
rect 6181 2499 6239 2505
rect 6181 2496 6193 2499
rect 6104 2468 6193 2496
rect 6181 2465 6193 2468
rect 6227 2465 6239 2499
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 6181 2459 6239 2465
rect 6294 2468 6377 2496
rect 1854 2439 1860 2440
rect 1305 2431 1363 2437
rect 1305 2397 1317 2431
rect 1351 2397 1363 2431
rect 1305 2391 1363 2397
rect 1811 2433 1860 2439
rect 1811 2399 1823 2433
rect 1857 2399 1860 2433
rect 1811 2393 1860 2399
rect 1320 2292 1348 2391
rect 1854 2388 1860 2393
rect 1912 2388 1918 2440
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 6018 2428 6046 2456
rect 6294 2428 6322 2468
rect 6365 2465 6377 2468
rect 6411 2496 6423 2499
rect 6454 2496 6460 2508
rect 6411 2468 6460 2496
rect 6411 2465 6423 2468
rect 6365 2459 6423 2465
rect 6454 2456 6460 2468
rect 6512 2456 6518 2508
rect 6822 2456 6828 2508
rect 6880 2496 6886 2508
rect 7098 2496 7104 2508
rect 6880 2468 7104 2496
rect 6880 2456 6886 2468
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 7653 2499 7711 2505
rect 7653 2465 7665 2499
rect 7699 2465 7711 2499
rect 7653 2459 7711 2465
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 4580 2400 5948 2428
rect 6018 2400 6322 2428
rect 6380 2400 7021 2428
rect 4580 2388 4586 2400
rect 4982 2360 4988 2372
rect 3252 2332 4988 2360
rect 3252 2304 3280 2332
rect 4982 2320 4988 2332
rect 5040 2320 5046 2372
rect 3050 2292 3056 2304
rect 1320 2264 3056 2292
rect 3050 2252 3056 2264
rect 3108 2252 3114 2304
rect 3234 2252 3240 2304
rect 3292 2252 3298 2304
rect 3329 2295 3387 2301
rect 3329 2261 3341 2295
rect 3375 2292 3387 2295
rect 4890 2292 4896 2304
rect 3375 2264 4896 2292
rect 3375 2261 3387 2264
rect 3329 2255 3387 2261
rect 4890 2252 4896 2264
rect 4948 2252 4954 2304
rect 5920 2292 5948 2400
rect 5994 2320 6000 2372
rect 6052 2320 6058 2372
rect 6380 2292 6408 2400
rect 7009 2397 7021 2400
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 7466 2388 7472 2440
rect 7524 2428 7530 2440
rect 7668 2428 7696 2459
rect 7834 2456 7840 2508
rect 7892 2496 7898 2508
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 7892 2468 8493 2496
rect 7892 2456 7898 2468
rect 8481 2465 8493 2468
rect 8527 2465 8539 2499
rect 8481 2459 8539 2465
rect 8570 2456 8576 2508
rect 8628 2496 8634 2508
rect 9490 2496 9496 2508
rect 8628 2468 9496 2496
rect 8628 2456 8634 2468
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 10229 2499 10287 2505
rect 10229 2496 10241 2499
rect 9784 2468 10241 2496
rect 9784 2440 9812 2468
rect 10229 2465 10241 2468
rect 10275 2465 10287 2499
rect 10229 2459 10287 2465
rect 10502 2456 10508 2508
rect 10560 2456 10566 2508
rect 10781 2499 10839 2505
rect 10781 2465 10793 2499
rect 10827 2465 10839 2499
rect 10781 2459 10839 2465
rect 7524 2400 7696 2428
rect 7524 2388 7530 2400
rect 7742 2388 7748 2440
rect 7800 2388 7806 2440
rect 8202 2388 8208 2440
rect 8260 2388 8266 2440
rect 8294 2388 8300 2440
rect 8352 2428 8358 2440
rect 9674 2428 9680 2440
rect 8352 2400 9680 2428
rect 8352 2388 8358 2400
rect 9646 2388 9680 2400
rect 9732 2388 9738 2440
rect 9766 2388 9772 2440
rect 9824 2388 9830 2440
rect 10796 2428 10824 2459
rect 11054 2456 11060 2508
rect 11112 2496 11118 2508
rect 11624 2496 11652 2604
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14191 2635 14249 2641
rect 14191 2632 14203 2635
rect 14056 2604 14203 2632
rect 14056 2592 14062 2604
rect 14191 2601 14203 2604
rect 14237 2601 14249 2635
rect 14191 2595 14249 2601
rect 16574 2592 16580 2644
rect 16632 2641 16638 2644
rect 16632 2632 16641 2641
rect 18791 2635 18849 2641
rect 16632 2604 16677 2632
rect 16632 2595 16641 2604
rect 18791 2601 18803 2635
rect 18837 2632 18849 2635
rect 18966 2632 18972 2644
rect 18837 2604 18972 2632
rect 18837 2601 18849 2604
rect 18791 2595 18849 2601
rect 16632 2592 16638 2595
rect 18966 2592 18972 2604
rect 19024 2592 19030 2644
rect 20809 2635 20867 2641
rect 20809 2632 20821 2635
rect 20640 2604 20821 2632
rect 13633 2499 13691 2505
rect 11112 2468 11560 2496
rect 11624 2468 12296 2496
rect 11112 2456 11118 2468
rect 11532 2437 11560 2468
rect 9876 2400 10824 2428
rect 11517 2431 11575 2437
rect 6454 2320 6460 2372
rect 6512 2360 6518 2372
rect 7760 2360 7788 2388
rect 6512 2332 7788 2360
rect 9646 2360 9674 2388
rect 9876 2360 9904 2400
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 11844 2431 11902 2437
rect 11844 2428 11856 2431
rect 11756 2400 11856 2428
rect 11756 2388 11762 2400
rect 11844 2397 11856 2400
rect 11890 2397 11902 2431
rect 11844 2391 11902 2397
rect 12023 2431 12081 2437
rect 12023 2397 12035 2431
rect 12069 2428 12081 2431
rect 12158 2428 12164 2440
rect 12069 2400 12164 2428
rect 12069 2397 12081 2400
rect 12023 2391 12081 2397
rect 12158 2388 12164 2400
rect 12216 2388 12222 2440
rect 12268 2437 12296 2468
rect 13633 2465 13645 2499
rect 13679 2496 13691 2499
rect 13679 2468 13860 2496
rect 13679 2465 13691 2468
rect 13633 2459 13691 2465
rect 12253 2431 12311 2437
rect 12253 2397 12265 2431
rect 12299 2397 12311 2431
rect 12253 2391 12311 2397
rect 13722 2388 13728 2440
rect 13780 2388 13786 2440
rect 13832 2428 13860 2468
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 14424 2468 15148 2496
rect 14424 2456 14430 2468
rect 14231 2433 14289 2439
rect 14231 2428 14243 2433
rect 13832 2400 14243 2428
rect 14231 2399 14243 2400
rect 14277 2399 14289 2433
rect 14231 2393 14289 2399
rect 14458 2388 14464 2440
rect 14516 2388 14522 2440
rect 9646 2332 9904 2360
rect 6512 2320 6518 2332
rect 10042 2320 10048 2372
rect 10100 2360 10106 2372
rect 15120 2360 15148 2468
rect 16114 2456 16120 2508
rect 16172 2456 16178 2508
rect 16206 2456 16212 2508
rect 16264 2496 16270 2508
rect 16853 2499 16911 2505
rect 16853 2496 16865 2499
rect 16264 2468 16865 2496
rect 16264 2456 16270 2468
rect 16853 2465 16865 2468
rect 16899 2465 16911 2499
rect 20530 2496 20536 2508
rect 16853 2459 16911 2465
rect 17512 2468 20536 2496
rect 16022 2388 16028 2440
rect 16080 2428 16086 2440
rect 16580 2431 16638 2437
rect 16580 2428 16592 2431
rect 16080 2400 16592 2428
rect 16080 2388 16086 2400
rect 16580 2397 16592 2400
rect 16626 2397 16638 2431
rect 16580 2391 16638 2397
rect 10100 2332 11284 2360
rect 15120 2332 16068 2360
rect 10100 2320 10106 2332
rect 5920 2264 6408 2292
rect 8846 2252 8852 2304
rect 8904 2292 8910 2304
rect 11149 2295 11207 2301
rect 11149 2292 11161 2295
rect 8904 2264 11161 2292
rect 8904 2252 8910 2264
rect 11149 2261 11161 2264
rect 11195 2261 11207 2295
rect 11256 2292 11284 2332
rect 14182 2292 14188 2304
rect 11256 2264 14188 2292
rect 11149 2255 11207 2261
rect 14182 2252 14188 2264
rect 14240 2252 14246 2304
rect 15749 2295 15807 2301
rect 15749 2261 15761 2295
rect 15795 2292 15807 2295
rect 15930 2292 15936 2304
rect 15795 2264 15936 2292
rect 15795 2261 15807 2264
rect 15749 2255 15807 2261
rect 15930 2252 15936 2264
rect 15988 2252 15994 2304
rect 16040 2292 16068 2332
rect 17512 2292 17540 2468
rect 20530 2456 20536 2468
rect 20588 2456 20594 2508
rect 20640 2496 20668 2604
rect 20809 2601 20821 2604
rect 20855 2632 20867 2635
rect 20898 2632 20904 2644
rect 20855 2604 20904 2632
rect 20855 2601 20867 2604
rect 20809 2595 20867 2601
rect 20898 2592 20904 2604
rect 20956 2592 20962 2644
rect 21542 2592 21548 2644
rect 21600 2632 21606 2644
rect 21735 2635 21793 2641
rect 21735 2632 21747 2635
rect 21600 2604 21747 2632
rect 21600 2592 21606 2604
rect 21735 2601 21747 2604
rect 21781 2601 21793 2635
rect 21735 2595 21793 2601
rect 24136 2604 25544 2632
rect 20717 2567 20775 2573
rect 20717 2533 20729 2567
rect 20763 2564 20775 2567
rect 20763 2536 21404 2564
rect 20763 2533 20775 2536
rect 20717 2527 20775 2533
rect 21376 2508 21404 2536
rect 23842 2524 23848 2576
rect 23900 2564 23906 2576
rect 24136 2564 24164 2604
rect 23900 2536 24164 2564
rect 25516 2564 25544 2604
rect 25958 2592 25964 2644
rect 26016 2592 26022 2644
rect 26605 2635 26663 2641
rect 26605 2632 26617 2635
rect 26068 2604 26617 2632
rect 26068 2564 26096 2604
rect 26605 2601 26617 2604
rect 26651 2601 26663 2635
rect 26605 2595 26663 2601
rect 27341 2635 27399 2641
rect 27341 2601 27353 2635
rect 27387 2601 27399 2635
rect 27341 2595 27399 2601
rect 25516 2536 26096 2564
rect 23900 2524 23906 2536
rect 21174 2496 21180 2508
rect 20640 2468 21180 2496
rect 21174 2456 21180 2468
rect 21232 2496 21238 2508
rect 21269 2499 21327 2505
rect 21269 2496 21281 2499
rect 21232 2468 21281 2496
rect 21232 2456 21238 2468
rect 21269 2465 21281 2468
rect 21315 2465 21327 2499
rect 21269 2459 21327 2465
rect 21358 2456 21364 2508
rect 21416 2456 21422 2508
rect 21652 2480 21772 2496
rect 21652 2468 21791 2480
rect 18325 2431 18383 2437
rect 18325 2397 18337 2431
rect 18371 2430 18383 2431
rect 18506 2430 18512 2440
rect 18371 2402 18512 2430
rect 18371 2397 18383 2402
rect 18325 2391 18383 2397
rect 18506 2388 18512 2402
rect 18564 2388 18570 2440
rect 18782 2388 18788 2440
rect 18840 2388 18846 2440
rect 19061 2431 19119 2437
rect 19061 2397 19073 2431
rect 19107 2428 19119 2431
rect 19242 2428 19248 2440
rect 19107 2400 19248 2428
rect 19107 2397 19119 2400
rect 19061 2391 19119 2397
rect 19242 2388 19248 2400
rect 19300 2388 19306 2440
rect 20441 2431 20499 2437
rect 20441 2397 20453 2431
rect 20487 2428 20499 2431
rect 21652 2428 21680 2468
rect 21744 2455 21791 2468
rect 23658 2456 23664 2508
rect 23716 2456 23722 2508
rect 23934 2456 23940 2508
rect 23992 2456 23998 2508
rect 24136 2505 24164 2536
rect 26234 2524 26240 2576
rect 26292 2564 26298 2576
rect 26513 2567 26571 2573
rect 26513 2564 26525 2567
rect 26292 2536 26525 2564
rect 26292 2524 26298 2536
rect 26513 2533 26525 2536
rect 26559 2564 26571 2567
rect 27356 2564 27384 2595
rect 27706 2592 27712 2644
rect 27764 2632 27770 2644
rect 28077 2635 28135 2641
rect 28077 2632 28089 2635
rect 27764 2604 28089 2632
rect 27764 2592 27770 2604
rect 28077 2601 28089 2604
rect 28123 2601 28135 2635
rect 28077 2595 28135 2601
rect 30006 2592 30012 2644
rect 30064 2592 30070 2644
rect 26559 2536 27384 2564
rect 26559 2533 26571 2536
rect 26513 2527 26571 2533
rect 24121 2499 24179 2505
rect 24121 2465 24133 2499
rect 24167 2496 24179 2499
rect 24210 2496 24216 2508
rect 24167 2468 24216 2496
rect 24167 2465 24179 2468
rect 24121 2459 24179 2465
rect 24210 2456 24216 2468
rect 24268 2456 24274 2508
rect 25314 2496 25320 2508
rect 24780 2468 25320 2496
rect 21744 2452 21823 2455
rect 20487 2400 21680 2428
rect 21763 2449 21823 2452
rect 21763 2418 21777 2449
rect 21765 2415 21777 2418
rect 21811 2415 21823 2449
rect 24617 2449 24675 2455
rect 24617 2446 24629 2449
rect 21765 2409 21823 2415
rect 20487 2397 20499 2400
rect 20441 2391 20499 2397
rect 22002 2388 22008 2440
rect 22060 2388 22066 2440
rect 24486 2437 24492 2440
rect 24448 2431 24492 2437
rect 24448 2397 24460 2431
rect 24448 2391 24492 2397
rect 24486 2388 24492 2391
rect 24544 2388 24550 2440
rect 24596 2415 24629 2446
rect 24663 2428 24675 2449
rect 24780 2428 24808 2468
rect 25314 2456 25320 2468
rect 25372 2456 25378 2508
rect 27249 2499 27307 2505
rect 27249 2465 27261 2499
rect 27295 2496 27307 2499
rect 27338 2496 27344 2508
rect 27295 2468 27344 2496
rect 27295 2465 27307 2468
rect 27249 2459 27307 2465
rect 27338 2456 27344 2468
rect 27396 2456 27402 2508
rect 27522 2456 27528 2508
rect 27580 2496 27586 2508
rect 27893 2499 27951 2505
rect 27893 2496 27905 2499
rect 27580 2468 27905 2496
rect 27580 2456 27586 2468
rect 24663 2415 24808 2428
rect 24596 2400 24808 2415
rect 24857 2431 24915 2437
rect 24857 2397 24869 2431
rect 24903 2428 24915 2431
rect 26418 2428 26424 2440
rect 24903 2400 26424 2428
rect 24903 2397 24915 2400
rect 24857 2391 24915 2397
rect 26418 2388 26424 2400
rect 26476 2388 26482 2440
rect 22922 2320 22928 2372
rect 22980 2360 22986 2372
rect 23477 2363 23535 2369
rect 23477 2360 23489 2363
rect 22980 2332 23489 2360
rect 22980 2320 22986 2332
rect 23477 2329 23489 2332
rect 23523 2329 23535 2363
rect 23477 2323 23535 2329
rect 16040 2264 17540 2292
rect 18141 2295 18199 2301
rect 18141 2261 18153 2295
rect 18187 2292 18199 2295
rect 18782 2292 18788 2304
rect 18187 2264 18788 2292
rect 18187 2261 18199 2264
rect 18141 2255 18199 2261
rect 18782 2252 18788 2264
rect 18840 2252 18846 2304
rect 20162 2252 20168 2304
rect 20220 2292 20226 2304
rect 21450 2292 21456 2304
rect 20220 2264 21456 2292
rect 20220 2252 20226 2264
rect 21450 2252 21456 2264
rect 21508 2252 21514 2304
rect 22186 2252 22192 2304
rect 22244 2292 22250 2304
rect 23109 2295 23167 2301
rect 23109 2292 23121 2295
rect 22244 2264 23121 2292
rect 22244 2252 22250 2264
rect 23109 2261 23121 2264
rect 23155 2261 23167 2295
rect 23109 2255 23167 2261
rect 23753 2295 23811 2301
rect 23753 2261 23765 2295
rect 23799 2292 23811 2295
rect 23842 2292 23848 2304
rect 23799 2264 23848 2292
rect 23799 2261 23811 2264
rect 23753 2255 23811 2261
rect 23842 2252 23848 2264
rect 23900 2252 23906 2304
rect 27816 2292 27844 2468
rect 27893 2465 27905 2468
rect 27939 2465 27951 2499
rect 27893 2459 27951 2465
rect 27982 2456 27988 2508
rect 28040 2496 28046 2508
rect 28169 2499 28227 2505
rect 28169 2496 28181 2499
rect 28040 2468 28181 2496
rect 28040 2456 28046 2468
rect 28169 2465 28181 2468
rect 28215 2465 28227 2499
rect 28169 2459 28227 2465
rect 28258 2456 28264 2508
rect 28316 2496 28322 2508
rect 28496 2499 28554 2505
rect 28496 2496 28508 2499
rect 28316 2468 28508 2496
rect 28316 2456 28322 2468
rect 28496 2465 28508 2468
rect 28542 2465 28554 2499
rect 28496 2459 28554 2465
rect 28902 2456 28908 2508
rect 28960 2456 28966 2508
rect 28632 2431 28690 2437
rect 28632 2428 28644 2431
rect 27908 2400 28644 2428
rect 27908 2372 27936 2400
rect 28632 2397 28644 2400
rect 28678 2397 28690 2431
rect 28632 2391 28690 2397
rect 27890 2320 27896 2372
rect 27948 2320 27954 2372
rect 29638 2292 29644 2304
rect 27816 2264 29644 2292
rect 29638 2252 29644 2264
rect 29696 2252 29702 2304
rect 552 2202 30912 2224
rect 552 2150 4193 2202
rect 4245 2150 4257 2202
rect 4309 2150 4321 2202
rect 4373 2150 4385 2202
rect 4437 2150 4449 2202
rect 4501 2150 11783 2202
rect 11835 2150 11847 2202
rect 11899 2150 11911 2202
rect 11963 2150 11975 2202
rect 12027 2150 12039 2202
rect 12091 2150 19373 2202
rect 19425 2150 19437 2202
rect 19489 2150 19501 2202
rect 19553 2150 19565 2202
rect 19617 2150 19629 2202
rect 19681 2150 26963 2202
rect 27015 2150 27027 2202
rect 27079 2150 27091 2202
rect 27143 2150 27155 2202
rect 27207 2150 27219 2202
rect 27271 2150 30912 2202
rect 552 2128 30912 2150
rect 2961 2091 3019 2097
rect 2961 2057 2973 2091
rect 3007 2088 3019 2091
rect 3326 2088 3332 2100
rect 3007 2060 3332 2088
rect 3007 2057 3019 2060
rect 2961 2051 3019 2057
rect 3326 2048 3332 2060
rect 3384 2048 3390 2100
rect 5534 2048 5540 2100
rect 5592 2048 5598 2100
rect 7837 2091 7895 2097
rect 5828 2060 7788 2088
rect 3234 1980 3240 2032
rect 3292 1980 3298 2032
rect 5258 1980 5264 2032
rect 5316 2020 5322 2032
rect 5828 2020 5856 2060
rect 5316 1992 5856 2020
rect 5316 1980 5322 1992
rect 1486 1952 1492 1964
rect 1418 1937 1492 1952
rect 1418 1906 1445 1937
rect 1433 1903 1445 1906
rect 1479 1912 1492 1937
rect 1544 1912 1550 1964
rect 1670 1912 1676 1964
rect 1728 1912 1734 1964
rect 3513 1955 3571 1961
rect 3513 1921 3525 1955
rect 3559 1921 3571 1955
rect 3513 1915 3571 1921
rect 1479 1903 1491 1912
rect 1433 1897 1491 1903
rect 937 1887 995 1893
rect 937 1853 949 1887
rect 983 1884 995 1887
rect 1302 1884 1308 1896
rect 983 1856 1308 1884
rect 983 1853 995 1856
rect 937 1847 995 1853
rect 1302 1844 1308 1856
rect 1360 1844 1366 1896
rect 3418 1844 3424 1896
rect 3476 1844 3482 1896
rect 3528 1884 3556 1915
rect 3970 1912 3976 1964
rect 4028 1912 4034 1964
rect 6178 1961 6184 1964
rect 6140 1955 6184 1961
rect 6140 1952 6152 1955
rect 4178 1924 6152 1952
rect 3602 1884 3608 1896
rect 3528 1856 3608 1884
rect 3602 1844 3608 1856
rect 3660 1844 3666 1896
rect 3840 1887 3898 1893
rect 3840 1853 3852 1887
rect 3886 1884 3898 1887
rect 4178 1884 4206 1924
rect 6140 1921 6152 1924
rect 6140 1915 6184 1921
rect 6178 1912 6184 1915
rect 6236 1912 6242 1964
rect 6276 1953 6334 1959
rect 6276 1919 6288 1953
rect 6322 1952 6334 1953
rect 6362 1952 6368 1964
rect 6322 1924 6368 1952
rect 6322 1919 6334 1924
rect 6276 1913 6334 1919
rect 6362 1912 6368 1924
rect 6420 1912 6426 1964
rect 6549 1955 6607 1961
rect 6549 1921 6561 1955
rect 6595 1952 6607 1955
rect 7282 1952 7288 1964
rect 6595 1924 7288 1952
rect 6595 1921 6607 1924
rect 6549 1915 6607 1921
rect 7282 1912 7288 1924
rect 7340 1912 7346 1964
rect 7760 1952 7788 2060
rect 7837 2057 7849 2091
rect 7883 2088 7895 2091
rect 8202 2088 8208 2100
rect 7883 2060 8208 2088
rect 7883 2057 7895 2060
rect 7837 2051 7895 2057
rect 8202 2048 8208 2060
rect 8260 2048 8266 2100
rect 10870 2088 10876 2100
rect 9048 2060 10876 2088
rect 8021 2023 8079 2029
rect 8021 1989 8033 2023
rect 8067 2020 8079 2023
rect 9048 2020 9076 2060
rect 10870 2048 10876 2060
rect 10928 2048 10934 2100
rect 11146 2048 11152 2100
rect 11204 2088 11210 2100
rect 12158 2088 12164 2100
rect 11204 2060 12164 2088
rect 11204 2048 11210 2060
rect 12158 2048 12164 2060
rect 12216 2048 12222 2100
rect 13170 2048 13176 2100
rect 13228 2088 13234 2100
rect 16758 2088 16764 2100
rect 13228 2060 16764 2088
rect 13228 2048 13234 2060
rect 16758 2048 16764 2060
rect 16816 2048 16822 2100
rect 17865 2091 17923 2097
rect 17865 2057 17877 2091
rect 17911 2088 17923 2091
rect 17954 2088 17960 2100
rect 17911 2060 17960 2088
rect 17911 2057 17923 2060
rect 17865 2051 17923 2057
rect 17954 2048 17960 2060
rect 18012 2048 18018 2100
rect 20714 2088 20720 2100
rect 18708 2060 20720 2088
rect 8067 1992 9076 2020
rect 18049 2023 18107 2029
rect 8067 1989 8079 1992
rect 8021 1983 8079 1989
rect 18049 1989 18061 2023
rect 18095 1989 18107 2023
rect 18049 1983 18107 1989
rect 7760 1924 8624 1952
rect 3886 1856 4206 1884
rect 4249 1887 4307 1893
rect 3886 1853 3898 1856
rect 3840 1847 3898 1853
rect 4249 1853 4261 1887
rect 4295 1884 4307 1887
rect 5718 1884 5724 1896
rect 4295 1856 5724 1884
rect 4295 1853 4307 1856
rect 4249 1847 4307 1853
rect 5718 1844 5724 1856
rect 5776 1844 5782 1896
rect 5810 1844 5816 1896
rect 5868 1844 5874 1896
rect 5902 1844 5908 1896
rect 5960 1884 5966 1896
rect 8205 1887 8263 1893
rect 8205 1884 8217 1887
rect 5960 1856 8217 1884
rect 5960 1844 5966 1856
rect 8205 1853 8217 1856
rect 8251 1884 8263 1887
rect 8294 1884 8300 1896
rect 8251 1856 8300 1884
rect 8251 1853 8263 1856
rect 8205 1847 8263 1853
rect 8294 1844 8300 1856
rect 8352 1844 8358 1896
rect 8596 1884 8624 1924
rect 8846 1912 8852 1964
rect 8904 1952 8910 1964
rect 9033 1955 9091 1961
rect 9033 1952 9045 1955
rect 8904 1924 9045 1952
rect 8904 1912 8910 1924
rect 9033 1921 9045 1924
rect 9079 1921 9091 1955
rect 9033 1915 9091 1921
rect 9496 1953 9554 1959
rect 9496 1919 9508 1953
rect 9542 1919 9554 1953
rect 9496 1913 9554 1919
rect 8662 1884 8668 1896
rect 8596 1856 8668 1884
rect 8662 1844 8668 1856
rect 8720 1884 8726 1896
rect 8941 1887 8999 1893
rect 8941 1884 8953 1887
rect 8720 1856 8953 1884
rect 8720 1844 8726 1856
rect 8941 1853 8953 1856
rect 8987 1853 8999 1887
rect 9514 1884 9542 1913
rect 9582 1912 9588 1964
rect 9640 1952 9646 1964
rect 9769 1955 9827 1961
rect 9769 1952 9781 1955
rect 9640 1924 9781 1952
rect 9640 1912 9646 1924
rect 9769 1921 9781 1924
rect 9815 1921 9827 1955
rect 9769 1915 9827 1921
rect 11149 1955 11207 1961
rect 11149 1921 11161 1955
rect 11195 1952 11207 1955
rect 11704 1955 11762 1961
rect 11704 1952 11716 1955
rect 11195 1924 11716 1952
rect 11195 1921 11207 1924
rect 11149 1915 11207 1921
rect 11704 1921 11716 1924
rect 11750 1921 11762 1955
rect 12342 1952 12348 1964
rect 11704 1915 11762 1921
rect 11808 1924 12348 1952
rect 8941 1847 8999 1853
rect 9146 1880 9447 1884
rect 9511 1880 9542 1884
rect 9146 1856 9542 1880
rect 1403 1751 1461 1757
rect 1403 1717 1415 1751
rect 1449 1748 1461 1751
rect 1670 1748 1676 1760
rect 1449 1720 1676 1748
rect 1449 1717 1461 1720
rect 1403 1711 1461 1717
rect 1670 1708 1676 1720
rect 1728 1708 1734 1760
rect 3620 1748 3648 1844
rect 5828 1816 5856 1844
rect 9146 1816 9174 1856
rect 9419 1852 9539 1856
rect 10778 1844 10784 1896
rect 10836 1884 10842 1896
rect 11054 1884 11060 1896
rect 10836 1856 11060 1884
rect 10836 1844 10842 1856
rect 11054 1844 11060 1856
rect 11112 1884 11118 1896
rect 11241 1887 11299 1893
rect 11241 1884 11253 1887
rect 11112 1856 11253 1884
rect 11112 1844 11118 1856
rect 11241 1853 11253 1856
rect 11287 1853 11299 1887
rect 11241 1847 11299 1853
rect 11514 1844 11520 1896
rect 11572 1884 11578 1896
rect 11808 1884 11836 1924
rect 12342 1912 12348 1924
rect 12400 1912 12406 1964
rect 13357 1955 13415 1961
rect 13357 1921 13369 1955
rect 13403 1952 13415 1955
rect 14096 1955 14154 1961
rect 14096 1952 14108 1955
rect 13403 1924 14108 1952
rect 13403 1921 13415 1924
rect 13357 1915 13415 1921
rect 14096 1921 14108 1924
rect 14142 1921 14154 1955
rect 14096 1915 14154 1921
rect 14182 1912 14188 1964
rect 14240 1952 14246 1964
rect 14369 1955 14427 1961
rect 14369 1952 14381 1955
rect 14240 1924 14381 1952
rect 14240 1912 14246 1924
rect 14369 1921 14381 1924
rect 14415 1921 14427 1955
rect 14369 1915 14427 1921
rect 15749 1955 15807 1961
rect 15749 1921 15761 1955
rect 15795 1952 15807 1955
rect 16304 1955 16362 1961
rect 16304 1952 16316 1955
rect 15795 1924 16316 1952
rect 15795 1921 15807 1924
rect 15749 1915 15807 1921
rect 16304 1921 16316 1924
rect 16350 1921 16362 1955
rect 16304 1915 16362 1921
rect 16577 1955 16635 1961
rect 16577 1921 16589 1955
rect 16623 1952 16635 1955
rect 18064 1952 18092 1983
rect 18322 1980 18328 2032
rect 18380 2020 18386 2032
rect 18708 2020 18736 2060
rect 20714 2048 20720 2060
rect 20772 2048 20778 2100
rect 21082 2048 21088 2100
rect 21140 2088 21146 2100
rect 21140 2060 22330 2088
rect 21140 2048 21146 2060
rect 18380 1992 18736 2020
rect 22302 2020 22330 2060
rect 22370 2048 22376 2100
rect 22428 2088 22434 2100
rect 23385 2091 23443 2097
rect 23385 2088 23397 2091
rect 22428 2060 23397 2088
rect 22428 2048 22434 2060
rect 23385 2057 23397 2060
rect 23431 2057 23443 2091
rect 23385 2051 23443 2057
rect 23474 2048 23480 2100
rect 23532 2088 23538 2100
rect 28169 2091 28227 2097
rect 28169 2088 28181 2091
rect 23532 2060 28181 2088
rect 23532 2048 23538 2060
rect 28169 2057 28181 2060
rect 28215 2057 28227 2091
rect 28169 2051 28227 2057
rect 28718 2048 28724 2100
rect 28776 2048 28782 2100
rect 23658 2020 23664 2032
rect 22302 1992 23664 2020
rect 18380 1980 18386 1992
rect 16623 1924 18092 1952
rect 16623 1921 16635 1924
rect 16577 1915 16635 1921
rect 11572 1856 11836 1884
rect 11572 1844 11578 1856
rect 11882 1844 11888 1896
rect 11940 1884 11946 1896
rect 11977 1887 12035 1893
rect 11977 1884 11989 1887
rect 11940 1856 11989 1884
rect 11940 1844 11946 1856
rect 11977 1853 11989 1856
rect 12023 1853 12035 1887
rect 11977 1847 12035 1853
rect 13633 1887 13691 1893
rect 13633 1853 13645 1887
rect 13679 1884 13691 1887
rect 13722 1884 13728 1896
rect 13679 1856 13728 1884
rect 13679 1853 13691 1856
rect 13633 1847 13691 1853
rect 13722 1844 13728 1856
rect 13780 1844 13786 1896
rect 13998 1893 14004 1896
rect 13960 1887 14004 1893
rect 13960 1853 13972 1887
rect 13960 1847 14004 1853
rect 13998 1844 14004 1847
rect 14056 1844 14062 1896
rect 15841 1887 15899 1893
rect 15841 1853 15853 1887
rect 15887 1884 15899 1887
rect 16114 1884 16120 1896
rect 15887 1856 16120 1884
rect 15887 1853 15899 1856
rect 15841 1847 15899 1853
rect 16114 1844 16120 1856
rect 16172 1844 16178 1896
rect 18230 1844 18236 1896
rect 18288 1844 18294 1896
rect 18524 1893 18552 1992
rect 18598 1912 18604 1964
rect 18656 1952 18662 1964
rect 18693 1955 18751 1961
rect 18693 1952 18705 1955
rect 18656 1924 18705 1952
rect 18656 1912 18662 1924
rect 18693 1921 18705 1924
rect 18739 1921 18751 1955
rect 19156 1955 19214 1961
rect 19156 1952 19168 1955
rect 18693 1915 18751 1921
rect 18800 1924 19168 1952
rect 18509 1887 18567 1893
rect 18509 1853 18521 1887
rect 18555 1853 18567 1887
rect 18509 1847 18567 1853
rect 5644 1788 5856 1816
rect 8956 1788 9174 1816
rect 5644 1748 5672 1788
rect 8956 1760 8984 1788
rect 18138 1776 18144 1828
rect 18196 1816 18202 1828
rect 18800 1816 18828 1924
rect 19156 1921 19168 1924
rect 19202 1921 19214 1955
rect 19156 1915 19214 1921
rect 20809 1955 20867 1961
rect 20809 1921 20821 1955
rect 20855 1950 20867 1955
rect 21364 1955 21422 1961
rect 21364 1952 21376 1955
rect 21008 1950 21376 1952
rect 20855 1924 21376 1950
rect 20855 1922 21036 1924
rect 20855 1921 20867 1922
rect 20809 1915 20867 1921
rect 21364 1921 21376 1924
rect 21410 1921 21422 1955
rect 21364 1915 21422 1921
rect 21450 1912 21456 1964
rect 21508 1912 21514 1964
rect 21637 1955 21695 1961
rect 21637 1921 21649 1955
rect 21683 1952 21695 1955
rect 23474 1952 23480 1964
rect 21683 1924 23480 1952
rect 21683 1921 21695 1924
rect 21637 1915 21695 1921
rect 23474 1912 23480 1924
rect 23532 1912 23538 1964
rect 19429 1887 19487 1893
rect 19429 1853 19441 1887
rect 19475 1884 19487 1887
rect 20438 1884 20444 1896
rect 19475 1856 20444 1884
rect 19475 1853 19487 1856
rect 19429 1847 19487 1853
rect 20438 1844 20444 1856
rect 20496 1844 20502 1896
rect 20927 1887 20985 1893
rect 20927 1853 20939 1887
rect 20973 1884 20985 1887
rect 21174 1884 21180 1896
rect 20973 1856 21180 1884
rect 20973 1853 20985 1856
rect 20927 1847 20985 1853
rect 21174 1844 21180 1856
rect 21232 1844 21238 1896
rect 21468 1884 21496 1912
rect 22646 1884 22652 1896
rect 21468 1856 22652 1884
rect 22646 1844 22652 1856
rect 22704 1884 22710 1896
rect 23584 1893 23612 1992
rect 23658 1980 23664 1992
rect 23716 1980 23722 2032
rect 26050 1980 26056 2032
rect 26108 2020 26114 2032
rect 26108 1992 26372 2020
rect 26108 1980 26114 1992
rect 24308 1955 24366 1961
rect 24308 1952 24320 1955
rect 24228 1924 24320 1952
rect 23293 1887 23351 1893
rect 23293 1884 23305 1887
rect 22704 1856 23305 1884
rect 22704 1844 22710 1856
rect 23293 1853 23305 1856
rect 23339 1853 23351 1887
rect 23293 1847 23351 1853
rect 23569 1887 23627 1893
rect 23569 1853 23581 1887
rect 23615 1853 23627 1887
rect 23750 1884 23756 1896
rect 23569 1847 23627 1853
rect 23676 1856 23756 1884
rect 18196 1788 18828 1816
rect 18196 1776 18202 1788
rect 23014 1776 23020 1828
rect 23072 1776 23078 1828
rect 23676 1816 23704 1856
rect 23750 1844 23756 1856
rect 23808 1884 23814 1896
rect 23845 1887 23903 1893
rect 23845 1884 23857 1887
rect 23808 1856 23857 1884
rect 23808 1844 23814 1856
rect 23845 1853 23857 1856
rect 23891 1853 23903 1887
rect 24228 1884 24256 1924
rect 24308 1921 24320 1924
rect 24354 1921 24366 1955
rect 24308 1915 24366 1921
rect 26234 1912 26240 1964
rect 26292 1912 26298 1964
rect 26344 1952 26372 1992
rect 26792 1955 26850 1961
rect 26792 1952 26804 1955
rect 26344 1924 26804 1952
rect 26792 1921 26804 1924
rect 26838 1921 26850 1955
rect 26792 1915 26850 1921
rect 26970 1912 26976 1964
rect 27028 1952 27034 1964
rect 27065 1955 27123 1961
rect 27065 1952 27077 1955
rect 27028 1924 27077 1952
rect 27028 1912 27034 1924
rect 27065 1921 27077 1924
rect 27111 1921 27123 1955
rect 27065 1915 27123 1921
rect 27172 1924 29040 1952
rect 23845 1847 23903 1853
rect 23971 1856 24256 1884
rect 24581 1887 24639 1893
rect 23971 1816 23999 1856
rect 24581 1853 24593 1887
rect 24627 1884 24639 1887
rect 26050 1884 26056 1896
rect 24627 1856 26056 1884
rect 24627 1853 24639 1856
rect 24581 1847 24639 1853
rect 26050 1844 26056 1856
rect 26108 1844 26114 1896
rect 26252 1884 26280 1912
rect 26329 1887 26387 1893
rect 26329 1884 26341 1887
rect 26252 1856 26341 1884
rect 26329 1853 26341 1856
rect 26375 1853 26387 1887
rect 26329 1847 26387 1853
rect 26418 1844 26424 1896
rect 26476 1884 26482 1896
rect 27172 1884 27200 1924
rect 29012 1893 29040 1924
rect 29270 1912 29276 1964
rect 29328 1912 29334 1964
rect 29546 1912 29552 1964
rect 29604 1912 29610 1964
rect 28537 1887 28595 1893
rect 28537 1884 28549 1887
rect 26476 1856 27200 1884
rect 27724 1856 28549 1884
rect 26476 1844 26482 1856
rect 23584 1788 23704 1816
rect 23768 1788 23999 1816
rect 23584 1760 23612 1788
rect 23768 1760 23796 1788
rect 27724 1760 27752 1856
rect 28537 1853 28549 1856
rect 28583 1853 28595 1887
rect 28537 1847 28595 1853
rect 28997 1887 29055 1893
rect 28997 1853 29009 1887
rect 29043 1884 29055 1887
rect 29288 1884 29316 1912
rect 29043 1856 29316 1884
rect 29043 1853 29055 1856
rect 28997 1847 29055 1853
rect 28552 1816 28580 1847
rect 29564 1816 29592 1912
rect 28552 1788 29592 1816
rect 3620 1720 5672 1748
rect 8481 1751 8539 1757
rect 8481 1717 8493 1751
rect 8527 1748 8539 1751
rect 8662 1748 8668 1760
rect 8527 1720 8668 1748
rect 8527 1717 8539 1720
rect 8481 1711 8539 1717
rect 8662 1708 8668 1720
rect 8720 1708 8726 1760
rect 8754 1708 8760 1760
rect 8812 1708 8818 1760
rect 8938 1708 8944 1760
rect 8996 1708 9002 1760
rect 9398 1708 9404 1760
rect 9456 1748 9462 1760
rect 9499 1751 9557 1757
rect 9499 1748 9511 1751
rect 9456 1720 9511 1748
rect 9456 1708 9462 1720
rect 9499 1717 9511 1720
rect 9545 1717 9557 1751
rect 9499 1711 9557 1717
rect 10870 1708 10876 1760
rect 10928 1748 10934 1760
rect 11698 1748 11704 1760
rect 11756 1757 11762 1760
rect 10928 1720 11704 1748
rect 10928 1708 10934 1720
rect 11698 1708 11704 1720
rect 11756 1711 11765 1757
rect 11756 1708 11762 1711
rect 11882 1708 11888 1760
rect 11940 1748 11946 1760
rect 13630 1748 13636 1760
rect 11940 1720 13636 1748
rect 11940 1708 11946 1720
rect 13630 1708 13636 1720
rect 13688 1708 13694 1760
rect 16307 1751 16365 1757
rect 16307 1717 16319 1751
rect 16353 1748 16365 1751
rect 16574 1748 16580 1760
rect 16353 1720 16580 1748
rect 16353 1717 16365 1720
rect 16307 1711 16365 1717
rect 16574 1708 16580 1720
rect 16632 1708 16638 1760
rect 17954 1708 17960 1760
rect 18012 1748 18018 1760
rect 18325 1751 18383 1757
rect 18325 1748 18337 1751
rect 18012 1720 18337 1748
rect 18012 1708 18018 1720
rect 18325 1717 18337 1720
rect 18371 1717 18383 1751
rect 18325 1711 18383 1717
rect 18966 1708 18972 1760
rect 19024 1748 19030 1760
rect 19159 1751 19217 1757
rect 19159 1748 19171 1751
rect 19024 1720 19171 1748
rect 19024 1708 19030 1720
rect 19159 1717 19171 1720
rect 19205 1717 19217 1751
rect 19159 1711 19217 1717
rect 19334 1708 19340 1760
rect 19392 1748 19398 1760
rect 20806 1748 20812 1760
rect 19392 1720 20812 1748
rect 19392 1708 19398 1720
rect 20806 1708 20812 1720
rect 20864 1708 20870 1760
rect 21367 1751 21425 1757
rect 21367 1717 21379 1751
rect 21413 1748 21425 1751
rect 21542 1748 21548 1760
rect 21413 1720 21548 1748
rect 21413 1717 21425 1720
rect 21367 1711 21425 1717
rect 21542 1708 21548 1720
rect 21600 1708 21606 1760
rect 22830 1708 22836 1760
rect 22888 1748 22894 1760
rect 23109 1751 23167 1757
rect 23109 1748 23121 1751
rect 22888 1720 23121 1748
rect 22888 1708 22894 1720
rect 23109 1717 23121 1720
rect 23155 1717 23167 1751
rect 23109 1711 23167 1717
rect 23566 1708 23572 1760
rect 23624 1708 23630 1760
rect 23750 1708 23756 1760
rect 23808 1708 23814 1760
rect 23934 1708 23940 1760
rect 23992 1748 23998 1760
rect 24118 1748 24124 1760
rect 23992 1720 24124 1748
rect 23992 1708 23998 1720
rect 24118 1708 24124 1720
rect 24176 1748 24182 1760
rect 24311 1751 24369 1757
rect 24311 1748 24323 1751
rect 24176 1720 24323 1748
rect 24176 1708 24182 1720
rect 24311 1717 24323 1720
rect 24357 1717 24369 1751
rect 24311 1711 24369 1717
rect 24854 1708 24860 1760
rect 24912 1748 24918 1760
rect 25685 1751 25743 1757
rect 25685 1748 25697 1751
rect 24912 1720 25697 1748
rect 24912 1708 24918 1720
rect 25685 1717 25697 1720
rect 25731 1717 25743 1751
rect 25685 1711 25743 1717
rect 26326 1708 26332 1760
rect 26384 1748 26390 1760
rect 26602 1748 26608 1760
rect 26384 1720 26608 1748
rect 26384 1708 26390 1720
rect 26602 1708 26608 1720
rect 26660 1748 26666 1760
rect 26795 1751 26853 1757
rect 26795 1748 26807 1751
rect 26660 1720 26807 1748
rect 26660 1708 26666 1720
rect 26795 1717 26807 1720
rect 26841 1717 26853 1751
rect 26795 1711 26853 1717
rect 26970 1708 26976 1760
rect 27028 1748 27034 1760
rect 27522 1748 27528 1760
rect 27028 1720 27528 1748
rect 27028 1708 27034 1720
rect 27522 1708 27528 1720
rect 27580 1708 27586 1760
rect 27706 1708 27712 1760
rect 27764 1708 27770 1760
rect 29178 1708 29184 1760
rect 29236 1708 29242 1760
rect 552 1658 31072 1680
rect 552 1606 7988 1658
rect 8040 1606 8052 1658
rect 8104 1606 8116 1658
rect 8168 1606 8180 1658
rect 8232 1606 8244 1658
rect 8296 1606 15578 1658
rect 15630 1606 15642 1658
rect 15694 1606 15706 1658
rect 15758 1606 15770 1658
rect 15822 1606 15834 1658
rect 15886 1606 23168 1658
rect 23220 1606 23232 1658
rect 23284 1606 23296 1658
rect 23348 1606 23360 1658
rect 23412 1606 23424 1658
rect 23476 1606 30758 1658
rect 30810 1606 30822 1658
rect 30874 1606 30886 1658
rect 30938 1606 30950 1658
rect 31002 1606 31014 1658
rect 31066 1606 31072 1658
rect 552 1584 31072 1606
rect 845 1547 903 1553
rect 845 1513 857 1547
rect 891 1544 903 1547
rect 1210 1544 1216 1556
rect 891 1516 1216 1544
rect 891 1513 903 1516
rect 845 1507 903 1513
rect 1210 1504 1216 1516
rect 1268 1504 1274 1556
rect 1762 1504 1768 1556
rect 1820 1544 1826 1556
rect 3329 1547 3387 1553
rect 1820 1516 2912 1544
rect 1820 1504 1826 1516
rect 1029 1411 1087 1417
rect 1029 1377 1041 1411
rect 1075 1377 1087 1411
rect 2884 1408 2912 1516
rect 3329 1513 3341 1547
rect 3375 1544 3387 1547
rect 3878 1544 3884 1556
rect 3375 1516 3884 1544
rect 3375 1513 3387 1516
rect 3329 1507 3387 1513
rect 3878 1504 3884 1516
rect 3936 1504 3942 1556
rect 3979 1547 4037 1553
rect 3979 1513 3991 1547
rect 4025 1544 4037 1547
rect 4522 1544 4528 1556
rect 4025 1516 4528 1544
rect 4025 1513 4037 1516
rect 3979 1507 4037 1513
rect 4522 1504 4528 1516
rect 4580 1504 4586 1556
rect 6914 1504 6920 1556
rect 6972 1553 6978 1556
rect 6972 1544 6981 1553
rect 8481 1547 8539 1553
rect 6972 1516 7017 1544
rect 6972 1507 6981 1516
rect 8481 1513 8493 1547
rect 8527 1544 8539 1547
rect 8938 1544 8944 1556
rect 8527 1516 8944 1544
rect 8527 1513 8539 1516
rect 8481 1507 8539 1513
rect 6972 1504 6978 1507
rect 8938 1504 8944 1516
rect 8996 1504 9002 1556
rect 9131 1547 9189 1553
rect 9131 1513 9143 1547
rect 9177 1544 9189 1547
rect 10870 1544 10876 1556
rect 9177 1516 10876 1544
rect 9177 1513 9189 1516
rect 9131 1507 9189 1513
rect 10870 1504 10876 1516
rect 10928 1504 10934 1556
rect 10962 1504 10968 1556
rect 11020 1504 11026 1556
rect 11054 1504 11060 1556
rect 11112 1544 11118 1556
rect 11241 1547 11299 1553
rect 11241 1544 11253 1547
rect 11112 1516 11253 1544
rect 11112 1504 11118 1516
rect 11241 1513 11253 1516
rect 11287 1513 11299 1547
rect 11241 1507 11299 1513
rect 11983 1547 12041 1553
rect 11983 1513 11995 1547
rect 12029 1544 12041 1547
rect 13814 1544 13820 1556
rect 12029 1516 13820 1544
rect 12029 1513 12041 1516
rect 11983 1507 12041 1513
rect 13814 1504 13820 1516
rect 13872 1504 13878 1556
rect 13998 1504 14004 1556
rect 14056 1544 14062 1556
rect 14191 1547 14249 1553
rect 14191 1544 14203 1547
rect 14056 1516 14203 1544
rect 14056 1504 14062 1516
rect 14191 1513 14203 1516
rect 14237 1513 14249 1547
rect 14191 1507 14249 1513
rect 15749 1547 15807 1553
rect 15749 1513 15761 1547
rect 15795 1544 15807 1547
rect 16022 1544 16028 1556
rect 15795 1516 16028 1544
rect 15795 1513 15807 1516
rect 15749 1507 15807 1513
rect 16022 1504 16028 1516
rect 16080 1504 16086 1556
rect 16574 1504 16580 1556
rect 16632 1553 16638 1556
rect 16632 1544 16641 1553
rect 16632 1516 16677 1544
rect 16632 1507 16641 1516
rect 16632 1504 16638 1507
rect 18138 1504 18144 1556
rect 18196 1504 18202 1556
rect 18791 1547 18849 1553
rect 18791 1513 18803 1547
rect 18837 1544 18849 1547
rect 18966 1544 18972 1556
rect 18837 1516 18972 1544
rect 18837 1513 18849 1516
rect 18791 1507 18849 1513
rect 18966 1504 18972 1516
rect 19024 1504 19030 1556
rect 20990 1544 20996 1556
rect 20088 1516 20996 1544
rect 10502 1436 10508 1488
rect 10560 1476 10566 1488
rect 10781 1479 10839 1485
rect 10560 1448 10732 1476
rect 10560 1436 10566 1448
rect 5813 1411 5871 1417
rect 1029 1371 1087 1377
rect 1964 1380 2176 1408
rect 2884 1380 4844 1408
rect 1044 1204 1072 1371
rect 1302 1300 1308 1352
rect 1360 1300 1366 1352
rect 1670 1349 1676 1352
rect 1632 1343 1676 1349
rect 1632 1309 1644 1343
rect 1632 1303 1676 1309
rect 1670 1300 1676 1303
rect 1728 1300 1734 1352
rect 1811 1343 1869 1349
rect 1811 1309 1823 1343
rect 1857 1340 1869 1343
rect 1964 1340 1992 1380
rect 1857 1312 1992 1340
rect 1857 1309 1869 1312
rect 1811 1303 1869 1309
rect 2038 1300 2044 1352
rect 2096 1300 2102 1352
rect 2148 1340 2176 1380
rect 2148 1312 2774 1340
rect 2498 1204 2504 1216
rect 1044 1176 2504 1204
rect 2498 1164 2504 1176
rect 2556 1164 2562 1216
rect 2746 1204 2774 1312
rect 3510 1300 3516 1352
rect 3568 1300 3574 1352
rect 3970 1300 3976 1352
rect 4028 1351 4034 1352
rect 4028 1345 4067 1351
rect 4055 1311 4067 1345
rect 4028 1305 4067 1311
rect 4249 1343 4307 1349
rect 4249 1309 4261 1343
rect 4295 1340 4307 1343
rect 4706 1340 4712 1352
rect 4295 1312 4712 1340
rect 4295 1309 4307 1312
rect 4028 1300 4034 1305
rect 4249 1303 4307 1309
rect 4706 1300 4712 1312
rect 4764 1300 4770 1352
rect 4816 1340 4844 1380
rect 5813 1377 5825 1411
rect 5859 1408 5871 1411
rect 6822 1408 6828 1420
rect 5859 1380 6828 1408
rect 5859 1377 5871 1380
rect 5813 1371 5871 1377
rect 6822 1368 6828 1380
rect 6880 1368 6886 1420
rect 8754 1368 8760 1420
rect 8812 1408 8818 1420
rect 9401 1411 9459 1417
rect 9401 1408 9413 1411
rect 8812 1380 9413 1408
rect 8812 1368 8818 1380
rect 9401 1377 9413 1380
rect 9447 1377 9459 1411
rect 9401 1371 9459 1377
rect 9490 1368 9496 1420
rect 9548 1408 9554 1420
rect 10704 1408 10732 1448
rect 10781 1445 10793 1479
rect 10827 1476 10839 1479
rect 10827 1448 11284 1476
rect 10827 1445 10839 1448
rect 10781 1439 10839 1445
rect 11149 1411 11207 1417
rect 11149 1408 11161 1411
rect 9548 1380 9674 1408
rect 10704 1380 11161 1408
rect 9548 1368 9554 1380
rect 6953 1361 7011 1367
rect 6953 1358 6965 1361
rect 5997 1343 6055 1349
rect 5997 1340 6009 1343
rect 4816 1312 6009 1340
rect 5997 1309 6009 1312
rect 6043 1309 6055 1343
rect 5997 1303 6055 1309
rect 6454 1300 6460 1352
rect 6512 1300 6518 1352
rect 6932 1327 6965 1358
rect 6999 1352 7011 1361
rect 6999 1327 7012 1352
rect 6932 1312 7012 1327
rect 7006 1300 7012 1312
rect 7064 1300 7070 1352
rect 7190 1300 7196 1352
rect 7248 1300 7254 1352
rect 8665 1343 8723 1349
rect 8665 1309 8677 1343
rect 8711 1309 8723 1343
rect 8665 1303 8723 1309
rect 5537 1275 5595 1281
rect 5537 1241 5549 1275
rect 5583 1272 5595 1275
rect 6362 1272 6368 1284
rect 5583 1244 6368 1272
rect 5583 1241 5595 1244
rect 5537 1235 5595 1241
rect 6362 1232 6368 1244
rect 6420 1232 6426 1284
rect 5074 1204 5080 1216
rect 2746 1176 5080 1204
rect 5074 1164 5080 1176
rect 5132 1164 5138 1216
rect 5718 1164 5724 1216
rect 5776 1204 5782 1216
rect 7558 1204 7564 1216
rect 5776 1176 7564 1204
rect 5776 1164 5782 1176
rect 7558 1164 7564 1176
rect 7616 1164 7622 1216
rect 8680 1204 8708 1303
rect 9122 1300 9128 1352
rect 9180 1300 9186 1352
rect 9646 1340 9674 1380
rect 11149 1377 11161 1380
rect 11195 1377 11207 1411
rect 11149 1371 11207 1377
rect 9646 1312 10916 1340
rect 10778 1204 10784 1216
rect 8680 1176 10784 1204
rect 10778 1164 10784 1176
rect 10836 1164 10842 1216
rect 10888 1204 10916 1312
rect 11256 1272 11284 1448
rect 18230 1436 18236 1488
rect 18288 1436 18294 1488
rect 11330 1368 11336 1420
rect 11388 1408 11394 1420
rect 11425 1411 11483 1417
rect 11425 1408 11437 1411
rect 11388 1380 11437 1408
rect 11388 1368 11394 1380
rect 11425 1377 11437 1380
rect 11471 1377 11483 1411
rect 11425 1371 11483 1377
rect 11606 1368 11612 1420
rect 11664 1408 11670 1420
rect 11664 1380 13860 1408
rect 11664 1368 11670 1380
rect 11517 1343 11575 1349
rect 11517 1309 11529 1343
rect 11563 1340 11575 1343
rect 11882 1340 11888 1352
rect 11563 1312 11888 1340
rect 11563 1309 11575 1312
rect 11517 1303 11575 1309
rect 11882 1300 11888 1312
rect 11940 1300 11946 1352
rect 12023 1343 12081 1349
rect 12023 1309 12035 1343
rect 12069 1340 12081 1343
rect 12158 1340 12164 1352
rect 12069 1312 12164 1340
rect 12069 1309 12081 1312
rect 12023 1303 12081 1309
rect 12158 1300 12164 1312
rect 12216 1300 12222 1352
rect 12253 1343 12311 1349
rect 12253 1309 12265 1343
rect 12299 1340 12311 1343
rect 12299 1312 13676 1340
rect 12299 1309 12311 1312
rect 12253 1303 12311 1309
rect 11422 1272 11428 1284
rect 11256 1244 11428 1272
rect 11422 1232 11428 1244
rect 11480 1232 11486 1284
rect 12342 1204 12348 1216
rect 10888 1176 12348 1204
rect 12342 1164 12348 1176
rect 12400 1164 12406 1216
rect 13354 1164 13360 1216
rect 13412 1164 13418 1216
rect 13648 1204 13676 1312
rect 13722 1300 13728 1352
rect 13780 1300 13786 1352
rect 13832 1340 13860 1380
rect 15930 1368 15936 1420
rect 15988 1368 15994 1420
rect 16114 1368 16120 1420
rect 16172 1368 16178 1420
rect 18248 1408 18276 1436
rect 20088 1408 20116 1516
rect 20990 1504 20996 1516
rect 21048 1504 21054 1556
rect 21542 1504 21548 1556
rect 21600 1544 21606 1556
rect 21735 1547 21793 1553
rect 21735 1544 21747 1547
rect 21600 1516 21747 1544
rect 21600 1504 21606 1516
rect 21735 1513 21747 1516
rect 21781 1513 21793 1547
rect 21735 1507 21793 1513
rect 23014 1504 23020 1556
rect 23072 1504 23078 1556
rect 23293 1547 23351 1553
rect 23293 1513 23305 1547
rect 23339 1544 23351 1547
rect 23750 1544 23756 1556
rect 23339 1516 23756 1544
rect 23339 1513 23351 1516
rect 23293 1507 23351 1513
rect 23750 1504 23756 1516
rect 23808 1504 23814 1556
rect 23842 1504 23848 1556
rect 23900 1544 23906 1556
rect 24118 1544 24124 1556
rect 23900 1516 24124 1544
rect 23900 1504 23906 1516
rect 24118 1504 24124 1516
rect 24176 1504 24182 1556
rect 24302 1504 24308 1556
rect 24360 1544 24366 1556
rect 26605 1547 26663 1553
rect 26605 1544 26617 1547
rect 24360 1516 26617 1544
rect 24360 1504 24366 1516
rect 26605 1513 26617 1516
rect 26651 1513 26663 1547
rect 26605 1507 26663 1513
rect 26878 1504 26884 1556
rect 26936 1504 26942 1556
rect 27157 1547 27215 1553
rect 27157 1513 27169 1547
rect 27203 1513 27215 1547
rect 27157 1507 27215 1513
rect 20162 1436 20168 1488
rect 20220 1436 20226 1488
rect 20441 1479 20499 1485
rect 20441 1445 20453 1479
rect 20487 1476 20499 1479
rect 20487 1448 21404 1476
rect 20487 1445 20499 1448
rect 20441 1439 20499 1445
rect 18248 1380 20116 1408
rect 20180 1408 20208 1436
rect 20717 1411 20775 1417
rect 20717 1408 20729 1411
rect 20180 1380 20729 1408
rect 20717 1377 20729 1380
rect 20763 1377 20775 1411
rect 20717 1371 20775 1377
rect 20806 1368 20812 1420
rect 20864 1368 20870 1420
rect 20990 1368 20996 1420
rect 21048 1368 21054 1420
rect 21174 1368 21180 1420
rect 21232 1408 21238 1420
rect 21232 1380 21312 1408
rect 21232 1368 21238 1380
rect 14188 1343 14246 1349
rect 14188 1340 14200 1343
rect 13832 1312 14200 1340
rect 14188 1309 14200 1312
rect 14234 1309 14246 1343
rect 14188 1303 14246 1309
rect 14458 1300 14464 1352
rect 14516 1300 14522 1352
rect 15948 1340 15976 1368
rect 16580 1343 16638 1349
rect 16580 1340 16592 1343
rect 15948 1312 16592 1340
rect 16580 1309 16592 1312
rect 16626 1309 16638 1343
rect 16580 1303 16638 1309
rect 16853 1343 16911 1349
rect 16853 1309 16865 1343
rect 16899 1340 16911 1343
rect 17954 1340 17960 1352
rect 16899 1312 17960 1340
rect 16899 1309 16911 1312
rect 16853 1303 16911 1309
rect 17954 1300 17960 1312
rect 18012 1300 18018 1352
rect 18325 1343 18383 1349
rect 18325 1309 18337 1343
rect 18371 1340 18383 1343
rect 18598 1340 18604 1352
rect 18371 1312 18604 1340
rect 18371 1309 18383 1312
rect 18325 1303 18383 1309
rect 18598 1300 18604 1312
rect 18656 1300 18662 1352
rect 18782 1300 18788 1352
rect 18840 1340 18846 1352
rect 19061 1343 19119 1349
rect 18840 1312 18885 1340
rect 18840 1300 18846 1312
rect 19061 1309 19073 1343
rect 19107 1340 19119 1343
rect 19107 1312 20576 1340
rect 19107 1309 19119 1312
rect 19061 1303 19119 1309
rect 20548 1281 20576 1312
rect 20824 1281 20852 1368
rect 21284 1349 21312 1380
rect 21269 1343 21327 1349
rect 21269 1309 21281 1343
rect 21315 1309 21327 1343
rect 21376 1340 21404 1448
rect 23032 1408 23060 1504
rect 25792 1448 26096 1476
rect 21928 1380 22968 1408
rect 23032 1380 23612 1408
rect 21732 1361 21790 1367
rect 21732 1340 21744 1361
rect 21376 1327 21744 1340
rect 21778 1327 21790 1361
rect 21928 1352 21956 1380
rect 21376 1321 21790 1327
rect 21376 1312 21775 1321
rect 21269 1303 21327 1309
rect 21910 1300 21916 1352
rect 21968 1300 21974 1352
rect 22005 1343 22063 1349
rect 22005 1309 22017 1343
rect 22051 1340 22063 1343
rect 22830 1340 22836 1352
rect 22051 1312 22836 1340
rect 22051 1309 22063 1312
rect 22005 1303 22063 1309
rect 22830 1300 22836 1312
rect 22888 1300 22894 1352
rect 22940 1340 22968 1380
rect 23474 1340 23480 1352
rect 22940 1312 23480 1340
rect 23474 1300 23480 1312
rect 23532 1300 23538 1352
rect 23584 1340 23612 1380
rect 23750 1368 23756 1420
rect 23808 1417 23814 1420
rect 23808 1411 23862 1417
rect 23808 1377 23816 1411
rect 23850 1377 23862 1411
rect 23808 1371 23862 1377
rect 23808 1368 23814 1371
rect 24118 1368 24124 1420
rect 24176 1408 24182 1420
rect 24213 1411 24271 1417
rect 24213 1408 24225 1411
rect 24176 1380 24225 1408
rect 24176 1368 24182 1380
rect 24213 1377 24225 1380
rect 24259 1377 24271 1411
rect 24213 1371 24271 1377
rect 24302 1368 24308 1420
rect 24360 1408 24366 1420
rect 25792 1412 25820 1448
rect 25869 1412 25927 1417
rect 25792 1411 25927 1412
rect 25792 1408 25881 1411
rect 24360 1384 25881 1408
rect 24360 1380 25820 1384
rect 24360 1368 24366 1380
rect 25869 1377 25881 1384
rect 25915 1377 25927 1411
rect 25869 1371 25927 1377
rect 25958 1368 25964 1420
rect 26016 1368 26022 1420
rect 26068 1408 26096 1448
rect 26234 1436 26240 1488
rect 26292 1476 26298 1488
rect 27172 1476 27200 1507
rect 27430 1504 27436 1556
rect 27488 1504 27494 1556
rect 27798 1504 27804 1556
rect 27856 1544 27862 1556
rect 27991 1547 28049 1553
rect 27991 1544 28003 1547
rect 27856 1516 28003 1544
rect 27856 1504 27862 1516
rect 27991 1513 28003 1516
rect 28037 1513 28049 1547
rect 27991 1507 28049 1513
rect 28994 1504 29000 1556
rect 29052 1544 29058 1556
rect 29365 1547 29423 1553
rect 29365 1544 29377 1547
rect 29052 1516 29377 1544
rect 29052 1504 29058 1516
rect 29365 1513 29377 1516
rect 29411 1513 29423 1547
rect 29365 1507 29423 1513
rect 26292 1448 27200 1476
rect 26292 1436 26298 1448
rect 26421 1411 26479 1417
rect 26068 1380 26372 1408
rect 23940 1343 23998 1349
rect 23940 1340 23952 1343
rect 23584 1312 23952 1340
rect 23940 1309 23952 1312
rect 23986 1309 23998 1343
rect 23940 1303 23998 1309
rect 25130 1300 25136 1352
rect 25188 1340 25194 1352
rect 26344 1340 26372 1380
rect 26421 1377 26433 1411
rect 26467 1408 26479 1411
rect 26510 1408 26516 1420
rect 26467 1380 26516 1408
rect 26467 1377 26479 1380
rect 26421 1371 26479 1377
rect 26510 1368 26516 1380
rect 26568 1408 26574 1420
rect 26697 1411 26755 1417
rect 26697 1408 26709 1411
rect 26568 1380 26709 1408
rect 26568 1368 26574 1380
rect 26697 1377 26709 1380
rect 26743 1377 26755 1411
rect 26697 1371 26755 1377
rect 26970 1368 26976 1420
rect 27028 1368 27034 1420
rect 27249 1411 27307 1417
rect 27249 1377 27261 1411
rect 27295 1377 27307 1411
rect 27249 1371 27307 1377
rect 27264 1340 27292 1371
rect 27338 1368 27344 1420
rect 27396 1408 27402 1420
rect 27525 1411 27583 1417
rect 27525 1408 27537 1411
rect 27396 1380 27537 1408
rect 27396 1368 27402 1380
rect 27525 1377 27537 1380
rect 27571 1377 27583 1411
rect 27525 1371 27583 1377
rect 28021 1361 28079 1367
rect 28021 1358 28033 1361
rect 27706 1340 27712 1352
rect 25188 1312 26280 1340
rect 26344 1312 27712 1340
rect 25188 1300 25194 1312
rect 20533 1275 20591 1281
rect 20533 1241 20545 1275
rect 20579 1241 20591 1275
rect 20533 1235 20591 1241
rect 20809 1275 20867 1281
rect 20809 1241 20821 1275
rect 20855 1241 20867 1275
rect 20809 1235 20867 1241
rect 23032 1244 23244 1272
rect 23032 1204 23060 1244
rect 13648 1176 23060 1204
rect 23216 1204 23244 1244
rect 24872 1244 26188 1272
rect 24872 1204 24900 1244
rect 23216 1176 24900 1204
rect 25314 1164 25320 1216
rect 25372 1164 25378 1216
rect 25682 1164 25688 1216
rect 25740 1164 25746 1216
rect 26160 1213 26188 1244
rect 26145 1207 26203 1213
rect 26145 1173 26157 1207
rect 26191 1173 26203 1207
rect 26252 1204 26280 1312
rect 27706 1300 27712 1312
rect 27764 1300 27770 1352
rect 28000 1327 28033 1358
rect 28067 1352 28079 1361
rect 28067 1327 28080 1352
rect 28000 1312 28080 1327
rect 28074 1300 28080 1312
rect 28132 1300 28138 1352
rect 28166 1300 28172 1352
rect 28224 1340 28230 1352
rect 28261 1343 28319 1349
rect 28261 1340 28273 1343
rect 28224 1312 28273 1340
rect 28224 1300 28230 1312
rect 28261 1309 28273 1312
rect 28307 1309 28319 1343
rect 28261 1303 28319 1309
rect 28166 1204 28172 1216
rect 26252 1176 28172 1204
rect 26145 1167 26203 1173
rect 28166 1164 28172 1176
rect 28224 1164 28230 1216
rect 552 1114 30912 1136
rect 552 1062 4193 1114
rect 4245 1062 4257 1114
rect 4309 1062 4321 1114
rect 4373 1062 4385 1114
rect 4437 1062 4449 1114
rect 4501 1062 11783 1114
rect 11835 1062 11847 1114
rect 11899 1062 11911 1114
rect 11963 1062 11975 1114
rect 12027 1062 12039 1114
rect 12091 1062 19373 1114
rect 19425 1062 19437 1114
rect 19489 1062 19501 1114
rect 19553 1062 19565 1114
rect 19617 1062 19629 1114
rect 19681 1062 26963 1114
rect 27015 1062 27027 1114
rect 27079 1062 27091 1114
rect 27143 1062 27155 1114
rect 27207 1062 27219 1114
rect 27271 1062 30912 1114
rect 552 1040 30912 1062
rect 1302 1000 1308 1012
rect 952 972 1308 1000
rect 952 873 980 972
rect 1302 960 1308 972
rect 1360 1000 1366 1012
rect 1360 972 2774 1000
rect 1360 960 1366 972
rect 2498 892 2504 944
rect 2556 892 2562 944
rect 2746 932 2774 972
rect 2958 960 2964 1012
rect 3016 960 3022 1012
rect 3513 1003 3571 1009
rect 3513 969 3525 1003
rect 3559 1000 3571 1003
rect 4157 1003 4215 1009
rect 4157 1000 4169 1003
rect 3559 972 4169 1000
rect 3559 969 3571 972
rect 3513 963 3571 969
rect 4157 969 4169 972
rect 4203 1000 4215 1003
rect 4798 1000 4804 1012
rect 4203 972 4804 1000
rect 4203 969 4215 972
rect 4157 963 4215 969
rect 3528 932 3556 963
rect 4798 960 4804 972
rect 4856 960 4862 1012
rect 5166 960 5172 1012
rect 5224 960 5230 1012
rect 5445 1003 5503 1009
rect 5445 969 5457 1003
rect 5491 1000 5503 1003
rect 5491 972 7512 1000
rect 5491 969 5503 972
rect 5445 963 5503 969
rect 2746 904 3556 932
rect 3605 935 3663 941
rect 3605 901 3617 935
rect 3651 932 3663 935
rect 6086 932 6092 944
rect 3651 904 6092 932
rect 3651 901 3663 904
rect 3605 895 3663 901
rect 6086 892 6092 904
rect 6144 892 6150 944
rect 937 867 995 873
rect 937 833 949 867
rect 983 833 995 867
rect 1578 864 1584 876
rect 937 827 995 833
rect 1418 849 1584 864
rect 1418 818 1445 849
rect 1433 815 1445 818
rect 1479 836 1584 849
rect 1479 815 1491 836
rect 1578 824 1584 836
rect 1636 824 1642 876
rect 1670 824 1676 876
rect 1728 824 1734 876
rect 2516 864 2544 892
rect 2516 836 4844 864
rect 1433 809 1491 815
rect 3789 799 3847 805
rect 3789 765 3801 799
rect 3835 796 3847 799
rect 4706 796 4712 808
rect 3835 768 4712 796
rect 3835 765 3847 768
rect 3789 759 3847 765
rect 4706 756 4712 768
rect 4764 756 4770 808
rect 4816 796 4844 836
rect 4890 824 4896 876
rect 4948 864 4954 876
rect 6552 867 6610 873
rect 6552 864 6564 867
rect 4948 836 6564 864
rect 4948 824 4954 836
rect 6552 833 6564 836
rect 6598 833 6610 867
rect 6552 827 6610 833
rect 6638 824 6644 876
rect 6696 864 6702 876
rect 7484 864 7512 972
rect 7558 960 7564 1012
rect 7616 960 7622 1012
rect 8113 1003 8171 1009
rect 8113 969 8125 1003
rect 8159 1000 8171 1003
rect 9122 1000 9128 1012
rect 8159 972 9128 1000
rect 8159 969 8171 972
rect 8113 963 8171 969
rect 9122 960 9128 972
rect 9180 960 9186 1012
rect 9306 960 9312 1012
rect 9364 1000 9370 1012
rect 10689 1003 10747 1009
rect 9364 972 10180 1000
rect 9364 960 9370 972
rect 7576 932 7604 960
rect 8389 935 8447 941
rect 8389 932 8401 935
rect 7576 904 8401 932
rect 8389 901 8401 904
rect 8435 901 8447 935
rect 10152 932 10180 972
rect 10689 969 10701 1003
rect 10735 1000 10747 1003
rect 11054 1000 11060 1012
rect 10735 972 11060 1000
rect 10735 969 10747 972
rect 10689 963 10747 969
rect 11054 960 11060 972
rect 11112 960 11118 1012
rect 11974 960 11980 1012
rect 12032 1000 12038 1012
rect 13170 1000 13176 1012
rect 12032 972 13176 1000
rect 12032 960 12038 972
rect 13170 960 13176 972
rect 13228 960 13234 1012
rect 13262 960 13268 1012
rect 13320 960 13326 1012
rect 15286 960 15292 1012
rect 15344 1000 15350 1012
rect 15749 1003 15807 1009
rect 15749 1000 15761 1003
rect 15344 972 15761 1000
rect 15344 960 15350 972
rect 15749 969 15761 972
rect 15795 969 15807 1003
rect 15749 963 15807 969
rect 16117 1003 16175 1009
rect 16117 969 16129 1003
rect 16163 1000 16175 1003
rect 16206 1000 16212 1012
rect 16163 972 16212 1000
rect 16163 969 16175 972
rect 16117 963 16175 969
rect 16206 960 16212 972
rect 16264 960 16270 1012
rect 16316 972 17816 1000
rect 10965 935 11023 941
rect 10965 932 10977 935
rect 10152 904 10977 932
rect 8389 895 8447 901
rect 10965 901 10977 904
rect 11011 901 11023 935
rect 10965 895 11023 901
rect 15378 892 15384 944
rect 15436 892 15442 944
rect 15470 892 15476 944
rect 15528 932 15534 944
rect 16316 932 16344 972
rect 15528 904 16344 932
rect 15528 892 15534 904
rect 9171 867 9229 873
rect 6696 836 7420 864
rect 7484 836 8800 864
rect 6696 824 6702 836
rect 5077 799 5135 805
rect 5077 796 5089 799
rect 4816 768 5089 796
rect 5077 765 5089 768
rect 5123 796 5135 799
rect 5258 796 5264 808
rect 5123 768 5264 796
rect 5123 765 5135 768
rect 5077 759 5135 765
rect 5258 756 5264 768
rect 5316 756 5322 808
rect 5350 756 5356 808
rect 5408 756 5414 808
rect 5629 799 5687 805
rect 5629 765 5641 799
rect 5675 796 5687 799
rect 5902 796 5908 808
rect 5675 768 5908 796
rect 5675 765 5687 768
rect 5629 759 5687 765
rect 3418 688 3424 740
rect 3476 728 3482 740
rect 5644 728 5672 759
rect 5902 756 5908 768
rect 5960 756 5966 808
rect 5997 799 6055 805
rect 5997 765 6009 799
rect 6043 765 6055 799
rect 5997 759 6055 765
rect 6089 799 6147 805
rect 6089 765 6101 799
rect 6135 765 6147 799
rect 6089 759 6147 765
rect 3476 700 5672 728
rect 3476 688 3482 700
rect 6012 672 6040 759
rect 1403 663 1461 669
rect 1403 629 1415 663
rect 1449 660 1461 663
rect 1762 660 1768 672
rect 1449 632 1768 660
rect 1449 629 1461 632
rect 1403 623 1461 629
rect 1762 620 1768 632
rect 1820 660 1826 672
rect 2682 660 2688 672
rect 1820 632 2688 660
rect 1820 620 1826 632
rect 2682 620 2688 632
rect 2740 620 2746 672
rect 4798 620 4804 672
rect 4856 620 4862 672
rect 4890 620 4896 672
rect 4948 620 4954 672
rect 5810 620 5816 672
rect 5868 620 5874 672
rect 5994 620 6000 672
rect 6052 620 6058 672
rect 6104 660 6132 759
rect 6178 756 6184 808
rect 6236 796 6242 808
rect 6825 799 6883 805
rect 6825 796 6837 799
rect 6236 768 6837 796
rect 6236 756 6242 768
rect 6825 765 6837 768
rect 6871 765 6883 799
rect 7392 796 7420 836
rect 7392 768 8524 796
rect 6825 759 6883 765
rect 8496 728 8524 768
rect 8570 756 8576 808
rect 8628 756 8634 808
rect 8665 799 8723 805
rect 8665 765 8677 799
rect 8711 765 8723 799
rect 8772 796 8800 836
rect 9171 833 9183 867
rect 9217 864 9229 867
rect 9217 836 11100 864
rect 9217 833 9229 836
rect 9171 827 9229 833
rect 9401 799 9459 805
rect 9401 796 9413 799
rect 8772 768 9413 796
rect 8665 759 8723 765
rect 9401 765 9413 768
rect 9447 765 9459 799
rect 9401 759 9459 765
rect 8680 728 8708 759
rect 8754 728 8760 740
rect 8496 700 8760 728
rect 8754 688 8760 700
rect 8812 688 8818 740
rect 6454 660 6460 672
rect 6104 632 6460 660
rect 6454 620 6460 632
rect 6512 620 6518 672
rect 6555 663 6613 669
rect 6555 629 6567 663
rect 6601 660 6613 663
rect 9131 663 9189 669
rect 9131 660 9143 663
rect 6601 632 9143 660
rect 6601 629 6613 632
rect 6555 623 6613 629
rect 9131 629 9143 632
rect 9177 660 9189 663
rect 9398 660 9404 672
rect 9177 632 9404 660
rect 9177 629 9189 632
rect 9131 623 9189 629
rect 9398 620 9404 632
rect 9456 620 9462 672
rect 11072 660 11100 836
rect 11238 824 11244 876
rect 11296 824 11302 876
rect 11790 871 11796 876
rect 11747 865 11796 871
rect 11747 831 11759 865
rect 11793 831 11796 865
rect 11747 825 11796 831
rect 11790 824 11796 825
rect 11848 824 11854 876
rect 12342 824 12348 876
rect 12400 864 12406 876
rect 14090 873 14096 876
rect 13541 867 13599 873
rect 13541 864 13553 867
rect 12400 836 13553 864
rect 12400 824 12406 836
rect 13541 833 13553 836
rect 13587 833 13599 867
rect 13541 827 13599 833
rect 14047 867 14096 873
rect 14047 833 14059 867
rect 14093 833 14096 867
rect 14047 827 14096 833
rect 14090 824 14096 827
rect 14148 824 14154 876
rect 14200 836 16436 864
rect 11149 799 11207 805
rect 11149 765 11161 799
rect 11195 796 11207 799
rect 11330 796 11336 808
rect 11195 768 11336 796
rect 11195 765 11207 768
rect 11149 759 11207 765
rect 11330 756 11336 768
rect 11388 756 11394 808
rect 11974 756 11980 808
rect 12032 756 12038 808
rect 13630 756 13636 808
rect 13688 796 13694 808
rect 14200 796 14228 836
rect 13688 768 14228 796
rect 13688 756 13694 768
rect 14274 756 14280 808
rect 14332 756 14338 808
rect 14550 756 14556 808
rect 14608 796 14614 808
rect 15933 799 15991 805
rect 15933 796 15945 799
rect 14608 768 15945 796
rect 14608 756 14614 768
rect 15933 765 15945 768
rect 15979 765 15991 799
rect 15933 759 15991 765
rect 16298 756 16304 808
rect 16356 756 16362 808
rect 16408 805 16436 836
rect 16850 824 16856 876
rect 16908 855 16914 876
rect 17788 864 17816 972
rect 18690 960 18696 1012
rect 18748 960 18754 1012
rect 19334 960 19340 1012
rect 19392 1000 19398 1012
rect 20070 1000 20076 1012
rect 19392 972 20076 1000
rect 19392 960 19398 972
rect 20070 960 20076 972
rect 20128 960 20134 1012
rect 22646 1000 22652 1012
rect 20732 972 22652 1000
rect 19475 867 19533 873
rect 16908 849 16947 855
rect 16868 818 16901 824
rect 16889 815 16901 818
rect 16935 815 16947 849
rect 17788 836 18920 864
rect 16889 809 16947 815
rect 16393 799 16451 805
rect 16393 765 16405 799
rect 16439 796 16451 799
rect 16482 796 16488 808
rect 16439 768 16488 796
rect 16439 765 16451 768
rect 16393 759 16451 765
rect 16482 756 16488 768
rect 16540 756 16546 808
rect 17126 756 17132 808
rect 17184 756 17190 808
rect 18892 805 18920 836
rect 19475 833 19487 867
rect 19521 864 19533 867
rect 20732 864 20760 972
rect 22646 960 22652 972
rect 22704 960 22710 1012
rect 22738 960 22744 1012
rect 22796 1000 22802 1012
rect 23385 1003 23443 1009
rect 23385 1000 23397 1003
rect 22796 972 23397 1000
rect 22796 960 22802 972
rect 23385 969 23397 972
rect 23431 969 23443 1003
rect 25961 1003 26019 1009
rect 25961 1000 25973 1003
rect 23385 963 23443 969
rect 23492 972 25973 1000
rect 19521 836 20760 864
rect 19521 833 19533 836
rect 19475 827 19533 833
rect 21358 824 21364 876
rect 21416 864 21422 876
rect 21545 867 21603 873
rect 21545 864 21557 867
rect 21416 836 21557 864
rect 21416 824 21422 836
rect 21545 833 21557 836
rect 21591 864 21603 867
rect 21910 864 21916 876
rect 21591 836 21916 864
rect 21591 833 21603 836
rect 21545 827 21603 833
rect 21910 824 21916 836
rect 21968 824 21974 876
rect 22051 867 22109 873
rect 22051 833 22063 867
rect 22097 864 22109 867
rect 22186 864 22192 876
rect 22097 836 22192 864
rect 22097 833 22109 836
rect 22051 827 22109 833
rect 22186 824 22192 836
rect 22244 824 22250 876
rect 22281 867 22339 873
rect 22281 833 22293 867
rect 22327 864 22339 867
rect 22922 864 22928 876
rect 22327 836 22928 864
rect 22327 833 22339 836
rect 22281 827 22339 833
rect 22922 824 22928 836
rect 22980 824 22986 876
rect 18877 799 18935 805
rect 18877 765 18889 799
rect 18923 765 18935 799
rect 18877 759 18935 765
rect 18969 799 19027 805
rect 18969 765 18981 799
rect 19015 796 19027 799
rect 19058 796 19064 808
rect 19015 768 19064 796
rect 19015 765 19027 768
rect 18969 759 19027 765
rect 19058 756 19064 768
rect 19116 756 19122 808
rect 19334 805 19340 808
rect 19296 799 19340 805
rect 19296 765 19308 799
rect 19296 759 19340 765
rect 19334 756 19340 759
rect 19392 756 19398 808
rect 19705 799 19763 805
rect 19705 765 19717 799
rect 19751 796 19763 799
rect 20622 796 20628 808
rect 19751 768 20628 796
rect 19751 765 19763 768
rect 19705 759 19763 765
rect 20622 756 20628 768
rect 20680 756 20686 808
rect 20714 756 20720 808
rect 20772 796 20778 808
rect 21450 796 21456 808
rect 20772 768 21456 796
rect 20772 756 20778 768
rect 21450 756 21456 768
rect 21508 756 21514 808
rect 22646 756 22652 808
rect 22704 796 22710 808
rect 23492 796 23520 972
rect 25961 969 25973 972
rect 26007 969 26019 1003
rect 25961 963 26019 969
rect 26050 960 26056 1012
rect 26108 1000 26114 1012
rect 26421 1003 26479 1009
rect 26421 1000 26433 1003
rect 26108 972 26433 1000
rect 26108 960 26114 972
rect 26421 969 26433 972
rect 26467 969 26479 1003
rect 29914 1000 29920 1012
rect 26421 963 26479 969
rect 26620 972 29920 1000
rect 23658 892 23664 944
rect 23716 932 23722 944
rect 23845 935 23903 941
rect 23845 932 23857 935
rect 23716 904 23857 932
rect 23716 892 23722 904
rect 23845 901 23857 904
rect 23891 901 23903 935
rect 23845 895 23903 901
rect 24026 892 24032 944
rect 24084 892 24090 944
rect 24044 864 24072 892
rect 24670 873 24676 876
rect 24627 867 24676 873
rect 24044 836 24532 864
rect 22704 768 23520 796
rect 22704 756 22710 768
rect 23934 756 23940 808
rect 23992 796 23998 808
rect 24029 799 24087 805
rect 24029 796 24041 799
rect 23992 768 24041 796
rect 23992 756 23998 768
rect 24029 765 24041 768
rect 24075 765 24087 799
rect 24029 759 24087 765
rect 24118 756 24124 808
rect 24176 756 24182 808
rect 24504 796 24532 836
rect 24627 833 24639 867
rect 24673 833 24676 867
rect 24627 827 24676 833
rect 24670 824 24676 827
rect 24728 824 24734 876
rect 26620 805 26648 972
rect 29914 960 29920 972
rect 29972 960 29978 1012
rect 28166 892 28172 944
rect 28224 932 28230 944
rect 28537 935 28595 941
rect 28537 932 28549 935
rect 28224 904 28549 932
rect 28224 892 28230 904
rect 28537 901 28549 904
rect 28583 901 28595 935
rect 28537 895 28595 901
rect 27203 867 27261 873
rect 27203 833 27215 867
rect 27249 864 27261 867
rect 27614 864 27620 876
rect 27249 836 27620 864
rect 27249 833 27261 836
rect 27203 827 27261 833
rect 27614 824 27620 836
rect 27672 824 27678 876
rect 24857 799 24915 805
rect 24857 796 24869 799
rect 24504 768 24869 796
rect 24857 765 24869 768
rect 24903 765 24915 799
rect 24857 759 24915 765
rect 26605 799 26663 805
rect 26605 765 26617 799
rect 26651 765 26663 799
rect 26605 759 26663 765
rect 26697 799 26755 805
rect 26697 765 26709 799
rect 26743 796 26755 799
rect 27338 796 27344 808
rect 26743 768 27344 796
rect 26743 765 26755 768
rect 26697 759 26755 765
rect 27338 756 27344 768
rect 27396 756 27402 808
rect 27433 799 27491 805
rect 27433 765 27445 799
rect 27479 796 27491 799
rect 29086 796 29092 808
rect 27479 768 29092 796
rect 27479 765 27491 768
rect 27433 759 27491 765
rect 29086 756 29092 768
rect 29144 756 29150 808
rect 20438 688 20444 740
rect 20496 728 20502 740
rect 20496 700 21312 728
rect 20496 688 20502 700
rect 11606 660 11612 672
rect 11072 632 11612 660
rect 11606 620 11612 632
rect 11664 620 11670 672
rect 11707 663 11765 669
rect 11707 629 11719 663
rect 11753 660 11765 663
rect 12250 660 12256 672
rect 11753 632 12256 660
rect 11753 629 11765 632
rect 11707 623 11765 629
rect 12250 620 12256 632
rect 12308 620 12314 672
rect 13814 620 13820 672
rect 13872 660 13878 672
rect 14007 663 14065 669
rect 14007 660 14019 663
rect 13872 632 14019 660
rect 13872 620 13878 632
rect 14007 629 14019 632
rect 14053 629 14065 663
rect 14007 623 14065 629
rect 15010 620 15016 672
rect 15068 660 15074 672
rect 16859 663 16917 669
rect 16859 660 16871 663
rect 15068 632 16871 660
rect 15068 620 15074 632
rect 16859 629 16871 632
rect 16905 660 16917 663
rect 17954 660 17960 672
rect 16905 632 17960 660
rect 16905 629 16917 632
rect 16859 623 16917 629
rect 17954 620 17960 632
rect 18012 620 18018 672
rect 18230 620 18236 672
rect 18288 620 18294 672
rect 18322 620 18328 672
rect 18380 660 18386 672
rect 21284 669 21312 700
rect 20809 663 20867 669
rect 20809 660 20821 663
rect 18380 632 20821 660
rect 18380 620 18386 632
rect 20809 629 20821 632
rect 20855 629 20867 663
rect 20809 623 20867 629
rect 21269 663 21327 669
rect 21269 629 21281 663
rect 21315 629 21327 663
rect 21269 623 21327 629
rect 22011 663 22069 669
rect 22011 629 22023 663
rect 22057 660 22069 663
rect 23750 660 23756 672
rect 22057 632 23756 660
rect 22057 629 22069 632
rect 22011 623 22069 629
rect 23750 620 23756 632
rect 23808 620 23814 672
rect 23934 620 23940 672
rect 23992 660 23998 672
rect 24486 660 24492 672
rect 23992 632 24492 660
rect 23992 620 23998 632
rect 24486 620 24492 632
rect 24544 660 24550 672
rect 24587 663 24645 669
rect 24587 660 24599 663
rect 24544 632 24599 660
rect 24544 620 24550 632
rect 24587 629 24599 632
rect 24633 629 24645 663
rect 24587 623 24645 629
rect 27163 663 27221 669
rect 27163 629 27175 663
rect 27209 660 27221 663
rect 27798 660 27804 672
rect 27209 632 27804 660
rect 27209 629 27221 632
rect 27163 623 27221 629
rect 27798 620 27804 632
rect 27856 620 27862 672
rect 552 570 31072 592
rect 552 518 7988 570
rect 8040 518 8052 570
rect 8104 518 8116 570
rect 8168 518 8180 570
rect 8232 518 8244 570
rect 8296 518 15578 570
rect 15630 518 15642 570
rect 15694 518 15706 570
rect 15758 518 15770 570
rect 15822 518 15834 570
rect 15886 518 23168 570
rect 23220 518 23232 570
rect 23284 518 23296 570
rect 23348 518 23360 570
rect 23412 518 23424 570
rect 23476 518 30758 570
rect 30810 518 30822 570
rect 30874 518 30886 570
rect 30938 518 30950 570
rect 31002 518 31014 570
rect 31066 518 31072 570
rect 552 496 31072 518
rect 1578 416 1584 468
rect 1636 416 1642 468
rect 5810 416 5816 468
rect 5868 456 5874 468
rect 11698 456 11704 468
rect 5868 428 11704 456
rect 5868 416 5874 428
rect 11698 416 11704 428
rect 11756 416 11762 468
rect 14274 456 14280 468
rect 12406 428 14280 456
rect 1596 252 1624 416
rect 9122 348 9128 400
rect 9180 388 9186 400
rect 12406 388 12434 428
rect 14274 416 14280 428
rect 14332 416 14338 468
rect 16850 416 16856 468
rect 16908 416 16914 468
rect 17126 416 17132 468
rect 17184 456 17190 468
rect 25682 456 25688 468
rect 17184 428 25688 456
rect 17184 416 17190 428
rect 25682 416 25688 428
rect 25740 416 25746 468
rect 9180 360 12434 388
rect 16868 388 16896 416
rect 24854 388 24860 400
rect 16868 360 24860 388
rect 9180 348 9186 360
rect 24854 348 24860 360
rect 24912 348 24918 400
rect 2682 280 2688 332
rect 2740 320 2746 332
rect 17034 320 17040 332
rect 2740 292 17040 320
rect 2740 280 2746 292
rect 17034 280 17040 292
rect 17092 280 17098 332
rect 17954 280 17960 332
rect 18012 320 18018 332
rect 23934 320 23940 332
rect 18012 292 23940 320
rect 18012 280 18018 292
rect 23934 280 23940 292
rect 23992 280 23998 332
rect 13354 252 13360 264
rect 1596 224 13360 252
rect 13354 212 13360 224
rect 13412 212 13418 264
rect 17052 252 17080 280
rect 19334 252 19340 264
rect 17052 224 19340 252
rect 19334 212 19340 224
rect 19392 212 19398 264
rect 4982 144 4988 196
rect 5040 144 5046 196
rect 5074 144 5080 196
rect 5132 184 5138 196
rect 15102 184 15108 196
rect 5132 156 15108 184
rect 5132 144 5138 156
rect 15102 144 15108 156
rect 15160 144 15166 196
rect 16482 144 16488 196
rect 16540 184 16546 196
rect 24118 184 24124 196
rect 16540 156 24124 184
rect 16540 144 16546 156
rect 24118 144 24124 156
rect 24176 144 24182 196
rect 5000 116 5028 144
rect 9122 116 9128 128
rect 5000 88 9128 116
rect 9122 76 9128 88
rect 9180 76 9186 128
rect 11790 76 11796 128
rect 11848 116 11854 128
rect 18322 116 18328 128
rect 11848 88 18328 116
rect 11848 76 11854 88
rect 18322 76 18328 88
rect 18380 76 18386 128
rect 4706 8 4712 60
rect 4764 48 4770 60
rect 5994 48 6000 60
rect 4764 20 6000 48
rect 4764 8 4770 20
rect 5994 8 6000 20
rect 6052 48 6058 60
rect 9766 48 9772 60
rect 6052 20 9772 48
rect 6052 8 6058 20
rect 9766 8 9772 20
rect 9824 8 9830 60
<< via1 >>
rect 10968 22244 11020 22296
rect 18880 22244 18932 22296
rect 24216 22244 24268 22296
rect 25044 22244 25096 22296
rect 31208 22244 31260 22296
rect 9128 22176 9180 22228
rect 15752 22176 15804 22228
rect 7564 22108 7616 22160
rect 16764 22176 16816 22228
rect 16856 22176 16908 22228
rect 27620 22176 27672 22228
rect 15936 22108 15988 22160
rect 25872 22108 25924 22160
rect 10508 22040 10560 22092
rect 16120 22040 16172 22092
rect 10140 21972 10192 22024
rect 10600 21972 10652 22024
rect 15568 21972 15620 22024
rect 18696 22040 18748 22092
rect 19248 22040 19300 22092
rect 24124 22040 24176 22092
rect 28724 22040 28776 22092
rect 5448 21904 5500 21956
rect 7748 21904 7800 21956
rect 11428 21904 11480 21956
rect 4804 21836 4856 21888
rect 10324 21836 10376 21888
rect 10416 21836 10468 21888
rect 30288 21972 30340 22024
rect 17500 21836 17552 21888
rect 19708 21836 19760 21888
rect 20628 21836 20680 21888
rect 23388 21836 23440 21888
rect 24584 21836 24636 21888
rect 25964 21836 26016 21888
rect 27804 21836 27856 21888
rect 4193 21734 4245 21786
rect 4257 21734 4309 21786
rect 4321 21734 4373 21786
rect 4385 21734 4437 21786
rect 4449 21734 4501 21786
rect 11783 21734 11835 21786
rect 11847 21734 11899 21786
rect 11911 21734 11963 21786
rect 11975 21734 12027 21786
rect 12039 21734 12091 21786
rect 19373 21734 19425 21786
rect 19437 21734 19489 21786
rect 19501 21734 19553 21786
rect 19565 21734 19617 21786
rect 19629 21734 19681 21786
rect 26963 21734 27015 21786
rect 27027 21734 27079 21786
rect 27091 21734 27143 21786
rect 27155 21734 27207 21786
rect 27219 21734 27271 21786
rect 848 21428 900 21480
rect 7564 21632 7616 21684
rect 11704 21632 11756 21684
rect 12532 21632 12584 21684
rect 2780 21428 2832 21480
rect 3240 21471 3292 21480
rect 3240 21437 3249 21471
rect 3249 21437 3283 21471
rect 3283 21437 3292 21471
rect 3240 21428 3292 21437
rect 2872 21360 2924 21412
rect 4068 21428 4120 21480
rect 5448 21428 5500 21480
rect 5356 21403 5408 21412
rect 5356 21369 5365 21403
rect 5365 21369 5399 21403
rect 5399 21369 5408 21403
rect 5356 21360 5408 21369
rect 5724 21360 5776 21412
rect 6184 21428 6236 21480
rect 8668 21496 8720 21548
rect 9128 21539 9180 21548
rect 9128 21505 9137 21539
rect 9137 21505 9171 21539
rect 9171 21505 9180 21539
rect 9128 21496 9180 21505
rect 9588 21496 9640 21548
rect 7380 21428 7432 21480
rect 8300 21428 8352 21480
rect 8392 21471 8444 21480
rect 8392 21437 8401 21471
rect 8401 21437 8435 21471
rect 8435 21437 8444 21471
rect 8392 21428 8444 21437
rect 7288 21360 7340 21412
rect 9772 21428 9824 21480
rect 11060 21496 11112 21548
rect 11244 21428 11296 21480
rect 11428 21428 11480 21480
rect 16856 21632 16908 21684
rect 18880 21675 18932 21684
rect 18880 21641 18889 21675
rect 18889 21641 18923 21675
rect 18923 21641 18932 21675
rect 18880 21632 18932 21641
rect 15568 21564 15620 21616
rect 1400 21335 1452 21344
rect 1400 21301 1415 21335
rect 1415 21301 1449 21335
rect 1449 21301 1452 21335
rect 1400 21292 1452 21301
rect 3608 21292 3660 21344
rect 3884 21292 3936 21344
rect 5908 21292 5960 21344
rect 6092 21292 6144 21344
rect 6460 21292 6512 21344
rect 8668 21292 8720 21344
rect 10232 21335 10284 21344
rect 10232 21301 10241 21335
rect 10241 21301 10275 21335
rect 10275 21301 10284 21335
rect 10232 21292 10284 21301
rect 10968 21292 11020 21344
rect 11612 21335 11664 21344
rect 11612 21301 11627 21335
rect 11627 21301 11661 21335
rect 11661 21301 11664 21335
rect 11612 21292 11664 21301
rect 12348 21292 12400 21344
rect 13820 21360 13872 21412
rect 23388 21675 23440 21684
rect 23388 21641 23397 21675
rect 23397 21641 23431 21675
rect 23431 21641 23440 21675
rect 23388 21632 23440 21641
rect 15936 21403 15988 21412
rect 15936 21369 15945 21403
rect 15945 21369 15979 21403
rect 15979 21369 15988 21403
rect 15936 21360 15988 21369
rect 12992 21335 13044 21344
rect 12992 21301 13001 21335
rect 13001 21301 13035 21335
rect 13035 21301 13044 21335
rect 12992 21292 13044 21301
rect 14188 21292 14240 21344
rect 15476 21292 15528 21344
rect 16120 21471 16172 21480
rect 16120 21437 16129 21471
rect 16129 21437 16163 21471
rect 16163 21437 16172 21471
rect 16120 21428 16172 21437
rect 16856 21471 16908 21480
rect 16856 21437 16865 21471
rect 16865 21437 16899 21471
rect 16899 21437 16908 21471
rect 16856 21428 16908 21437
rect 22100 21496 22152 21548
rect 24216 21564 24268 21616
rect 24492 21632 24544 21684
rect 25964 21632 26016 21684
rect 27804 21675 27856 21684
rect 27804 21641 27813 21675
rect 27813 21641 27847 21675
rect 27847 21641 27856 21675
rect 27804 21632 27856 21641
rect 23940 21496 23992 21548
rect 24400 21496 24452 21548
rect 25688 21496 25740 21548
rect 26792 21496 26844 21548
rect 30564 21564 30616 21616
rect 19248 21428 19300 21480
rect 19708 21471 19760 21480
rect 19708 21437 19717 21471
rect 19717 21437 19751 21471
rect 19751 21437 19760 21471
rect 19708 21428 19760 21437
rect 18512 21403 18564 21412
rect 18512 21369 18521 21403
rect 18521 21369 18555 21403
rect 18555 21369 18564 21403
rect 18512 21360 18564 21369
rect 21456 21428 21508 21480
rect 22284 21471 22336 21480
rect 22284 21437 22293 21471
rect 22293 21437 22327 21471
rect 22327 21437 22336 21471
rect 22284 21428 22336 21437
rect 23664 21428 23716 21480
rect 18604 21292 18656 21344
rect 21364 21292 21416 21344
rect 23020 21292 23072 21344
rect 24860 21471 24912 21480
rect 24860 21437 24894 21471
rect 24894 21437 24912 21471
rect 24860 21428 24912 21437
rect 25044 21471 25096 21480
rect 25044 21437 25053 21471
rect 25053 21437 25087 21471
rect 25087 21437 25096 21471
rect 25044 21428 25096 21437
rect 26332 21428 26384 21480
rect 27344 21428 27396 21480
rect 27620 21428 27672 21480
rect 28356 21428 28408 21480
rect 29092 21471 29144 21480
rect 29092 21437 29101 21471
rect 29101 21437 29135 21471
rect 29135 21437 29144 21471
rect 29092 21428 29144 21437
rect 29276 21471 29328 21480
rect 29276 21437 29285 21471
rect 29285 21437 29319 21471
rect 29319 21437 29328 21471
rect 29276 21428 29328 21437
rect 31116 21428 31168 21480
rect 25320 21292 25372 21344
rect 25780 21292 25832 21344
rect 29828 21360 29880 21412
rect 29920 21403 29972 21412
rect 29920 21369 29929 21403
rect 29929 21369 29963 21403
rect 29963 21369 29972 21403
rect 29920 21360 29972 21369
rect 28724 21292 28776 21344
rect 29736 21292 29788 21344
rect 7988 21190 8040 21242
rect 8052 21190 8104 21242
rect 8116 21190 8168 21242
rect 8180 21190 8232 21242
rect 8244 21190 8296 21242
rect 15578 21190 15630 21242
rect 15642 21190 15694 21242
rect 15706 21190 15758 21242
rect 15770 21190 15822 21242
rect 15834 21190 15886 21242
rect 23168 21190 23220 21242
rect 23232 21190 23284 21242
rect 23296 21190 23348 21242
rect 23360 21190 23412 21242
rect 23424 21190 23476 21242
rect 30758 21190 30810 21242
rect 30822 21190 30874 21242
rect 30886 21190 30938 21242
rect 30950 21190 31002 21242
rect 31014 21190 31066 21242
rect 1400 21131 1452 21140
rect 1400 21097 1415 21131
rect 1415 21097 1449 21131
rect 1449 21097 1452 21131
rect 1400 21088 1452 21097
rect 3608 21131 3660 21140
rect 3608 21097 3623 21131
rect 3623 21097 3657 21131
rect 3657 21097 3660 21131
rect 3608 21088 3660 21097
rect 5816 21088 5868 21140
rect 6552 21088 6604 21140
rect 10232 21088 10284 21140
rect 14464 21088 14516 21140
rect 14832 21088 14884 21140
rect 15384 21088 15436 21140
rect 15660 21131 15712 21140
rect 15660 21097 15669 21131
rect 15669 21097 15703 21131
rect 15703 21097 15712 21131
rect 15660 21088 15712 21097
rect 16580 21088 16632 21140
rect 1676 20995 1728 21004
rect 1676 20961 1685 20995
rect 1685 20961 1719 20995
rect 1719 20961 1728 20995
rect 1676 20952 1728 20961
rect 5448 20952 5500 21004
rect 5540 20952 5592 21004
rect 940 20927 992 20936
rect 940 20893 949 20927
rect 949 20893 983 20927
rect 983 20893 992 20927
rect 940 20884 992 20893
rect 1860 20884 1912 20936
rect 3332 20884 3384 20936
rect 3608 20927 3660 20936
rect 3608 20893 3620 20927
rect 3620 20893 3654 20927
rect 3654 20893 3660 20927
rect 3608 20884 3660 20893
rect 2964 20791 3016 20800
rect 2964 20757 2973 20791
rect 2973 20757 3007 20791
rect 3007 20757 3016 20791
rect 2964 20748 3016 20757
rect 5540 20791 5592 20800
rect 5540 20757 5549 20791
rect 5549 20757 5583 20791
rect 5583 20757 5592 20791
rect 5540 20748 5592 20757
rect 6736 20884 6788 20936
rect 7656 20748 7708 20800
rect 7840 20791 7892 20800
rect 7840 20757 7849 20791
rect 7849 20757 7883 20791
rect 7883 20757 7892 20791
rect 7840 20748 7892 20757
rect 8392 20884 8444 20936
rect 8760 20952 8812 21004
rect 9128 20952 9180 21004
rect 10416 21063 10468 21072
rect 10416 21029 10425 21063
rect 10425 21029 10459 21063
rect 10459 21029 10468 21063
rect 10416 21020 10468 21029
rect 17132 21131 17184 21140
rect 17132 21097 17141 21131
rect 17141 21097 17175 21131
rect 17175 21097 17184 21131
rect 17132 21088 17184 21097
rect 17868 21088 17920 21140
rect 18604 21131 18656 21140
rect 18604 21097 18613 21131
rect 18613 21097 18647 21131
rect 18647 21097 18656 21131
rect 18604 21088 18656 21097
rect 19248 21088 19300 21140
rect 21364 21088 21416 21140
rect 22284 21088 22336 21140
rect 23388 21088 23440 21140
rect 24768 21088 24820 21140
rect 25320 21131 25372 21140
rect 25320 21097 25329 21131
rect 25329 21097 25363 21131
rect 25363 21097 25372 21131
rect 25320 21088 25372 21097
rect 29920 21088 29972 21140
rect 10324 20952 10376 21004
rect 12624 20952 12676 21004
rect 16120 20952 16172 21004
rect 16672 20995 16724 21004
rect 16672 20961 16681 20995
rect 16681 20961 16715 20995
rect 16715 20961 16724 20995
rect 16672 20952 16724 20961
rect 17500 20995 17552 21004
rect 17500 20961 17509 20995
rect 17509 20961 17543 20995
rect 17543 20961 17552 20995
rect 17500 20952 17552 20961
rect 25136 21020 25188 21072
rect 26056 21063 26108 21072
rect 26056 21029 26065 21063
rect 26065 21029 26099 21063
rect 26099 21029 26108 21063
rect 26056 21020 26108 21029
rect 8668 20884 8720 20936
rect 8944 20884 8996 20936
rect 9036 20884 9088 20936
rect 11152 20884 11204 20936
rect 11428 20927 11480 20936
rect 11428 20893 11440 20927
rect 11440 20893 11474 20927
rect 11474 20893 11480 20927
rect 11428 20884 11480 20893
rect 20720 20952 20772 21004
rect 8484 20748 8536 20800
rect 9588 20748 9640 20800
rect 10784 20748 10836 20800
rect 11428 20748 11480 20800
rect 12716 20748 12768 20800
rect 13176 20748 13228 20800
rect 19708 20884 19760 20936
rect 23112 20952 23164 21004
rect 21272 20927 21324 20936
rect 21272 20893 21281 20927
rect 21281 20893 21315 20927
rect 21315 20893 21324 20927
rect 21272 20884 21324 20893
rect 21732 20748 21784 20800
rect 22192 20748 22244 20800
rect 25596 20952 25648 21004
rect 26148 20995 26200 21004
rect 26148 20961 26157 20995
rect 26157 20961 26191 20995
rect 26191 20961 26200 20995
rect 26148 20952 26200 20961
rect 26976 20952 27028 21004
rect 26240 20884 26292 20936
rect 27436 20884 27488 20936
rect 27528 20884 27580 20936
rect 29000 20884 29052 20936
rect 29828 20884 29880 20936
rect 28264 20748 28316 20800
rect 28540 20748 28592 20800
rect 4193 20646 4245 20698
rect 4257 20646 4309 20698
rect 4321 20646 4373 20698
rect 4385 20646 4437 20698
rect 4449 20646 4501 20698
rect 11783 20646 11835 20698
rect 11847 20646 11899 20698
rect 11911 20646 11963 20698
rect 11975 20646 12027 20698
rect 12039 20646 12091 20698
rect 19373 20646 19425 20698
rect 19437 20646 19489 20698
rect 19501 20646 19553 20698
rect 19565 20646 19617 20698
rect 19629 20646 19681 20698
rect 26963 20646 27015 20698
rect 27027 20646 27079 20698
rect 27091 20646 27143 20698
rect 27155 20646 27207 20698
rect 27219 20646 27271 20698
rect 848 20340 900 20392
rect 1308 20451 1360 20460
rect 1308 20417 1310 20451
rect 1310 20417 1360 20451
rect 1308 20408 1360 20417
rect 1584 20408 1636 20460
rect 1676 20451 1728 20460
rect 1676 20417 1685 20451
rect 1685 20417 1719 20451
rect 1719 20417 1728 20451
rect 1676 20408 1728 20417
rect 3608 20544 3660 20596
rect 4712 20544 4764 20596
rect 6276 20408 6328 20460
rect 6644 20408 6696 20460
rect 6736 20408 6788 20460
rect 9128 20544 9180 20596
rect 10232 20408 10284 20460
rect 3424 20340 3476 20392
rect 4528 20340 4580 20392
rect 4896 20340 4948 20392
rect 5724 20340 5776 20392
rect 6184 20340 6236 20392
rect 6920 20340 6972 20392
rect 7564 20340 7616 20392
rect 8760 20340 8812 20392
rect 10692 20340 10744 20392
rect 12992 20544 13044 20596
rect 14004 20544 14056 20596
rect 21916 20544 21968 20596
rect 23848 20544 23900 20596
rect 25780 20544 25832 20596
rect 10876 20476 10928 20528
rect 20720 20476 20772 20528
rect 21364 20476 21416 20528
rect 14188 20408 14240 20460
rect 18696 20451 18748 20460
rect 18696 20417 18705 20451
rect 18705 20417 18739 20451
rect 18739 20417 18748 20451
rect 18696 20408 18748 20417
rect 19708 20408 19760 20460
rect 19984 20408 20036 20460
rect 27528 20544 27580 20596
rect 28172 20544 28224 20596
rect 28356 20544 28408 20596
rect 28908 20476 28960 20528
rect 29460 20476 29512 20528
rect 10876 20340 10928 20392
rect 11244 20383 11296 20392
rect 11244 20349 11253 20383
rect 11253 20349 11287 20383
rect 11287 20349 11296 20383
rect 11244 20340 11296 20349
rect 3700 20315 3752 20324
rect 3700 20281 3709 20315
rect 3709 20281 3743 20315
rect 3743 20281 3752 20315
rect 3700 20272 3752 20281
rect 11060 20272 11112 20324
rect 5816 20204 5868 20256
rect 7288 20204 7340 20256
rect 7472 20204 7524 20256
rect 9128 20204 9180 20256
rect 10508 20204 10560 20256
rect 12072 20340 12124 20392
rect 14004 20272 14056 20324
rect 16672 20340 16724 20392
rect 18052 20340 18104 20392
rect 18880 20383 18932 20392
rect 18880 20349 18889 20383
rect 18889 20349 18923 20383
rect 18923 20349 18932 20383
rect 18880 20340 18932 20349
rect 14832 20272 14884 20324
rect 11612 20204 11664 20256
rect 13084 20247 13136 20256
rect 13084 20213 13093 20247
rect 13093 20213 13127 20247
rect 13127 20213 13136 20247
rect 13084 20204 13136 20213
rect 14464 20204 14516 20256
rect 15384 20204 15436 20256
rect 16120 20272 16172 20324
rect 17500 20247 17552 20256
rect 17500 20213 17509 20247
rect 17509 20213 17543 20247
rect 17543 20213 17552 20247
rect 17500 20204 17552 20213
rect 17868 20204 17920 20256
rect 21272 20340 21324 20392
rect 21548 20383 21600 20392
rect 21548 20349 21557 20383
rect 21557 20349 21591 20383
rect 21591 20349 21600 20383
rect 21548 20340 21600 20349
rect 23388 20383 23440 20392
rect 23388 20349 23410 20383
rect 23410 20349 23440 20383
rect 23388 20340 23440 20349
rect 25136 20340 25188 20392
rect 26700 20451 26752 20460
rect 26700 20417 26709 20451
rect 26709 20417 26743 20451
rect 26743 20417 26752 20451
rect 26700 20408 26752 20417
rect 26884 20408 26936 20460
rect 22100 20272 22152 20324
rect 23112 20272 23164 20324
rect 23756 20272 23808 20324
rect 21364 20204 21416 20256
rect 24768 20204 24820 20256
rect 25688 20247 25740 20256
rect 25688 20213 25697 20247
rect 25697 20213 25731 20247
rect 25731 20213 25740 20247
rect 25688 20204 25740 20213
rect 26332 20204 26384 20256
rect 27528 20204 27580 20256
rect 29276 20340 29328 20392
rect 29460 20383 29512 20392
rect 29460 20349 29469 20383
rect 29469 20349 29503 20383
rect 29503 20349 29512 20383
rect 29460 20340 29512 20349
rect 29920 20340 29972 20392
rect 29092 20315 29144 20324
rect 29092 20281 29101 20315
rect 29101 20281 29135 20315
rect 29135 20281 29144 20315
rect 29092 20272 29144 20281
rect 30104 20315 30156 20324
rect 30104 20281 30113 20315
rect 30113 20281 30147 20315
rect 30147 20281 30156 20315
rect 30104 20272 30156 20281
rect 29460 20204 29512 20256
rect 29552 20204 29604 20256
rect 7988 20102 8040 20154
rect 8052 20102 8104 20154
rect 8116 20102 8168 20154
rect 8180 20102 8232 20154
rect 8244 20102 8296 20154
rect 15578 20102 15630 20154
rect 15642 20102 15694 20154
rect 15706 20102 15758 20154
rect 15770 20102 15822 20154
rect 15834 20102 15886 20154
rect 23168 20102 23220 20154
rect 23232 20102 23284 20154
rect 23296 20102 23348 20154
rect 23360 20102 23412 20154
rect 23424 20102 23476 20154
rect 30758 20102 30810 20154
rect 30822 20102 30874 20154
rect 30886 20102 30938 20154
rect 30950 20102 31002 20154
rect 31014 20102 31066 20154
rect 1308 20000 1360 20052
rect 1768 20000 1820 20052
rect 4068 20000 4120 20052
rect 5816 20000 5868 20052
rect 7472 20000 7524 20052
rect 848 19796 900 19848
rect 3148 19864 3200 19916
rect 3608 19864 3660 19916
rect 3884 19907 3936 19916
rect 3884 19873 3886 19907
rect 3886 19873 3936 19907
rect 5908 19932 5960 19984
rect 13084 20000 13136 20052
rect 17500 20000 17552 20052
rect 18880 20000 18932 20052
rect 21272 20000 21324 20052
rect 21824 20043 21876 20052
rect 21824 20009 21833 20043
rect 21833 20009 21867 20043
rect 21867 20009 21876 20043
rect 21824 20000 21876 20009
rect 23940 20000 23992 20052
rect 8392 19932 8444 19984
rect 10600 19975 10652 19984
rect 10600 19941 10609 19975
rect 10609 19941 10643 19975
rect 10643 19941 10652 19975
rect 10600 19932 10652 19941
rect 3884 19864 3936 19873
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 3332 19796 3384 19848
rect 4068 19796 4120 19848
rect 5172 19796 5224 19848
rect 5448 19796 5500 19848
rect 6460 19796 6512 19848
rect 8392 19796 8444 19848
rect 8484 19839 8536 19848
rect 8484 19805 8493 19839
rect 8493 19805 8527 19839
rect 8527 19805 8536 19839
rect 8484 19796 8536 19805
rect 9036 19864 9088 19916
rect 11336 19864 11388 19916
rect 12072 19932 12124 19984
rect 8944 19839 8996 19848
rect 8944 19805 8956 19839
rect 8956 19805 8990 19839
rect 8990 19805 8996 19839
rect 8944 19796 8996 19805
rect 9220 19839 9272 19848
rect 9220 19805 9229 19839
rect 9229 19805 9263 19839
rect 9263 19805 9272 19839
rect 9220 19796 9272 19805
rect 11980 19796 12032 19848
rect 12440 19839 12492 19848
rect 12440 19805 12442 19839
rect 12442 19805 12492 19839
rect 12440 19796 12492 19805
rect 12716 19796 12768 19848
rect 12808 19839 12860 19848
rect 12808 19805 12817 19839
rect 12817 19805 12851 19839
rect 12851 19805 12860 19839
rect 12808 19796 12860 19805
rect 14188 19864 14240 19916
rect 15384 19864 15436 19916
rect 20996 19932 21048 19984
rect 21916 19932 21968 19984
rect 23756 19932 23808 19984
rect 25136 20000 25188 20052
rect 27344 20000 27396 20052
rect 17960 19864 18012 19916
rect 20628 19864 20680 19916
rect 20904 19864 20956 19916
rect 21364 19907 21416 19916
rect 21364 19873 21373 19907
rect 21373 19873 21407 19907
rect 21407 19873 21416 19907
rect 21364 19864 21416 19873
rect 21456 19864 21508 19916
rect 21548 19864 21600 19916
rect 22192 19907 22244 19916
rect 22192 19873 22201 19907
rect 22201 19873 22235 19907
rect 22235 19873 22244 19907
rect 22192 19864 22244 19873
rect 15936 19796 15988 19848
rect 17224 19796 17276 19848
rect 17868 19839 17920 19848
rect 17868 19805 17877 19839
rect 17877 19805 17911 19839
rect 17911 19805 17920 19839
rect 17868 19796 17920 19805
rect 18236 19796 18288 19848
rect 8300 19703 8352 19712
rect 8300 19669 8309 19703
rect 8309 19669 8343 19703
rect 8343 19669 8352 19703
rect 8300 19660 8352 19669
rect 23480 19728 23532 19780
rect 26240 19864 26292 19916
rect 27896 19932 27948 19984
rect 28356 19907 28408 19916
rect 28356 19873 28365 19907
rect 28365 19873 28399 19907
rect 28399 19873 28408 19907
rect 28356 19864 28408 19873
rect 24400 19839 24452 19848
rect 24400 19805 24409 19839
rect 24409 19805 24443 19839
rect 24443 19805 24452 19839
rect 24400 19796 24452 19805
rect 25964 19796 26016 19848
rect 26424 19728 26476 19780
rect 8668 19660 8720 19712
rect 13728 19660 13780 19712
rect 13912 19703 13964 19712
rect 13912 19669 13921 19703
rect 13921 19669 13955 19703
rect 13955 19669 13964 19703
rect 13912 19660 13964 19669
rect 15844 19703 15896 19712
rect 15844 19669 15853 19703
rect 15853 19669 15887 19703
rect 15887 19669 15896 19703
rect 15844 19660 15896 19669
rect 18144 19660 18196 19712
rect 19156 19660 19208 19712
rect 21272 19660 21324 19712
rect 21548 19660 21600 19712
rect 22652 19660 22704 19712
rect 23572 19660 23624 19712
rect 28448 19839 28500 19848
rect 28448 19805 28457 19839
rect 28457 19805 28491 19839
rect 28491 19805 28500 19839
rect 28448 19796 28500 19805
rect 28816 19839 28868 19848
rect 28816 19805 28818 19839
rect 28818 19805 28868 19839
rect 28816 19796 28868 19805
rect 29644 19796 29696 19848
rect 4193 19558 4245 19610
rect 4257 19558 4309 19610
rect 4321 19558 4373 19610
rect 4385 19558 4437 19610
rect 4449 19558 4501 19610
rect 11783 19558 11835 19610
rect 11847 19558 11899 19610
rect 11911 19558 11963 19610
rect 11975 19558 12027 19610
rect 12039 19558 12091 19610
rect 19373 19558 19425 19610
rect 19437 19558 19489 19610
rect 19501 19558 19553 19610
rect 19565 19558 19617 19610
rect 19629 19558 19681 19610
rect 26963 19558 27015 19610
rect 27027 19558 27079 19610
rect 27091 19558 27143 19610
rect 27155 19558 27207 19610
rect 27219 19558 27271 19610
rect 2780 19499 2832 19508
rect 2780 19465 2789 19499
rect 2789 19465 2823 19499
rect 2823 19465 2832 19499
rect 2780 19456 2832 19465
rect 3332 19456 3384 19508
rect 5632 19456 5684 19508
rect 5724 19456 5776 19508
rect 5356 19388 5408 19440
rect 3056 19320 3108 19372
rect 3884 19363 3936 19372
rect 3884 19329 3893 19363
rect 3893 19329 3927 19363
rect 3927 19329 3936 19363
rect 3884 19320 3936 19329
rect 6000 19320 6052 19372
rect 8300 19456 8352 19508
rect 9588 19456 9640 19508
rect 10232 19499 10284 19508
rect 10232 19465 10241 19499
rect 10241 19465 10275 19499
rect 10275 19465 10284 19499
rect 10232 19456 10284 19465
rect 10692 19456 10744 19508
rect 13452 19456 13504 19508
rect 14004 19499 14056 19508
rect 14004 19465 14013 19499
rect 14013 19465 14047 19499
rect 14047 19465 14056 19499
rect 14004 19456 14056 19465
rect 6920 19388 6972 19440
rect 1032 19252 1084 19304
rect 2136 19252 2188 19304
rect 3608 19295 3660 19304
rect 3608 19261 3617 19295
rect 3617 19261 3651 19295
rect 3651 19261 3660 19295
rect 3608 19252 3660 19261
rect 4528 19252 4580 19304
rect 5448 19252 5500 19304
rect 6460 19252 6512 19304
rect 3884 19184 3936 19236
rect 1768 19116 1820 19168
rect 4804 19184 4856 19236
rect 7288 19252 7340 19304
rect 5724 19116 5776 19168
rect 5816 19159 5868 19168
rect 5816 19125 5831 19159
rect 5831 19125 5865 19159
rect 5865 19125 5868 19159
rect 5816 19116 5868 19125
rect 6736 19116 6788 19168
rect 7840 19184 7892 19236
rect 8576 19320 8628 19372
rect 8944 19320 8996 19372
rect 8668 19252 8720 19304
rect 9404 19252 9456 19304
rect 11060 19320 11112 19372
rect 14188 19363 14240 19372
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 14832 19320 14884 19372
rect 8484 19184 8536 19236
rect 9956 19184 10008 19236
rect 11980 19252 12032 19304
rect 13268 19252 13320 19304
rect 16120 19456 16172 19508
rect 15844 19320 15896 19372
rect 17776 19320 17828 19372
rect 15936 19295 15988 19304
rect 15936 19261 15945 19295
rect 15945 19261 15979 19295
rect 15979 19261 15988 19295
rect 15936 19252 15988 19261
rect 17224 19252 17276 19304
rect 17684 19252 17736 19304
rect 18236 19320 18288 19372
rect 23480 19456 23532 19508
rect 24400 19456 24452 19508
rect 26516 19456 26568 19508
rect 30104 19456 30156 19508
rect 21548 19388 21600 19440
rect 9128 19116 9180 19168
rect 11152 19116 11204 19168
rect 11428 19116 11480 19168
rect 12164 19116 12216 19168
rect 12532 19116 12584 19168
rect 12992 19159 13044 19168
rect 12992 19125 13001 19159
rect 13001 19125 13035 19159
rect 13035 19125 13044 19159
rect 12992 19116 13044 19125
rect 20444 19295 20496 19304
rect 20444 19261 20453 19295
rect 20453 19261 20487 19295
rect 20487 19261 20496 19295
rect 20444 19252 20496 19261
rect 20536 19252 20588 19304
rect 23572 19363 23624 19372
rect 23572 19329 23581 19363
rect 23581 19329 23615 19363
rect 23615 19329 23624 19363
rect 23572 19320 23624 19329
rect 26700 19363 26752 19372
rect 26700 19329 26709 19363
rect 26709 19329 26743 19363
rect 26743 19329 26752 19363
rect 26700 19320 26752 19329
rect 27344 19320 27396 19372
rect 28908 19320 28960 19372
rect 22836 19184 22888 19236
rect 23020 19252 23072 19304
rect 24492 19252 24544 19304
rect 27068 19295 27120 19304
rect 27068 19261 27070 19295
rect 27070 19261 27120 19295
rect 27068 19252 27120 19261
rect 23572 19184 23624 19236
rect 24124 19227 24176 19236
rect 24124 19193 24133 19227
rect 24133 19193 24167 19227
rect 24167 19193 24176 19227
rect 24124 19184 24176 19193
rect 24216 19184 24268 19236
rect 26516 19184 26568 19236
rect 16028 19116 16080 19168
rect 16304 19116 16356 19168
rect 20076 19159 20128 19168
rect 20076 19125 20085 19159
rect 20085 19125 20119 19159
rect 20119 19125 20128 19159
rect 20076 19116 20128 19125
rect 24492 19116 24544 19168
rect 25136 19116 25188 19168
rect 25504 19116 25556 19168
rect 26056 19116 26108 19168
rect 26608 19116 26660 19168
rect 29092 19184 29144 19236
rect 29920 19252 29972 19304
rect 29552 19184 29604 19236
rect 27712 19116 27764 19168
rect 28540 19159 28592 19168
rect 28540 19125 28549 19159
rect 28549 19125 28583 19159
rect 28583 19125 28592 19159
rect 28540 19116 28592 19125
rect 30012 19116 30064 19168
rect 30104 19159 30156 19168
rect 30104 19125 30113 19159
rect 30113 19125 30147 19159
rect 30147 19125 30156 19159
rect 30104 19116 30156 19125
rect 30656 19116 30708 19168
rect 7988 19014 8040 19066
rect 8052 19014 8104 19066
rect 8116 19014 8168 19066
rect 8180 19014 8232 19066
rect 8244 19014 8296 19066
rect 15578 19014 15630 19066
rect 15642 19014 15694 19066
rect 15706 19014 15758 19066
rect 15770 19014 15822 19066
rect 15834 19014 15886 19066
rect 23168 19014 23220 19066
rect 23232 19014 23284 19066
rect 23296 19014 23348 19066
rect 23360 19014 23412 19066
rect 23424 19014 23476 19066
rect 30758 19014 30810 19066
rect 30822 19014 30874 19066
rect 30886 19014 30938 19066
rect 30950 19014 31002 19066
rect 31014 19014 31066 19066
rect 1676 18912 1728 18964
rect 3148 18955 3200 18964
rect 3148 18921 3157 18955
rect 3157 18921 3191 18955
rect 3191 18921 3200 18955
rect 3148 18912 3200 18921
rect 1216 18819 1268 18828
rect 1216 18785 1225 18819
rect 1225 18785 1259 18819
rect 1259 18785 1268 18819
rect 1216 18776 1268 18785
rect 1124 18708 1176 18760
rect 2320 18776 2372 18828
rect 1032 18615 1084 18624
rect 1032 18581 1041 18615
rect 1041 18581 1075 18615
rect 1075 18581 1084 18615
rect 1032 18572 1084 18581
rect 1768 18572 1820 18624
rect 4712 18887 4764 18896
rect 4712 18853 4721 18887
rect 4721 18853 4755 18887
rect 4755 18853 4764 18887
rect 4712 18844 4764 18853
rect 5080 18887 5132 18896
rect 5080 18853 5089 18887
rect 5089 18853 5123 18887
rect 5123 18853 5132 18887
rect 5080 18844 5132 18853
rect 6828 18912 6880 18964
rect 11980 18912 12032 18964
rect 12348 18955 12400 18964
rect 12348 18921 12363 18955
rect 12363 18921 12397 18955
rect 12397 18921 12400 18955
rect 12348 18912 12400 18921
rect 13820 18912 13872 18964
rect 16028 18912 16080 18964
rect 17960 18912 18012 18964
rect 8576 18844 8628 18896
rect 10416 18844 10468 18896
rect 3884 18819 3936 18828
rect 3884 18785 3893 18819
rect 3893 18785 3927 18819
rect 3927 18785 3936 18819
rect 3884 18776 3936 18785
rect 5908 18776 5960 18828
rect 6092 18776 6144 18828
rect 8760 18776 8812 18828
rect 9036 18819 9088 18828
rect 9036 18785 9038 18819
rect 9038 18785 9088 18819
rect 9036 18776 9088 18785
rect 10876 18844 10928 18896
rect 6460 18751 6512 18760
rect 6460 18717 6472 18751
rect 6472 18717 6506 18751
rect 6506 18717 6512 18751
rect 6460 18708 6512 18717
rect 6736 18751 6788 18760
rect 6736 18717 6745 18751
rect 6745 18717 6779 18751
rect 6779 18717 6788 18751
rect 6736 18708 6788 18717
rect 3792 18615 3844 18624
rect 3792 18581 3801 18615
rect 3801 18581 3835 18615
rect 3835 18581 3844 18615
rect 3792 18572 3844 18581
rect 8484 18708 8536 18760
rect 8576 18708 8628 18760
rect 11336 18776 11388 18828
rect 9404 18751 9456 18760
rect 9404 18717 9413 18751
rect 9413 18717 9447 18751
rect 9447 18717 9456 18751
rect 9404 18708 9456 18717
rect 9496 18708 9548 18760
rect 8392 18640 8444 18692
rect 10508 18708 10560 18760
rect 11152 18751 11204 18760
rect 11152 18717 11161 18751
rect 11161 18717 11195 18751
rect 11195 18717 11204 18751
rect 11152 18708 11204 18717
rect 12532 18776 12584 18828
rect 12992 18776 13044 18828
rect 14556 18819 14608 18828
rect 14556 18785 14565 18819
rect 14565 18785 14599 18819
rect 14599 18785 14608 18819
rect 14556 18776 14608 18785
rect 15936 18776 15988 18828
rect 17224 18776 17276 18828
rect 18144 18819 18196 18828
rect 18144 18785 18153 18819
rect 18153 18785 18187 18819
rect 18187 18785 18196 18819
rect 18144 18776 18196 18785
rect 19892 18819 19944 18828
rect 19892 18785 19901 18819
rect 19901 18785 19935 18819
rect 19935 18785 19944 18819
rect 19892 18776 19944 18785
rect 20628 18912 20680 18964
rect 22836 18912 22888 18964
rect 23664 18912 23716 18964
rect 25228 18912 25280 18964
rect 25320 18912 25372 18964
rect 28540 18912 28592 18964
rect 28816 18912 28868 18964
rect 29276 18912 29328 18964
rect 25596 18844 25648 18896
rect 20444 18776 20496 18828
rect 20628 18776 20680 18828
rect 11796 18640 11848 18692
rect 9404 18572 9456 18624
rect 15844 18708 15896 18760
rect 12624 18572 12676 18624
rect 19708 18708 19760 18760
rect 24400 18776 24452 18828
rect 21272 18751 21324 18760
rect 21272 18717 21281 18751
rect 21281 18717 21315 18751
rect 21315 18717 21324 18751
rect 21272 18708 21324 18717
rect 21548 18751 21600 18760
rect 21548 18717 21557 18751
rect 21557 18717 21591 18751
rect 21591 18717 21600 18751
rect 21548 18708 21600 18717
rect 24124 18751 24176 18760
rect 24124 18717 24133 18751
rect 24133 18717 24167 18751
rect 24167 18717 24176 18751
rect 24124 18708 24176 18717
rect 24308 18708 24360 18760
rect 25964 18776 26016 18828
rect 26516 18776 26568 18828
rect 24860 18751 24912 18760
rect 24860 18717 24869 18751
rect 24869 18717 24903 18751
rect 24903 18717 24912 18751
rect 24860 18708 24912 18717
rect 25228 18708 25280 18760
rect 26240 18708 26292 18760
rect 18880 18640 18932 18692
rect 19064 18572 19116 18624
rect 20444 18640 20496 18692
rect 20996 18572 21048 18624
rect 25596 18640 25648 18692
rect 27620 18708 27672 18760
rect 24768 18572 24820 18624
rect 24860 18572 24912 18624
rect 25872 18572 25924 18624
rect 25964 18615 26016 18624
rect 25964 18581 25973 18615
rect 25973 18581 26007 18615
rect 26007 18581 26016 18615
rect 25964 18572 26016 18581
rect 26056 18572 26108 18624
rect 28448 18819 28500 18828
rect 28448 18785 28457 18819
rect 28457 18785 28491 18819
rect 28491 18785 28500 18819
rect 28448 18776 28500 18785
rect 29276 18776 29328 18828
rect 30012 18776 30064 18828
rect 28908 18751 28960 18760
rect 28908 18717 28920 18751
rect 28920 18717 28954 18751
rect 28954 18717 28960 18751
rect 28908 18708 28960 18717
rect 29184 18751 29236 18760
rect 29184 18717 29193 18751
rect 29193 18717 29227 18751
rect 29227 18717 29236 18751
rect 29184 18708 29236 18717
rect 28356 18615 28408 18624
rect 28356 18581 28365 18615
rect 28365 18581 28399 18615
rect 28399 18581 28408 18615
rect 28356 18572 28408 18581
rect 4193 18470 4245 18522
rect 4257 18470 4309 18522
rect 4321 18470 4373 18522
rect 4385 18470 4437 18522
rect 4449 18470 4501 18522
rect 11783 18470 11835 18522
rect 11847 18470 11899 18522
rect 11911 18470 11963 18522
rect 11975 18470 12027 18522
rect 12039 18470 12091 18522
rect 19373 18470 19425 18522
rect 19437 18470 19489 18522
rect 19501 18470 19553 18522
rect 19565 18470 19617 18522
rect 19629 18470 19681 18522
rect 26963 18470 27015 18522
rect 27027 18470 27079 18522
rect 27091 18470 27143 18522
rect 27155 18470 27207 18522
rect 27219 18470 27271 18522
rect 1124 18368 1176 18420
rect 848 18232 900 18284
rect 2688 18232 2740 18284
rect 4068 18368 4120 18420
rect 4160 18368 4212 18420
rect 3424 18300 3476 18352
rect 4068 18232 4120 18284
rect 3332 18207 3384 18216
rect 3332 18173 3341 18207
rect 3341 18173 3375 18207
rect 3375 18173 3384 18207
rect 3332 18164 3384 18173
rect 3700 18164 3752 18216
rect 4620 18207 4672 18216
rect 4620 18173 4629 18207
rect 4629 18173 4663 18207
rect 4663 18173 4672 18207
rect 4620 18164 4672 18173
rect 5632 18164 5684 18216
rect 6460 18368 6512 18420
rect 9772 18368 9824 18420
rect 11060 18368 11112 18420
rect 8208 18300 8260 18352
rect 13360 18368 13412 18420
rect 13544 18300 13596 18352
rect 6000 18232 6052 18284
rect 9036 18275 9088 18284
rect 9036 18241 9048 18275
rect 9048 18241 9082 18275
rect 9082 18241 9088 18275
rect 9036 18232 9088 18241
rect 11060 18232 11112 18284
rect 5908 18164 5960 18216
rect 5356 18096 5408 18148
rect 8576 18207 8628 18216
rect 8576 18173 8585 18207
rect 8585 18173 8619 18207
rect 8619 18173 8628 18207
rect 8576 18164 8628 18173
rect 9312 18207 9364 18216
rect 9312 18173 9321 18207
rect 9321 18173 9355 18207
rect 9355 18173 9364 18207
rect 9312 18164 9364 18173
rect 10968 18207 11020 18216
rect 10968 18173 10977 18207
rect 10977 18173 11011 18207
rect 11011 18173 11020 18207
rect 10968 18164 11020 18173
rect 11244 18207 11296 18216
rect 11244 18173 11253 18207
rect 11253 18173 11287 18207
rect 11287 18173 11296 18207
rect 11244 18164 11296 18173
rect 11520 18164 11572 18216
rect 13820 18164 13872 18216
rect 13912 18164 13964 18216
rect 15016 18232 15068 18284
rect 15384 18232 15436 18284
rect 15844 18232 15896 18284
rect 17040 18232 17092 18284
rect 20076 18368 20128 18420
rect 20536 18368 20588 18420
rect 19708 18300 19760 18352
rect 21180 18368 21232 18420
rect 21732 18368 21784 18420
rect 26884 18368 26936 18420
rect 8392 18096 8444 18148
rect 11152 18139 11204 18148
rect 11152 18105 11161 18139
rect 11161 18105 11195 18139
rect 11195 18105 11204 18139
rect 11152 18096 11204 18105
rect 13176 18096 13228 18148
rect 15292 18164 15344 18216
rect 18052 18164 18104 18216
rect 18880 18232 18932 18284
rect 19064 18232 19116 18284
rect 20812 18232 20864 18284
rect 20720 18164 20772 18216
rect 24584 18343 24636 18352
rect 24584 18309 24593 18343
rect 24593 18309 24627 18343
rect 24627 18309 24636 18343
rect 24584 18300 24636 18309
rect 27068 18300 27120 18352
rect 22652 18232 22704 18284
rect 22928 18164 22980 18216
rect 24492 18232 24544 18284
rect 25044 18232 25096 18284
rect 25964 18232 26016 18284
rect 26240 18232 26292 18284
rect 26516 18232 26568 18284
rect 29552 18300 29604 18352
rect 23664 18164 23716 18216
rect 24860 18207 24912 18216
rect 24860 18173 24869 18207
rect 24869 18173 24903 18207
rect 24903 18173 24912 18207
rect 24860 18164 24912 18173
rect 1676 18028 1728 18080
rect 3148 18028 3200 18080
rect 4528 18028 4580 18080
rect 6092 18028 6144 18080
rect 6828 18028 6880 18080
rect 9036 18071 9088 18080
rect 9036 18037 9051 18071
rect 9051 18037 9085 18071
rect 9085 18037 9088 18071
rect 9036 18028 9088 18037
rect 9588 18028 9640 18080
rect 11336 18028 11388 18080
rect 11612 18028 11664 18080
rect 12072 18028 12124 18080
rect 12716 18028 12768 18080
rect 12992 18028 13044 18080
rect 14280 18028 14332 18080
rect 15108 18028 15160 18080
rect 24400 18139 24452 18148
rect 24400 18105 24409 18139
rect 24409 18105 24443 18139
rect 24443 18105 24452 18139
rect 24400 18096 24452 18105
rect 24768 18096 24820 18148
rect 19340 18028 19392 18080
rect 21456 18028 21508 18080
rect 21824 18028 21876 18080
rect 24032 18028 24084 18080
rect 25504 18164 25556 18216
rect 25228 18028 25280 18080
rect 26700 18071 26752 18080
rect 26700 18037 26709 18071
rect 26709 18037 26743 18071
rect 26743 18037 26752 18071
rect 26700 18028 26752 18037
rect 27068 18207 27120 18216
rect 27068 18173 27077 18207
rect 27077 18173 27111 18207
rect 27111 18173 27120 18207
rect 27068 18164 27120 18173
rect 27160 18164 27212 18216
rect 27620 18164 27672 18216
rect 28448 18071 28500 18080
rect 28448 18037 28457 18071
rect 28457 18037 28491 18071
rect 28491 18037 28500 18071
rect 28448 18028 28500 18037
rect 29368 18096 29420 18148
rect 29920 18096 29972 18148
rect 30104 18071 30156 18080
rect 30104 18037 30113 18071
rect 30113 18037 30147 18071
rect 30147 18037 30156 18071
rect 30104 18028 30156 18037
rect 30196 18028 30248 18080
rect 30380 18071 30432 18080
rect 30380 18037 30389 18071
rect 30389 18037 30423 18071
rect 30423 18037 30432 18071
rect 30380 18028 30432 18037
rect 30656 18028 30708 18080
rect 7988 17926 8040 17978
rect 8052 17926 8104 17978
rect 8116 17926 8168 17978
rect 8180 17926 8232 17978
rect 8244 17926 8296 17978
rect 15578 17926 15630 17978
rect 15642 17926 15694 17978
rect 15706 17926 15758 17978
rect 15770 17926 15822 17978
rect 15834 17926 15886 17978
rect 23168 17926 23220 17978
rect 23232 17926 23284 17978
rect 23296 17926 23348 17978
rect 23360 17926 23412 17978
rect 23424 17926 23476 17978
rect 30758 17926 30810 17978
rect 30822 17926 30874 17978
rect 30886 17926 30938 17978
rect 30950 17926 31002 17978
rect 31014 17926 31066 17978
rect 1124 17756 1176 17808
rect 3148 17867 3200 17876
rect 3148 17833 3157 17867
rect 3157 17833 3191 17867
rect 3191 17833 3200 17867
rect 3148 17824 3200 17833
rect 4528 17824 4580 17876
rect 6828 17824 6880 17876
rect 1676 17731 1728 17740
rect 1676 17697 1678 17731
rect 1678 17697 1728 17731
rect 1676 17688 1728 17697
rect 3148 17688 3200 17740
rect 2044 17663 2096 17672
rect 2044 17629 2053 17663
rect 2053 17629 2087 17663
rect 2087 17629 2096 17663
rect 2044 17620 2096 17629
rect 3240 17484 3292 17536
rect 6000 17756 6052 17808
rect 3700 17620 3752 17672
rect 6552 17688 6604 17740
rect 12072 17824 12124 17876
rect 12256 17824 12308 17876
rect 12808 17824 12860 17876
rect 14280 17867 14332 17876
rect 14280 17833 14295 17867
rect 14295 17833 14329 17867
rect 14329 17833 14332 17867
rect 14280 17824 14332 17833
rect 15384 17824 15436 17876
rect 16120 17824 16172 17876
rect 10784 17799 10836 17808
rect 10784 17765 10793 17799
rect 10793 17765 10827 17799
rect 10827 17765 10836 17799
rect 10784 17756 10836 17765
rect 15568 17756 15620 17808
rect 16580 17824 16632 17876
rect 5264 17620 5316 17672
rect 5816 17620 5868 17672
rect 6368 17620 6420 17672
rect 6460 17663 6512 17672
rect 6460 17629 6469 17663
rect 6469 17629 6503 17663
rect 6503 17629 6512 17663
rect 6460 17620 6512 17629
rect 6920 17663 6972 17672
rect 6920 17629 6932 17663
rect 6932 17629 6966 17663
rect 6966 17629 6972 17663
rect 6920 17620 6972 17629
rect 8668 17663 8720 17672
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 9036 17663 9088 17672
rect 9036 17629 9038 17663
rect 9038 17629 9088 17663
rect 9036 17620 9088 17629
rect 10324 17688 10376 17740
rect 11612 17731 11664 17740
rect 11612 17697 11614 17731
rect 11614 17697 11664 17731
rect 9404 17663 9456 17672
rect 9404 17629 9413 17663
rect 9413 17629 9447 17663
rect 9447 17629 9456 17663
rect 9404 17620 9456 17629
rect 9864 17484 9916 17536
rect 10968 17527 11020 17536
rect 10968 17493 10977 17527
rect 10977 17493 11011 17527
rect 11011 17493 11020 17527
rect 10968 17484 11020 17493
rect 11612 17688 11664 17697
rect 11244 17663 11296 17672
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 11888 17620 11940 17672
rect 12072 17620 12124 17672
rect 12900 17620 12952 17672
rect 13268 17688 13320 17740
rect 12992 17484 13044 17536
rect 13084 17527 13136 17536
rect 13084 17493 13093 17527
rect 13093 17493 13127 17527
rect 13127 17493 13136 17527
rect 13084 17484 13136 17493
rect 13636 17527 13688 17536
rect 13636 17493 13645 17527
rect 13645 17493 13679 17527
rect 13679 17493 13688 17527
rect 13636 17484 13688 17493
rect 13820 17663 13872 17672
rect 13820 17629 13829 17663
rect 13829 17629 13863 17663
rect 13863 17629 13872 17663
rect 13820 17620 13872 17629
rect 16120 17688 16172 17740
rect 16580 17731 16632 17740
rect 16580 17697 16589 17731
rect 16589 17697 16623 17731
rect 16623 17697 16632 17731
rect 16580 17688 16632 17697
rect 17776 17824 17828 17876
rect 21640 17824 21692 17876
rect 23020 17824 23072 17876
rect 24584 17824 24636 17876
rect 24768 17824 24820 17876
rect 27436 17824 27488 17876
rect 28816 17867 28868 17876
rect 16672 17620 16724 17672
rect 17040 17620 17092 17672
rect 17500 17663 17552 17672
rect 17500 17629 17502 17663
rect 17502 17629 17552 17663
rect 17500 17620 17552 17629
rect 19340 17688 19392 17740
rect 23664 17731 23716 17740
rect 23664 17697 23673 17731
rect 23673 17697 23707 17731
rect 23707 17697 23716 17731
rect 23664 17688 23716 17697
rect 23756 17688 23808 17740
rect 17868 17663 17920 17672
rect 17868 17629 17877 17663
rect 17877 17629 17911 17663
rect 17911 17629 17920 17663
rect 17868 17620 17920 17629
rect 20444 17620 20496 17672
rect 20720 17620 20772 17672
rect 15476 17484 15528 17536
rect 17592 17484 17644 17536
rect 21456 17620 21508 17672
rect 21916 17620 21968 17672
rect 23572 17620 23624 17672
rect 24492 17663 24544 17672
rect 24492 17629 24494 17663
rect 24494 17629 24544 17663
rect 24492 17620 24544 17629
rect 24676 17620 24728 17672
rect 24860 17663 24912 17672
rect 24860 17629 24869 17663
rect 24869 17629 24903 17663
rect 24903 17629 24912 17663
rect 24860 17620 24912 17629
rect 25044 17620 25096 17672
rect 26424 17663 26476 17672
rect 26424 17629 26433 17663
rect 26433 17629 26467 17663
rect 26467 17629 26476 17663
rect 26424 17620 26476 17629
rect 27344 17620 27396 17672
rect 28816 17833 28831 17867
rect 28831 17833 28865 17867
rect 28865 17833 28868 17867
rect 28816 17824 28868 17833
rect 29000 17824 29052 17876
rect 28540 17620 28592 17672
rect 29736 17620 29788 17672
rect 29920 17620 29972 17672
rect 22008 17484 22060 17536
rect 22744 17484 22796 17536
rect 25504 17484 25556 17536
rect 26424 17484 26476 17536
rect 29276 17484 29328 17536
rect 30104 17484 30156 17536
rect 4193 17382 4245 17434
rect 4257 17382 4309 17434
rect 4321 17382 4373 17434
rect 4385 17382 4437 17434
rect 4449 17382 4501 17434
rect 11783 17382 11835 17434
rect 11847 17382 11899 17434
rect 11911 17382 11963 17434
rect 11975 17382 12027 17434
rect 12039 17382 12091 17434
rect 19373 17382 19425 17434
rect 19437 17382 19489 17434
rect 19501 17382 19553 17434
rect 19565 17382 19617 17434
rect 19629 17382 19681 17434
rect 26963 17382 27015 17434
rect 27027 17382 27079 17434
rect 27091 17382 27143 17434
rect 27155 17382 27207 17434
rect 27219 17382 27271 17434
rect 1584 17280 1636 17332
rect 3240 17280 3292 17332
rect 3700 17212 3752 17264
rect 1124 17144 1176 17196
rect 2780 17144 2832 17196
rect 4068 17144 4120 17196
rect 5540 17144 5592 17196
rect 2412 17076 2464 17128
rect 3240 17119 3292 17128
rect 3240 17085 3249 17119
rect 3249 17085 3283 17119
rect 3283 17085 3292 17119
rect 3240 17076 3292 17085
rect 5080 17076 5132 17128
rect 6920 17280 6972 17332
rect 8484 17280 8536 17332
rect 5908 17144 5960 17196
rect 6460 17144 6512 17196
rect 6552 17187 6604 17196
rect 6552 17153 6564 17187
rect 6564 17153 6598 17187
rect 6598 17153 6604 17187
rect 6552 17144 6604 17153
rect 8392 17144 8444 17196
rect 7472 17076 7524 17128
rect 10232 17280 10284 17332
rect 10508 17323 10560 17332
rect 10508 17289 10517 17323
rect 10517 17289 10551 17323
rect 10551 17289 10560 17323
rect 10508 17280 10560 17289
rect 8668 17187 8720 17196
rect 8668 17153 8677 17187
rect 8677 17153 8711 17187
rect 8711 17153 8720 17187
rect 8668 17144 8720 17153
rect 9036 17187 9088 17196
rect 9036 17153 9038 17187
rect 9038 17153 9088 17187
rect 9036 17144 9088 17153
rect 9128 17144 9180 17196
rect 9588 17144 9640 17196
rect 11520 17280 11572 17332
rect 11704 17280 11756 17332
rect 15200 17280 15252 17332
rect 13268 17212 13320 17264
rect 14464 17212 14516 17264
rect 15384 17212 15436 17264
rect 11796 17144 11848 17196
rect 1768 16940 1820 16992
rect 4528 16940 4580 16992
rect 4988 16940 5040 16992
rect 6828 16940 6880 16992
rect 10968 17119 11020 17128
rect 10968 17085 10977 17119
rect 10977 17085 11011 17119
rect 11011 17085 11020 17119
rect 10968 17076 11020 17085
rect 11244 17119 11296 17128
rect 11244 17085 11253 17119
rect 11253 17085 11287 17119
rect 11287 17085 11296 17119
rect 11244 17076 11296 17085
rect 11980 17119 12032 17128
rect 11980 17085 11989 17119
rect 11989 17085 12023 17119
rect 12023 17085 12032 17119
rect 11980 17076 12032 17085
rect 14004 17076 14056 17128
rect 14096 17076 14148 17128
rect 21548 17280 21600 17332
rect 22100 17280 22152 17332
rect 10140 17008 10192 17060
rect 10784 17008 10836 17060
rect 9496 16940 9548 16992
rect 11060 16940 11112 16992
rect 11612 16940 11664 16992
rect 12072 16940 12124 16992
rect 14648 17008 14700 17060
rect 15016 17076 15068 17128
rect 14924 17008 14976 17060
rect 15936 17076 15988 17128
rect 15200 17008 15252 17060
rect 17040 17076 17092 17128
rect 17132 17119 17184 17128
rect 17132 17085 17141 17119
rect 17141 17085 17175 17119
rect 17175 17085 17184 17119
rect 17132 17076 17184 17085
rect 18788 17076 18840 17128
rect 19156 17144 19208 17196
rect 12716 16940 12768 16992
rect 13268 16940 13320 16992
rect 15568 16940 15620 16992
rect 16488 17008 16540 17060
rect 20720 17076 20772 17128
rect 21272 17144 21324 17196
rect 23664 17212 23716 17264
rect 24124 17212 24176 17264
rect 24216 17212 24268 17264
rect 22284 17144 22336 17196
rect 23020 17144 23072 17196
rect 23756 17144 23808 17196
rect 21824 17076 21876 17128
rect 22008 17076 22060 17128
rect 23664 17076 23716 17128
rect 24676 17212 24728 17264
rect 28356 17212 28408 17264
rect 29552 17212 29604 17264
rect 24492 17144 24544 17196
rect 25228 17187 25280 17196
rect 25228 17153 25230 17187
rect 25230 17153 25280 17187
rect 25228 17144 25280 17153
rect 25320 17187 25372 17196
rect 25320 17153 25332 17187
rect 25332 17153 25366 17187
rect 25366 17153 25372 17187
rect 25320 17144 25372 17153
rect 25504 17144 25556 17196
rect 28448 17144 28500 17196
rect 24860 17119 24912 17128
rect 24860 17085 24869 17119
rect 24869 17085 24903 17119
rect 24903 17085 24912 17119
rect 24860 17076 24912 17085
rect 26424 17076 26476 17128
rect 28724 17051 28776 17060
rect 28724 17017 28733 17051
rect 28733 17017 28767 17051
rect 28767 17017 28776 17051
rect 28724 17008 28776 17017
rect 17500 16940 17552 16992
rect 19892 16940 19944 16992
rect 21456 16940 21508 16992
rect 21824 16940 21876 16992
rect 22008 16940 22060 16992
rect 22468 16983 22520 16992
rect 22468 16949 22477 16983
rect 22477 16949 22511 16983
rect 22511 16949 22520 16983
rect 22468 16940 22520 16949
rect 23572 16940 23624 16992
rect 23848 16983 23900 16992
rect 23848 16949 23857 16983
rect 23857 16949 23891 16983
rect 23891 16949 23900 16983
rect 23848 16940 23900 16949
rect 25596 16940 25648 16992
rect 27988 16940 28040 16992
rect 28632 16940 28684 16992
rect 30012 17008 30064 17060
rect 29276 16940 29328 16992
rect 29552 16940 29604 16992
rect 30380 16983 30432 16992
rect 30380 16949 30389 16983
rect 30389 16949 30423 16983
rect 30423 16949 30432 16983
rect 30380 16940 30432 16949
rect 7988 16838 8040 16890
rect 8052 16838 8104 16890
rect 8116 16838 8168 16890
rect 8180 16838 8232 16890
rect 8244 16838 8296 16890
rect 15578 16838 15630 16890
rect 15642 16838 15694 16890
rect 15706 16838 15758 16890
rect 15770 16838 15822 16890
rect 15834 16838 15886 16890
rect 23168 16838 23220 16890
rect 23232 16838 23284 16890
rect 23296 16838 23348 16890
rect 23360 16838 23412 16890
rect 23424 16838 23476 16890
rect 30758 16838 30810 16890
rect 30822 16838 30874 16890
rect 30886 16838 30938 16890
rect 30950 16838 31002 16890
rect 31014 16838 31066 16890
rect 1032 16736 1084 16788
rect 1860 16736 1912 16788
rect 3056 16779 3108 16788
rect 3056 16745 3065 16779
rect 3065 16745 3099 16779
rect 3099 16745 3108 16779
rect 3056 16736 3108 16745
rect 6552 16736 6604 16788
rect 9956 16736 10008 16788
rect 10876 16736 10928 16788
rect 11888 16779 11940 16788
rect 1308 16668 1360 16720
rect 5632 16711 5684 16720
rect 5632 16677 5641 16711
rect 5641 16677 5675 16711
rect 5675 16677 5684 16711
rect 5632 16668 5684 16677
rect 7380 16668 7432 16720
rect 7840 16668 7892 16720
rect 1124 16643 1176 16652
rect 1124 16609 1133 16643
rect 1133 16609 1167 16643
rect 1167 16609 1176 16643
rect 1124 16600 1176 16609
rect 4068 16600 4120 16652
rect 1216 16575 1268 16584
rect 1216 16541 1225 16575
rect 1225 16541 1259 16575
rect 1259 16541 1268 16575
rect 1216 16532 1268 16541
rect 1584 16575 1636 16584
rect 1584 16541 1586 16575
rect 1586 16541 1636 16575
rect 1584 16532 1636 16541
rect 1768 16532 1820 16584
rect 1860 16532 1912 16584
rect 3516 16575 3568 16584
rect 3516 16541 3525 16575
rect 3525 16541 3559 16575
rect 3559 16541 3568 16575
rect 3516 16532 3568 16541
rect 3884 16575 3936 16584
rect 3884 16541 3886 16575
rect 3886 16541 3936 16575
rect 3884 16532 3936 16541
rect 3976 16575 4028 16584
rect 3976 16541 3988 16575
rect 3988 16541 4022 16575
rect 4022 16541 4028 16575
rect 4712 16600 4764 16652
rect 4988 16600 5040 16652
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 7472 16600 7524 16652
rect 3976 16532 4028 16541
rect 6368 16532 6420 16584
rect 7012 16532 7064 16584
rect 8116 16532 8168 16584
rect 8668 16600 8720 16652
rect 9220 16600 9272 16652
rect 9956 16600 10008 16652
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 12900 16736 12952 16788
rect 15200 16736 15252 16788
rect 15476 16736 15528 16788
rect 15936 16736 15988 16788
rect 16672 16779 16724 16788
rect 16672 16745 16681 16779
rect 16681 16745 16715 16779
rect 16715 16745 16724 16779
rect 16672 16736 16724 16745
rect 11336 16668 11388 16720
rect 12440 16668 12492 16720
rect 11980 16600 12032 16652
rect 12072 16643 12124 16652
rect 12072 16609 12081 16643
rect 12081 16609 12115 16643
rect 12115 16609 12124 16643
rect 12072 16600 12124 16609
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 12992 16600 13044 16652
rect 13268 16600 13320 16652
rect 16120 16668 16172 16720
rect 15568 16600 15620 16652
rect 16304 16600 16356 16652
rect 16856 16643 16908 16652
rect 8944 16575 8996 16584
rect 8944 16541 8946 16575
rect 8946 16541 8996 16575
rect 8944 16532 8996 16541
rect 9496 16532 9548 16584
rect 9680 16532 9732 16584
rect 10048 16532 10100 16584
rect 11704 16532 11756 16584
rect 13820 16575 13872 16584
rect 13820 16541 13837 16575
rect 13837 16541 13871 16575
rect 13871 16541 13872 16575
rect 14188 16575 14240 16584
rect 13820 16532 13872 16541
rect 14188 16541 14190 16575
rect 14190 16541 14240 16575
rect 14188 16532 14240 16541
rect 15016 16532 15068 16584
rect 16856 16609 16865 16643
rect 16865 16609 16899 16643
rect 16899 16609 16908 16643
rect 16856 16600 16908 16609
rect 17040 16600 17092 16652
rect 17224 16600 17276 16652
rect 22468 16736 22520 16788
rect 22652 16736 22704 16788
rect 21088 16711 21140 16720
rect 21088 16677 21097 16711
rect 21097 16677 21131 16711
rect 21131 16677 21140 16711
rect 21088 16668 21140 16677
rect 17500 16575 17552 16584
rect 17500 16541 17502 16575
rect 17502 16541 17552 16575
rect 17500 16532 17552 16541
rect 20628 16600 20680 16652
rect 18052 16532 18104 16584
rect 20904 16600 20956 16652
rect 23848 16736 23900 16788
rect 24216 16736 24268 16788
rect 24492 16736 24544 16788
rect 21272 16575 21324 16584
rect 21272 16541 21281 16575
rect 21281 16541 21315 16575
rect 21315 16541 21324 16575
rect 21272 16532 21324 16541
rect 21456 16532 21508 16584
rect 24952 16668 25004 16720
rect 25228 16668 25280 16720
rect 21824 16532 21876 16584
rect 21916 16532 21968 16584
rect 22376 16532 22428 16584
rect 23020 16532 23072 16584
rect 23480 16575 23532 16584
rect 23480 16541 23489 16575
rect 23489 16541 23523 16575
rect 23523 16541 23532 16575
rect 23480 16532 23532 16541
rect 23664 16532 23716 16584
rect 27988 16736 28040 16788
rect 29368 16736 29420 16788
rect 30288 16711 30340 16720
rect 30288 16677 30297 16711
rect 30297 16677 30331 16711
rect 30331 16677 30340 16711
rect 30288 16668 30340 16677
rect 25688 16532 25740 16584
rect 27528 16600 27580 16652
rect 27804 16600 27856 16652
rect 28264 16600 28316 16652
rect 30104 16600 30156 16652
rect 30472 16600 30524 16652
rect 26976 16532 27028 16584
rect 28632 16575 28684 16584
rect 28632 16541 28641 16575
rect 28641 16541 28675 16575
rect 28675 16541 28684 16575
rect 28632 16532 28684 16541
rect 8484 16464 8536 16516
rect 16028 16464 16080 16516
rect 16396 16464 16448 16516
rect 16672 16464 16724 16516
rect 25964 16507 26016 16516
rect 2044 16396 2096 16448
rect 3792 16396 3844 16448
rect 4068 16396 4120 16448
rect 7196 16396 7248 16448
rect 9220 16396 9272 16448
rect 10416 16439 10468 16448
rect 10416 16405 10425 16439
rect 10425 16405 10459 16439
rect 10459 16405 10468 16439
rect 10416 16396 10468 16405
rect 10968 16396 11020 16448
rect 12440 16396 12492 16448
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 14464 16396 14516 16448
rect 17592 16396 17644 16448
rect 17684 16396 17736 16448
rect 25964 16473 25973 16507
rect 25973 16473 26007 16507
rect 26007 16473 26016 16507
rect 25964 16464 26016 16473
rect 22928 16396 22980 16448
rect 23020 16396 23072 16448
rect 26700 16396 26752 16448
rect 28080 16396 28132 16448
rect 30104 16396 30156 16448
rect 4193 16294 4245 16346
rect 4257 16294 4309 16346
rect 4321 16294 4373 16346
rect 4385 16294 4437 16346
rect 4449 16294 4501 16346
rect 11783 16294 11835 16346
rect 11847 16294 11899 16346
rect 11911 16294 11963 16346
rect 11975 16294 12027 16346
rect 12039 16294 12091 16346
rect 19373 16294 19425 16346
rect 19437 16294 19489 16346
rect 19501 16294 19553 16346
rect 19565 16294 19617 16346
rect 19629 16294 19681 16346
rect 26963 16294 27015 16346
rect 27027 16294 27079 16346
rect 27091 16294 27143 16346
rect 27155 16294 27207 16346
rect 27219 16294 27271 16346
rect 2320 16192 2372 16244
rect 848 16056 900 16108
rect 5632 16192 5684 16244
rect 3700 16124 3752 16176
rect 3792 16124 3844 16176
rect 5816 16167 5868 16176
rect 5816 16133 5825 16167
rect 5825 16133 5859 16167
rect 5859 16133 5868 16167
rect 5816 16124 5868 16133
rect 1308 15852 1360 15904
rect 1584 15852 1636 15904
rect 3516 15852 3568 15904
rect 8116 16192 8168 16244
rect 10508 16192 10560 16244
rect 6460 16099 6512 16108
rect 6460 16065 6462 16099
rect 6462 16065 6512 16099
rect 6460 16056 6512 16065
rect 8484 16056 8536 16108
rect 9220 16056 9272 16108
rect 4436 15988 4488 16040
rect 4988 15988 5040 16040
rect 6092 16031 6144 16040
rect 6092 15997 6101 16031
rect 6101 15997 6135 16031
rect 6135 15997 6144 16031
rect 6092 15988 6144 15997
rect 5448 15920 5500 15972
rect 8668 15988 8720 16040
rect 8944 16031 8996 16040
rect 8944 15997 8946 16031
rect 8946 15997 8996 16031
rect 8944 15988 8996 15997
rect 13452 16192 13504 16244
rect 15292 16192 15344 16244
rect 15476 16192 15528 16244
rect 16672 16192 16724 16244
rect 17132 16192 17184 16244
rect 17868 16192 17920 16244
rect 19892 16192 19944 16244
rect 16304 16124 16356 16176
rect 11060 16056 11112 16108
rect 11612 16099 11664 16108
rect 11612 16065 11614 16099
rect 11614 16065 11664 16099
rect 11612 16056 11664 16065
rect 13544 16056 13596 16108
rect 11244 16031 11296 16040
rect 11244 15997 11253 16031
rect 11253 15997 11287 16031
rect 11287 15997 11296 16031
rect 11244 15988 11296 15997
rect 3884 15852 3936 15904
rect 4436 15852 4488 15904
rect 10692 15920 10744 15972
rect 10416 15895 10468 15904
rect 10416 15861 10425 15895
rect 10425 15861 10459 15895
rect 10459 15861 10468 15895
rect 10416 15852 10468 15861
rect 13820 15988 13872 16040
rect 13912 15988 13964 16040
rect 13544 15920 13596 15972
rect 14004 15920 14056 15972
rect 16120 15988 16172 16040
rect 16948 16031 17000 16040
rect 16948 15997 16957 16031
rect 16957 15997 16991 16031
rect 16991 15997 17000 16031
rect 16948 15988 17000 15997
rect 17592 15988 17644 16040
rect 17684 16031 17736 16040
rect 17684 15997 17693 16031
rect 17693 15997 17727 16031
rect 17727 15997 17736 16031
rect 17684 15988 17736 15997
rect 18604 15988 18656 16040
rect 22744 16192 22796 16244
rect 22928 16192 22980 16244
rect 25872 16192 25924 16244
rect 29000 16192 29052 16244
rect 27712 16124 27764 16176
rect 28448 16124 28500 16176
rect 20812 16099 20864 16108
rect 20812 16065 20821 16099
rect 20821 16065 20855 16099
rect 20855 16065 20864 16099
rect 20812 16056 20864 16065
rect 21824 16056 21876 16108
rect 22008 16056 22060 16108
rect 24216 16099 24268 16108
rect 17868 15920 17920 15972
rect 22284 16031 22336 16040
rect 22284 15997 22293 16031
rect 22293 15997 22327 16031
rect 22327 15997 22336 16031
rect 22284 15988 22336 15997
rect 23480 15988 23532 16040
rect 23848 16031 23900 16040
rect 23848 15997 23857 16031
rect 23857 15997 23891 16031
rect 23891 15997 23900 16031
rect 23848 15988 23900 15997
rect 11520 15852 11572 15904
rect 13084 15852 13136 15904
rect 13728 15895 13780 15904
rect 13728 15861 13737 15895
rect 13737 15861 13771 15895
rect 13771 15861 13780 15895
rect 13728 15852 13780 15861
rect 14740 15852 14792 15904
rect 14832 15852 14884 15904
rect 16580 15895 16632 15904
rect 16580 15861 16589 15895
rect 16589 15861 16623 15895
rect 16623 15861 16632 15895
rect 16580 15852 16632 15861
rect 17132 15895 17184 15904
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17132 15852 17184 15861
rect 17224 15852 17276 15904
rect 21456 15920 21508 15972
rect 23756 15920 23808 15972
rect 18972 15852 19024 15904
rect 19524 15852 19576 15904
rect 21916 15852 21968 15904
rect 22652 15852 22704 15904
rect 24216 16065 24218 16099
rect 24218 16065 24268 16099
rect 24216 16056 24268 16065
rect 24400 16056 24452 16108
rect 25872 16056 25924 16108
rect 25964 16056 26016 16108
rect 24492 15988 24544 16040
rect 25964 15920 26016 15972
rect 26332 15988 26384 16040
rect 27712 15920 27764 15972
rect 29092 16031 29144 16040
rect 29092 15997 29101 16031
rect 29101 15997 29135 16031
rect 29135 15997 29144 16031
rect 29092 15988 29144 15997
rect 29184 16031 29236 16040
rect 29184 15997 29193 16031
rect 29193 15997 29227 16031
rect 29227 15997 29236 16031
rect 29184 15988 29236 15997
rect 30012 16124 30064 16176
rect 30012 15988 30064 16040
rect 29000 15920 29052 15972
rect 30104 15963 30156 15972
rect 30104 15929 30113 15963
rect 30113 15929 30147 15963
rect 30147 15929 30156 15963
rect 30104 15920 30156 15929
rect 26700 15852 26752 15904
rect 27528 15852 27580 15904
rect 27896 15895 27948 15904
rect 27896 15861 27905 15895
rect 27905 15861 27939 15895
rect 27939 15861 27948 15895
rect 27896 15852 27948 15861
rect 29368 15852 29420 15904
rect 7988 15750 8040 15802
rect 8052 15750 8104 15802
rect 8116 15750 8168 15802
rect 8180 15750 8232 15802
rect 8244 15750 8296 15802
rect 15578 15750 15630 15802
rect 15642 15750 15694 15802
rect 15706 15750 15758 15802
rect 15770 15750 15822 15802
rect 15834 15750 15886 15802
rect 23168 15750 23220 15802
rect 23232 15750 23284 15802
rect 23296 15750 23348 15802
rect 23360 15750 23412 15802
rect 23424 15750 23476 15802
rect 30758 15750 30810 15802
rect 30822 15750 30874 15802
rect 30886 15750 30938 15802
rect 30950 15750 31002 15802
rect 31014 15750 31066 15802
rect 3056 15648 3108 15700
rect 3148 15691 3200 15700
rect 3148 15657 3157 15691
rect 3157 15657 3191 15691
rect 3191 15657 3200 15691
rect 3148 15648 3200 15657
rect 5540 15691 5592 15700
rect 5540 15657 5549 15691
rect 5549 15657 5583 15691
rect 5583 15657 5592 15691
rect 5540 15648 5592 15657
rect 1676 15487 1728 15496
rect 1676 15453 1678 15487
rect 1678 15453 1728 15487
rect 1676 15444 1728 15453
rect 2044 15487 2096 15496
rect 2044 15453 2053 15487
rect 2053 15453 2087 15487
rect 2087 15453 2096 15487
rect 2044 15444 2096 15453
rect 3516 15487 3568 15496
rect 3516 15453 3525 15487
rect 3525 15453 3559 15487
rect 3559 15453 3568 15487
rect 3516 15444 3568 15453
rect 3884 15487 3936 15496
rect 3884 15453 3886 15487
rect 3886 15453 3936 15487
rect 3884 15444 3936 15453
rect 4068 15444 4120 15496
rect 4528 15512 4580 15564
rect 10416 15648 10468 15700
rect 1032 15351 1084 15360
rect 1032 15317 1041 15351
rect 1041 15317 1075 15351
rect 1075 15317 1084 15351
rect 1032 15308 1084 15317
rect 1308 15308 1360 15360
rect 3792 15308 3844 15360
rect 6460 15512 6512 15564
rect 8300 15512 8352 15564
rect 8668 15512 8720 15564
rect 11520 15648 11572 15700
rect 11612 15648 11664 15700
rect 13452 15691 13504 15700
rect 13452 15657 13461 15691
rect 13461 15657 13495 15691
rect 13495 15657 13504 15691
rect 13452 15648 13504 15657
rect 7104 15487 7156 15496
rect 7104 15453 7113 15487
rect 7113 15453 7147 15487
rect 7147 15453 7156 15487
rect 7104 15444 7156 15453
rect 8208 15444 8260 15496
rect 8944 15487 8996 15496
rect 8944 15453 8946 15487
rect 8946 15453 8996 15487
rect 6184 15351 6236 15360
rect 6184 15317 6193 15351
rect 6193 15317 6227 15351
rect 6227 15317 6236 15351
rect 6184 15308 6236 15317
rect 6276 15308 6328 15360
rect 8944 15444 8996 15453
rect 16580 15648 16632 15700
rect 16948 15648 17000 15700
rect 17040 15648 17092 15700
rect 17592 15648 17644 15700
rect 20720 15648 20772 15700
rect 22836 15648 22888 15700
rect 23020 15648 23072 15700
rect 24216 15648 24268 15700
rect 24492 15648 24544 15700
rect 15936 15623 15988 15632
rect 15936 15589 15945 15623
rect 15945 15589 15979 15623
rect 15979 15589 15988 15623
rect 15936 15580 15988 15589
rect 14188 15555 14240 15564
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 14188 15521 14190 15555
rect 14190 15521 14240 15555
rect 14188 15512 14240 15521
rect 14832 15512 14884 15564
rect 11244 15419 11296 15428
rect 11244 15385 11253 15419
rect 11253 15385 11287 15419
rect 11287 15385 11296 15419
rect 12348 15487 12400 15496
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 12348 15444 12400 15453
rect 13820 15487 13872 15496
rect 13820 15453 13829 15487
rect 13829 15453 13863 15487
rect 13863 15453 13872 15487
rect 13820 15444 13872 15453
rect 14464 15444 14516 15496
rect 15384 15444 15436 15496
rect 16028 15444 16080 15496
rect 16764 15444 16816 15496
rect 17500 15512 17552 15564
rect 17224 15487 17276 15496
rect 17224 15453 17233 15487
rect 17233 15453 17267 15487
rect 17267 15453 17276 15487
rect 17224 15444 17276 15453
rect 17960 15487 18012 15496
rect 17960 15453 17969 15487
rect 17969 15453 18003 15487
rect 18003 15453 18012 15487
rect 17960 15444 18012 15453
rect 18604 15512 18656 15564
rect 19524 15580 19576 15632
rect 19708 15555 19760 15564
rect 19708 15521 19717 15555
rect 19717 15521 19751 15555
rect 19751 15521 19760 15555
rect 19708 15512 19760 15521
rect 19800 15512 19852 15564
rect 21364 15512 21416 15564
rect 26240 15623 26292 15632
rect 26240 15589 26249 15623
rect 26249 15589 26283 15623
rect 26283 15589 26292 15623
rect 26240 15580 26292 15589
rect 29736 15580 29788 15632
rect 11244 15376 11296 15385
rect 10416 15351 10468 15360
rect 10416 15317 10425 15351
rect 10425 15317 10459 15351
rect 10459 15317 10468 15351
rect 10416 15308 10468 15317
rect 10508 15308 10560 15360
rect 16856 15419 16908 15428
rect 16856 15385 16865 15419
rect 16865 15385 16899 15419
rect 16899 15385 16908 15419
rect 16856 15376 16908 15385
rect 15568 15308 15620 15360
rect 16396 15308 16448 15360
rect 16580 15308 16632 15360
rect 19064 15351 19116 15360
rect 19064 15317 19073 15351
rect 19073 15317 19107 15351
rect 19107 15317 19116 15351
rect 19064 15308 19116 15317
rect 19432 15487 19484 15496
rect 19432 15453 19441 15487
rect 19441 15453 19475 15487
rect 19475 15453 19484 15487
rect 19432 15444 19484 15453
rect 21272 15487 21324 15496
rect 21272 15453 21281 15487
rect 21281 15453 21315 15487
rect 21315 15453 21324 15487
rect 21272 15444 21324 15453
rect 21456 15444 21508 15496
rect 23756 15512 23808 15564
rect 21916 15444 21968 15496
rect 23848 15444 23900 15496
rect 24676 15512 24728 15564
rect 25872 15555 25924 15564
rect 25872 15521 25881 15555
rect 25881 15521 25915 15555
rect 25915 15521 25924 15555
rect 25872 15512 25924 15521
rect 25964 15512 26016 15564
rect 24216 15487 24268 15496
rect 24216 15453 24225 15487
rect 24225 15453 24259 15487
rect 24259 15453 24268 15487
rect 24216 15444 24268 15453
rect 19708 15308 19760 15360
rect 19800 15308 19852 15360
rect 23664 15308 23716 15360
rect 26700 15512 26752 15564
rect 26976 15512 27028 15564
rect 28724 15512 28776 15564
rect 29000 15512 29052 15564
rect 26884 15487 26936 15496
rect 26884 15453 26896 15487
rect 26896 15453 26930 15487
rect 26930 15453 26936 15487
rect 26884 15444 26936 15453
rect 28816 15444 28868 15496
rect 29368 15444 29420 15496
rect 30288 15444 30340 15496
rect 30656 15444 30708 15496
rect 28816 15308 28868 15360
rect 30012 15351 30064 15360
rect 30012 15317 30021 15351
rect 30021 15317 30055 15351
rect 30055 15317 30064 15351
rect 30012 15308 30064 15317
rect 4193 15206 4245 15258
rect 4257 15206 4309 15258
rect 4321 15206 4373 15258
rect 4385 15206 4437 15258
rect 4449 15206 4501 15258
rect 11783 15206 11835 15258
rect 11847 15206 11899 15258
rect 11911 15206 11963 15258
rect 11975 15206 12027 15258
rect 12039 15206 12091 15258
rect 19373 15206 19425 15258
rect 19437 15206 19489 15258
rect 19501 15206 19553 15258
rect 19565 15206 19617 15258
rect 19629 15206 19681 15258
rect 26963 15206 27015 15258
rect 27027 15206 27079 15258
rect 27091 15206 27143 15258
rect 27155 15206 27207 15258
rect 27219 15206 27271 15258
rect 2780 15147 2832 15156
rect 2780 15113 2789 15147
rect 2789 15113 2823 15147
rect 2823 15113 2832 15147
rect 2780 15104 2832 15113
rect 2504 15036 2556 15088
rect 3516 15036 3568 15088
rect 1308 14968 1360 15020
rect 2136 14968 2188 15020
rect 1768 14900 1820 14952
rect 3240 14943 3292 14952
rect 3240 14909 3249 14943
rect 3249 14909 3283 14943
rect 3283 14909 3292 14943
rect 6368 15104 6420 15156
rect 6736 15104 6788 15156
rect 6092 15036 6144 15088
rect 3792 15011 3844 15020
rect 3792 14977 3801 15011
rect 3801 14977 3835 15011
rect 3835 14977 3844 15011
rect 3792 14968 3844 14977
rect 6276 14968 6328 15020
rect 10508 15104 10560 15156
rect 10140 15036 10192 15088
rect 10600 15036 10652 15088
rect 8208 14968 8260 15020
rect 3240 14900 3292 14909
rect 3884 14900 3936 14952
rect 4528 14943 4580 14952
rect 4528 14909 4537 14943
rect 4537 14909 4571 14943
rect 4571 14909 4580 14943
rect 4528 14900 4580 14909
rect 1676 14764 1728 14816
rect 6368 14900 6420 14952
rect 9680 14900 9732 14952
rect 10232 14968 10284 15020
rect 13728 15104 13780 15156
rect 11612 15011 11664 15020
rect 11612 14977 11614 15011
rect 11614 14977 11664 15011
rect 11612 14968 11664 14977
rect 11888 14968 11940 15020
rect 11980 15011 12032 15018
rect 11980 14977 11989 15011
rect 11989 14977 12023 15011
rect 12023 14977 12032 15011
rect 11980 14966 12032 14977
rect 12072 14968 12124 15020
rect 18052 15104 18104 15156
rect 21916 15104 21968 15156
rect 17868 15036 17920 15088
rect 22468 15079 22520 15088
rect 22468 15045 22477 15079
rect 22477 15045 22511 15079
rect 22511 15045 22520 15079
rect 22468 15036 22520 15045
rect 24216 15104 24268 15156
rect 24952 15104 25004 15156
rect 27528 15104 27580 15156
rect 27804 15104 27856 15156
rect 23572 15036 23624 15088
rect 10876 14900 10928 14952
rect 11152 14943 11204 14952
rect 11152 14909 11161 14943
rect 11161 14909 11195 14943
rect 11195 14909 11204 14943
rect 11152 14900 11204 14909
rect 11244 14943 11296 14952
rect 11244 14909 11253 14943
rect 11253 14909 11287 14943
rect 11287 14909 11296 14943
rect 11244 14900 11296 14909
rect 13820 14900 13872 14952
rect 3608 14764 3660 14816
rect 4620 14764 4672 14816
rect 5540 14764 5592 14816
rect 5908 14764 5960 14816
rect 6092 14764 6144 14816
rect 6460 14764 6512 14816
rect 8944 14764 8996 14816
rect 9772 14764 9824 14816
rect 13636 14764 13688 14816
rect 13820 14764 13872 14816
rect 14832 14764 14884 14816
rect 16580 14968 16632 15020
rect 19800 14968 19852 15020
rect 19892 15011 19944 15020
rect 19892 14977 19901 15011
rect 19901 14977 19935 15011
rect 19935 14977 19944 15011
rect 19892 14968 19944 14977
rect 20536 14968 20588 15020
rect 20628 15011 20680 15020
rect 20628 14977 20637 15011
rect 20637 14977 20671 15011
rect 20671 14977 20680 15011
rect 20628 14968 20680 14977
rect 20720 14968 20772 15020
rect 18696 14943 18748 14952
rect 18696 14909 18705 14943
rect 18705 14909 18739 14943
rect 18739 14909 18748 14943
rect 18696 14900 18748 14909
rect 18880 14832 18932 14884
rect 18972 14875 19024 14884
rect 18972 14841 18981 14875
rect 18981 14841 19015 14875
rect 19015 14841 19024 14875
rect 18972 14832 19024 14841
rect 19708 14943 19760 14952
rect 19708 14909 19717 14943
rect 19717 14909 19751 14943
rect 19751 14909 19760 14943
rect 22836 14968 22888 15020
rect 23756 14968 23808 15020
rect 24216 15011 24268 15020
rect 24216 14977 24218 15011
rect 24218 14977 24268 15011
rect 24216 14968 24268 14977
rect 26056 15036 26108 15088
rect 25964 14968 26016 15020
rect 19708 14900 19760 14909
rect 19984 14832 20036 14884
rect 23204 14943 23256 14952
rect 23204 14909 23213 14943
rect 23213 14909 23247 14943
rect 23247 14909 23256 14943
rect 23204 14900 23256 14909
rect 16396 14764 16448 14816
rect 16764 14764 16816 14816
rect 23020 14832 23072 14884
rect 23848 14943 23900 14952
rect 23848 14909 23857 14943
rect 23857 14909 23891 14943
rect 23891 14909 23900 14943
rect 23848 14900 23900 14909
rect 20260 14764 20312 14816
rect 21456 14764 21508 14816
rect 21732 14807 21784 14816
rect 21732 14773 21741 14807
rect 21741 14773 21775 14807
rect 21775 14773 21784 14807
rect 21732 14764 21784 14773
rect 22652 14764 22704 14816
rect 24216 14764 24268 14816
rect 25688 14807 25740 14816
rect 25688 14773 25697 14807
rect 25697 14773 25731 14807
rect 25731 14773 25740 14807
rect 25688 14764 25740 14773
rect 26056 14764 26108 14816
rect 26608 14968 26660 15020
rect 28172 14968 28224 15020
rect 30104 15104 30156 15156
rect 27988 14832 28040 14884
rect 28540 14968 28592 15020
rect 26700 14764 26752 14816
rect 26792 14764 26844 14816
rect 27528 14764 27580 14816
rect 28724 14943 28776 14952
rect 28724 14909 28733 14943
rect 28733 14909 28767 14943
rect 28767 14909 28776 14943
rect 28724 14900 28776 14909
rect 28816 14832 28868 14884
rect 29552 14943 29604 14952
rect 29552 14909 29561 14943
rect 29561 14909 29595 14943
rect 29595 14909 29604 14943
rect 29552 14900 29604 14909
rect 29736 14832 29788 14884
rect 29276 14764 29328 14816
rect 31116 14764 31168 14816
rect 7988 14662 8040 14714
rect 8052 14662 8104 14714
rect 8116 14662 8168 14714
rect 8180 14662 8232 14714
rect 8244 14662 8296 14714
rect 15578 14662 15630 14714
rect 15642 14662 15694 14714
rect 15706 14662 15758 14714
rect 15770 14662 15822 14714
rect 15834 14662 15886 14714
rect 23168 14662 23220 14714
rect 23232 14662 23284 14714
rect 23296 14662 23348 14714
rect 23360 14662 23412 14714
rect 23424 14662 23476 14714
rect 30758 14662 30810 14714
rect 30822 14662 30874 14714
rect 30886 14662 30938 14714
rect 30950 14662 31002 14714
rect 31014 14662 31066 14714
rect 2504 14560 2556 14612
rect 2596 14560 2648 14612
rect 3056 14492 3108 14544
rect 3424 14560 3476 14612
rect 4436 14603 4488 14612
rect 4436 14569 4445 14603
rect 4445 14569 4479 14603
rect 4479 14569 4488 14603
rect 4436 14560 4488 14569
rect 4528 14560 4580 14612
rect 4988 14603 5040 14612
rect 4988 14569 4997 14603
rect 4997 14569 5031 14603
rect 5031 14569 5040 14603
rect 4988 14560 5040 14569
rect 5448 14603 5500 14612
rect 5448 14569 5457 14603
rect 5457 14569 5491 14603
rect 5491 14569 5500 14603
rect 5448 14560 5500 14569
rect 6368 14603 6420 14612
rect 6368 14569 6377 14603
rect 6377 14569 6411 14603
rect 6411 14569 6420 14603
rect 6368 14560 6420 14569
rect 7104 14560 7156 14612
rect 7288 14560 7340 14612
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2596 14424 2648 14476
rect 1676 14356 1728 14408
rect 2044 14356 2096 14408
rect 3148 14356 3200 14408
rect 3792 14356 3844 14408
rect 4436 14424 4488 14476
rect 4620 14467 4672 14476
rect 4620 14433 4629 14467
rect 4629 14433 4663 14467
rect 4663 14433 4672 14467
rect 4620 14424 4672 14433
rect 4712 14424 4764 14476
rect 4988 14424 5040 14476
rect 5356 14356 5408 14408
rect 5908 14424 5960 14476
rect 6276 14467 6328 14476
rect 6276 14433 6285 14467
rect 6285 14433 6319 14467
rect 6319 14433 6328 14467
rect 6276 14424 6328 14433
rect 6368 14424 6420 14476
rect 6644 14467 6696 14476
rect 6644 14433 6653 14467
rect 6653 14433 6687 14467
rect 6687 14433 6696 14467
rect 6644 14424 6696 14433
rect 8944 14560 8996 14612
rect 9036 14560 9088 14612
rect 9312 14560 9364 14612
rect 9680 14603 9732 14612
rect 9680 14569 9689 14603
rect 9689 14569 9723 14603
rect 9723 14569 9732 14603
rect 9680 14560 9732 14569
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 10048 14560 10100 14612
rect 11980 14560 12032 14612
rect 13452 14603 13504 14612
rect 13452 14569 13461 14603
rect 13461 14569 13495 14603
rect 13495 14569 13504 14603
rect 13452 14560 13504 14569
rect 14832 14560 14884 14612
rect 14924 14560 14976 14612
rect 18328 14560 18380 14612
rect 20628 14560 20680 14612
rect 7012 14399 7064 14408
rect 7012 14365 7014 14399
rect 7014 14365 7064 14399
rect 7012 14356 7064 14365
rect 7288 14356 7340 14408
rect 7380 14399 7432 14408
rect 7380 14365 7389 14399
rect 7389 14365 7423 14399
rect 7423 14365 7432 14399
rect 7380 14356 7432 14365
rect 7564 14356 7616 14408
rect 4712 14288 4764 14340
rect 5724 14288 5776 14340
rect 6368 14288 6420 14340
rect 4804 14220 4856 14272
rect 5816 14263 5868 14272
rect 5816 14229 5825 14263
rect 5825 14229 5859 14263
rect 5859 14229 5868 14263
rect 5816 14220 5868 14229
rect 6000 14220 6052 14272
rect 6644 14220 6696 14272
rect 9312 14424 9364 14476
rect 9956 14424 10008 14476
rect 10968 14492 11020 14544
rect 11520 14492 11572 14544
rect 10232 14424 10284 14476
rect 10324 14424 10376 14476
rect 10784 14467 10836 14476
rect 10784 14433 10793 14467
rect 10793 14433 10827 14467
rect 10827 14433 10836 14467
rect 10784 14424 10836 14433
rect 11244 14424 11296 14476
rect 11796 14356 11848 14408
rect 12256 14356 12308 14408
rect 13820 14399 13872 14408
rect 13820 14365 13829 14399
rect 13829 14365 13863 14399
rect 13863 14365 13872 14399
rect 13820 14356 13872 14365
rect 14464 14356 14516 14408
rect 14556 14399 14608 14408
rect 14556 14365 14565 14399
rect 14565 14365 14599 14399
rect 14599 14365 14608 14399
rect 14556 14356 14608 14365
rect 14648 14356 14700 14408
rect 15384 14356 15436 14408
rect 8392 14288 8444 14340
rect 10140 14288 10192 14340
rect 10876 14288 10928 14340
rect 10048 14220 10100 14272
rect 10232 14220 10284 14272
rect 10416 14220 10468 14272
rect 10600 14263 10652 14272
rect 10600 14229 10609 14263
rect 10609 14229 10643 14263
rect 10643 14229 10652 14263
rect 10600 14220 10652 14229
rect 12716 14220 12768 14272
rect 14188 14220 14240 14272
rect 16672 14467 16724 14476
rect 16672 14433 16681 14467
rect 16681 14433 16715 14467
rect 16715 14433 16724 14467
rect 16672 14424 16724 14433
rect 16764 14424 16816 14476
rect 20168 14424 20220 14476
rect 20536 14424 20588 14476
rect 20720 14467 20772 14476
rect 20720 14433 20737 14467
rect 20737 14433 20771 14467
rect 20771 14433 20772 14467
rect 20720 14424 20772 14433
rect 21732 14560 21784 14612
rect 22652 14560 22704 14612
rect 23664 14560 23716 14612
rect 23848 14560 23900 14612
rect 24032 14560 24084 14612
rect 24400 14560 24452 14612
rect 26056 14603 26108 14612
rect 26056 14569 26065 14603
rect 26065 14569 26099 14603
rect 26099 14569 26108 14603
rect 26056 14560 26108 14569
rect 18972 14331 19024 14340
rect 18972 14297 18981 14331
rect 18981 14297 19015 14331
rect 19015 14297 19024 14331
rect 18972 14288 19024 14297
rect 16580 14220 16632 14272
rect 18696 14220 18748 14272
rect 19800 14220 19852 14272
rect 20812 14220 20864 14272
rect 20996 14220 21048 14272
rect 22100 14424 22152 14476
rect 22836 14424 22888 14476
rect 23664 14467 23716 14476
rect 23664 14433 23673 14467
rect 23673 14433 23707 14467
rect 23707 14433 23716 14467
rect 23664 14424 23716 14433
rect 23756 14424 23808 14476
rect 26792 14492 26844 14544
rect 27344 14560 27396 14612
rect 28724 14560 28776 14612
rect 29920 14603 29972 14612
rect 29920 14569 29929 14603
rect 29929 14569 29963 14603
rect 29963 14569 29972 14603
rect 29920 14560 29972 14569
rect 27528 14535 27580 14544
rect 27528 14501 27537 14535
rect 27537 14501 27571 14535
rect 27571 14501 27580 14535
rect 27528 14492 27580 14501
rect 24860 14424 24912 14476
rect 26424 14424 26476 14476
rect 27068 14424 27120 14476
rect 21272 14399 21324 14408
rect 21272 14365 21281 14399
rect 21281 14365 21315 14399
rect 21315 14365 21324 14399
rect 21272 14356 21324 14365
rect 21456 14356 21508 14408
rect 22928 14356 22980 14408
rect 24032 14399 24084 14408
rect 24032 14365 24041 14399
rect 24041 14365 24075 14399
rect 24075 14365 24084 14399
rect 24032 14356 24084 14365
rect 24492 14399 24544 14408
rect 24492 14365 24504 14399
rect 24504 14365 24538 14399
rect 24538 14365 24544 14399
rect 24492 14356 24544 14365
rect 23940 14288 23992 14340
rect 28724 14356 28776 14408
rect 28816 14399 28868 14408
rect 28816 14365 28825 14399
rect 28825 14365 28859 14399
rect 28859 14365 28868 14399
rect 28816 14356 28868 14365
rect 29920 14424 29972 14476
rect 30564 14424 30616 14476
rect 31116 14424 31168 14476
rect 29920 14288 29972 14340
rect 23296 14263 23348 14272
rect 23296 14229 23305 14263
rect 23305 14229 23339 14263
rect 23339 14229 23348 14263
rect 23296 14220 23348 14229
rect 24676 14220 24728 14272
rect 26516 14220 26568 14272
rect 27344 14220 27396 14272
rect 27712 14220 27764 14272
rect 30564 14220 30616 14272
rect 4193 14118 4245 14170
rect 4257 14118 4309 14170
rect 4321 14118 4373 14170
rect 4385 14118 4437 14170
rect 4449 14118 4501 14170
rect 11783 14118 11835 14170
rect 11847 14118 11899 14170
rect 11911 14118 11963 14170
rect 11975 14118 12027 14170
rect 12039 14118 12091 14170
rect 19373 14118 19425 14170
rect 19437 14118 19489 14170
rect 19501 14118 19553 14170
rect 19565 14118 19617 14170
rect 19629 14118 19681 14170
rect 26963 14118 27015 14170
rect 27027 14118 27079 14170
rect 27091 14118 27143 14170
rect 27155 14118 27207 14170
rect 27219 14118 27271 14170
rect 1124 14016 1176 14068
rect 940 13923 992 13932
rect 940 13889 949 13923
rect 949 13889 983 13923
rect 983 13889 992 13923
rect 940 13880 992 13889
rect 1308 13923 1360 13932
rect 1308 13889 1310 13923
rect 1310 13889 1360 13923
rect 1308 13880 1360 13889
rect 2320 13880 2372 13932
rect 2596 13812 2648 13864
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 4988 14016 5040 14068
rect 5816 14016 5868 14068
rect 7196 14016 7248 14068
rect 3792 13948 3844 14000
rect 3792 13855 3844 13864
rect 3792 13821 3801 13855
rect 3801 13821 3835 13855
rect 3835 13821 3844 13855
rect 3792 13812 3844 13821
rect 4620 13880 4672 13932
rect 4712 13880 4764 13932
rect 5908 13855 5960 13864
rect 5908 13821 5917 13855
rect 5917 13821 5951 13855
rect 5951 13821 5960 13855
rect 5908 13812 5960 13821
rect 6092 13855 6144 13864
rect 6092 13821 6101 13855
rect 6101 13821 6135 13855
rect 6135 13821 6144 13855
rect 6092 13812 6144 13821
rect 9772 14016 9824 14068
rect 10140 14016 10192 14068
rect 10508 14016 10560 14068
rect 13636 14059 13688 14068
rect 13636 14025 13645 14059
rect 13645 14025 13679 14059
rect 13679 14025 13688 14059
rect 13636 14016 13688 14025
rect 8944 13880 8996 13932
rect 9312 13880 9364 13932
rect 10140 13880 10192 13932
rect 10600 13880 10652 13932
rect 11612 13923 11664 13932
rect 7564 13812 7616 13864
rect 8760 13812 8812 13864
rect 10876 13812 10928 13864
rect 10968 13812 11020 13864
rect 11244 13855 11296 13864
rect 11244 13821 11253 13855
rect 11253 13821 11287 13855
rect 11287 13821 11296 13855
rect 11244 13812 11296 13821
rect 11612 13889 11614 13923
rect 11614 13889 11664 13923
rect 11612 13880 11664 13889
rect 16396 14016 16448 14068
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 14096 13855 14148 13864
rect 14096 13821 14105 13855
rect 14105 13821 14139 13855
rect 14139 13821 14148 13855
rect 14096 13812 14148 13821
rect 14188 13855 14240 13864
rect 14188 13821 14197 13855
rect 14197 13821 14231 13855
rect 14231 13821 14240 13855
rect 14188 13812 14240 13821
rect 15108 13880 15160 13932
rect 16580 13880 16632 13932
rect 16764 13923 16816 13932
rect 16764 13889 16766 13923
rect 16766 13889 16816 13923
rect 16764 13880 16816 13889
rect 23296 14016 23348 14068
rect 23848 14016 23900 14068
rect 24032 14016 24084 14068
rect 18880 13948 18932 14000
rect 19156 13948 19208 14000
rect 19800 13948 19852 14000
rect 21364 13948 21416 14000
rect 18972 13812 19024 13864
rect 19432 13923 19484 13932
rect 19432 13889 19441 13923
rect 19441 13889 19475 13923
rect 19475 13889 19484 13923
rect 19432 13880 19484 13889
rect 19892 13812 19944 13864
rect 20628 13880 20680 13932
rect 21180 13880 21232 13932
rect 21824 13880 21876 13932
rect 20812 13812 20864 13864
rect 3240 13719 3292 13728
rect 3240 13685 3249 13719
rect 3249 13685 3283 13719
rect 3283 13685 3292 13719
rect 3240 13676 3292 13685
rect 3884 13676 3936 13728
rect 6460 13676 6512 13728
rect 7196 13676 7248 13728
rect 9864 13744 9916 13796
rect 10692 13744 10744 13796
rect 9128 13676 9180 13728
rect 11244 13676 11296 13728
rect 15936 13744 15988 13796
rect 16212 13744 16264 13796
rect 23848 13880 23900 13932
rect 24400 13923 24452 13932
rect 24400 13889 24402 13923
rect 24402 13889 24452 13923
rect 24400 13880 24452 13889
rect 24584 13880 24636 13932
rect 24676 13880 24728 13932
rect 24952 13880 25004 13932
rect 25872 14016 25924 14068
rect 26332 14016 26384 14068
rect 27436 14016 27488 14068
rect 28172 13948 28224 14000
rect 29000 13948 29052 14000
rect 29276 13991 29328 14000
rect 29276 13957 29285 13991
rect 29285 13957 29319 13991
rect 29319 13957 29328 13991
rect 29276 13948 29328 13957
rect 26700 13923 26752 13932
rect 26700 13889 26709 13923
rect 26709 13889 26743 13923
rect 26743 13889 26752 13923
rect 26700 13880 26752 13889
rect 23664 13812 23716 13864
rect 26792 13812 26844 13864
rect 30472 14016 30524 14068
rect 30288 13991 30340 14000
rect 30288 13957 30297 13991
rect 30297 13957 30331 13991
rect 30331 13957 30340 13991
rect 30288 13948 30340 13957
rect 30380 13880 30432 13932
rect 11888 13676 11940 13728
rect 14832 13676 14884 13728
rect 20260 13719 20312 13728
rect 20260 13685 20275 13719
rect 20275 13685 20309 13719
rect 20309 13685 20312 13719
rect 20260 13676 20312 13685
rect 20996 13676 21048 13728
rect 26608 13744 26660 13796
rect 29000 13812 29052 13864
rect 29184 13812 29236 13864
rect 29276 13812 29328 13864
rect 29368 13812 29420 13864
rect 28540 13744 28592 13796
rect 27712 13676 27764 13728
rect 28264 13676 28316 13728
rect 28632 13676 28684 13728
rect 30564 13676 30616 13728
rect 7988 13574 8040 13626
rect 8052 13574 8104 13626
rect 8116 13574 8168 13626
rect 8180 13574 8232 13626
rect 8244 13574 8296 13626
rect 15578 13574 15630 13626
rect 15642 13574 15694 13626
rect 15706 13574 15758 13626
rect 15770 13574 15822 13626
rect 15834 13574 15886 13626
rect 23168 13574 23220 13626
rect 23232 13574 23284 13626
rect 23296 13574 23348 13626
rect 23360 13574 23412 13626
rect 23424 13574 23476 13626
rect 30758 13574 30810 13626
rect 30822 13574 30874 13626
rect 30886 13574 30938 13626
rect 30950 13574 31002 13626
rect 31014 13574 31066 13626
rect 756 13472 808 13524
rect 1768 13472 1820 13524
rect 1124 13404 1176 13456
rect 1308 13311 1360 13320
rect 1308 13277 1317 13311
rect 1317 13277 1351 13311
rect 1351 13277 1360 13311
rect 1308 13268 1360 13277
rect 1492 13268 1544 13320
rect 1676 13311 1728 13320
rect 1676 13277 1678 13311
rect 1678 13277 1728 13311
rect 1676 13268 1728 13277
rect 1952 13268 2004 13320
rect 2044 13311 2096 13320
rect 2044 13277 2053 13311
rect 2053 13277 2087 13311
rect 2087 13277 2096 13311
rect 2044 13268 2096 13277
rect 5264 13472 5316 13524
rect 5356 13472 5408 13524
rect 6092 13472 6144 13524
rect 7380 13472 7432 13524
rect 8576 13515 8628 13524
rect 8576 13481 8585 13515
rect 8585 13481 8619 13515
rect 8619 13481 8628 13515
rect 8576 13472 8628 13481
rect 8668 13472 8720 13524
rect 8944 13515 8996 13524
rect 8944 13481 8953 13515
rect 8953 13481 8987 13515
rect 8987 13481 8996 13515
rect 8944 13472 8996 13481
rect 9220 13515 9272 13524
rect 9220 13481 9229 13515
rect 9229 13481 9263 13515
rect 9263 13481 9272 13515
rect 9220 13472 9272 13481
rect 9404 13472 9456 13524
rect 9588 13472 9640 13524
rect 11152 13472 11204 13524
rect 11428 13515 11480 13524
rect 11428 13481 11437 13515
rect 11437 13481 11471 13515
rect 11471 13481 11480 13515
rect 11428 13472 11480 13481
rect 11888 13515 11940 13524
rect 11888 13481 11897 13515
rect 11897 13481 11931 13515
rect 11931 13481 11940 13515
rect 11888 13472 11940 13481
rect 12164 13472 12216 13524
rect 6276 13404 6328 13456
rect 3884 13311 3936 13320
rect 3884 13277 3886 13311
rect 3886 13277 3936 13311
rect 3884 13268 3936 13277
rect 6368 13379 6420 13388
rect 5816 13268 5868 13320
rect 4988 13200 5040 13252
rect 6368 13345 6377 13379
rect 6377 13345 6411 13379
rect 6411 13345 6420 13379
rect 6368 13336 6420 13345
rect 6092 13268 6144 13320
rect 9312 13336 9364 13388
rect 9680 13379 9732 13388
rect 9680 13345 9689 13379
rect 9689 13345 9723 13379
rect 9723 13345 9732 13379
rect 9680 13336 9732 13345
rect 9864 13336 9916 13388
rect 11612 13404 11664 13456
rect 10232 13379 10284 13388
rect 10232 13345 10241 13379
rect 10241 13345 10275 13379
rect 10275 13345 10284 13379
rect 10232 13336 10284 13345
rect 10324 13336 10376 13388
rect 10784 13379 10836 13388
rect 10784 13345 10793 13379
rect 10793 13345 10827 13379
rect 10827 13345 10836 13379
rect 10784 13336 10836 13345
rect 11060 13336 11112 13388
rect 11428 13336 11480 13388
rect 12532 13472 12584 13524
rect 13268 13472 13320 13524
rect 14556 13472 14608 13524
rect 14832 13472 14884 13524
rect 15108 13472 15160 13524
rect 19156 13472 19208 13524
rect 24032 13472 24084 13524
rect 15384 13404 15436 13456
rect 6736 13311 6788 13320
rect 6736 13277 6753 13311
rect 6753 13277 6787 13311
rect 6787 13277 6788 13311
rect 6736 13268 6788 13277
rect 7012 13268 7064 13320
rect 7196 13311 7248 13320
rect 7196 13277 7208 13311
rect 7208 13277 7242 13311
rect 7242 13277 7248 13311
rect 7196 13268 7248 13277
rect 7472 13311 7524 13320
rect 7472 13277 7481 13311
rect 7481 13277 7515 13311
rect 7515 13277 7524 13311
rect 7472 13268 7524 13277
rect 9496 13268 9548 13320
rect 8392 13200 8444 13252
rect 9220 13200 9272 13252
rect 3792 13132 3844 13184
rect 5448 13132 5500 13184
rect 6644 13132 6696 13184
rect 7932 13132 7984 13184
rect 9680 13132 9732 13184
rect 10232 13132 10284 13184
rect 10416 13132 10468 13184
rect 10600 13175 10652 13184
rect 10600 13141 10609 13175
rect 10609 13141 10643 13175
rect 10643 13141 10652 13175
rect 10600 13132 10652 13141
rect 14924 13379 14976 13388
rect 14924 13345 14933 13379
rect 14933 13345 14967 13379
rect 14967 13345 14976 13379
rect 14924 13336 14976 13345
rect 12716 13268 12768 13320
rect 13176 13268 13228 13320
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 13636 13268 13688 13320
rect 12256 13132 12308 13184
rect 16028 13336 16080 13388
rect 15108 13268 15160 13320
rect 16304 13268 16356 13320
rect 16580 13311 16632 13320
rect 16580 13277 16592 13311
rect 16592 13277 16626 13311
rect 16626 13277 16632 13311
rect 16580 13268 16632 13277
rect 16856 13311 16908 13320
rect 16856 13277 16865 13311
rect 16865 13277 16899 13311
rect 16899 13277 16908 13311
rect 16856 13268 16908 13277
rect 18604 13268 18656 13320
rect 18788 13311 18840 13320
rect 18788 13277 18800 13311
rect 18800 13277 18834 13311
rect 18834 13277 18840 13311
rect 18788 13268 18840 13277
rect 19708 13268 19760 13320
rect 20168 13268 20220 13320
rect 23664 13336 23716 13388
rect 26884 13472 26936 13524
rect 27620 13472 27672 13524
rect 29276 13472 29328 13524
rect 30288 13472 30340 13524
rect 30472 13404 30524 13456
rect 26792 13379 26844 13388
rect 26792 13345 26794 13379
rect 26794 13345 26844 13379
rect 26792 13336 26844 13345
rect 28356 13336 28408 13388
rect 30012 13336 30064 13388
rect 22100 13268 22152 13320
rect 22468 13268 22520 13320
rect 22652 13311 22704 13320
rect 22652 13277 22661 13311
rect 22661 13277 22695 13311
rect 22695 13277 22704 13311
rect 22652 13268 22704 13277
rect 24124 13311 24176 13320
rect 24124 13277 24133 13311
rect 24133 13277 24167 13311
rect 24167 13277 24176 13311
rect 24124 13268 24176 13277
rect 25044 13268 25096 13320
rect 26608 13268 26660 13320
rect 26884 13311 26936 13320
rect 26884 13277 26896 13311
rect 26896 13277 26930 13311
rect 26930 13277 26936 13311
rect 26884 13268 26936 13277
rect 27344 13268 27396 13320
rect 14372 13175 14424 13184
rect 14372 13141 14381 13175
rect 14381 13141 14415 13175
rect 14415 13141 14424 13175
rect 14372 13132 14424 13141
rect 14464 13132 14516 13184
rect 15752 13175 15804 13184
rect 15752 13141 15761 13175
rect 15761 13141 15795 13175
rect 15795 13141 15804 13175
rect 15752 13132 15804 13141
rect 18696 13132 18748 13184
rect 20352 13175 20404 13184
rect 20352 13141 20361 13175
rect 20361 13141 20395 13175
rect 20395 13141 20404 13175
rect 20352 13132 20404 13141
rect 24124 13132 24176 13184
rect 24308 13132 24360 13184
rect 29552 13132 29604 13184
rect 30288 13132 30340 13184
rect 31208 13132 31260 13184
rect 4193 13030 4245 13082
rect 4257 13030 4309 13082
rect 4321 13030 4373 13082
rect 4385 13030 4437 13082
rect 4449 13030 4501 13082
rect 11783 13030 11835 13082
rect 11847 13030 11899 13082
rect 11911 13030 11963 13082
rect 11975 13030 12027 13082
rect 12039 13030 12091 13082
rect 19373 13030 19425 13082
rect 19437 13030 19489 13082
rect 19501 13030 19553 13082
rect 19565 13030 19617 13082
rect 19629 13030 19681 13082
rect 26963 13030 27015 13082
rect 27027 13030 27079 13082
rect 27091 13030 27143 13082
rect 27155 13030 27207 13082
rect 27219 13030 27271 13082
rect 3148 12928 3200 12980
rect 3608 12928 3660 12980
rect 5724 12928 5776 12980
rect 7196 12928 7248 12980
rect 7472 12928 7524 12980
rect 9312 12928 9364 12980
rect 1308 12792 1360 12844
rect 2136 12792 2188 12844
rect 4620 12835 4672 12844
rect 4620 12801 4629 12835
rect 4629 12801 4663 12835
rect 4663 12801 4672 12835
rect 4620 12792 4672 12801
rect 7840 12860 7892 12912
rect 9496 12860 9548 12912
rect 3240 12724 3292 12776
rect 3608 12724 3660 12776
rect 3792 12724 3844 12776
rect 5356 12724 5408 12776
rect 6644 12792 6696 12844
rect 6736 12792 6788 12844
rect 8852 12724 8904 12776
rect 11428 12928 11480 12980
rect 11336 12860 11388 12912
rect 12808 12928 12860 12980
rect 16212 12928 16264 12980
rect 16856 12928 16908 12980
rect 17960 12928 18012 12980
rect 1676 12588 1728 12640
rect 3240 12631 3292 12640
rect 3240 12597 3249 12631
rect 3249 12597 3283 12631
rect 3283 12597 3292 12631
rect 3240 12588 3292 12597
rect 3976 12588 4028 12640
rect 6000 12588 6052 12640
rect 6460 12588 6512 12640
rect 7104 12588 7156 12640
rect 7472 12588 7524 12640
rect 8852 12588 8904 12640
rect 9588 12767 9640 12776
rect 9588 12733 9597 12767
rect 9597 12733 9631 12767
rect 9631 12733 9640 12767
rect 9588 12724 9640 12733
rect 9680 12774 9732 12826
rect 9772 12792 9824 12844
rect 10508 12792 10560 12844
rect 11152 12792 11204 12844
rect 11520 12792 11572 12844
rect 13452 12860 13504 12912
rect 10784 12724 10836 12776
rect 11336 12724 11388 12776
rect 11704 12767 11756 12776
rect 11704 12733 11713 12767
rect 11713 12733 11747 12767
rect 11747 12733 11756 12767
rect 11704 12724 11756 12733
rect 12624 12792 12676 12844
rect 13912 12792 13964 12844
rect 15200 12792 15252 12844
rect 16396 12792 16448 12844
rect 16672 12792 16724 12844
rect 12164 12724 12216 12776
rect 12992 12724 13044 12776
rect 13176 12724 13228 12776
rect 13360 12767 13412 12776
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 9220 12588 9272 12640
rect 9312 12631 9364 12640
rect 9312 12597 9321 12631
rect 9321 12597 9355 12631
rect 9355 12597 9364 12631
rect 9312 12588 9364 12597
rect 11336 12588 11388 12640
rect 12532 12656 12584 12708
rect 14648 12724 14700 12776
rect 15108 12724 15160 12776
rect 15200 12656 15252 12708
rect 16764 12724 16816 12776
rect 18144 12767 18196 12776
rect 18144 12733 18153 12767
rect 18153 12733 18187 12767
rect 18187 12733 18196 12767
rect 18144 12724 18196 12733
rect 18604 12792 18656 12844
rect 18972 12928 19024 12980
rect 20352 12928 20404 12980
rect 22652 12928 22704 12980
rect 23572 12928 23624 12980
rect 23848 12928 23900 12980
rect 24492 12928 24544 12980
rect 28908 12928 28960 12980
rect 29092 12928 29144 12980
rect 29460 12928 29512 12980
rect 29644 12971 29696 12980
rect 29644 12937 29653 12971
rect 29653 12937 29687 12971
rect 29687 12937 29696 12971
rect 29644 12928 29696 12937
rect 29828 12928 29880 12980
rect 22928 12792 22980 12844
rect 24952 12792 25004 12844
rect 26608 12792 26660 12844
rect 31208 12792 31260 12844
rect 19064 12767 19116 12776
rect 19064 12733 19066 12767
rect 19066 12733 19116 12767
rect 13084 12588 13136 12640
rect 13176 12631 13228 12640
rect 13176 12597 13185 12631
rect 13185 12597 13219 12631
rect 13219 12597 13228 12631
rect 13176 12588 13228 12597
rect 13636 12588 13688 12640
rect 15108 12588 15160 12640
rect 17592 12631 17644 12640
rect 17592 12597 17601 12631
rect 17601 12597 17635 12631
rect 17635 12597 17644 12631
rect 17592 12588 17644 12597
rect 17960 12631 18012 12640
rect 17960 12597 17969 12631
rect 17969 12597 18003 12631
rect 18003 12597 18012 12631
rect 17960 12588 18012 12597
rect 19064 12724 19116 12733
rect 19432 12767 19484 12776
rect 19432 12733 19441 12767
rect 19441 12733 19475 12767
rect 19475 12733 19484 12767
rect 19432 12724 19484 12733
rect 19524 12724 19576 12776
rect 20720 12724 20772 12776
rect 21272 12724 21324 12776
rect 21640 12767 21692 12776
rect 21640 12733 21649 12767
rect 21649 12733 21683 12767
rect 21683 12733 21692 12767
rect 21640 12724 21692 12733
rect 23020 12724 23072 12776
rect 23480 12724 23532 12776
rect 20812 12699 20864 12708
rect 20812 12665 20821 12699
rect 20821 12665 20855 12699
rect 20855 12665 20864 12699
rect 20812 12656 20864 12665
rect 23664 12724 23716 12776
rect 23756 12656 23808 12708
rect 20996 12588 21048 12640
rect 21732 12588 21784 12640
rect 22744 12631 22796 12640
rect 22744 12597 22753 12631
rect 22753 12597 22787 12631
rect 22787 12597 22796 12631
rect 22744 12588 22796 12597
rect 24860 12724 24912 12776
rect 26516 12724 26568 12776
rect 28448 12724 28500 12776
rect 29184 12724 29236 12776
rect 24124 12588 24176 12640
rect 24676 12588 24728 12640
rect 29276 12656 29328 12708
rect 26792 12588 26844 12640
rect 27804 12588 27856 12640
rect 29000 12588 29052 12640
rect 29920 12724 29972 12776
rect 30012 12724 30064 12776
rect 30564 12724 30616 12776
rect 30656 12656 30708 12708
rect 7988 12486 8040 12538
rect 8052 12486 8104 12538
rect 8116 12486 8168 12538
rect 8180 12486 8232 12538
rect 8244 12486 8296 12538
rect 15578 12486 15630 12538
rect 15642 12486 15694 12538
rect 15706 12486 15758 12538
rect 15770 12486 15822 12538
rect 15834 12486 15886 12538
rect 23168 12486 23220 12538
rect 23232 12486 23284 12538
rect 23296 12486 23348 12538
rect 23360 12486 23412 12538
rect 23424 12486 23476 12538
rect 30758 12486 30810 12538
rect 30822 12486 30874 12538
rect 30886 12486 30938 12538
rect 30950 12486 31002 12538
rect 31014 12486 31066 12538
rect 1032 12384 1084 12436
rect 2136 12384 2188 12436
rect 5816 12427 5868 12436
rect 5816 12393 5825 12427
rect 5825 12393 5859 12427
rect 5859 12393 5868 12427
rect 5816 12384 5868 12393
rect 6276 12384 6328 12436
rect 6828 12384 6880 12436
rect 7104 12384 7156 12436
rect 9772 12384 9824 12436
rect 11244 12427 11296 12436
rect 11244 12393 11253 12427
rect 11253 12393 11287 12427
rect 11287 12393 11296 12427
rect 11244 12384 11296 12393
rect 11704 12384 11756 12436
rect 1216 12291 1268 12300
rect 1216 12257 1225 12291
rect 1225 12257 1259 12291
rect 1259 12257 1268 12291
rect 1216 12248 1268 12257
rect 1676 12291 1728 12300
rect 1676 12257 1678 12291
rect 1678 12257 1728 12291
rect 1676 12248 1728 12257
rect 1308 12223 1360 12232
rect 1308 12189 1317 12223
rect 1317 12189 1351 12223
rect 1351 12189 1360 12223
rect 1308 12180 1360 12189
rect 1768 12223 1820 12232
rect 1768 12189 1780 12223
rect 1780 12189 1814 12223
rect 1814 12189 1820 12223
rect 1768 12180 1820 12189
rect 2136 12180 2188 12232
rect 3516 12223 3568 12232
rect 3516 12189 3525 12223
rect 3525 12189 3559 12223
rect 3559 12189 3568 12223
rect 3516 12180 3568 12189
rect 3884 12223 3936 12232
rect 3884 12189 3886 12223
rect 3886 12189 3936 12223
rect 3884 12180 3936 12189
rect 4712 12248 4764 12300
rect 5540 12248 5592 12300
rect 8576 12316 8628 12368
rect 6000 12112 6052 12164
rect 6828 12180 6880 12232
rect 2136 12044 2188 12096
rect 6736 12044 6788 12096
rect 7012 12044 7064 12096
rect 8484 12044 8536 12096
rect 8852 12180 8904 12232
rect 9312 12248 9364 12300
rect 11520 12291 11572 12300
rect 11520 12257 11529 12291
rect 11529 12257 11563 12291
rect 11563 12257 11572 12291
rect 11520 12248 11572 12257
rect 12440 12291 12492 12300
rect 10784 12180 10836 12232
rect 12440 12257 12449 12291
rect 12449 12257 12483 12291
rect 12483 12257 12492 12291
rect 12440 12248 12492 12257
rect 12808 12384 12860 12436
rect 13636 12384 13688 12436
rect 14280 12384 14332 12436
rect 16120 12427 16172 12436
rect 16120 12393 16129 12427
rect 16129 12393 16163 12427
rect 16163 12393 16172 12427
rect 16120 12384 16172 12393
rect 17224 12384 17276 12436
rect 18788 12427 18840 12436
rect 18788 12393 18797 12427
rect 18797 12393 18831 12427
rect 18831 12393 18840 12427
rect 18788 12384 18840 12393
rect 18880 12316 18932 12368
rect 19708 12427 19760 12436
rect 19708 12393 19717 12427
rect 19717 12393 19751 12427
rect 19751 12393 19760 12427
rect 19708 12384 19760 12393
rect 21640 12384 21692 12436
rect 21732 12427 21784 12436
rect 21732 12393 21747 12427
rect 21747 12393 21781 12427
rect 21781 12393 21784 12427
rect 21732 12384 21784 12393
rect 21916 12384 21968 12436
rect 22468 12384 22520 12436
rect 24124 12384 24176 12436
rect 24584 12384 24636 12436
rect 26792 12384 26844 12436
rect 28264 12427 28316 12436
rect 28264 12393 28273 12427
rect 28273 12393 28307 12427
rect 28307 12393 28316 12427
rect 28264 12384 28316 12393
rect 30196 12384 30248 12436
rect 13176 12248 13228 12300
rect 14004 12248 14056 12300
rect 12716 12180 12768 12232
rect 13452 12180 13504 12232
rect 10324 12112 10376 12164
rect 14280 12180 14332 12232
rect 17500 12180 17552 12232
rect 17960 12248 18012 12300
rect 18052 12248 18104 12300
rect 19524 12272 19576 12324
rect 19800 12248 19852 12300
rect 20168 12248 20220 12300
rect 20628 12248 20680 12300
rect 21088 12291 21140 12300
rect 21088 12257 21097 12291
rect 21097 12257 21131 12291
rect 21131 12257 21140 12291
rect 21088 12248 21140 12257
rect 22744 12316 22796 12368
rect 26424 12316 26476 12368
rect 29920 12316 29972 12368
rect 21272 12291 21324 12300
rect 21272 12257 21281 12291
rect 21281 12257 21315 12291
rect 21315 12257 21324 12291
rect 21272 12248 21324 12257
rect 21732 12223 21784 12232
rect 21732 12189 21744 12223
rect 21744 12189 21778 12223
rect 21778 12189 21784 12223
rect 21732 12180 21784 12189
rect 19248 12112 19300 12164
rect 20536 12112 20588 12164
rect 9312 12044 9364 12096
rect 9588 12044 9640 12096
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 10968 12087 11020 12096
rect 10968 12053 10977 12087
rect 10977 12053 11011 12087
rect 11011 12053 11020 12087
rect 10968 12044 11020 12053
rect 11060 12044 11112 12096
rect 13268 12044 13320 12096
rect 14556 12087 14608 12096
rect 14556 12053 14565 12087
rect 14565 12053 14599 12087
rect 14599 12053 14608 12087
rect 14556 12044 14608 12053
rect 15568 12087 15620 12096
rect 15568 12053 15577 12087
rect 15577 12053 15611 12087
rect 15611 12053 15620 12087
rect 15568 12044 15620 12053
rect 16672 12087 16724 12096
rect 16672 12053 16681 12087
rect 16681 12053 16715 12087
rect 16715 12053 16724 12087
rect 16672 12044 16724 12053
rect 16764 12044 16816 12096
rect 17500 12044 17552 12096
rect 18420 12044 18472 12096
rect 19064 12044 19116 12096
rect 19432 12087 19484 12096
rect 19432 12053 19441 12087
rect 19441 12053 19475 12087
rect 19475 12053 19484 12087
rect 19432 12044 19484 12053
rect 21456 12044 21508 12096
rect 22376 12044 22428 12096
rect 23296 12044 23348 12096
rect 23664 12180 23716 12232
rect 24216 12291 24268 12300
rect 24216 12257 24225 12291
rect 24225 12257 24259 12291
rect 24259 12257 24268 12291
rect 24216 12248 24268 12257
rect 24216 12044 24268 12096
rect 26516 12248 26568 12300
rect 28080 12248 28132 12300
rect 28908 12291 28960 12300
rect 28908 12257 28917 12291
rect 28917 12257 28951 12291
rect 28951 12257 28960 12291
rect 28908 12248 28960 12257
rect 26884 12223 26936 12232
rect 26884 12189 26896 12223
rect 26896 12189 26930 12223
rect 26930 12189 26936 12223
rect 26884 12180 26936 12189
rect 27804 12180 27856 12232
rect 28632 12223 28684 12232
rect 28632 12189 28641 12223
rect 28641 12189 28675 12223
rect 28675 12189 28684 12223
rect 28632 12180 28684 12189
rect 25504 12044 25556 12096
rect 4193 11942 4245 11994
rect 4257 11942 4309 11994
rect 4321 11942 4373 11994
rect 4385 11942 4437 11994
rect 4449 11942 4501 11994
rect 11783 11942 11835 11994
rect 11847 11942 11899 11994
rect 11911 11942 11963 11994
rect 11975 11942 12027 11994
rect 12039 11942 12091 11994
rect 19373 11942 19425 11994
rect 19437 11942 19489 11994
rect 19501 11942 19553 11994
rect 19565 11942 19617 11994
rect 19629 11942 19681 11994
rect 26963 11942 27015 11994
rect 27027 11942 27079 11994
rect 27091 11942 27143 11994
rect 27155 11942 27207 11994
rect 27219 11942 27271 11994
rect 2780 11883 2832 11892
rect 2780 11849 2789 11883
rect 2789 11849 2823 11883
rect 2823 11849 2832 11883
rect 2780 11840 2832 11849
rect 3700 11772 3752 11824
rect 7288 11840 7340 11892
rect 940 11679 992 11688
rect 940 11645 949 11679
rect 949 11645 983 11679
rect 983 11645 992 11679
rect 940 11636 992 11645
rect 1216 11636 1268 11688
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 1400 11543 1452 11552
rect 1400 11509 1415 11543
rect 1415 11509 1449 11543
rect 1449 11509 1452 11543
rect 1400 11500 1452 11509
rect 1584 11500 1636 11552
rect 2964 11500 3016 11552
rect 3516 11704 3568 11756
rect 4252 11747 4304 11756
rect 4252 11713 4264 11747
rect 4264 11713 4298 11747
rect 4298 11713 4304 11747
rect 4252 11704 4304 11713
rect 5448 11704 5500 11756
rect 4160 11636 4212 11688
rect 5172 11636 5224 11688
rect 3424 11500 3476 11552
rect 3516 11543 3568 11552
rect 3516 11509 3525 11543
rect 3525 11509 3559 11543
rect 3559 11509 3568 11543
rect 3516 11500 3568 11509
rect 4068 11500 4120 11552
rect 4528 11500 4580 11552
rect 5908 11704 5960 11756
rect 7840 11704 7892 11756
rect 6000 11636 6052 11688
rect 10140 11840 10192 11892
rect 10692 11840 10744 11892
rect 11612 11772 11664 11824
rect 12164 11772 12216 11824
rect 9036 11704 9088 11756
rect 9496 11704 9548 11756
rect 7840 11568 7892 11620
rect 8484 11568 8536 11620
rect 8944 11568 8996 11620
rect 6460 11500 6512 11552
rect 6920 11500 6972 11552
rect 9312 11500 9364 11552
rect 9864 11704 9916 11756
rect 10232 11704 10284 11756
rect 11152 11636 11204 11688
rect 12532 11772 12584 11824
rect 12716 11840 12768 11892
rect 13268 11840 13320 11892
rect 13820 11840 13872 11892
rect 12992 11772 13044 11824
rect 13452 11772 13504 11824
rect 15936 11883 15988 11892
rect 15936 11849 15945 11883
rect 15945 11849 15979 11883
rect 15979 11849 15988 11883
rect 15936 11840 15988 11849
rect 17960 11840 18012 11892
rect 9956 11500 10008 11552
rect 11704 11568 11756 11620
rect 13176 11679 13228 11688
rect 13176 11645 13185 11679
rect 13185 11645 13219 11679
rect 13219 11645 13228 11679
rect 13176 11636 13228 11645
rect 13268 11636 13320 11688
rect 13544 11679 13596 11688
rect 13544 11645 13553 11679
rect 13553 11645 13587 11679
rect 13587 11645 13596 11679
rect 13544 11636 13596 11645
rect 14096 11636 14148 11688
rect 19800 11840 19852 11892
rect 21732 11840 21784 11892
rect 22928 11883 22980 11892
rect 22928 11849 22937 11883
rect 22937 11849 22971 11883
rect 22971 11849 22980 11883
rect 22928 11840 22980 11849
rect 23296 11840 23348 11892
rect 23940 11840 23992 11892
rect 26792 11840 26844 11892
rect 26884 11840 26936 11892
rect 28448 11840 28500 11892
rect 28816 11840 28868 11892
rect 30288 11883 30340 11892
rect 30288 11849 30297 11883
rect 30297 11849 30331 11883
rect 30331 11849 30340 11883
rect 30288 11840 30340 11849
rect 20812 11704 20864 11756
rect 21456 11704 21508 11756
rect 30380 11815 30432 11824
rect 30380 11781 30389 11815
rect 30389 11781 30423 11815
rect 30423 11781 30432 11815
rect 30380 11772 30432 11781
rect 24400 11704 24452 11756
rect 25964 11704 26016 11756
rect 12164 11500 12216 11552
rect 12348 11543 12400 11552
rect 12348 11509 12357 11543
rect 12357 11509 12391 11543
rect 12391 11509 12400 11543
rect 12348 11500 12400 11509
rect 13176 11500 13228 11552
rect 13268 11500 13320 11552
rect 14924 11500 14976 11552
rect 18696 11679 18748 11688
rect 18696 11645 18705 11679
rect 18705 11645 18739 11679
rect 18739 11645 18748 11679
rect 18696 11636 18748 11645
rect 19064 11636 19116 11688
rect 21272 11636 21324 11688
rect 22928 11636 22980 11688
rect 23296 11636 23348 11688
rect 23848 11679 23900 11688
rect 23848 11645 23857 11679
rect 23857 11645 23891 11679
rect 23891 11645 23900 11679
rect 23848 11636 23900 11645
rect 23940 11636 23992 11688
rect 24216 11679 24268 11688
rect 24216 11645 24225 11679
rect 24225 11645 24259 11679
rect 24259 11645 24268 11679
rect 24216 11636 24268 11645
rect 25320 11636 25372 11688
rect 26424 11679 26476 11688
rect 26424 11645 26433 11679
rect 26433 11645 26467 11679
rect 26467 11645 26476 11679
rect 26424 11636 26476 11645
rect 27160 11679 27212 11688
rect 27160 11645 27169 11679
rect 27169 11645 27203 11679
rect 27203 11645 27212 11679
rect 27160 11636 27212 11645
rect 28908 11704 28960 11756
rect 29184 11704 29236 11756
rect 29276 11704 29328 11756
rect 30472 11704 30524 11756
rect 31116 11704 31168 11756
rect 29092 11679 29144 11688
rect 29092 11645 29101 11679
rect 29101 11645 29135 11679
rect 29135 11645 29144 11679
rect 29092 11636 29144 11645
rect 29460 11636 29512 11688
rect 29828 11679 29880 11688
rect 29828 11645 29837 11679
rect 29837 11645 29871 11679
rect 29871 11645 29880 11679
rect 29828 11636 29880 11645
rect 29920 11636 29972 11688
rect 30564 11679 30616 11688
rect 30564 11645 30573 11679
rect 30573 11645 30607 11679
rect 30607 11645 30616 11679
rect 30564 11636 30616 11645
rect 16764 11500 16816 11552
rect 17224 11500 17276 11552
rect 19156 11543 19208 11552
rect 19156 11509 19171 11543
rect 19171 11509 19205 11543
rect 19205 11509 19208 11543
rect 19156 11500 19208 11509
rect 21916 11500 21968 11552
rect 22376 11500 22428 11552
rect 22560 11500 22612 11552
rect 23940 11500 23992 11552
rect 24676 11543 24728 11552
rect 24676 11509 24691 11543
rect 24691 11509 24725 11543
rect 24725 11509 24728 11543
rect 24676 11500 24728 11509
rect 26700 11500 26752 11552
rect 28816 11500 28868 11552
rect 29092 11500 29144 11552
rect 29460 11500 29512 11552
rect 29644 11543 29696 11552
rect 29644 11509 29653 11543
rect 29653 11509 29687 11543
rect 29687 11509 29696 11543
rect 29644 11500 29696 11509
rect 7988 11398 8040 11450
rect 8052 11398 8104 11450
rect 8116 11398 8168 11450
rect 8180 11398 8232 11450
rect 8244 11398 8296 11450
rect 15578 11398 15630 11450
rect 15642 11398 15694 11450
rect 15706 11398 15758 11450
rect 15770 11398 15822 11450
rect 15834 11398 15886 11450
rect 23168 11398 23220 11450
rect 23232 11398 23284 11450
rect 23296 11398 23348 11450
rect 23360 11398 23412 11450
rect 23424 11398 23476 11450
rect 30758 11398 30810 11450
rect 30822 11398 30874 11450
rect 30886 11398 30938 11450
rect 30950 11398 31002 11450
rect 31014 11398 31066 11450
rect 1308 11339 1360 11348
rect 1308 11305 1317 11339
rect 1317 11305 1351 11339
rect 1351 11305 1360 11339
rect 1308 11296 1360 11305
rect 1768 11296 1820 11348
rect 1584 11160 1636 11212
rect 2136 11160 2188 11212
rect 4068 11228 4120 11280
rect 1952 11119 1997 11144
rect 1997 11119 2004 11144
rect 1952 11092 2004 11119
rect 4252 11160 4304 11212
rect 3976 11092 4028 11144
rect 4620 11024 4672 11076
rect 5172 11160 5224 11212
rect 8392 11296 8444 11348
rect 8484 11296 8536 11348
rect 8576 11296 8628 11348
rect 11428 11296 11480 11348
rect 11520 11339 11572 11348
rect 11520 11305 11529 11339
rect 11529 11305 11563 11339
rect 11563 11305 11572 11339
rect 11520 11296 11572 11305
rect 5540 11092 5592 11144
rect 6000 11092 6052 11144
rect 6368 11160 6420 11212
rect 6828 11160 6880 11212
rect 7472 11160 7524 11212
rect 12808 11296 12860 11348
rect 13268 11296 13320 11348
rect 14188 11296 14240 11348
rect 15108 11296 15160 11348
rect 16396 11296 16448 11348
rect 16672 11296 16724 11348
rect 6276 11135 6328 11144
rect 6276 11101 6288 11135
rect 6288 11101 6322 11135
rect 6322 11101 6328 11135
rect 6276 11092 6328 11101
rect 6460 11092 6512 11144
rect 7656 11092 7708 11144
rect 7840 11024 7892 11076
rect 8300 11092 8352 11144
rect 8852 11092 8904 11144
rect 9036 11135 9088 11144
rect 9036 11101 9038 11135
rect 9038 11101 9088 11135
rect 9036 11092 9088 11101
rect 10600 11160 10652 11212
rect 9496 11092 9548 11144
rect 12072 11228 12124 11280
rect 11060 11160 11112 11212
rect 5172 10956 5224 11008
rect 6552 10956 6604 11008
rect 11244 11067 11296 11076
rect 11244 11033 11253 11067
rect 11253 11033 11287 11067
rect 11287 11033 11296 11067
rect 11244 11024 11296 11033
rect 11336 11024 11388 11076
rect 11520 11160 11572 11212
rect 12164 11092 12216 11144
rect 12716 11092 12768 11144
rect 13084 11160 13136 11212
rect 13360 11160 13412 11212
rect 13176 11092 13228 11144
rect 14740 11092 14792 11144
rect 16304 11271 16356 11280
rect 16304 11237 16313 11271
rect 16313 11237 16347 11271
rect 16347 11237 16356 11271
rect 16304 11228 16356 11237
rect 15200 11203 15252 11212
rect 15200 11169 15209 11203
rect 15209 11169 15243 11203
rect 15243 11169 15252 11203
rect 16856 11228 16908 11280
rect 15200 11160 15252 11169
rect 18972 11296 19024 11348
rect 20352 11296 20404 11348
rect 22008 11296 22060 11348
rect 22376 11296 22428 11348
rect 19156 11228 19208 11280
rect 21364 11228 21416 11280
rect 23020 11228 23072 11280
rect 25320 11339 25372 11348
rect 25320 11305 25329 11339
rect 25329 11305 25363 11339
rect 25363 11305 25372 11339
rect 25320 11296 25372 11305
rect 26424 11296 26476 11348
rect 26700 11271 26752 11280
rect 16764 11092 16816 11144
rect 17224 11135 17276 11144
rect 17224 11101 17226 11135
rect 17226 11101 17276 11135
rect 11520 11024 11572 11076
rect 11796 11024 11848 11076
rect 12256 11024 12308 11076
rect 12440 11067 12492 11076
rect 12440 11033 12449 11067
rect 12449 11033 12483 11067
rect 12483 11033 12492 11067
rect 12440 11024 12492 11033
rect 14832 11024 14884 11076
rect 9864 10956 9916 11008
rect 10600 10956 10652 11008
rect 11704 10956 11756 11008
rect 12532 10956 12584 11008
rect 13728 10956 13780 11008
rect 14740 10999 14792 11008
rect 14740 10965 14749 10999
rect 14749 10965 14783 10999
rect 14783 10965 14792 10999
rect 14740 10956 14792 10965
rect 15476 10999 15528 11008
rect 15476 10965 15485 10999
rect 15485 10965 15519 10999
rect 15519 10965 15528 10999
rect 15476 10956 15528 10965
rect 17224 11092 17276 11101
rect 20812 11092 20864 11144
rect 21088 11092 21140 11144
rect 21548 11092 21600 11144
rect 22652 11160 22704 11212
rect 26700 11237 26709 11271
rect 26709 11237 26743 11271
rect 26743 11237 26752 11271
rect 26700 11228 26752 11237
rect 27160 11296 27212 11348
rect 27712 11296 27764 11348
rect 27804 11339 27856 11348
rect 27804 11305 27813 11339
rect 27813 11305 27847 11339
rect 27847 11305 27856 11339
rect 27804 11296 27856 11305
rect 27896 11296 27948 11348
rect 30472 11339 30524 11348
rect 30472 11305 30481 11339
rect 30481 11305 30515 11339
rect 30515 11305 30524 11339
rect 30472 11296 30524 11305
rect 25596 11160 25648 11212
rect 26148 11160 26200 11212
rect 26332 11160 26384 11212
rect 29644 11228 29696 11280
rect 22008 11135 22060 11144
rect 22008 11101 22017 11135
rect 22017 11101 22051 11135
rect 22051 11101 22060 11135
rect 22008 11092 22060 11101
rect 22928 11092 22980 11144
rect 23848 11092 23900 11144
rect 23940 11135 23992 11144
rect 23940 11101 23952 11135
rect 23952 11101 23986 11135
rect 23986 11101 23992 11135
rect 23940 11092 23992 11101
rect 24032 11092 24084 11144
rect 19064 10956 19116 11008
rect 26332 11024 26384 11076
rect 23756 10956 23808 11008
rect 25872 10999 25924 11008
rect 25872 10965 25881 10999
rect 25881 10965 25915 10999
rect 25915 10965 25924 10999
rect 25872 10956 25924 10965
rect 26240 10956 26292 11008
rect 30288 11203 30340 11212
rect 30288 11169 30297 11203
rect 30297 11169 30331 11203
rect 30331 11169 30340 11203
rect 30288 11160 30340 11169
rect 28080 11135 28132 11144
rect 28080 11101 28089 11135
rect 28089 11101 28123 11135
rect 28123 11101 28132 11135
rect 28080 11092 28132 11101
rect 29552 11092 29604 11144
rect 29460 10956 29512 11008
rect 30656 10956 30708 11008
rect 4193 10854 4245 10906
rect 4257 10854 4309 10906
rect 4321 10854 4373 10906
rect 4385 10854 4437 10906
rect 4449 10854 4501 10906
rect 11783 10854 11835 10906
rect 11847 10854 11899 10906
rect 11911 10854 11963 10906
rect 11975 10854 12027 10906
rect 12039 10854 12091 10906
rect 19373 10854 19425 10906
rect 19437 10854 19489 10906
rect 19501 10854 19553 10906
rect 19565 10854 19617 10906
rect 19629 10854 19681 10906
rect 26963 10854 27015 10906
rect 27027 10854 27079 10906
rect 27091 10854 27143 10906
rect 27155 10854 27207 10906
rect 27219 10854 27271 10906
rect 1308 10616 1360 10668
rect 15476 10752 15528 10804
rect 21364 10752 21416 10804
rect 11704 10684 11756 10736
rect 11980 10684 12032 10736
rect 12716 10684 12768 10736
rect 13820 10727 13872 10736
rect 13820 10693 13829 10727
rect 13829 10693 13863 10727
rect 13863 10693 13872 10727
rect 13820 10684 13872 10693
rect 5356 10616 5408 10668
rect 6368 10616 6420 10668
rect 7840 10616 7892 10668
rect 664 10548 716 10600
rect 3148 10548 3200 10600
rect 3608 10548 3660 10600
rect 5264 10548 5316 10600
rect 5540 10591 5592 10600
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 5540 10548 5592 10557
rect 3056 10523 3108 10532
rect 3056 10489 3065 10523
rect 3065 10489 3099 10523
rect 3099 10489 3108 10523
rect 3056 10480 3108 10489
rect 5356 10523 5408 10532
rect 5356 10489 5365 10523
rect 5365 10489 5399 10523
rect 5399 10489 5408 10523
rect 5356 10480 5408 10489
rect 1768 10412 1820 10464
rect 3332 10412 3384 10464
rect 3976 10412 4028 10464
rect 6092 10548 6144 10600
rect 6184 10548 6236 10600
rect 8852 10616 8904 10668
rect 9956 10659 10008 10668
rect 9956 10625 9958 10659
rect 9958 10625 10008 10659
rect 9956 10616 10008 10625
rect 10048 10659 10100 10668
rect 10048 10625 10060 10659
rect 10060 10625 10094 10659
rect 10094 10625 10100 10659
rect 10048 10616 10100 10625
rect 10968 10616 11020 10668
rect 11520 10616 11572 10668
rect 14280 10659 14332 10668
rect 14280 10625 14282 10659
rect 14282 10625 14332 10659
rect 14280 10616 14332 10625
rect 14556 10616 14608 10668
rect 14740 10616 14792 10668
rect 16580 10616 16632 10668
rect 8668 10548 8720 10600
rect 9036 10591 9088 10600
rect 9036 10557 9045 10591
rect 9045 10557 9079 10591
rect 9079 10557 9088 10591
rect 9036 10548 9088 10557
rect 7104 10480 7156 10532
rect 7564 10480 7616 10532
rect 8300 10480 8352 10532
rect 9312 10548 9364 10600
rect 9220 10455 9272 10464
rect 9220 10421 9229 10455
rect 9229 10421 9263 10455
rect 9263 10421 9272 10455
rect 9220 10412 9272 10421
rect 10692 10548 10744 10600
rect 11152 10480 11204 10532
rect 9864 10412 9916 10464
rect 11980 10455 12032 10464
rect 11980 10421 11989 10455
rect 11989 10421 12023 10455
rect 12023 10421 12032 10455
rect 11980 10412 12032 10421
rect 12348 10412 12400 10464
rect 12808 10523 12860 10532
rect 12808 10489 12817 10523
rect 12817 10489 12851 10523
rect 12851 10489 12860 10523
rect 12808 10480 12860 10489
rect 13084 10480 13136 10532
rect 13912 10591 13964 10600
rect 13912 10557 13921 10591
rect 13921 10557 13955 10591
rect 13955 10557 13964 10591
rect 13912 10548 13964 10557
rect 16396 10591 16448 10600
rect 16396 10557 16405 10591
rect 16405 10557 16439 10591
rect 16439 10557 16448 10591
rect 16396 10548 16448 10557
rect 16948 10548 17000 10600
rect 17132 10591 17184 10600
rect 17132 10557 17141 10591
rect 17141 10557 17175 10591
rect 17175 10557 17184 10591
rect 17132 10548 17184 10557
rect 18696 10548 18748 10600
rect 19064 10548 19116 10600
rect 20536 10548 20588 10600
rect 21180 10548 21232 10600
rect 21364 10548 21416 10600
rect 22560 10591 22612 10600
rect 22560 10557 22569 10591
rect 22569 10557 22603 10591
rect 22603 10557 22612 10591
rect 22560 10548 22612 10557
rect 14004 10480 14056 10532
rect 18512 10523 18564 10532
rect 18512 10489 18521 10523
rect 18521 10489 18555 10523
rect 18555 10489 18564 10523
rect 18512 10480 18564 10489
rect 22284 10480 22336 10532
rect 13544 10412 13596 10464
rect 14648 10412 14700 10464
rect 15292 10412 15344 10464
rect 17224 10412 17276 10464
rect 21548 10412 21600 10464
rect 21916 10412 21968 10464
rect 22376 10455 22428 10464
rect 22376 10421 22385 10455
rect 22385 10421 22419 10455
rect 22419 10421 22428 10455
rect 22376 10412 22428 10421
rect 23020 10795 23072 10804
rect 23020 10761 23029 10795
rect 23029 10761 23063 10795
rect 23063 10761 23072 10795
rect 23020 10752 23072 10761
rect 23756 10616 23808 10668
rect 24400 10616 24452 10668
rect 25964 10752 26016 10804
rect 26148 10752 26200 10804
rect 28172 10752 28224 10804
rect 29644 10752 29696 10804
rect 29736 10752 29788 10804
rect 28448 10727 28500 10736
rect 28448 10693 28457 10727
rect 28457 10693 28491 10727
rect 28491 10693 28500 10727
rect 28448 10684 28500 10693
rect 29184 10727 29236 10736
rect 29184 10693 29193 10727
rect 29193 10693 29227 10727
rect 29227 10693 29236 10727
rect 29184 10684 29236 10693
rect 25320 10616 25372 10668
rect 26516 10616 26568 10668
rect 26240 10591 26292 10600
rect 26240 10557 26249 10591
rect 26249 10557 26283 10591
rect 26283 10557 26292 10591
rect 26240 10548 26292 10557
rect 23664 10480 23716 10532
rect 23756 10480 23808 10532
rect 27988 10548 28040 10600
rect 27804 10480 27856 10532
rect 28816 10548 28868 10600
rect 29092 10548 29144 10600
rect 30104 10752 30156 10804
rect 30104 10616 30156 10668
rect 28356 10523 28408 10532
rect 28356 10489 28365 10523
rect 28365 10489 28399 10523
rect 28399 10489 28408 10523
rect 28356 10480 28408 10489
rect 25320 10412 25372 10464
rect 26148 10412 26200 10464
rect 26332 10412 26384 10464
rect 29276 10480 29328 10532
rect 28540 10412 28592 10464
rect 29828 10412 29880 10464
rect 29920 10412 29972 10464
rect 7988 10310 8040 10362
rect 8052 10310 8104 10362
rect 8116 10310 8168 10362
rect 8180 10310 8232 10362
rect 8244 10310 8296 10362
rect 15578 10310 15630 10362
rect 15642 10310 15694 10362
rect 15706 10310 15758 10362
rect 15770 10310 15822 10362
rect 15834 10310 15886 10362
rect 23168 10310 23220 10362
rect 23232 10310 23284 10362
rect 23296 10310 23348 10362
rect 23360 10310 23412 10362
rect 23424 10310 23476 10362
rect 30758 10310 30810 10362
rect 30822 10310 30874 10362
rect 30886 10310 30938 10362
rect 30950 10310 31002 10362
rect 31014 10310 31066 10362
rect 940 10072 992 10124
rect 1308 10208 1360 10260
rect 1768 10208 1820 10260
rect 3056 10208 3108 10260
rect 4068 10208 4120 10260
rect 4896 10208 4948 10260
rect 2964 10072 3016 10124
rect 1492 10031 1537 10056
rect 1537 10031 1544 10056
rect 1492 10004 1544 10031
rect 1860 10004 1912 10056
rect 3240 10047 3292 10056
rect 3240 10013 3249 10047
rect 3249 10013 3283 10047
rect 3283 10013 3292 10047
rect 3240 10004 3292 10013
rect 3792 10072 3844 10124
rect 9036 10208 9088 10260
rect 9312 10208 9364 10260
rect 9680 10208 9732 10260
rect 13544 10208 13596 10260
rect 14280 10251 14332 10260
rect 14280 10217 14295 10251
rect 14295 10217 14329 10251
rect 14329 10217 14332 10251
rect 14280 10208 14332 10217
rect 17868 10251 17920 10260
rect 17868 10217 17883 10251
rect 17883 10217 17917 10251
rect 17917 10217 17920 10251
rect 17868 10208 17920 10217
rect 18420 10208 18472 10260
rect 20352 10251 20404 10260
rect 20352 10217 20361 10251
rect 20361 10217 20395 10251
rect 20395 10217 20404 10251
rect 20352 10208 20404 10217
rect 6552 10140 6604 10192
rect 13452 10140 13504 10192
rect 4620 10004 4672 10056
rect 6092 10072 6144 10124
rect 2596 9936 2648 9988
rect 6368 10004 6420 10056
rect 3056 9911 3108 9920
rect 3056 9877 3065 9911
rect 3065 9877 3099 9911
rect 3099 9877 3108 9911
rect 3056 9868 3108 9877
rect 5908 9868 5960 9920
rect 6644 10004 6696 10056
rect 6828 10047 6880 10056
rect 6828 10013 6830 10047
rect 6830 10013 6880 10047
rect 6828 10004 6880 10013
rect 7656 10072 7708 10124
rect 10600 10072 10652 10124
rect 8392 10004 8444 10056
rect 8668 10047 8720 10056
rect 8668 10013 8677 10047
rect 8677 10013 8711 10047
rect 8711 10013 8720 10047
rect 8668 10004 8720 10013
rect 8944 10004 8996 10056
rect 13084 10072 13136 10124
rect 13912 10072 13964 10124
rect 16856 10115 16908 10124
rect 16856 10081 16865 10115
rect 16865 10081 16899 10115
rect 16899 10081 16908 10115
rect 16856 10072 16908 10081
rect 9588 10004 9640 10056
rect 10784 10004 10836 10056
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 11520 10047 11572 10056
rect 11520 10013 11522 10047
rect 11522 10013 11572 10047
rect 11520 10004 11572 10013
rect 11612 10047 11664 10056
rect 11612 10013 11624 10047
rect 11624 10013 11658 10047
rect 11658 10013 11664 10047
rect 11612 10004 11664 10013
rect 11704 10004 11756 10056
rect 14556 10047 14608 10056
rect 14556 10013 14565 10047
rect 14565 10013 14599 10047
rect 14599 10013 14608 10047
rect 14556 10004 14608 10013
rect 16672 10004 16724 10056
rect 13728 9936 13780 9988
rect 7656 9868 7708 9920
rect 9036 9868 9088 9920
rect 9588 9868 9640 9920
rect 11060 9868 11112 9920
rect 12348 9868 12400 9920
rect 14556 9868 14608 9920
rect 16488 9911 16540 9920
rect 16488 9877 16497 9911
rect 16497 9877 16531 9911
rect 16531 9877 16540 9911
rect 16488 9868 16540 9877
rect 20444 10140 20496 10192
rect 17132 10072 17184 10124
rect 18788 10072 18840 10124
rect 19892 10072 19944 10124
rect 17224 10004 17276 10056
rect 17408 10047 17460 10056
rect 17408 10013 17417 10047
rect 17417 10013 17451 10047
rect 17451 10013 17460 10047
rect 17408 10004 17460 10013
rect 19248 10004 19300 10056
rect 20628 10072 20680 10124
rect 22284 10208 22336 10260
rect 23940 10208 23992 10260
rect 24216 10208 24268 10260
rect 26148 10251 26200 10260
rect 26148 10217 26157 10251
rect 26157 10217 26191 10251
rect 26191 10217 26200 10251
rect 26148 10208 26200 10217
rect 26516 10208 26568 10260
rect 26332 10140 26384 10192
rect 20996 10072 21048 10124
rect 21272 10115 21324 10124
rect 21272 10081 21281 10115
rect 21281 10081 21315 10115
rect 21315 10081 21324 10115
rect 21272 10072 21324 10081
rect 21916 10072 21968 10124
rect 22376 10072 22428 10124
rect 21180 10004 21232 10056
rect 21456 10004 21508 10056
rect 19156 9868 19208 9920
rect 19708 9868 19760 9920
rect 20904 9911 20956 9920
rect 20904 9877 20913 9911
rect 20913 9877 20947 9911
rect 20947 9877 20956 9911
rect 20904 9868 20956 9877
rect 21548 9868 21600 9920
rect 24124 10047 24176 10056
rect 24124 10013 24133 10047
rect 24133 10013 24167 10047
rect 24167 10013 24176 10047
rect 24124 10004 24176 10013
rect 25780 10072 25832 10124
rect 24860 10047 24912 10056
rect 24860 10013 24869 10047
rect 24869 10013 24903 10047
rect 24903 10013 24912 10047
rect 24860 10004 24912 10013
rect 25044 10004 25096 10056
rect 26056 10004 26108 10056
rect 26240 10004 26292 10056
rect 26884 10047 26936 10056
rect 26884 10013 26896 10047
rect 26896 10013 26930 10047
rect 26930 10013 26936 10047
rect 26884 10004 26936 10013
rect 27620 10004 27672 10056
rect 28632 10115 28684 10124
rect 28632 10081 28641 10115
rect 28641 10081 28675 10115
rect 28675 10081 28684 10115
rect 28632 10072 28684 10081
rect 29644 10072 29696 10124
rect 24952 9868 25004 9920
rect 28172 9868 28224 9920
rect 30012 9911 30064 9920
rect 30012 9877 30021 9911
rect 30021 9877 30055 9911
rect 30055 9877 30064 9911
rect 30012 9868 30064 9877
rect 4193 9766 4245 9818
rect 4257 9766 4309 9818
rect 4321 9766 4373 9818
rect 4385 9766 4437 9818
rect 4449 9766 4501 9818
rect 11783 9766 11835 9818
rect 11847 9766 11899 9818
rect 11911 9766 11963 9818
rect 11975 9766 12027 9818
rect 12039 9766 12091 9818
rect 19373 9766 19425 9818
rect 19437 9766 19489 9818
rect 19501 9766 19553 9818
rect 19565 9766 19617 9818
rect 19629 9766 19681 9818
rect 26963 9766 27015 9818
rect 27027 9766 27079 9818
rect 27091 9766 27143 9818
rect 27155 9766 27207 9818
rect 27219 9766 27271 9818
rect 940 9571 992 9580
rect 940 9537 949 9571
rect 949 9537 983 9571
rect 983 9537 992 9571
rect 940 9528 992 9537
rect 5172 9596 5224 9648
rect 6644 9664 6696 9716
rect 6828 9664 6880 9716
rect 7012 9664 7064 9716
rect 8944 9664 8996 9716
rect 10692 9664 10744 9716
rect 3056 9528 3108 9580
rect 3976 9528 4028 9580
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 3240 9460 3292 9512
rect 3608 9460 3660 9512
rect 4988 9528 5040 9580
rect 5816 9528 5868 9580
rect 11612 9664 11664 9716
rect 17132 9664 17184 9716
rect 20720 9664 20772 9716
rect 21088 9664 21140 9716
rect 21364 9664 21416 9716
rect 24860 9664 24912 9716
rect 6368 9528 6420 9580
rect 8668 9528 8720 9580
rect 9312 9571 9364 9580
rect 9312 9537 9314 9571
rect 9314 9537 9364 9571
rect 1768 9324 1820 9376
rect 3608 9324 3660 9376
rect 4068 9324 4120 9376
rect 4344 9324 4396 9376
rect 5356 9392 5408 9444
rect 4804 9324 4856 9376
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 6920 9460 6972 9512
rect 8484 9460 8536 9512
rect 9312 9528 9364 9537
rect 9496 9528 9548 9580
rect 11060 9528 11112 9580
rect 9680 9503 9732 9512
rect 9680 9469 9689 9503
rect 9689 9469 9723 9503
rect 9723 9469 9732 9503
rect 9680 9460 9732 9469
rect 9772 9460 9824 9512
rect 11152 9503 11204 9512
rect 11152 9469 11161 9503
rect 11161 9469 11195 9503
rect 11195 9469 11204 9503
rect 11152 9460 11204 9469
rect 11520 9503 11572 9512
rect 11520 9469 11522 9503
rect 11522 9469 11572 9503
rect 11520 9460 11572 9469
rect 12164 9460 12216 9512
rect 6184 9392 6236 9444
rect 7564 9392 7616 9444
rect 6368 9324 6420 9376
rect 7104 9324 7156 9376
rect 7748 9324 7800 9376
rect 9036 9392 9088 9444
rect 13912 9460 13964 9512
rect 14372 9528 14424 9580
rect 16396 9571 16448 9580
rect 16396 9537 16405 9571
rect 16405 9537 16439 9571
rect 16439 9537 16448 9571
rect 16396 9528 16448 9537
rect 16580 9528 16632 9580
rect 16028 9460 16080 9512
rect 16948 9460 17000 9512
rect 17776 9528 17828 9580
rect 20720 9528 20772 9580
rect 20812 9571 20864 9580
rect 20812 9537 20821 9571
rect 20821 9537 20855 9571
rect 20855 9537 20864 9571
rect 20812 9528 20864 9537
rect 22744 9528 22796 9580
rect 17408 9460 17460 9512
rect 19340 9460 19392 9512
rect 19708 9460 19760 9512
rect 8668 9324 8720 9376
rect 12992 9367 13044 9376
rect 12992 9333 13001 9367
rect 13001 9333 13035 9367
rect 13035 9333 13044 9367
rect 12992 9324 13044 9333
rect 13728 9324 13780 9376
rect 14280 9367 14332 9376
rect 14280 9333 14295 9367
rect 14295 9333 14329 9367
rect 14329 9333 14332 9367
rect 14280 9324 14332 9333
rect 14648 9324 14700 9376
rect 15384 9324 15436 9376
rect 17868 9392 17920 9444
rect 17960 9324 18012 9376
rect 18144 9324 18196 9376
rect 18788 9392 18840 9444
rect 20812 9392 20864 9444
rect 21640 9503 21692 9512
rect 21640 9469 21649 9503
rect 21649 9469 21683 9503
rect 21683 9469 21692 9503
rect 21640 9460 21692 9469
rect 21916 9460 21968 9512
rect 24492 9596 24544 9648
rect 26884 9664 26936 9716
rect 27620 9664 27672 9716
rect 27988 9707 28040 9716
rect 27988 9673 27997 9707
rect 27997 9673 28031 9707
rect 28031 9673 28040 9707
rect 27988 9664 28040 9673
rect 27252 9571 27304 9580
rect 27252 9537 27261 9571
rect 27261 9537 27295 9571
rect 27295 9537 27304 9571
rect 27252 9528 27304 9537
rect 24124 9460 24176 9512
rect 24308 9503 24360 9512
rect 24308 9469 24317 9503
rect 24317 9469 24351 9503
rect 24351 9469 24360 9503
rect 24952 9503 25004 9512
rect 24308 9460 24360 9469
rect 24584 9392 24636 9444
rect 22008 9324 22060 9376
rect 23572 9324 23624 9376
rect 23940 9324 23992 9376
rect 24400 9324 24452 9376
rect 24952 9469 24954 9503
rect 24954 9469 25004 9503
rect 24952 9460 25004 9469
rect 25228 9460 25280 9512
rect 25688 9460 25740 9512
rect 25964 9460 26016 9512
rect 26332 9460 26384 9512
rect 29184 9528 29236 9580
rect 26792 9392 26844 9444
rect 27804 9392 27856 9444
rect 27252 9324 27304 9376
rect 28540 9460 28592 9512
rect 27988 9324 28040 9376
rect 28080 9324 28132 9376
rect 7988 9222 8040 9274
rect 8052 9222 8104 9274
rect 8116 9222 8168 9274
rect 8180 9222 8232 9274
rect 8244 9222 8296 9274
rect 15578 9222 15630 9274
rect 15642 9222 15694 9274
rect 15706 9222 15758 9274
rect 15770 9222 15822 9274
rect 15834 9222 15886 9274
rect 23168 9222 23220 9274
rect 23232 9222 23284 9274
rect 23296 9222 23348 9274
rect 23360 9222 23412 9274
rect 23424 9222 23476 9274
rect 30758 9222 30810 9274
rect 30822 9222 30874 9274
rect 30886 9222 30938 9274
rect 30950 9222 31002 9274
rect 31014 9222 31066 9274
rect 1308 9120 1360 9172
rect 2228 9120 2280 9172
rect 4068 9120 4120 9172
rect 6276 9120 6328 9172
rect 6368 9120 6420 9172
rect 7104 9120 7156 9172
rect 7196 9120 7248 9172
rect 3148 9095 3200 9104
rect 3148 9061 3157 9095
rect 3157 9061 3191 9095
rect 3191 9061 3200 9095
rect 3148 9052 3200 9061
rect 7748 9120 7800 9172
rect 9496 9163 9548 9172
rect 9496 9129 9505 9163
rect 9505 9129 9539 9163
rect 9539 9129 9548 9163
rect 9496 9120 9548 9129
rect 9680 9120 9732 9172
rect 11520 9120 11572 9172
rect 13728 9120 13780 9172
rect 16488 9120 16540 9172
rect 17868 9163 17920 9172
rect 1400 9027 1452 9036
rect 1400 8993 1402 9027
rect 1402 8993 1452 9027
rect 1400 8984 1452 8993
rect 1768 9027 1820 9036
rect 1768 8993 1777 9027
rect 1777 8993 1811 9027
rect 1811 8993 1820 9027
rect 1768 8984 1820 8993
rect 3792 8984 3844 9036
rect 1216 8916 1268 8968
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3608 8916 3660 8968
rect 3884 8916 3936 8968
rect 5632 9027 5684 9036
rect 5632 8993 5641 9027
rect 5641 8993 5675 9027
rect 5675 8993 5684 9027
rect 5632 8984 5684 8993
rect 5816 9027 5868 9036
rect 5816 8993 5825 9027
rect 5825 8993 5859 9027
rect 5859 8993 5868 9027
rect 5816 8984 5868 8993
rect 6644 8984 6696 9036
rect 7012 8984 7064 9036
rect 7288 8984 7340 9036
rect 7564 9027 7616 9036
rect 7564 8993 7573 9027
rect 7573 8993 7607 9027
rect 7607 8993 7616 9027
rect 7564 8984 7616 8993
rect 7656 9027 7708 9036
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 9312 8984 9364 9036
rect 4436 8916 4488 8968
rect 5540 8916 5592 8968
rect 6368 8916 6420 8968
rect 7472 8916 7524 8968
rect 6736 8891 6788 8900
rect 6736 8857 6745 8891
rect 6745 8857 6779 8891
rect 6779 8857 6788 8891
rect 6736 8848 6788 8857
rect 10600 8984 10652 9036
rect 10692 8984 10744 9036
rect 11152 9027 11204 9036
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11152 8984 11204 8993
rect 12808 9052 12860 9104
rect 17868 9129 17883 9163
rect 17883 9129 17917 9163
rect 17917 9129 17920 9163
rect 17868 9120 17920 9129
rect 19340 9120 19392 9172
rect 21640 9120 21692 9172
rect 22008 9120 22060 9172
rect 22652 9120 22704 9172
rect 23572 9120 23624 9172
rect 23756 9120 23808 9172
rect 24124 9120 24176 9172
rect 14372 8984 14424 9036
rect 14832 8984 14884 9036
rect 14924 8984 14976 9036
rect 16856 9027 16908 9036
rect 16856 8993 16865 9027
rect 16865 8993 16899 9027
rect 16899 8993 16908 9027
rect 16856 8984 16908 8993
rect 17316 8984 17368 9036
rect 17408 9027 17460 9036
rect 17408 8993 17417 9027
rect 17417 8993 17451 9027
rect 17451 8993 17460 9027
rect 17408 8984 17460 8993
rect 19800 9052 19852 9104
rect 20628 9052 20680 9104
rect 21088 9052 21140 9104
rect 8116 8959 8168 8968
rect 8116 8925 8128 8959
rect 8128 8925 8162 8959
rect 8162 8925 8168 8959
rect 8116 8916 8168 8925
rect 9036 8916 9088 8968
rect 3884 8780 3936 8832
rect 6184 8780 6236 8832
rect 6276 8780 6328 8832
rect 7104 8780 7156 8832
rect 7656 8848 7708 8900
rect 9772 8916 9824 8968
rect 11520 8916 11572 8968
rect 11704 8916 11756 8968
rect 13728 8959 13780 8968
rect 13728 8925 13737 8959
rect 13737 8925 13771 8959
rect 13771 8925 13780 8959
rect 13728 8916 13780 8925
rect 13912 8916 13964 8968
rect 18144 8959 18196 8968
rect 18144 8925 18153 8959
rect 18153 8925 18187 8959
rect 18187 8925 18196 8959
rect 18144 8916 18196 8925
rect 20168 8916 20220 8968
rect 20444 8984 20496 9036
rect 20904 8984 20956 9036
rect 25228 9120 25280 9172
rect 25688 9163 25740 9172
rect 25688 9129 25697 9163
rect 25697 9129 25731 9163
rect 25731 9129 25740 9163
rect 25688 9120 25740 9129
rect 24492 8984 24544 9036
rect 26056 8984 26108 9036
rect 29000 9120 29052 9172
rect 29368 9120 29420 9172
rect 30012 8984 30064 9036
rect 20812 8916 20864 8968
rect 11152 8848 11204 8900
rect 19064 8848 19116 8900
rect 21180 8848 21232 8900
rect 8852 8780 8904 8832
rect 9496 8780 9548 8832
rect 9864 8780 9916 8832
rect 11612 8780 11664 8832
rect 12716 8780 12768 8832
rect 14280 8780 14332 8832
rect 15108 8780 15160 8832
rect 16304 8823 16356 8832
rect 16304 8789 16313 8823
rect 16313 8789 16347 8823
rect 16347 8789 16356 8823
rect 16304 8780 16356 8789
rect 16764 8823 16816 8832
rect 16764 8789 16773 8823
rect 16773 8789 16807 8823
rect 16807 8789 16816 8823
rect 16764 8780 16816 8789
rect 18788 8780 18840 8832
rect 19708 8780 19760 8832
rect 22652 8916 22704 8968
rect 25320 8916 25372 8968
rect 25964 8916 26016 8968
rect 24952 8848 25004 8900
rect 26884 8959 26936 8968
rect 26884 8925 26896 8959
rect 26896 8925 26930 8959
rect 26930 8925 26936 8959
rect 26884 8916 26936 8925
rect 23480 8780 23532 8832
rect 24584 8780 24636 8832
rect 26056 8780 26108 8832
rect 26792 8780 26844 8832
rect 27988 8780 28040 8832
rect 28264 8823 28316 8832
rect 28264 8789 28273 8823
rect 28273 8789 28307 8823
rect 28307 8789 28316 8823
rect 28264 8780 28316 8789
rect 4193 8678 4245 8730
rect 4257 8678 4309 8730
rect 4321 8678 4373 8730
rect 4385 8678 4437 8730
rect 4449 8678 4501 8730
rect 11783 8678 11835 8730
rect 11847 8678 11899 8730
rect 11911 8678 11963 8730
rect 11975 8678 12027 8730
rect 12039 8678 12091 8730
rect 19373 8678 19425 8730
rect 19437 8678 19489 8730
rect 19501 8678 19553 8730
rect 19565 8678 19617 8730
rect 19629 8678 19681 8730
rect 26963 8678 27015 8730
rect 27027 8678 27079 8730
rect 27091 8678 27143 8730
rect 27155 8678 27207 8730
rect 27219 8678 27271 8730
rect 1216 8576 1268 8628
rect 2872 8576 2924 8628
rect 2412 8508 2464 8560
rect 3792 8576 3844 8628
rect 3884 8576 3936 8628
rect 6920 8576 6972 8628
rect 8392 8619 8444 8628
rect 8392 8585 8401 8619
rect 8401 8585 8435 8619
rect 8435 8585 8444 8619
rect 8392 8576 8444 8585
rect 7748 8508 7800 8560
rect 8760 8508 8812 8560
rect 11428 8576 11480 8628
rect 11704 8619 11756 8628
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 12164 8576 12216 8628
rect 4068 8440 4120 8492
rect 1032 8372 1084 8424
rect 2136 8372 2188 8424
rect 2504 8372 2556 8424
rect 1584 8236 1636 8288
rect 2780 8279 2832 8288
rect 2780 8245 2789 8279
rect 2789 8245 2823 8279
rect 2823 8245 2832 8279
rect 2780 8236 2832 8245
rect 5448 8372 5500 8424
rect 5908 8440 5960 8492
rect 6184 8440 6236 8492
rect 7012 8440 7064 8492
rect 7288 8440 7340 8492
rect 9864 8440 9916 8492
rect 11244 8440 11296 8492
rect 11520 8440 11572 8492
rect 13728 8576 13780 8628
rect 16304 8576 16356 8628
rect 18144 8619 18196 8628
rect 18144 8585 18153 8619
rect 18153 8585 18187 8619
rect 18187 8585 18196 8619
rect 18144 8576 18196 8585
rect 19248 8576 19300 8628
rect 12900 8508 12952 8560
rect 3792 8236 3844 8288
rect 3884 8236 3936 8288
rect 5540 8236 5592 8288
rect 6000 8279 6052 8288
rect 6000 8245 6015 8279
rect 6015 8245 6049 8279
rect 6049 8245 6052 8279
rect 6000 8236 6052 8245
rect 6184 8236 6236 8288
rect 6552 8236 6604 8288
rect 7012 8236 7064 8288
rect 7840 8236 7892 8288
rect 9036 8372 9088 8424
rect 8392 8236 8444 8288
rect 8576 8236 8628 8288
rect 8852 8236 8904 8288
rect 9128 8236 9180 8288
rect 9496 8372 9548 8424
rect 9680 8415 9732 8440
rect 9680 8388 9689 8415
rect 9689 8388 9723 8415
rect 9723 8388 9732 8415
rect 9312 8304 9364 8356
rect 9772 8372 9824 8424
rect 11336 8372 11388 8424
rect 14188 8483 14240 8492
rect 14188 8449 14200 8483
rect 14200 8449 14234 8483
rect 14234 8449 14240 8483
rect 14188 8440 14240 8449
rect 14280 8440 14332 8492
rect 21548 8576 21600 8628
rect 9404 8279 9456 8288
rect 9404 8245 9413 8279
rect 9413 8245 9447 8279
rect 9447 8245 9456 8279
rect 9404 8236 9456 8245
rect 9956 8236 10008 8288
rect 10692 8236 10744 8288
rect 12164 8304 12216 8356
rect 12256 8304 12308 8356
rect 13820 8372 13872 8424
rect 14372 8372 14424 8424
rect 15936 8415 15988 8424
rect 15936 8381 15945 8415
rect 15945 8381 15979 8415
rect 15979 8381 15988 8415
rect 15936 8372 15988 8381
rect 16580 8372 16632 8424
rect 18696 8415 18748 8424
rect 18696 8381 18705 8415
rect 18705 8381 18739 8415
rect 18739 8381 18748 8415
rect 18696 8372 18748 8381
rect 19064 8372 19116 8424
rect 19432 8415 19484 8424
rect 19432 8381 19441 8415
rect 19441 8381 19475 8415
rect 19475 8381 19484 8415
rect 19432 8372 19484 8381
rect 21180 8372 21232 8424
rect 25412 8576 25464 8628
rect 26884 8576 26936 8628
rect 28264 8576 28316 8628
rect 23480 8440 23532 8492
rect 26240 8440 26292 8492
rect 26516 8440 26568 8492
rect 21824 8372 21876 8424
rect 22284 8415 22336 8424
rect 22284 8381 22293 8415
rect 22293 8381 22327 8415
rect 22327 8381 22336 8415
rect 22284 8372 22336 8381
rect 23848 8415 23900 8424
rect 23848 8381 23857 8415
rect 23857 8381 23891 8415
rect 23891 8381 23900 8415
rect 23848 8372 23900 8381
rect 23940 8372 23992 8424
rect 25964 8372 26016 8424
rect 26976 8372 27028 8424
rect 28080 8372 28132 8424
rect 23756 8304 23808 8356
rect 27988 8304 28040 8356
rect 29460 8372 29512 8424
rect 31392 8372 31444 8424
rect 30012 8304 30064 8356
rect 12808 8279 12860 8288
rect 12808 8245 12817 8279
rect 12817 8245 12851 8279
rect 12851 8245 12860 8279
rect 12808 8236 12860 8245
rect 14924 8236 14976 8288
rect 16396 8279 16448 8288
rect 16396 8245 16411 8279
rect 16411 8245 16445 8279
rect 16445 8245 16448 8279
rect 16396 8236 16448 8245
rect 18328 8236 18380 8288
rect 19156 8279 19208 8288
rect 19156 8245 19171 8279
rect 19171 8245 19205 8279
rect 19205 8245 19208 8279
rect 19156 8236 19208 8245
rect 21364 8236 21416 8288
rect 21456 8236 21508 8288
rect 23572 8236 23624 8288
rect 24216 8236 24268 8288
rect 25228 8236 25280 8288
rect 26608 8236 26660 8288
rect 27068 8236 27120 8288
rect 27804 8236 27856 8288
rect 28540 8279 28592 8288
rect 28540 8245 28549 8279
rect 28549 8245 28583 8279
rect 28583 8245 28592 8279
rect 28540 8236 28592 8245
rect 29276 8236 29328 8288
rect 29736 8279 29788 8288
rect 29736 8245 29745 8279
rect 29745 8245 29779 8279
rect 29779 8245 29788 8279
rect 29736 8236 29788 8245
rect 30104 8236 30156 8288
rect 7988 8134 8040 8186
rect 8052 8134 8104 8186
rect 8116 8134 8168 8186
rect 8180 8134 8232 8186
rect 8244 8134 8296 8186
rect 15578 8134 15630 8186
rect 15642 8134 15694 8186
rect 15706 8134 15758 8186
rect 15770 8134 15822 8186
rect 15834 8134 15886 8186
rect 23168 8134 23220 8186
rect 23232 8134 23284 8186
rect 23296 8134 23348 8186
rect 23360 8134 23412 8186
rect 23424 8134 23476 8186
rect 30758 8134 30810 8186
rect 30822 8134 30874 8186
rect 30886 8134 30938 8186
rect 30950 8134 31002 8186
rect 31014 8134 31066 8186
rect 1584 8032 1636 8084
rect 3516 8032 3568 8084
rect 3608 7964 3660 8016
rect 5448 8032 5500 8084
rect 8392 8032 8444 8084
rect 9496 8032 9548 8084
rect 10876 8032 10928 8084
rect 11704 8032 11756 8084
rect 14924 8032 14976 8084
rect 15292 8032 15344 8084
rect 16396 8032 16448 8084
rect 18144 8032 18196 8084
rect 19892 8032 19944 8084
rect 20168 8075 20220 8084
rect 20168 8041 20177 8075
rect 20177 8041 20211 8075
rect 20211 8041 20220 8075
rect 20168 8032 20220 8041
rect 6368 7964 6420 8016
rect 10416 7964 10468 8016
rect 11612 7964 11664 8016
rect 1124 7939 1176 7948
rect 1124 7905 1133 7939
rect 1133 7905 1167 7939
rect 1167 7905 1176 7939
rect 1124 7896 1176 7905
rect 1032 7828 1084 7880
rect 1492 7828 1544 7880
rect 5448 7896 5500 7948
rect 6000 7896 6052 7948
rect 1952 7871 2004 7880
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 3516 7871 3568 7880
rect 3516 7837 3525 7871
rect 3525 7837 3559 7871
rect 3559 7837 3568 7871
rect 3516 7828 3568 7837
rect 3700 7828 3752 7880
rect 3884 7871 3936 7880
rect 3884 7837 3886 7871
rect 3886 7837 3936 7871
rect 3884 7828 3936 7837
rect 4160 7828 4212 7880
rect 6368 7828 6420 7880
rect 7104 7896 7156 7948
rect 9036 7896 9088 7948
rect 12808 7896 12860 7948
rect 20996 7964 21048 8016
rect 6644 7828 6696 7880
rect 6828 7871 6880 7880
rect 6828 7837 6830 7871
rect 6830 7837 6880 7871
rect 6828 7828 6880 7837
rect 6920 7855 6965 7880
rect 6965 7855 6972 7880
rect 6920 7828 6972 7855
rect 9128 7828 9180 7880
rect 9404 7871 9456 7880
rect 9404 7837 9413 7871
rect 9413 7837 9447 7871
rect 9447 7837 9456 7871
rect 9404 7828 9456 7837
rect 11244 7828 11296 7880
rect 940 7735 992 7744
rect 940 7701 949 7735
rect 949 7701 983 7735
rect 983 7701 992 7735
rect 940 7692 992 7701
rect 1492 7692 1544 7744
rect 3148 7692 3200 7744
rect 5540 7735 5592 7744
rect 5540 7701 5549 7735
rect 5549 7701 5583 7735
rect 5583 7701 5592 7735
rect 5540 7692 5592 7701
rect 12716 7828 12768 7880
rect 13820 7871 13872 7880
rect 13820 7837 13829 7871
rect 13829 7837 13863 7871
rect 13863 7837 13872 7871
rect 13820 7828 13872 7837
rect 15936 7896 15988 7948
rect 14556 7871 14608 7880
rect 14556 7837 14565 7871
rect 14565 7837 14599 7871
rect 14599 7837 14608 7871
rect 14556 7828 14608 7837
rect 14740 7828 14792 7880
rect 16396 7828 16448 7880
rect 22468 8032 22520 8084
rect 22652 8032 22704 8084
rect 23572 8032 23624 8084
rect 25320 8075 25372 8084
rect 25320 8041 25329 8075
rect 25329 8041 25363 8075
rect 25363 8041 25372 8075
rect 25320 8032 25372 8041
rect 26700 8032 26752 8084
rect 28080 8032 28132 8084
rect 29552 8075 29604 8084
rect 29552 8041 29561 8075
rect 29561 8041 29595 8075
rect 29595 8041 29604 8075
rect 29552 8032 29604 8041
rect 16856 7871 16908 7880
rect 16856 7837 16865 7871
rect 16865 7837 16899 7871
rect 16899 7837 16908 7871
rect 16856 7828 16908 7837
rect 12256 7692 12308 7744
rect 15660 7803 15712 7812
rect 15660 7769 15669 7803
rect 15669 7769 15703 7803
rect 15703 7769 15712 7803
rect 15660 7760 15712 7769
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 14372 7692 14424 7744
rect 15016 7692 15068 7744
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 18972 7828 19024 7880
rect 19064 7871 19116 7880
rect 19064 7837 19073 7871
rect 19073 7837 19107 7871
rect 19107 7837 19116 7871
rect 19064 7828 19116 7837
rect 19156 7828 19208 7880
rect 26332 7896 26384 7948
rect 26424 7896 26476 7948
rect 26792 7896 26844 7948
rect 26884 7896 26936 7948
rect 27068 7896 27120 7948
rect 27528 7896 27580 7948
rect 27988 7896 28040 7948
rect 28448 7939 28500 7948
rect 28448 7905 28457 7939
rect 28457 7905 28491 7939
rect 28491 7905 28500 7939
rect 28448 7896 28500 7905
rect 29644 7896 29696 7948
rect 30104 7939 30156 7948
rect 30104 7905 30113 7939
rect 30113 7905 30147 7939
rect 30147 7905 30156 7939
rect 30104 7896 30156 7905
rect 21272 7871 21324 7880
rect 21272 7837 21281 7871
rect 21281 7837 21315 7871
rect 21315 7837 21324 7871
rect 21272 7828 21324 7837
rect 21456 7828 21508 7880
rect 22652 7828 22704 7880
rect 22836 7828 22888 7880
rect 23204 7828 23256 7880
rect 26056 7828 26108 7880
rect 27712 7871 27764 7880
rect 27712 7837 27721 7871
rect 27721 7837 27755 7871
rect 27755 7837 27764 7871
rect 27712 7828 27764 7837
rect 28172 7873 28224 7880
rect 28172 7839 28200 7873
rect 28200 7839 28224 7873
rect 28172 7828 28224 7839
rect 18696 7692 18748 7744
rect 18880 7692 18932 7744
rect 19432 7692 19484 7744
rect 22836 7692 22888 7744
rect 25688 7735 25740 7744
rect 25688 7701 25697 7735
rect 25697 7701 25731 7735
rect 25731 7701 25740 7735
rect 25688 7692 25740 7701
rect 25964 7735 26016 7744
rect 25964 7701 25973 7735
rect 25973 7701 26007 7735
rect 26007 7701 26016 7735
rect 25964 7692 26016 7701
rect 26792 7735 26844 7744
rect 26792 7701 26801 7735
rect 26801 7701 26835 7735
rect 26835 7701 26844 7735
rect 26792 7692 26844 7701
rect 28264 7692 28316 7744
rect 28816 7692 28868 7744
rect 4193 7590 4245 7642
rect 4257 7590 4309 7642
rect 4321 7590 4373 7642
rect 4385 7590 4437 7642
rect 4449 7590 4501 7642
rect 11783 7590 11835 7642
rect 11847 7590 11899 7642
rect 11911 7590 11963 7642
rect 11975 7590 12027 7642
rect 12039 7590 12091 7642
rect 19373 7590 19425 7642
rect 19437 7590 19489 7642
rect 19501 7590 19553 7642
rect 19565 7590 19617 7642
rect 19629 7590 19681 7642
rect 26963 7590 27015 7642
rect 27027 7590 27079 7642
rect 27091 7590 27143 7642
rect 27155 7590 27207 7642
rect 27219 7590 27271 7642
rect 940 7488 992 7540
rect 2136 7352 2188 7404
rect 3056 7488 3108 7540
rect 3516 7488 3568 7540
rect 3608 7488 3660 7540
rect 4068 7488 4120 7540
rect 5816 7531 5868 7540
rect 5816 7497 5825 7531
rect 5825 7497 5859 7531
rect 5859 7497 5868 7531
rect 5816 7488 5868 7497
rect 6000 7420 6052 7472
rect 1032 7284 1084 7336
rect 3700 7395 3752 7404
rect 3700 7361 3702 7395
rect 3702 7361 3752 7395
rect 3700 7352 3752 7361
rect 6828 7488 6880 7540
rect 7012 7488 7064 7540
rect 9680 7488 9732 7540
rect 7564 7420 7616 7472
rect 6276 7352 6328 7404
rect 6552 7395 6604 7404
rect 6552 7361 6564 7395
rect 6564 7361 6598 7395
rect 6598 7361 6604 7395
rect 6552 7352 6604 7361
rect 7748 7352 7800 7404
rect 9404 7395 9456 7404
rect 5724 7327 5776 7336
rect 5724 7293 5733 7327
rect 5733 7293 5767 7327
rect 5767 7293 5776 7327
rect 5724 7284 5776 7293
rect 5908 7284 5960 7336
rect 6644 7284 6696 7336
rect 3240 7216 3292 7268
rect 8576 7216 8628 7268
rect 1584 7148 1636 7200
rect 2964 7148 3016 7200
rect 6552 7191 6604 7200
rect 6552 7157 6567 7191
rect 6567 7157 6601 7191
rect 6601 7157 6604 7191
rect 6552 7148 6604 7157
rect 6920 7148 6972 7200
rect 7564 7148 7616 7200
rect 8484 7191 8536 7200
rect 8484 7157 8493 7191
rect 8493 7157 8527 7191
rect 8527 7157 8536 7191
rect 8484 7148 8536 7157
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 9404 7361 9406 7395
rect 9406 7361 9456 7395
rect 9404 7352 9456 7361
rect 13452 7488 13504 7540
rect 14004 7488 14056 7540
rect 14556 7488 14608 7540
rect 12808 7420 12860 7472
rect 13084 7420 13136 7472
rect 11244 7395 11296 7404
rect 11244 7361 11253 7395
rect 11253 7361 11287 7395
rect 11287 7361 11296 7395
rect 11244 7352 11296 7361
rect 12348 7352 12400 7404
rect 10968 7284 11020 7336
rect 11888 7284 11940 7336
rect 12716 7284 12768 7336
rect 16672 7420 16724 7472
rect 13820 7352 13872 7404
rect 14740 7395 14792 7404
rect 14740 7361 14749 7395
rect 14749 7361 14783 7395
rect 14783 7361 14792 7395
rect 14740 7352 14792 7361
rect 9128 7216 9180 7268
rect 14464 7327 14516 7336
rect 14464 7293 14473 7327
rect 14473 7293 14507 7327
rect 14507 7293 14516 7327
rect 14924 7352 14976 7404
rect 15384 7352 15436 7404
rect 15476 7395 15528 7404
rect 15476 7361 15485 7395
rect 15485 7361 15519 7395
rect 15519 7361 15528 7395
rect 15476 7352 15528 7361
rect 19064 7488 19116 7540
rect 18052 7463 18104 7472
rect 18052 7429 18061 7463
rect 18061 7429 18095 7463
rect 18095 7429 18104 7463
rect 18052 7420 18104 7429
rect 18236 7420 18288 7472
rect 18880 7352 18932 7404
rect 19064 7395 19116 7404
rect 19064 7361 19066 7395
rect 19066 7361 19116 7395
rect 19064 7352 19116 7361
rect 20720 7463 20772 7472
rect 20720 7429 20729 7463
rect 20729 7429 20763 7463
rect 20763 7429 20772 7463
rect 20720 7420 20772 7429
rect 22744 7531 22796 7540
rect 22744 7497 22753 7531
rect 22753 7497 22787 7531
rect 22787 7497 22796 7531
rect 22744 7488 22796 7497
rect 24676 7488 24728 7540
rect 25044 7488 25096 7540
rect 26700 7488 26752 7540
rect 28724 7531 28776 7540
rect 28724 7497 28733 7531
rect 28733 7497 28767 7531
rect 28767 7497 28776 7531
rect 28724 7488 28776 7497
rect 21180 7352 21232 7404
rect 14464 7284 14516 7293
rect 17408 7327 17460 7336
rect 17408 7293 17417 7327
rect 17417 7293 17451 7327
rect 17451 7293 17460 7327
rect 17408 7284 17460 7293
rect 14832 7216 14884 7268
rect 16488 7216 16540 7268
rect 17868 7284 17920 7336
rect 18052 7284 18104 7336
rect 18144 7284 18196 7336
rect 18328 7284 18380 7336
rect 18696 7327 18748 7336
rect 18696 7293 18705 7327
rect 18705 7293 18739 7327
rect 18739 7293 18748 7327
rect 18696 7284 18748 7293
rect 21640 7327 21692 7336
rect 21640 7293 21649 7327
rect 21649 7293 21683 7327
rect 21683 7293 21692 7327
rect 21640 7284 21692 7293
rect 23848 7327 23900 7336
rect 23848 7293 23857 7327
rect 23857 7293 23891 7327
rect 23891 7293 23900 7327
rect 23848 7284 23900 7293
rect 24032 7352 24084 7404
rect 24400 7352 24452 7404
rect 24952 7352 25004 7404
rect 26424 7352 26476 7404
rect 28908 7420 28960 7472
rect 27804 7352 27856 7404
rect 25044 7284 25096 7336
rect 25872 7284 25924 7336
rect 29920 7352 29972 7404
rect 10600 7148 10652 7200
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 12072 7148 12124 7200
rect 12624 7148 12676 7200
rect 13820 7148 13872 7200
rect 15384 7148 15436 7200
rect 17224 7191 17276 7200
rect 17224 7157 17233 7191
rect 17233 7157 17267 7191
rect 17267 7157 17276 7191
rect 17224 7148 17276 7157
rect 17500 7191 17552 7200
rect 17500 7157 17509 7191
rect 17509 7157 17543 7191
rect 17543 7157 17552 7191
rect 17500 7148 17552 7157
rect 23204 7259 23256 7268
rect 23204 7225 23213 7259
rect 23213 7225 23247 7259
rect 23247 7225 23256 7259
rect 23204 7216 23256 7225
rect 23572 7259 23624 7268
rect 23572 7225 23581 7259
rect 23581 7225 23615 7259
rect 23615 7225 23624 7259
rect 23572 7216 23624 7225
rect 26332 7259 26384 7268
rect 26332 7225 26341 7259
rect 26341 7225 26375 7259
rect 26375 7225 26384 7259
rect 26332 7216 26384 7225
rect 29276 7284 29328 7336
rect 18236 7148 18288 7200
rect 19248 7148 19300 7200
rect 21364 7191 21416 7200
rect 21364 7157 21379 7191
rect 21379 7157 21413 7191
rect 21413 7157 21416 7191
rect 21364 7148 21416 7157
rect 21916 7148 21968 7200
rect 29736 7216 29788 7268
rect 24216 7148 24268 7200
rect 24676 7148 24728 7200
rect 28448 7148 28500 7200
rect 29000 7191 29052 7200
rect 29000 7157 29009 7191
rect 29009 7157 29043 7191
rect 29043 7157 29052 7191
rect 29000 7148 29052 7157
rect 29552 7148 29604 7200
rect 7988 7046 8040 7098
rect 8052 7046 8104 7098
rect 8116 7046 8168 7098
rect 8180 7046 8232 7098
rect 8244 7046 8296 7098
rect 15578 7046 15630 7098
rect 15642 7046 15694 7098
rect 15706 7046 15758 7098
rect 15770 7046 15822 7098
rect 15834 7046 15886 7098
rect 23168 7046 23220 7098
rect 23232 7046 23284 7098
rect 23296 7046 23348 7098
rect 23360 7046 23412 7098
rect 23424 7046 23476 7098
rect 30758 7046 30810 7098
rect 30822 7046 30874 7098
rect 30886 7046 30938 7098
rect 30950 7046 31002 7098
rect 31014 7046 31066 7098
rect 1584 6987 1636 6996
rect 1584 6953 1599 6987
rect 1599 6953 1633 6987
rect 1633 6953 1636 6987
rect 1584 6944 1636 6953
rect 2136 6944 2188 6996
rect 3148 6944 3200 6996
rect 3240 6944 3292 6996
rect 5448 6944 5500 6996
rect 6460 6944 6512 6996
rect 6920 6987 6972 6996
rect 6920 6953 6935 6987
rect 6935 6953 6969 6987
rect 6969 6953 6972 6987
rect 6920 6944 6972 6953
rect 9496 6944 9548 6996
rect 10508 6987 10560 6996
rect 10508 6953 10517 6987
rect 10517 6953 10551 6987
rect 10551 6953 10560 6987
rect 10508 6944 10560 6953
rect 10692 6944 10744 6996
rect 11704 6987 11756 6996
rect 11704 6953 11713 6987
rect 11713 6953 11747 6987
rect 11747 6953 11756 6987
rect 11704 6944 11756 6953
rect 2320 6808 2372 6860
rect 3608 6876 3660 6928
rect 6184 6876 6236 6928
rect 11612 6876 11664 6928
rect 12072 6944 12124 6996
rect 14464 6944 14516 6996
rect 15476 6944 15528 6996
rect 16856 6944 16908 6996
rect 18236 6944 18288 6996
rect 21272 6944 21324 6996
rect 21456 6944 21508 6996
rect 24860 6944 24912 6996
rect 24952 6944 25004 6996
rect 28080 6944 28132 6996
rect 24032 6876 24084 6928
rect 3516 6851 3568 6860
rect 3516 6817 3525 6851
rect 3525 6817 3559 6851
rect 3559 6817 3568 6851
rect 3516 6808 3568 6817
rect 4988 6808 5040 6860
rect 6092 6808 6144 6860
rect 1768 6740 1820 6792
rect 1032 6672 1084 6724
rect 2044 6604 2096 6656
rect 3700 6740 3752 6792
rect 5816 6715 5868 6724
rect 5816 6681 5825 6715
rect 5825 6681 5859 6715
rect 5859 6681 5868 6715
rect 5816 6672 5868 6681
rect 4896 6604 4948 6656
rect 5356 6647 5408 6656
rect 5356 6613 5365 6647
rect 5365 6613 5399 6647
rect 5399 6613 5408 6647
rect 5356 6604 5408 6613
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 6644 6740 6696 6792
rect 6920 6783 6972 6792
rect 6920 6749 6932 6783
rect 6932 6749 6966 6783
rect 6966 6749 6972 6783
rect 6920 6740 6972 6749
rect 8760 6808 8812 6860
rect 9036 6808 9088 6860
rect 10968 6808 11020 6860
rect 11152 6851 11204 6860
rect 11152 6817 11161 6851
rect 11161 6817 11195 6851
rect 11195 6817 11204 6851
rect 11152 6808 11204 6817
rect 11336 6808 11388 6860
rect 8484 6672 8536 6724
rect 11704 6808 11756 6860
rect 12256 6808 12308 6860
rect 12808 6808 12860 6860
rect 12900 6851 12952 6860
rect 12900 6817 12909 6851
rect 12909 6817 12943 6851
rect 12943 6817 12952 6851
rect 12900 6808 12952 6817
rect 12992 6808 13044 6860
rect 13636 6808 13688 6860
rect 14648 6808 14700 6860
rect 15200 6851 15252 6860
rect 15200 6817 15209 6851
rect 15209 6817 15243 6851
rect 15243 6817 15252 6851
rect 15200 6808 15252 6817
rect 16488 6851 16540 6860
rect 16488 6817 16497 6851
rect 16497 6817 16531 6851
rect 16531 6817 16540 6851
rect 16488 6808 16540 6817
rect 16304 6740 16356 6792
rect 17960 6808 18012 6860
rect 19340 6851 19392 6860
rect 7932 6604 7984 6656
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 9312 6604 9364 6656
rect 9404 6604 9456 6656
rect 13820 6672 13872 6724
rect 11888 6604 11940 6656
rect 16672 6672 16724 6724
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 16396 6604 16448 6656
rect 16580 6604 16632 6656
rect 16948 6740 17000 6792
rect 17224 6783 17276 6792
rect 17224 6749 17236 6783
rect 17236 6749 17270 6783
rect 17270 6749 17276 6783
rect 17224 6740 17276 6749
rect 17500 6783 17552 6792
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 17684 6740 17736 6792
rect 19340 6817 19342 6851
rect 19342 6817 19392 6851
rect 19340 6808 19392 6817
rect 18972 6783 19024 6792
rect 18972 6749 18981 6783
rect 18981 6749 19015 6783
rect 19015 6749 19024 6783
rect 18972 6740 19024 6749
rect 20536 6808 20588 6860
rect 21180 6808 21232 6860
rect 21916 6808 21968 6860
rect 20628 6740 20680 6792
rect 21548 6783 21600 6792
rect 21548 6749 21557 6783
rect 21557 6749 21591 6783
rect 21591 6749 21600 6783
rect 21548 6740 21600 6749
rect 22560 6783 22612 6792
rect 22560 6749 22569 6783
rect 22569 6749 22603 6783
rect 22603 6749 22612 6783
rect 22560 6740 22612 6749
rect 23204 6740 23256 6792
rect 18788 6647 18840 6656
rect 18788 6613 18797 6647
rect 18797 6613 18831 6647
rect 18831 6613 18840 6647
rect 18788 6604 18840 6613
rect 19340 6604 19392 6656
rect 20076 6604 20128 6656
rect 23572 6740 23624 6792
rect 25688 6808 25740 6860
rect 26424 6808 26476 6860
rect 27712 6851 27764 6860
rect 27712 6817 27721 6851
rect 27721 6817 27755 6851
rect 27755 6817 27764 6851
rect 27712 6808 27764 6817
rect 28356 6808 28408 6860
rect 29828 6808 29880 6860
rect 26240 6740 26292 6792
rect 26700 6740 26752 6792
rect 25872 6672 25924 6724
rect 24492 6604 24544 6656
rect 26424 6604 26476 6656
rect 26516 6604 26568 6656
rect 26884 6604 26936 6656
rect 27344 6647 27396 6656
rect 27344 6613 27353 6647
rect 27353 6613 27387 6647
rect 27387 6613 27396 6647
rect 27344 6604 27396 6613
rect 29092 6604 29144 6656
rect 31208 6604 31260 6656
rect 4193 6502 4245 6554
rect 4257 6502 4309 6554
rect 4321 6502 4373 6554
rect 4385 6502 4437 6554
rect 4449 6502 4501 6554
rect 11783 6502 11835 6554
rect 11847 6502 11899 6554
rect 11911 6502 11963 6554
rect 11975 6502 12027 6554
rect 12039 6502 12091 6554
rect 19373 6502 19425 6554
rect 19437 6502 19489 6554
rect 19501 6502 19553 6554
rect 19565 6502 19617 6554
rect 19629 6502 19681 6554
rect 26963 6502 27015 6554
rect 27027 6502 27079 6554
rect 27091 6502 27143 6554
rect 27155 6502 27207 6554
rect 27219 6502 27271 6554
rect 5356 6400 5408 6452
rect 5448 6400 5500 6452
rect 4896 6332 4948 6384
rect 3516 6264 3568 6316
rect 3700 6307 3752 6316
rect 3700 6273 3702 6307
rect 3702 6273 3752 6307
rect 3700 6264 3752 6273
rect 8300 6400 8352 6452
rect 7932 6375 7984 6384
rect 7932 6341 7941 6375
rect 7941 6341 7975 6375
rect 7975 6341 7984 6375
rect 7932 6332 7984 6341
rect 9128 6443 9180 6452
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 9220 6400 9272 6452
rect 9680 6400 9732 6452
rect 11428 6400 11480 6452
rect 14464 6400 14516 6452
rect 16488 6400 16540 6452
rect 16672 6443 16724 6452
rect 16672 6409 16681 6443
rect 16681 6409 16715 6443
rect 16715 6409 16724 6443
rect 16672 6400 16724 6409
rect 16856 6400 16908 6452
rect 17684 6400 17736 6452
rect 17960 6400 18012 6452
rect 19892 6400 19944 6452
rect 6460 6264 6512 6316
rect 1584 6196 1636 6248
rect 2136 6196 2188 6248
rect 4804 6196 4856 6248
rect 5908 6196 5960 6248
rect 6736 6264 6788 6316
rect 7472 6264 7524 6316
rect 6920 6196 6972 6248
rect 7656 6196 7708 6248
rect 8668 6332 8720 6384
rect 9036 6264 9088 6316
rect 5632 6128 5684 6180
rect 8484 6128 8536 6180
rect 1308 6060 1360 6112
rect 1584 6060 1636 6112
rect 1768 6060 1820 6112
rect 2412 6060 2464 6112
rect 4528 6060 4580 6112
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 6552 6103 6604 6112
rect 6552 6069 6567 6103
rect 6567 6069 6601 6103
rect 6601 6069 6604 6103
rect 6552 6060 6604 6069
rect 6736 6060 6788 6112
rect 11060 6332 11112 6384
rect 9312 6264 9364 6316
rect 12624 6264 12676 6316
rect 12256 6239 12308 6248
rect 12256 6205 12265 6239
rect 12265 6205 12299 6239
rect 12299 6205 12308 6239
rect 12256 6196 12308 6205
rect 12532 6239 12584 6248
rect 12532 6205 12541 6239
rect 12541 6205 12575 6239
rect 12575 6205 12584 6239
rect 12532 6196 12584 6205
rect 14372 6332 14424 6384
rect 13820 6264 13872 6316
rect 14280 6264 14332 6316
rect 15108 6307 15160 6316
rect 15108 6273 15120 6307
rect 15120 6273 15154 6307
rect 15154 6273 15160 6307
rect 15108 6264 15160 6273
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 16396 6264 16448 6316
rect 19708 6332 19760 6384
rect 9404 6060 9456 6112
rect 9496 6060 9548 6112
rect 10140 6060 10192 6112
rect 11704 6060 11756 6112
rect 13636 6128 13688 6180
rect 14740 6196 14792 6248
rect 13912 6128 13964 6180
rect 17316 6196 17368 6248
rect 16948 6128 17000 6180
rect 17132 6171 17184 6180
rect 17132 6137 17141 6171
rect 17141 6137 17175 6171
rect 17175 6137 17184 6171
rect 17132 6128 17184 6137
rect 17960 6196 18012 6248
rect 19340 6307 19392 6316
rect 19340 6273 19349 6307
rect 19349 6273 19383 6307
rect 19383 6273 19392 6307
rect 19340 6264 19392 6273
rect 21640 6400 21692 6452
rect 22560 6400 22612 6452
rect 23204 6400 23256 6452
rect 22836 6332 22888 6384
rect 24308 6332 24360 6384
rect 24400 6332 24452 6384
rect 26056 6332 26108 6384
rect 19064 6196 19116 6248
rect 19248 6196 19300 6248
rect 19524 6128 19576 6180
rect 12164 6060 12216 6112
rect 12348 6103 12400 6112
rect 12348 6069 12357 6103
rect 12357 6069 12391 6103
rect 12391 6069 12400 6103
rect 12348 6060 12400 6069
rect 12624 6103 12676 6112
rect 12624 6069 12633 6103
rect 12633 6069 12667 6103
rect 12667 6069 12676 6103
rect 12624 6060 12676 6069
rect 12716 6060 12768 6112
rect 14556 6060 14608 6112
rect 14924 6060 14976 6112
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 17684 6103 17736 6112
rect 17684 6069 17693 6103
rect 17693 6069 17727 6103
rect 17727 6069 17736 6103
rect 17684 6060 17736 6069
rect 17960 6103 18012 6112
rect 17960 6069 17969 6103
rect 17969 6069 18003 6103
rect 18003 6069 18012 6103
rect 17960 6060 18012 6069
rect 18880 6060 18932 6112
rect 19892 6239 19944 6248
rect 19892 6205 19901 6239
rect 19901 6205 19935 6239
rect 19935 6205 19944 6239
rect 19892 6196 19944 6205
rect 19984 6239 20036 6248
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 19984 6196 20036 6205
rect 20260 6264 20312 6316
rect 24032 6264 24084 6316
rect 20352 6196 20404 6248
rect 20720 6239 20772 6248
rect 20720 6205 20729 6239
rect 20729 6205 20763 6239
rect 20763 6205 20772 6239
rect 20720 6196 20772 6205
rect 22836 6196 22888 6248
rect 24492 6307 24544 6316
rect 24492 6273 24501 6307
rect 24501 6273 24535 6307
rect 24535 6273 24544 6307
rect 24492 6264 24544 6273
rect 25044 6264 25096 6316
rect 25964 6264 26016 6316
rect 26240 6264 26292 6316
rect 27252 6264 27304 6316
rect 27528 6264 27580 6316
rect 25596 6196 25648 6248
rect 26424 6196 26476 6248
rect 26792 6196 26844 6248
rect 30564 6196 30616 6248
rect 20996 6060 21048 6112
rect 21456 6060 21508 6112
rect 22560 6103 22612 6112
rect 22560 6069 22569 6103
rect 22569 6069 22603 6103
rect 22603 6069 22612 6103
rect 22560 6060 22612 6069
rect 22744 6060 22796 6112
rect 23756 6060 23808 6112
rect 24492 6060 24544 6112
rect 24768 6060 24820 6112
rect 24860 6060 24912 6112
rect 26332 6060 26384 6112
rect 27896 6060 27948 6112
rect 28632 6060 28684 6112
rect 7988 5958 8040 6010
rect 8052 5958 8104 6010
rect 8116 5958 8168 6010
rect 8180 5958 8232 6010
rect 8244 5958 8296 6010
rect 15578 5958 15630 6010
rect 15642 5958 15694 6010
rect 15706 5958 15758 6010
rect 15770 5958 15822 6010
rect 15834 5958 15886 6010
rect 23168 5958 23220 6010
rect 23232 5958 23284 6010
rect 23296 5958 23348 6010
rect 23360 5958 23412 6010
rect 23424 5958 23476 6010
rect 30758 5958 30810 6010
rect 30822 5958 30874 6010
rect 30886 5958 30938 6010
rect 30950 5958 31002 6010
rect 31014 5958 31066 6010
rect 1860 5856 1912 5908
rect 3516 5856 3568 5908
rect 5080 5856 5132 5908
rect 5172 5856 5224 5908
rect 6276 5856 6328 5908
rect 6368 5899 6420 5908
rect 6368 5865 6377 5899
rect 6377 5865 6411 5899
rect 6411 5865 6420 5899
rect 6368 5856 6420 5865
rect 6460 5856 6512 5908
rect 7380 5856 7432 5908
rect 8484 5856 8536 5908
rect 10140 5856 10192 5908
rect 940 5652 992 5704
rect 1584 5720 1636 5772
rect 6092 5788 6144 5840
rect 1308 5695 1360 5704
rect 1308 5661 1317 5695
rect 1317 5661 1351 5695
rect 1351 5661 1360 5695
rect 1308 5652 1360 5661
rect 3884 5720 3936 5772
rect 3976 5763 4028 5772
rect 3976 5729 3985 5763
rect 3985 5729 4019 5763
rect 4019 5729 4028 5763
rect 3976 5720 4028 5729
rect 4160 5720 4212 5772
rect 4896 5763 4948 5772
rect 4896 5729 4905 5763
rect 4905 5729 4939 5763
rect 4939 5729 4948 5763
rect 4896 5720 4948 5729
rect 5540 5720 5592 5772
rect 2872 5584 2924 5636
rect 4712 5627 4764 5636
rect 4712 5593 4721 5627
rect 4721 5593 4755 5627
rect 4755 5593 4764 5627
rect 4712 5584 4764 5593
rect 6460 5720 6512 5772
rect 7012 5720 7064 5772
rect 7288 5720 7340 5772
rect 7564 5720 7616 5772
rect 7656 5763 7708 5772
rect 7656 5729 7665 5763
rect 7665 5729 7699 5763
rect 7699 5729 7708 5763
rect 7656 5720 7708 5729
rect 7932 5720 7984 5772
rect 8852 5720 8904 5772
rect 12440 5856 12492 5908
rect 13636 5856 13688 5908
rect 10600 5788 10652 5840
rect 11060 5788 11112 5840
rect 11152 5788 11204 5840
rect 16028 5856 16080 5908
rect 16488 5856 16540 5908
rect 16580 5899 16632 5908
rect 16580 5865 16595 5899
rect 16595 5865 16629 5899
rect 16629 5865 16632 5899
rect 16580 5856 16632 5865
rect 17132 5856 17184 5908
rect 17960 5856 18012 5908
rect 19064 5856 19116 5908
rect 6736 5652 6788 5704
rect 6920 5652 6972 5704
rect 8024 5652 8076 5704
rect 8392 5652 8444 5704
rect 8576 5695 8628 5704
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 10048 5652 10100 5704
rect 11428 5720 11480 5772
rect 11060 5652 11112 5704
rect 11796 5652 11848 5704
rect 12624 5720 12676 5772
rect 12440 5652 12492 5704
rect 13820 5695 13872 5704
rect 13820 5661 13829 5695
rect 13829 5661 13863 5695
rect 13863 5661 13872 5695
rect 13820 5652 13872 5661
rect 14188 5695 14240 5704
rect 14188 5661 14190 5695
rect 14190 5661 14240 5695
rect 14188 5652 14240 5661
rect 14372 5720 14424 5772
rect 16948 5720 17000 5772
rect 20352 5899 20404 5908
rect 20352 5865 20361 5899
rect 20361 5865 20395 5899
rect 20395 5865 20404 5899
rect 20352 5856 20404 5865
rect 20720 5856 20772 5908
rect 22928 5856 22980 5908
rect 23388 5856 23440 5908
rect 19524 5720 19576 5772
rect 20904 5720 20956 5772
rect 21456 5763 21508 5772
rect 21456 5729 21465 5763
rect 21465 5729 21499 5763
rect 21499 5729 21508 5763
rect 21456 5720 21508 5729
rect 21824 5763 21876 5772
rect 21824 5729 21833 5763
rect 21833 5729 21867 5763
rect 21867 5729 21876 5763
rect 21824 5720 21876 5729
rect 25596 5788 25648 5840
rect 16028 5652 16080 5704
rect 16672 5652 16724 5704
rect 18512 5652 18564 5704
rect 18696 5695 18748 5704
rect 18696 5661 18698 5695
rect 18698 5661 18748 5695
rect 18696 5652 18748 5661
rect 18788 5695 18840 5704
rect 18788 5661 18800 5695
rect 18800 5661 18834 5695
rect 18834 5661 18840 5695
rect 18788 5652 18840 5661
rect 20444 5652 20496 5704
rect 21916 5695 21968 5704
rect 21916 5661 21925 5695
rect 21925 5661 21959 5695
rect 21959 5661 21968 5695
rect 21916 5652 21968 5661
rect 22376 5695 22428 5704
rect 22376 5661 22388 5695
rect 22388 5661 22422 5695
rect 22422 5661 22428 5695
rect 22376 5652 22428 5661
rect 22560 5720 22612 5772
rect 23572 5652 23624 5704
rect 3332 5559 3384 5568
rect 3332 5525 3341 5559
rect 3341 5525 3375 5559
rect 3375 5525 3384 5559
rect 3332 5516 3384 5525
rect 3884 5516 3936 5568
rect 3976 5516 4028 5568
rect 6460 5584 6512 5636
rect 9404 5584 9456 5636
rect 10968 5584 11020 5636
rect 11244 5584 11296 5636
rect 11520 5627 11572 5636
rect 11520 5593 11529 5627
rect 11529 5593 11563 5627
rect 11563 5593 11572 5627
rect 11520 5584 11572 5593
rect 21456 5584 21508 5636
rect 24400 5720 24452 5772
rect 24768 5720 24820 5772
rect 26424 5720 26476 5772
rect 26792 5720 26844 5772
rect 27252 5720 27304 5772
rect 27620 5856 27672 5908
rect 24676 5652 24728 5704
rect 25872 5652 25924 5704
rect 27528 5695 27580 5704
rect 27528 5661 27537 5695
rect 27537 5661 27571 5695
rect 27571 5661 27580 5695
rect 27528 5652 27580 5661
rect 27896 5695 27948 5704
rect 27896 5661 27898 5695
rect 27898 5661 27948 5695
rect 27896 5652 27948 5661
rect 28540 5720 28592 5772
rect 24124 5584 24176 5636
rect 5172 5559 5224 5568
rect 5172 5525 5181 5559
rect 5181 5525 5215 5559
rect 5215 5525 5224 5559
rect 5172 5516 5224 5525
rect 6644 5559 6696 5568
rect 6644 5525 6653 5559
rect 6653 5525 6687 5559
rect 6687 5525 6696 5559
rect 6644 5516 6696 5525
rect 6920 5559 6972 5568
rect 6920 5525 6929 5559
rect 6929 5525 6963 5559
rect 6963 5525 6972 5559
rect 6920 5516 6972 5525
rect 7380 5516 7432 5568
rect 7840 5516 7892 5568
rect 9588 5516 9640 5568
rect 9772 5516 9824 5568
rect 10508 5516 10560 5568
rect 11336 5516 11388 5568
rect 16396 5516 16448 5568
rect 18144 5559 18196 5568
rect 18144 5525 18153 5559
rect 18153 5525 18187 5559
rect 18187 5525 18196 5559
rect 18144 5516 18196 5525
rect 18236 5516 18288 5568
rect 19248 5516 19300 5568
rect 19984 5516 20036 5568
rect 20720 5516 20772 5568
rect 20812 5559 20864 5568
rect 20812 5525 20821 5559
rect 20821 5525 20855 5559
rect 20855 5525 20864 5559
rect 20812 5516 20864 5525
rect 22560 5516 22612 5568
rect 22744 5516 22796 5568
rect 26240 5584 26292 5636
rect 26792 5584 26844 5636
rect 26148 5559 26200 5568
rect 26148 5525 26157 5559
rect 26157 5525 26191 5559
rect 26191 5525 26200 5559
rect 26148 5516 26200 5525
rect 26608 5516 26660 5568
rect 26884 5516 26936 5568
rect 28172 5516 28224 5568
rect 4193 5414 4245 5466
rect 4257 5414 4309 5466
rect 4321 5414 4373 5466
rect 4385 5414 4437 5466
rect 4449 5414 4501 5466
rect 11783 5414 11835 5466
rect 11847 5414 11899 5466
rect 11911 5414 11963 5466
rect 11975 5414 12027 5466
rect 12039 5414 12091 5466
rect 19373 5414 19425 5466
rect 19437 5414 19489 5466
rect 19501 5414 19553 5466
rect 19565 5414 19617 5466
rect 19629 5414 19681 5466
rect 26963 5414 27015 5466
rect 27027 5414 27079 5466
rect 27091 5414 27143 5466
rect 27155 5414 27207 5466
rect 27219 5414 27271 5466
rect 940 5312 992 5364
rect 2504 5312 2556 5364
rect 1308 5176 1360 5228
rect 2596 5176 2648 5228
rect 2320 5108 2372 5160
rect 4988 5312 5040 5364
rect 2872 5176 2924 5228
rect 3240 5176 3292 5228
rect 6552 5312 6604 5364
rect 6828 5312 6880 5364
rect 7012 5312 7064 5364
rect 8760 5312 8812 5364
rect 9220 5312 9272 5364
rect 11152 5312 11204 5364
rect 16672 5312 16724 5364
rect 16948 5312 17000 5364
rect 21364 5312 21416 5364
rect 21548 5312 21600 5364
rect 24676 5312 24728 5364
rect 24768 5312 24820 5364
rect 6276 5176 6328 5228
rect 6736 5176 6788 5228
rect 7472 5176 7524 5228
rect 7932 5176 7984 5228
rect 8484 5176 8536 5228
rect 4528 5108 4580 5160
rect 9772 5219 9824 5228
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 12164 5176 12216 5228
rect 14188 5176 14240 5228
rect 14556 5176 14608 5228
rect 16120 5176 16172 5228
rect 17408 5176 17460 5228
rect 18144 5176 18196 5228
rect 1584 4972 1636 5024
rect 1768 4972 1820 5024
rect 3976 5015 4028 5024
rect 3976 4981 3991 5015
rect 3991 4981 4025 5015
rect 4025 4981 4028 5015
rect 3976 4972 4028 4981
rect 5448 4972 5500 5024
rect 6920 4972 6972 5024
rect 8024 5040 8076 5092
rect 7840 4972 7892 5024
rect 8760 5040 8812 5092
rect 9588 5108 9640 5160
rect 11060 5108 11112 5160
rect 13452 5108 13504 5160
rect 13728 5108 13780 5160
rect 15844 5151 15896 5160
rect 15844 5117 15853 5151
rect 15853 5117 15887 5151
rect 15887 5117 15896 5151
rect 15844 5108 15896 5117
rect 17316 5108 17368 5160
rect 18236 5108 18288 5160
rect 18512 5108 18564 5160
rect 18972 5108 19024 5160
rect 19708 5108 19760 5160
rect 17960 5083 18012 5092
rect 17960 5049 17969 5083
rect 17969 5049 18003 5083
rect 18003 5049 18012 5083
rect 17960 5040 18012 5049
rect 8852 4972 8904 5024
rect 9036 4972 9088 5024
rect 11704 5015 11756 5024
rect 11704 4981 11719 5015
rect 11719 4981 11753 5015
rect 11753 4981 11756 5015
rect 11704 4972 11756 4981
rect 16580 4972 16632 5024
rect 18696 4972 18748 5024
rect 18972 4972 19024 5024
rect 20720 5176 20772 5228
rect 21456 5176 21508 5228
rect 23756 5176 23808 5228
rect 20996 5108 21048 5160
rect 21916 5108 21968 5160
rect 24032 5176 24084 5228
rect 24676 5176 24728 5228
rect 28448 5244 28500 5296
rect 29184 5244 29236 5296
rect 26332 5176 26384 5228
rect 29000 5176 29052 5228
rect 26240 5151 26292 5160
rect 26240 5117 26249 5151
rect 26249 5117 26283 5151
rect 26283 5117 26292 5151
rect 26240 5108 26292 5117
rect 26424 5108 26476 5160
rect 23664 5040 23716 5092
rect 23756 5040 23808 5092
rect 23940 5040 23992 5092
rect 26516 5040 26568 5092
rect 22468 4972 22520 5024
rect 22928 4972 22980 5024
rect 24952 4972 25004 5024
rect 27896 4972 27948 5024
rect 29000 5015 29052 5024
rect 29000 4981 29009 5015
rect 29009 4981 29043 5015
rect 29043 4981 29052 5015
rect 29000 4972 29052 4981
rect 7988 4870 8040 4922
rect 8052 4870 8104 4922
rect 8116 4870 8168 4922
rect 8180 4870 8232 4922
rect 8244 4870 8296 4922
rect 15578 4870 15630 4922
rect 15642 4870 15694 4922
rect 15706 4870 15758 4922
rect 15770 4870 15822 4922
rect 15834 4870 15886 4922
rect 23168 4870 23220 4922
rect 23232 4870 23284 4922
rect 23296 4870 23348 4922
rect 23360 4870 23412 4922
rect 23424 4870 23476 4922
rect 30758 4870 30810 4922
rect 30822 4870 30874 4922
rect 30886 4870 30938 4922
rect 30950 4870 31002 4922
rect 31014 4870 31066 4922
rect 848 4768 900 4820
rect 2872 4768 2924 4820
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 6276 4768 6328 4820
rect 6920 4811 6972 4820
rect 6920 4777 6935 4811
rect 6935 4777 6969 4811
rect 6969 4777 6972 4811
rect 6920 4768 6972 4777
rect 7840 4768 7892 4820
rect 8484 4768 8536 4820
rect 9220 4768 9272 4820
rect 11428 4768 11480 4820
rect 11704 4768 11756 4820
rect 14188 4768 14240 4820
rect 16580 4811 16632 4820
rect 16580 4777 16595 4811
rect 16595 4777 16629 4811
rect 16629 4777 16632 4811
rect 16580 4768 16632 4777
rect 17960 4768 18012 4820
rect 18696 4768 18748 4820
rect 18972 4768 19024 4820
rect 1308 4675 1360 4684
rect 1308 4641 1317 4675
rect 1317 4641 1351 4675
rect 1351 4641 1360 4675
rect 1308 4632 1360 4641
rect 1584 4632 1636 4684
rect 2780 4632 2832 4684
rect 3608 4632 3660 4684
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 16120 4700 16172 4752
rect 4896 4564 4948 4616
rect 5264 4564 5316 4616
rect 6000 4607 6052 4616
rect 3516 4496 3568 4548
rect 6000 4573 6009 4607
rect 6009 4573 6043 4607
rect 6043 4573 6052 4607
rect 6000 4564 6052 4573
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 6460 4564 6512 4573
rect 7104 4564 7156 4616
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 8852 4564 8904 4616
rect 9036 4607 9088 4616
rect 9036 4573 9038 4607
rect 9038 4573 9088 4607
rect 9036 4564 9088 4573
rect 9404 4675 9456 4684
rect 9404 4641 9413 4675
rect 9413 4641 9447 4675
rect 9447 4641 9456 4675
rect 9404 4632 9456 4641
rect 5816 4428 5868 4480
rect 7288 4428 7340 4480
rect 11060 4428 11112 4480
rect 12164 4564 12216 4616
rect 12348 4675 12400 4684
rect 12348 4641 12357 4675
rect 12357 4641 12391 4675
rect 12391 4641 12400 4675
rect 12348 4632 12400 4641
rect 12532 4564 12584 4616
rect 13820 4607 13872 4616
rect 13820 4573 13829 4607
rect 13829 4573 13863 4607
rect 13863 4573 13872 4607
rect 13820 4564 13872 4573
rect 14464 4632 14516 4684
rect 17684 4632 17736 4684
rect 16120 4607 16172 4616
rect 16120 4573 16129 4607
rect 16129 4573 16163 4607
rect 16163 4573 16172 4607
rect 16120 4564 16172 4573
rect 16396 4564 16448 4616
rect 18512 4564 18564 4616
rect 18880 4632 18932 4684
rect 13452 4428 13504 4480
rect 17868 4428 17920 4480
rect 27896 4768 27948 4820
rect 28356 4768 28408 4820
rect 20536 4700 20588 4752
rect 21640 4700 21692 4752
rect 26700 4700 26752 4752
rect 19800 4632 19852 4684
rect 20904 4632 20956 4684
rect 21272 4675 21324 4684
rect 21272 4641 21281 4675
rect 21281 4641 21315 4675
rect 21315 4641 21324 4675
rect 21272 4632 21324 4641
rect 21456 4632 21508 4684
rect 21916 4632 21968 4684
rect 22468 4632 22520 4684
rect 22560 4675 22612 4684
rect 22560 4641 22569 4675
rect 22569 4641 22603 4675
rect 22603 4641 22612 4675
rect 22560 4632 22612 4641
rect 22008 4564 22060 4616
rect 22192 4607 22244 4616
rect 22192 4573 22194 4607
rect 22194 4573 22244 4607
rect 22192 4564 22244 4573
rect 24032 4607 24084 4616
rect 24032 4573 24041 4607
rect 24041 4573 24075 4607
rect 24075 4573 24084 4607
rect 24032 4564 24084 4573
rect 24400 4607 24452 4616
rect 24400 4573 24402 4607
rect 24402 4573 24452 4607
rect 24400 4564 24452 4573
rect 24584 4632 24636 4684
rect 24860 4632 24912 4684
rect 25412 4564 25464 4616
rect 27528 4675 27580 4684
rect 27528 4641 27537 4675
rect 27537 4641 27571 4675
rect 27571 4641 27580 4675
rect 27528 4632 27580 4641
rect 27896 4632 27948 4684
rect 19800 4496 19852 4548
rect 20352 4471 20404 4480
rect 20352 4437 20361 4471
rect 20361 4437 20395 4471
rect 20395 4437 20404 4471
rect 20352 4428 20404 4437
rect 21272 4428 21324 4480
rect 21364 4428 21416 4480
rect 21824 4428 21876 4480
rect 22284 4428 22336 4480
rect 26056 4471 26108 4480
rect 26056 4437 26065 4471
rect 26065 4437 26099 4471
rect 26099 4437 26108 4471
rect 26056 4428 26108 4437
rect 27436 4564 27488 4616
rect 27804 4564 27856 4616
rect 29000 4632 29052 4684
rect 28264 4607 28316 4616
rect 28264 4573 28273 4607
rect 28273 4573 28307 4607
rect 28307 4573 28316 4607
rect 28264 4564 28316 4573
rect 4193 4326 4245 4378
rect 4257 4326 4309 4378
rect 4321 4326 4373 4378
rect 4385 4326 4437 4378
rect 4449 4326 4501 4378
rect 11783 4326 11835 4378
rect 11847 4326 11899 4378
rect 11911 4326 11963 4378
rect 11975 4326 12027 4378
rect 12039 4326 12091 4378
rect 19373 4326 19425 4378
rect 19437 4326 19489 4378
rect 19501 4326 19553 4378
rect 19565 4326 19617 4378
rect 19629 4326 19681 4378
rect 26963 4326 27015 4378
rect 27027 4326 27079 4378
rect 27091 4326 27143 4378
rect 27155 4326 27207 4378
rect 27219 4326 27271 4378
rect 1308 4088 1360 4140
rect 1492 4088 1544 4140
rect 2688 4088 2740 4140
rect 1032 4020 1084 4072
rect 5632 4224 5684 4276
rect 5356 4156 5408 4208
rect 6828 4224 6880 4276
rect 8760 4224 8812 4276
rect 9404 4156 9456 4208
rect 12164 4224 12216 4276
rect 12532 4267 12584 4276
rect 12532 4233 12541 4267
rect 12541 4233 12575 4267
rect 12575 4233 12584 4267
rect 12532 4224 12584 4233
rect 14556 4224 14608 4276
rect 17500 4224 17552 4276
rect 18512 4224 18564 4276
rect 21548 4224 21600 4276
rect 21640 4224 21692 4276
rect 23572 4224 23624 4276
rect 22192 4156 22244 4208
rect 3240 4088 3292 4140
rect 3332 4088 3384 4140
rect 4988 4088 5040 4140
rect 5540 4088 5592 4140
rect 8392 4088 8444 4140
rect 8852 4088 8904 4140
rect 3424 4063 3476 4072
rect 3424 4029 3433 4063
rect 3433 4029 3467 4063
rect 3467 4029 3476 4063
rect 3424 4020 3476 4029
rect 1768 3884 1820 3936
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 2780 3884 2832 3893
rect 5816 4020 5868 4072
rect 7656 4020 7708 4072
rect 8484 3952 8536 4004
rect 9036 4020 9088 4072
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 9404 4020 9456 4072
rect 10048 4088 10100 4140
rect 10508 4088 10560 4140
rect 11244 4088 11296 4140
rect 14004 4088 14056 4140
rect 14188 4131 14240 4140
rect 14188 4097 14190 4131
rect 14190 4097 14240 4131
rect 14188 4088 14240 4097
rect 3976 3927 4028 3936
rect 3976 3893 3991 3927
rect 3991 3893 4025 3927
rect 4025 3893 4028 3927
rect 3976 3884 4028 3893
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 6000 3884 6052 3936
rect 8576 3884 8628 3936
rect 9312 3884 9364 3936
rect 9680 3884 9732 3936
rect 9864 3884 9916 3936
rect 13452 3952 13504 4004
rect 13636 4020 13688 4072
rect 13820 4063 13872 4072
rect 13820 4029 13829 4063
rect 13829 4029 13863 4063
rect 13863 4029 13872 4063
rect 13820 4020 13872 4029
rect 14464 4088 14516 4140
rect 14372 4020 14424 4072
rect 14648 4020 14700 4072
rect 16212 4020 16264 4072
rect 16396 4063 16448 4072
rect 16396 4029 16405 4063
rect 16405 4029 16439 4063
rect 16439 4029 16448 4063
rect 16396 4020 16448 4029
rect 16948 4088 17000 4140
rect 17868 4088 17920 4140
rect 19616 4020 19668 4072
rect 20352 4131 20404 4140
rect 20352 4097 20364 4131
rect 20364 4097 20398 4131
rect 20398 4097 20404 4131
rect 20352 4088 20404 4097
rect 20812 4088 20864 4140
rect 22376 4088 22428 4140
rect 22836 4156 22888 4208
rect 19800 4063 19852 4072
rect 19800 4029 19801 4063
rect 19801 4029 19835 4063
rect 19835 4029 19852 4063
rect 19800 4020 19852 4029
rect 12072 3927 12124 3936
rect 12072 3893 12081 3927
rect 12081 3893 12115 3927
rect 12115 3893 12124 3927
rect 12072 3884 12124 3893
rect 13544 3927 13596 3936
rect 13544 3893 13553 3927
rect 13553 3893 13587 3927
rect 13587 3893 13596 3927
rect 13544 3884 13596 3893
rect 13912 3952 13964 4004
rect 19984 4020 20036 4072
rect 22652 4020 22704 4072
rect 22928 4020 22980 4072
rect 24216 4224 24268 4276
rect 24676 4088 24728 4140
rect 24768 4131 24820 4140
rect 24768 4097 24777 4131
rect 24777 4097 24811 4131
rect 24811 4097 24820 4131
rect 24768 4088 24820 4097
rect 26056 4088 26108 4140
rect 26792 4088 26844 4140
rect 25228 4020 25280 4072
rect 26240 4063 26292 4072
rect 14280 3884 14332 3936
rect 16028 3884 16080 3936
rect 16672 3884 16724 3936
rect 17040 3884 17092 3936
rect 17224 3884 17276 3936
rect 19340 3927 19392 3936
rect 19340 3893 19349 3927
rect 19349 3893 19383 3927
rect 19383 3893 19392 3927
rect 19340 3884 19392 3893
rect 19708 3884 19760 3936
rect 20996 3884 21048 3936
rect 22836 3927 22888 3936
rect 22836 3893 22845 3927
rect 22845 3893 22879 3927
rect 22879 3893 22888 3927
rect 22836 3884 22888 3893
rect 24032 3884 24084 3936
rect 24400 3884 24452 3936
rect 24492 3927 24544 3936
rect 24492 3893 24507 3927
rect 24507 3893 24541 3927
rect 24541 3893 24544 3927
rect 24492 3884 24544 3893
rect 25136 3884 25188 3936
rect 26240 4029 26249 4063
rect 26249 4029 26283 4063
rect 26283 4029 26292 4063
rect 26240 4020 26292 4029
rect 26056 3927 26108 3936
rect 26056 3893 26065 3927
rect 26065 3893 26099 3927
rect 26099 3893 26108 3927
rect 26056 3884 26108 3893
rect 26700 3927 26752 3936
rect 26700 3893 26715 3927
rect 26715 3893 26749 3927
rect 26749 3893 26752 3927
rect 26700 3884 26752 3893
rect 28080 3927 28132 3936
rect 28080 3893 28089 3927
rect 28089 3893 28123 3927
rect 28123 3893 28132 3927
rect 28080 3884 28132 3893
rect 7988 3782 8040 3834
rect 8052 3782 8104 3834
rect 8116 3782 8168 3834
rect 8180 3782 8232 3834
rect 8244 3782 8296 3834
rect 15578 3782 15630 3834
rect 15642 3782 15694 3834
rect 15706 3782 15758 3834
rect 15770 3782 15822 3834
rect 15834 3782 15886 3834
rect 23168 3782 23220 3834
rect 23232 3782 23284 3834
rect 23296 3782 23348 3834
rect 23360 3782 23412 3834
rect 23424 3782 23476 3834
rect 30758 3782 30810 3834
rect 30822 3782 30874 3834
rect 30886 3782 30938 3834
rect 30950 3782 31002 3834
rect 31014 3782 31066 3834
rect 756 3680 808 3732
rect 1124 3612 1176 3664
rect 4528 3680 4580 3732
rect 5540 3680 5592 3732
rect 6552 3680 6604 3732
rect 7104 3680 7156 3732
rect 9220 3680 9272 3732
rect 10508 3680 10560 3732
rect 10968 3680 11020 3732
rect 12072 3680 12124 3732
rect 1216 3587 1268 3596
rect 1216 3553 1225 3587
rect 1225 3553 1259 3587
rect 1259 3553 1268 3587
rect 1216 3544 1268 3553
rect 3240 3612 3292 3664
rect 3608 3612 3660 3664
rect 6000 3612 6052 3664
rect 940 3476 992 3528
rect 1676 3408 1728 3460
rect 3976 3519 4028 3528
rect 3976 3485 3988 3519
rect 3988 3485 4022 3519
rect 4022 3485 4028 3519
rect 3976 3476 4028 3485
rect 4252 3587 4304 3596
rect 4252 3553 4261 3587
rect 4261 3553 4295 3587
rect 4295 3553 4304 3587
rect 4252 3544 4304 3553
rect 6184 3544 6236 3596
rect 6552 3544 6604 3596
rect 6644 3587 6696 3596
rect 6644 3553 6653 3587
rect 6653 3553 6687 3587
rect 6687 3553 6696 3587
rect 6644 3544 6696 3553
rect 7104 3544 7156 3596
rect 7288 3544 7340 3596
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 9312 3544 9364 3596
rect 9496 3544 9548 3596
rect 14188 3680 14240 3732
rect 16212 3680 16264 3732
rect 16488 3680 16540 3732
rect 16580 3723 16632 3732
rect 16580 3689 16595 3723
rect 16595 3689 16629 3723
rect 16629 3689 16632 3723
rect 16580 3680 16632 3689
rect 18972 3680 19024 3732
rect 20996 3680 21048 3732
rect 21548 3680 21600 3732
rect 22836 3680 22888 3732
rect 22928 3680 22980 3732
rect 24124 3680 24176 3732
rect 24584 3680 24636 3732
rect 26516 3680 26568 3732
rect 13912 3612 13964 3664
rect 5448 3340 5500 3392
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 5632 3476 5684 3485
rect 5816 3476 5868 3528
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 8852 3476 8904 3528
rect 9036 3519 9088 3528
rect 9036 3485 9038 3519
rect 9038 3485 9088 3519
rect 9036 3476 9088 3485
rect 9772 3476 9824 3528
rect 11520 3476 11572 3528
rect 11060 3408 11112 3460
rect 11796 3476 11848 3528
rect 12348 3519 12400 3528
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 13544 3476 13596 3528
rect 13820 3519 13872 3528
rect 13820 3485 13829 3519
rect 13829 3485 13863 3519
rect 13863 3485 13872 3519
rect 13820 3476 13872 3485
rect 14280 3519 14332 3528
rect 14280 3485 14292 3519
rect 14292 3485 14326 3519
rect 14326 3485 14332 3519
rect 14280 3476 14332 3485
rect 16120 3519 16172 3528
rect 16120 3485 16129 3519
rect 16129 3485 16163 3519
rect 16163 3485 16172 3519
rect 16120 3476 16172 3485
rect 16672 3544 16724 3596
rect 18512 3476 18564 3528
rect 19340 3544 19392 3596
rect 19248 3476 19300 3528
rect 20996 3544 21048 3596
rect 21824 3544 21876 3596
rect 24492 3544 24544 3596
rect 25504 3544 25556 3596
rect 26700 3680 26752 3732
rect 27620 3655 27672 3664
rect 27620 3621 27629 3655
rect 27629 3621 27663 3655
rect 27663 3621 27672 3655
rect 27620 3612 27672 3621
rect 27804 3612 27856 3664
rect 9220 3340 9272 3392
rect 19984 3408 20036 3460
rect 20904 3408 20956 3460
rect 23756 3476 23808 3528
rect 23848 3476 23900 3528
rect 27896 3587 27948 3596
rect 27896 3553 27905 3587
rect 27905 3553 27939 3587
rect 27939 3553 27948 3587
rect 27896 3544 27948 3553
rect 28264 3519 28316 3528
rect 28264 3485 28266 3519
rect 28266 3485 28316 3519
rect 28264 3476 28316 3485
rect 28540 3476 28592 3528
rect 28816 3476 28868 3528
rect 25780 3408 25832 3460
rect 16396 3340 16448 3392
rect 16488 3340 16540 3392
rect 19524 3340 19576 3392
rect 23296 3383 23348 3392
rect 23296 3349 23305 3383
rect 23305 3349 23339 3383
rect 23339 3349 23348 3383
rect 23296 3340 23348 3349
rect 25320 3383 25372 3392
rect 25320 3349 25329 3383
rect 25329 3349 25363 3383
rect 25363 3349 25372 3383
rect 25320 3340 25372 3349
rect 26424 3383 26476 3392
rect 26424 3349 26433 3383
rect 26433 3349 26467 3383
rect 26467 3349 26476 3383
rect 26424 3340 26476 3349
rect 4193 3238 4245 3290
rect 4257 3238 4309 3290
rect 4321 3238 4373 3290
rect 4385 3238 4437 3290
rect 4449 3238 4501 3290
rect 11783 3238 11835 3290
rect 11847 3238 11899 3290
rect 11911 3238 11963 3290
rect 11975 3238 12027 3290
rect 12039 3238 12091 3290
rect 19373 3238 19425 3290
rect 19437 3238 19489 3290
rect 19501 3238 19553 3290
rect 19565 3238 19617 3290
rect 19629 3238 19681 3290
rect 26963 3238 27015 3290
rect 27027 3238 27079 3290
rect 27091 3238 27143 3290
rect 27155 3238 27207 3290
rect 27219 3238 27271 3290
rect 5264 3136 5316 3188
rect 5448 3068 5500 3120
rect 7288 3136 7340 3188
rect 8116 3136 8168 3188
rect 9864 3136 9916 3188
rect 10968 3136 11020 3188
rect 8852 3068 8904 3120
rect 1308 3000 1360 3052
rect 2964 3000 3016 3052
rect 4068 3000 4120 3052
rect 4620 3000 4672 3052
rect 6000 3000 6052 3052
rect 1676 2975 1728 2984
rect 1676 2941 1685 2975
rect 1685 2941 1719 2975
rect 1719 2941 1728 2975
rect 1676 2932 1728 2941
rect 3240 2932 3292 2984
rect 3516 2932 3568 2984
rect 5172 2932 5224 2984
rect 7748 3000 7800 3052
rect 8576 3000 8628 3052
rect 1768 2796 1820 2848
rect 4160 2839 4212 2848
rect 4160 2805 4175 2839
rect 4175 2805 4209 2839
rect 4209 2805 4212 2839
rect 4160 2796 4212 2805
rect 4528 2796 4580 2848
rect 5540 2796 5592 2848
rect 5724 2796 5776 2848
rect 6920 2796 6972 2848
rect 8852 2864 8904 2916
rect 9680 3000 9732 3052
rect 14280 3136 14332 3188
rect 16948 3136 17000 3188
rect 25964 3136 26016 3188
rect 23848 3068 23900 3120
rect 25504 3068 25556 3120
rect 25872 3068 25924 3120
rect 30012 3136 30064 3188
rect 11060 2932 11112 2984
rect 11336 2932 11388 2984
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 15108 3000 15160 3052
rect 16028 3000 16080 3052
rect 16396 3000 16448 3052
rect 23296 3000 23348 3052
rect 24400 3000 24452 3052
rect 14280 2932 14332 2984
rect 14372 2975 14424 2984
rect 14372 2941 14381 2975
rect 14381 2941 14415 2975
rect 14415 2941 14424 2975
rect 14372 2932 14424 2941
rect 16120 2932 16172 2984
rect 9312 2796 9364 2848
rect 9404 2796 9456 2848
rect 11704 2839 11756 2848
rect 11704 2805 11719 2839
rect 11719 2805 11753 2839
rect 11753 2805 11756 2839
rect 11704 2796 11756 2805
rect 13912 2796 13964 2848
rect 15016 2796 15068 2848
rect 15200 2796 15252 2848
rect 16580 2796 16632 2848
rect 18512 2932 18564 2984
rect 19708 2932 19760 2984
rect 20904 2975 20956 2984
rect 20904 2941 20913 2975
rect 20913 2941 20947 2975
rect 20947 2941 20956 2975
rect 20904 2932 20956 2941
rect 21272 2932 21324 2984
rect 22652 2932 22704 2984
rect 23756 2932 23808 2984
rect 26148 3000 26200 3052
rect 27068 3000 27120 3052
rect 26240 2975 26292 2984
rect 26240 2941 26249 2975
rect 26249 2941 26283 2975
rect 26283 2941 26292 2975
rect 26240 2932 26292 2941
rect 26608 2932 26660 2984
rect 27436 2932 27488 2984
rect 18972 2796 19024 2848
rect 21548 2796 21600 2848
rect 23848 2796 23900 2848
rect 24124 2796 24176 2848
rect 24676 2796 24728 2848
rect 26700 2839 26752 2848
rect 26700 2805 26715 2839
rect 26715 2805 26749 2839
rect 26749 2805 26752 2839
rect 26700 2796 26752 2805
rect 27620 2796 27672 2848
rect 7988 2694 8040 2746
rect 8052 2694 8104 2746
rect 8116 2694 8168 2746
rect 8180 2694 8232 2746
rect 8244 2694 8296 2746
rect 15578 2694 15630 2746
rect 15642 2694 15694 2746
rect 15706 2694 15758 2746
rect 15770 2694 15822 2746
rect 15834 2694 15886 2746
rect 23168 2694 23220 2746
rect 23232 2694 23284 2746
rect 23296 2694 23348 2746
rect 23360 2694 23412 2746
rect 23424 2694 23476 2746
rect 30758 2694 30810 2746
rect 30822 2694 30874 2746
rect 30886 2694 30938 2746
rect 30950 2694 31002 2746
rect 31014 2694 31066 2746
rect 664 2592 716 2644
rect 1400 2592 1452 2644
rect 1952 2592 2004 2644
rect 2044 2592 2096 2644
rect 5724 2592 5776 2644
rect 5816 2592 5868 2644
rect 6920 2592 6972 2644
rect 7196 2592 7248 2644
rect 3056 2524 3108 2576
rect 1032 2456 1084 2508
rect 1952 2456 2004 2508
rect 5080 2456 5132 2508
rect 6092 2524 6144 2576
rect 8392 2592 8444 2644
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 10600 2635 10652 2644
rect 10600 2601 10609 2635
rect 10609 2601 10643 2635
rect 10643 2601 10652 2635
rect 10600 2592 10652 2601
rect 10876 2592 10928 2644
rect 11520 2524 11572 2576
rect 6000 2456 6052 2508
rect 1860 2388 1912 2440
rect 4528 2388 4580 2440
rect 6460 2456 6512 2508
rect 6828 2499 6880 2508
rect 6828 2465 6837 2499
rect 6837 2465 6871 2499
rect 6871 2465 6880 2499
rect 6828 2456 6880 2465
rect 7104 2456 7156 2508
rect 4988 2320 5040 2372
rect 3056 2252 3108 2304
rect 3240 2252 3292 2304
rect 4896 2252 4948 2304
rect 6000 2363 6052 2372
rect 6000 2329 6009 2363
rect 6009 2329 6043 2363
rect 6043 2329 6052 2363
rect 6000 2320 6052 2329
rect 7472 2388 7524 2440
rect 7840 2456 7892 2508
rect 8576 2456 8628 2508
rect 9496 2456 9548 2508
rect 10508 2499 10560 2508
rect 10508 2465 10517 2499
rect 10517 2465 10551 2499
rect 10551 2465 10560 2499
rect 10508 2456 10560 2465
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 8208 2431 8260 2440
rect 8208 2397 8220 2431
rect 8220 2397 8254 2431
rect 8254 2397 8260 2431
rect 8208 2388 8260 2397
rect 8300 2388 8352 2440
rect 9680 2388 9732 2440
rect 9772 2388 9824 2440
rect 11060 2499 11112 2508
rect 11060 2465 11069 2499
rect 11069 2465 11103 2499
rect 11103 2465 11112 2499
rect 14004 2592 14056 2644
rect 16580 2635 16632 2644
rect 16580 2601 16595 2635
rect 16595 2601 16629 2635
rect 16629 2601 16632 2635
rect 16580 2592 16632 2601
rect 18972 2592 19024 2644
rect 11060 2456 11112 2465
rect 6460 2320 6512 2372
rect 11704 2388 11756 2440
rect 12164 2388 12216 2440
rect 13728 2431 13780 2440
rect 13728 2397 13737 2431
rect 13737 2397 13771 2431
rect 13771 2397 13780 2431
rect 13728 2388 13780 2397
rect 14372 2456 14424 2508
rect 14464 2431 14516 2440
rect 14464 2397 14473 2431
rect 14473 2397 14507 2431
rect 14507 2397 14516 2431
rect 14464 2388 14516 2397
rect 10048 2320 10100 2372
rect 16120 2499 16172 2508
rect 16120 2465 16129 2499
rect 16129 2465 16163 2499
rect 16163 2465 16172 2499
rect 16120 2456 16172 2465
rect 16212 2456 16264 2508
rect 16028 2388 16080 2440
rect 8852 2252 8904 2304
rect 14188 2252 14240 2304
rect 15936 2252 15988 2304
rect 20536 2456 20588 2508
rect 20904 2592 20956 2644
rect 21548 2592 21600 2644
rect 23848 2524 23900 2576
rect 25964 2635 26016 2644
rect 25964 2601 25973 2635
rect 25973 2601 26007 2635
rect 26007 2601 26016 2635
rect 25964 2592 26016 2601
rect 21180 2456 21232 2508
rect 21364 2456 21416 2508
rect 18512 2388 18564 2440
rect 18788 2431 18840 2440
rect 18788 2397 18800 2431
rect 18800 2397 18834 2431
rect 18834 2397 18840 2431
rect 18788 2388 18840 2397
rect 19248 2388 19300 2440
rect 23664 2499 23716 2508
rect 23664 2465 23673 2499
rect 23673 2465 23707 2499
rect 23707 2465 23716 2499
rect 23664 2456 23716 2465
rect 23940 2499 23992 2508
rect 23940 2465 23949 2499
rect 23949 2465 23983 2499
rect 23983 2465 23992 2499
rect 23940 2456 23992 2465
rect 26240 2524 26292 2576
rect 27712 2592 27764 2644
rect 30012 2635 30064 2644
rect 30012 2601 30021 2635
rect 30021 2601 30055 2635
rect 30055 2601 30064 2635
rect 30012 2592 30064 2601
rect 24216 2456 24268 2508
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 24492 2431 24544 2440
rect 24492 2397 24494 2431
rect 24494 2397 24544 2431
rect 24492 2388 24544 2397
rect 25320 2456 25372 2508
rect 27344 2456 27396 2508
rect 27528 2456 27580 2508
rect 26424 2388 26476 2440
rect 22928 2320 22980 2372
rect 18788 2252 18840 2304
rect 20168 2252 20220 2304
rect 21456 2252 21508 2304
rect 22192 2252 22244 2304
rect 23848 2252 23900 2304
rect 27988 2456 28040 2508
rect 28264 2456 28316 2508
rect 28908 2499 28960 2508
rect 28908 2465 28917 2499
rect 28917 2465 28951 2499
rect 28951 2465 28960 2499
rect 28908 2456 28960 2465
rect 27896 2320 27948 2372
rect 29644 2252 29696 2304
rect 4193 2150 4245 2202
rect 4257 2150 4309 2202
rect 4321 2150 4373 2202
rect 4385 2150 4437 2202
rect 4449 2150 4501 2202
rect 11783 2150 11835 2202
rect 11847 2150 11899 2202
rect 11911 2150 11963 2202
rect 11975 2150 12027 2202
rect 12039 2150 12091 2202
rect 19373 2150 19425 2202
rect 19437 2150 19489 2202
rect 19501 2150 19553 2202
rect 19565 2150 19617 2202
rect 19629 2150 19681 2202
rect 26963 2150 27015 2202
rect 27027 2150 27079 2202
rect 27091 2150 27143 2202
rect 27155 2150 27207 2202
rect 27219 2150 27271 2202
rect 3332 2048 3384 2100
rect 5540 2091 5592 2100
rect 5540 2057 5549 2091
rect 5549 2057 5583 2091
rect 5583 2057 5592 2091
rect 5540 2048 5592 2057
rect 3240 2023 3292 2032
rect 3240 1989 3249 2023
rect 3249 1989 3283 2023
rect 3283 1989 3292 2023
rect 3240 1980 3292 1989
rect 5264 1980 5316 2032
rect 1492 1912 1544 1964
rect 1676 1955 1728 1964
rect 1676 1921 1685 1955
rect 1685 1921 1719 1955
rect 1719 1921 1728 1955
rect 1676 1912 1728 1921
rect 1308 1844 1360 1896
rect 3424 1887 3476 1896
rect 3424 1853 3433 1887
rect 3433 1853 3467 1887
rect 3467 1853 3476 1887
rect 3424 1844 3476 1853
rect 3976 1953 4028 1964
rect 3976 1919 3988 1953
rect 3988 1919 4022 1953
rect 4022 1919 4028 1953
rect 3976 1912 4028 1919
rect 6184 1955 6236 1964
rect 3608 1844 3660 1896
rect 6184 1921 6186 1955
rect 6186 1921 6236 1955
rect 6184 1912 6236 1921
rect 6368 1912 6420 1964
rect 7288 1912 7340 1964
rect 8208 2048 8260 2100
rect 10876 2048 10928 2100
rect 11152 2048 11204 2100
rect 12164 2048 12216 2100
rect 13176 2048 13228 2100
rect 16764 2048 16816 2100
rect 17960 2048 18012 2100
rect 5724 1844 5776 1896
rect 5816 1887 5868 1896
rect 5816 1853 5825 1887
rect 5825 1853 5859 1887
rect 5859 1853 5868 1887
rect 5816 1844 5868 1853
rect 5908 1844 5960 1896
rect 8300 1844 8352 1896
rect 8852 1912 8904 1964
rect 8668 1887 8720 1896
rect 8668 1853 8677 1887
rect 8677 1853 8711 1887
rect 8711 1853 8720 1887
rect 8668 1844 8720 1853
rect 9588 1912 9640 1964
rect 1676 1708 1728 1760
rect 10784 1844 10836 1896
rect 11060 1844 11112 1896
rect 11520 1844 11572 1896
rect 12348 1912 12400 1964
rect 14188 1912 14240 1964
rect 18328 1980 18380 2032
rect 20720 2048 20772 2100
rect 21088 2048 21140 2100
rect 22376 2048 22428 2100
rect 23480 2048 23532 2100
rect 28724 2091 28776 2100
rect 28724 2057 28733 2091
rect 28733 2057 28767 2091
rect 28767 2057 28776 2091
rect 28724 2048 28776 2057
rect 11888 1844 11940 1896
rect 13728 1844 13780 1896
rect 14004 1887 14056 1896
rect 14004 1853 14006 1887
rect 14006 1853 14056 1887
rect 14004 1844 14056 1853
rect 16120 1844 16172 1896
rect 18236 1887 18288 1896
rect 18236 1853 18245 1887
rect 18245 1853 18279 1887
rect 18279 1853 18288 1887
rect 18236 1844 18288 1853
rect 18604 1912 18656 1964
rect 18144 1776 18196 1828
rect 21456 1912 21508 1964
rect 23480 1912 23532 1964
rect 20444 1844 20496 1896
rect 21180 1844 21232 1896
rect 22652 1844 22704 1896
rect 23664 1980 23716 2032
rect 26056 1980 26108 2032
rect 23020 1819 23072 1828
rect 23020 1785 23029 1819
rect 23029 1785 23063 1819
rect 23063 1785 23072 1819
rect 23020 1776 23072 1785
rect 23756 1844 23808 1896
rect 26240 1912 26292 1964
rect 26976 1912 27028 1964
rect 26056 1844 26108 1896
rect 26424 1844 26476 1896
rect 29276 1912 29328 1964
rect 29552 1912 29604 1964
rect 8668 1708 8720 1760
rect 8760 1751 8812 1760
rect 8760 1717 8769 1751
rect 8769 1717 8803 1751
rect 8803 1717 8812 1751
rect 8760 1708 8812 1717
rect 8944 1708 8996 1760
rect 9404 1708 9456 1760
rect 10876 1708 10928 1760
rect 11704 1751 11756 1760
rect 11704 1717 11719 1751
rect 11719 1717 11753 1751
rect 11753 1717 11756 1751
rect 11704 1708 11756 1717
rect 11888 1708 11940 1760
rect 13636 1708 13688 1760
rect 16580 1708 16632 1760
rect 17960 1708 18012 1760
rect 18972 1708 19024 1760
rect 19340 1708 19392 1760
rect 20812 1708 20864 1760
rect 21548 1708 21600 1760
rect 22836 1708 22888 1760
rect 23572 1708 23624 1760
rect 23756 1708 23808 1760
rect 23940 1708 23992 1760
rect 24124 1708 24176 1760
rect 24860 1708 24912 1760
rect 26332 1708 26384 1760
rect 26608 1708 26660 1760
rect 26976 1708 27028 1760
rect 27528 1708 27580 1760
rect 27712 1708 27764 1760
rect 29184 1751 29236 1760
rect 29184 1717 29193 1751
rect 29193 1717 29227 1751
rect 29227 1717 29236 1751
rect 29184 1708 29236 1717
rect 7988 1606 8040 1658
rect 8052 1606 8104 1658
rect 8116 1606 8168 1658
rect 8180 1606 8232 1658
rect 8244 1606 8296 1658
rect 15578 1606 15630 1658
rect 15642 1606 15694 1658
rect 15706 1606 15758 1658
rect 15770 1606 15822 1658
rect 15834 1606 15886 1658
rect 23168 1606 23220 1658
rect 23232 1606 23284 1658
rect 23296 1606 23348 1658
rect 23360 1606 23412 1658
rect 23424 1606 23476 1658
rect 30758 1606 30810 1658
rect 30822 1606 30874 1658
rect 30886 1606 30938 1658
rect 30950 1606 31002 1658
rect 31014 1606 31066 1658
rect 1216 1504 1268 1556
rect 1768 1504 1820 1556
rect 3884 1504 3936 1556
rect 4528 1504 4580 1556
rect 6920 1547 6972 1556
rect 6920 1513 6935 1547
rect 6935 1513 6969 1547
rect 6969 1513 6972 1547
rect 6920 1504 6972 1513
rect 8944 1504 8996 1556
rect 10876 1504 10928 1556
rect 10968 1547 11020 1556
rect 10968 1513 10977 1547
rect 10977 1513 11011 1547
rect 11011 1513 11020 1547
rect 10968 1504 11020 1513
rect 11060 1504 11112 1556
rect 13820 1504 13872 1556
rect 14004 1504 14056 1556
rect 16028 1504 16080 1556
rect 16580 1547 16632 1556
rect 16580 1513 16595 1547
rect 16595 1513 16629 1547
rect 16629 1513 16632 1547
rect 16580 1504 16632 1513
rect 18144 1547 18196 1556
rect 18144 1513 18153 1547
rect 18153 1513 18187 1547
rect 18187 1513 18196 1547
rect 18144 1504 18196 1513
rect 18972 1504 19024 1556
rect 10508 1436 10560 1488
rect 1308 1343 1360 1352
rect 1308 1309 1317 1343
rect 1317 1309 1351 1343
rect 1351 1309 1360 1343
rect 1308 1300 1360 1309
rect 1676 1343 1728 1352
rect 1676 1309 1678 1343
rect 1678 1309 1728 1343
rect 1676 1300 1728 1309
rect 2044 1343 2096 1352
rect 2044 1309 2053 1343
rect 2053 1309 2087 1343
rect 2087 1309 2096 1343
rect 2044 1300 2096 1309
rect 2504 1164 2556 1216
rect 3516 1343 3568 1352
rect 3516 1309 3525 1343
rect 3525 1309 3559 1343
rect 3559 1309 3568 1343
rect 3516 1300 3568 1309
rect 3976 1345 4028 1352
rect 3976 1311 4021 1345
rect 4021 1311 4028 1345
rect 3976 1300 4028 1311
rect 4712 1300 4764 1352
rect 6828 1368 6880 1420
rect 8760 1368 8812 1420
rect 9496 1368 9548 1420
rect 6460 1343 6512 1352
rect 6460 1309 6469 1343
rect 6469 1309 6503 1343
rect 6503 1309 6512 1343
rect 6460 1300 6512 1309
rect 7012 1300 7064 1352
rect 7196 1343 7248 1352
rect 7196 1309 7205 1343
rect 7205 1309 7239 1343
rect 7239 1309 7248 1343
rect 7196 1300 7248 1309
rect 6368 1232 6420 1284
rect 5080 1164 5132 1216
rect 5724 1164 5776 1216
rect 7564 1164 7616 1216
rect 9128 1343 9180 1352
rect 9128 1309 9140 1343
rect 9140 1309 9174 1343
rect 9174 1309 9180 1343
rect 9128 1300 9180 1309
rect 10784 1164 10836 1216
rect 18236 1436 18288 1488
rect 11336 1368 11388 1420
rect 11612 1368 11664 1420
rect 11888 1300 11940 1352
rect 12164 1300 12216 1352
rect 11428 1232 11480 1284
rect 12348 1164 12400 1216
rect 13360 1207 13412 1216
rect 13360 1173 13369 1207
rect 13369 1173 13403 1207
rect 13403 1173 13412 1207
rect 13360 1164 13412 1173
rect 13728 1343 13780 1352
rect 13728 1309 13737 1343
rect 13737 1309 13771 1343
rect 13771 1309 13780 1343
rect 13728 1300 13780 1309
rect 15936 1368 15988 1420
rect 16120 1411 16172 1420
rect 16120 1377 16129 1411
rect 16129 1377 16163 1411
rect 16163 1377 16172 1411
rect 16120 1368 16172 1377
rect 20996 1504 21048 1556
rect 21548 1504 21600 1556
rect 23020 1504 23072 1556
rect 23756 1504 23808 1556
rect 23848 1504 23900 1556
rect 24124 1504 24176 1556
rect 24308 1504 24360 1556
rect 26884 1547 26936 1556
rect 26884 1513 26893 1547
rect 26893 1513 26927 1547
rect 26927 1513 26936 1547
rect 26884 1504 26936 1513
rect 20168 1436 20220 1488
rect 20812 1368 20864 1420
rect 20996 1411 21048 1420
rect 20996 1377 21005 1411
rect 21005 1377 21039 1411
rect 21039 1377 21048 1411
rect 20996 1368 21048 1377
rect 21180 1368 21232 1420
rect 14464 1343 14516 1352
rect 14464 1309 14473 1343
rect 14473 1309 14507 1343
rect 14507 1309 14516 1343
rect 14464 1300 14516 1309
rect 17960 1300 18012 1352
rect 18604 1300 18656 1352
rect 18788 1343 18840 1352
rect 18788 1309 18800 1343
rect 18800 1309 18834 1343
rect 18834 1309 18840 1343
rect 18788 1300 18840 1309
rect 21916 1300 21968 1352
rect 22836 1300 22888 1352
rect 23480 1343 23532 1352
rect 23480 1309 23489 1343
rect 23489 1309 23523 1343
rect 23523 1309 23532 1343
rect 23480 1300 23532 1309
rect 23756 1368 23808 1420
rect 24124 1368 24176 1420
rect 24308 1368 24360 1420
rect 25964 1411 26016 1420
rect 25964 1377 25973 1411
rect 25973 1377 26007 1411
rect 26007 1377 26016 1411
rect 25964 1368 26016 1377
rect 26240 1436 26292 1488
rect 27436 1547 27488 1556
rect 27436 1513 27445 1547
rect 27445 1513 27479 1547
rect 27479 1513 27488 1547
rect 27436 1504 27488 1513
rect 27804 1504 27856 1556
rect 29000 1504 29052 1556
rect 25136 1300 25188 1352
rect 26516 1368 26568 1420
rect 26976 1411 27028 1420
rect 26976 1377 26985 1411
rect 26985 1377 27019 1411
rect 27019 1377 27028 1411
rect 26976 1368 27028 1377
rect 27344 1368 27396 1420
rect 25320 1207 25372 1216
rect 25320 1173 25329 1207
rect 25329 1173 25363 1207
rect 25363 1173 25372 1207
rect 25320 1164 25372 1173
rect 25688 1207 25740 1216
rect 25688 1173 25697 1207
rect 25697 1173 25731 1207
rect 25731 1173 25740 1207
rect 25688 1164 25740 1173
rect 27712 1300 27764 1352
rect 28080 1300 28132 1352
rect 28172 1300 28224 1352
rect 28172 1164 28224 1216
rect 4193 1062 4245 1114
rect 4257 1062 4309 1114
rect 4321 1062 4373 1114
rect 4385 1062 4437 1114
rect 4449 1062 4501 1114
rect 11783 1062 11835 1114
rect 11847 1062 11899 1114
rect 11911 1062 11963 1114
rect 11975 1062 12027 1114
rect 12039 1062 12091 1114
rect 19373 1062 19425 1114
rect 19437 1062 19489 1114
rect 19501 1062 19553 1114
rect 19565 1062 19617 1114
rect 19629 1062 19681 1114
rect 26963 1062 27015 1114
rect 27027 1062 27079 1114
rect 27091 1062 27143 1114
rect 27155 1062 27207 1114
rect 27219 1062 27271 1114
rect 1308 960 1360 1012
rect 2504 892 2556 944
rect 2964 1003 3016 1012
rect 2964 969 2973 1003
rect 2973 969 3007 1003
rect 3007 969 3016 1003
rect 2964 960 3016 969
rect 4804 960 4856 1012
rect 5172 1003 5224 1012
rect 5172 969 5181 1003
rect 5181 969 5215 1003
rect 5215 969 5224 1003
rect 5172 960 5224 969
rect 6092 892 6144 944
rect 1584 824 1636 876
rect 1676 867 1728 876
rect 1676 833 1685 867
rect 1685 833 1719 867
rect 1719 833 1728 867
rect 1676 824 1728 833
rect 4712 756 4764 808
rect 4896 824 4948 876
rect 6644 824 6696 876
rect 7564 960 7616 1012
rect 9128 960 9180 1012
rect 9312 960 9364 1012
rect 11060 960 11112 1012
rect 11980 960 12032 1012
rect 13176 960 13228 1012
rect 13268 1003 13320 1012
rect 13268 969 13277 1003
rect 13277 969 13311 1003
rect 13311 969 13320 1003
rect 13268 960 13320 969
rect 15292 960 15344 1012
rect 16212 960 16264 1012
rect 15384 935 15436 944
rect 15384 901 15393 935
rect 15393 901 15427 935
rect 15427 901 15436 935
rect 15384 892 15436 901
rect 15476 892 15528 944
rect 5264 756 5316 808
rect 5356 799 5408 808
rect 5356 765 5365 799
rect 5365 765 5399 799
rect 5399 765 5408 799
rect 5356 756 5408 765
rect 3424 688 3476 740
rect 5908 756 5960 808
rect 1768 620 1820 672
rect 2688 620 2740 672
rect 4804 663 4856 672
rect 4804 629 4813 663
rect 4813 629 4847 663
rect 4847 629 4856 663
rect 4804 620 4856 629
rect 4896 663 4948 672
rect 4896 629 4905 663
rect 4905 629 4939 663
rect 4939 629 4948 663
rect 4896 620 4948 629
rect 5816 663 5868 672
rect 5816 629 5825 663
rect 5825 629 5859 663
rect 5859 629 5868 663
rect 5816 620 5868 629
rect 6000 620 6052 672
rect 6184 756 6236 808
rect 8576 799 8628 808
rect 8576 765 8585 799
rect 8585 765 8619 799
rect 8619 765 8628 799
rect 8576 756 8628 765
rect 8760 688 8812 740
rect 6460 620 6512 672
rect 9404 620 9456 672
rect 11244 867 11296 876
rect 11244 833 11253 867
rect 11253 833 11287 867
rect 11287 833 11296 867
rect 11244 824 11296 833
rect 11796 824 11848 876
rect 12348 824 12400 876
rect 14096 824 14148 876
rect 11336 756 11388 808
rect 11980 799 12032 808
rect 11980 765 11989 799
rect 11989 765 12023 799
rect 12023 765 12032 799
rect 11980 756 12032 765
rect 13636 756 13688 808
rect 14280 799 14332 808
rect 14280 765 14289 799
rect 14289 765 14323 799
rect 14323 765 14332 799
rect 14280 756 14332 765
rect 14556 756 14608 808
rect 16304 799 16356 808
rect 16304 765 16313 799
rect 16313 765 16347 799
rect 16347 765 16356 799
rect 16304 756 16356 765
rect 16856 849 16908 876
rect 18696 1003 18748 1012
rect 18696 969 18705 1003
rect 18705 969 18739 1003
rect 18739 969 18748 1003
rect 18696 960 18748 969
rect 19340 960 19392 1012
rect 20076 960 20128 1012
rect 16856 824 16901 849
rect 16901 824 16908 849
rect 16488 756 16540 808
rect 17132 799 17184 808
rect 17132 765 17141 799
rect 17141 765 17175 799
rect 17175 765 17184 799
rect 17132 756 17184 765
rect 22652 960 22704 1012
rect 22744 960 22796 1012
rect 21364 824 21416 876
rect 21916 824 21968 876
rect 22192 824 22244 876
rect 22928 824 22980 876
rect 19064 756 19116 808
rect 19340 799 19392 808
rect 19340 765 19342 799
rect 19342 765 19392 799
rect 19340 756 19392 765
rect 20628 756 20680 808
rect 20720 756 20772 808
rect 21456 799 21508 808
rect 21456 765 21465 799
rect 21465 765 21499 799
rect 21499 765 21508 799
rect 21456 756 21508 765
rect 22652 756 22704 808
rect 26056 960 26108 1012
rect 23664 892 23716 944
rect 24032 892 24084 944
rect 23940 756 23992 808
rect 24124 799 24176 808
rect 24124 765 24133 799
rect 24133 765 24167 799
rect 24167 765 24176 799
rect 24124 756 24176 765
rect 24676 824 24728 876
rect 29920 960 29972 1012
rect 28172 892 28224 944
rect 27620 824 27672 876
rect 27344 756 27396 808
rect 29092 756 29144 808
rect 20444 688 20496 740
rect 11612 620 11664 672
rect 12256 620 12308 672
rect 13820 620 13872 672
rect 15016 620 15068 672
rect 17960 620 18012 672
rect 18236 663 18288 672
rect 18236 629 18245 663
rect 18245 629 18279 663
rect 18279 629 18288 663
rect 18236 620 18288 629
rect 18328 620 18380 672
rect 23756 620 23808 672
rect 23940 620 23992 672
rect 24492 620 24544 672
rect 27804 620 27856 672
rect 7988 518 8040 570
rect 8052 518 8104 570
rect 8116 518 8168 570
rect 8180 518 8232 570
rect 8244 518 8296 570
rect 15578 518 15630 570
rect 15642 518 15694 570
rect 15706 518 15758 570
rect 15770 518 15822 570
rect 15834 518 15886 570
rect 23168 518 23220 570
rect 23232 518 23284 570
rect 23296 518 23348 570
rect 23360 518 23412 570
rect 23424 518 23476 570
rect 30758 518 30810 570
rect 30822 518 30874 570
rect 30886 518 30938 570
rect 30950 518 31002 570
rect 31014 518 31066 570
rect 1584 416 1636 468
rect 5816 416 5868 468
rect 11704 416 11756 468
rect 9128 348 9180 400
rect 14280 416 14332 468
rect 16856 416 16908 468
rect 17132 416 17184 468
rect 25688 416 25740 468
rect 24860 348 24912 400
rect 2688 280 2740 332
rect 17040 280 17092 332
rect 17960 280 18012 332
rect 23940 280 23992 332
rect 13360 212 13412 264
rect 19340 212 19392 264
rect 4988 144 5040 196
rect 5080 144 5132 196
rect 15108 144 15160 196
rect 16488 144 16540 196
rect 24124 144 24176 196
rect 9128 76 9180 128
rect 11796 76 11848 128
rect 18328 76 18380 128
rect 4712 8 4764 60
rect 6000 8 6052 60
rect 9772 8 9824 60
<< metal2 >>
rect 10968 22296 11020 22302
rect 10966 22264 10968 22273
rect 18880 22296 18932 22302
rect 11020 22264 11022 22273
rect 9128 22228 9180 22234
rect 15764 22234 16252 22250
rect 18880 22238 18932 22244
rect 24216 22296 24268 22302
rect 24216 22238 24268 22244
rect 25044 22296 25096 22302
rect 25044 22238 25096 22244
rect 31208 22296 31260 22302
rect 31208 22238 31260 22244
rect 10966 22199 11022 22208
rect 15752 22228 16252 22234
rect 9128 22170 9180 22176
rect 15804 22222 16252 22228
rect 15752 22170 15804 22176
rect 7564 22160 7616 22166
rect 7564 22102 7616 22108
rect 5448 21956 5500 21962
rect 5448 21898 5500 21904
rect 4804 21888 4856 21894
rect 4804 21830 4856 21836
rect 4193 21788 4501 21797
rect 4193 21786 4199 21788
rect 4255 21786 4279 21788
rect 4335 21786 4359 21788
rect 4415 21786 4439 21788
rect 4495 21786 4501 21788
rect 4255 21734 4257 21786
rect 4437 21734 4439 21786
rect 4193 21732 4199 21734
rect 4255 21732 4279 21734
rect 4335 21732 4359 21734
rect 4415 21732 4439 21734
rect 4495 21732 4501 21734
rect 4193 21723 4501 21732
rect 848 21480 900 21486
rect 848 21422 900 21428
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 3240 21480 3292 21486
rect 3240 21422 3292 21428
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 860 20398 888 21422
rect 1400 21344 1452 21350
rect 1320 21292 1400 21298
rect 1320 21286 1452 21292
rect 1320 21270 1440 21286
rect 940 20936 992 20942
rect 940 20878 992 20884
rect 848 20392 900 20398
rect 848 20334 900 20340
rect 860 19854 888 20334
rect 848 19848 900 19854
rect 848 19790 900 19796
rect 860 18290 888 19790
rect 848 18284 900 18290
rect 848 18226 900 18232
rect 848 16108 900 16114
rect 848 16050 900 16056
rect 756 13524 808 13530
rect 756 13466 808 13472
rect 664 10600 716 10606
rect 664 10542 716 10548
rect 676 2650 704 10542
rect 768 3738 796 13466
rect 860 4826 888 16050
rect 952 13938 980 20878
rect 1320 20466 1348 21270
rect 1400 21140 1452 21146
rect 1400 21082 1452 21088
rect 1308 20460 1360 20466
rect 1308 20402 1360 20408
rect 1320 20058 1348 20402
rect 1308 20052 1360 20058
rect 1308 19994 1360 20000
rect 1032 19304 1084 19310
rect 1032 19246 1084 19252
rect 1044 18714 1072 19246
rect 1412 18952 1440 21082
rect 1674 21040 1730 21049
rect 1674 20975 1676 20984
rect 1728 20975 1730 20984
rect 1676 20946 1728 20952
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1674 20496 1730 20505
rect 1584 20460 1636 20466
rect 1674 20431 1676 20440
rect 1584 20402 1636 20408
rect 1728 20431 1730 20440
rect 1676 20402 1728 20408
rect 1412 18924 1532 18952
rect 1216 18828 1268 18834
rect 1268 18788 1440 18816
rect 1216 18770 1268 18776
rect 1124 18760 1176 18766
rect 1044 18708 1124 18714
rect 1412 18737 1440 18788
rect 1044 18702 1176 18708
rect 1398 18728 1454 18737
rect 1044 18686 1164 18702
rect 1032 18624 1084 18630
rect 1032 18566 1084 18572
rect 1044 16794 1072 18566
rect 1136 18426 1164 18686
rect 1398 18663 1454 18672
rect 1124 18420 1176 18426
rect 1124 18362 1176 18368
rect 1136 17814 1164 18362
rect 1306 18184 1362 18193
rect 1306 18119 1362 18128
rect 1124 17808 1176 17814
rect 1124 17750 1176 17756
rect 1136 17202 1164 17750
rect 1124 17196 1176 17202
rect 1124 17138 1176 17144
rect 1032 16788 1084 16794
rect 1032 16730 1084 16736
rect 1320 16726 1348 18119
rect 1308 16720 1360 16726
rect 1308 16662 1360 16668
rect 1124 16652 1176 16658
rect 1124 16594 1176 16600
rect 1032 15360 1084 15366
rect 1032 15302 1084 15308
rect 940 13932 992 13938
rect 940 13874 992 13880
rect 952 11694 980 13874
rect 1044 12442 1072 15302
rect 1136 14074 1164 16594
rect 1216 16584 1268 16590
rect 1216 16526 1268 16532
rect 1228 15994 1256 16526
rect 1228 15966 1348 15994
rect 1320 15910 1348 15966
rect 1308 15904 1360 15910
rect 1308 15846 1360 15852
rect 1320 15366 1348 15846
rect 1504 15688 1532 18924
rect 1596 17338 1624 20402
rect 1768 20052 1820 20058
rect 1768 19994 1820 20000
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 1688 19417 1716 19790
rect 1674 19408 1730 19417
rect 1674 19343 1730 19352
rect 1780 19258 1808 19994
rect 1688 19230 1808 19258
rect 1688 18970 1716 19230
rect 1768 19168 1820 19174
rect 1768 19110 1820 19116
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1688 18086 1716 18906
rect 1780 18630 1808 19110
rect 1768 18624 1820 18630
rect 1768 18566 1820 18572
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1676 17740 1728 17746
rect 1780 17728 1808 18566
rect 1728 17700 1808 17728
rect 1676 17682 1728 17688
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1780 16998 1808 17700
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1872 16946 1900 20878
rect 2792 19514 2820 21422
rect 2872 21412 2924 21418
rect 2872 21354 2924 21360
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2136 19304 2188 19310
rect 2136 19246 2188 19252
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 1872 16918 1992 16946
rect 1766 16824 1822 16833
rect 1766 16759 1822 16768
rect 1860 16788 1912 16794
rect 1780 16590 1808 16759
rect 1860 16730 1912 16736
rect 1872 16590 1900 16730
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1768 16584 1820 16590
rect 1768 16526 1820 16532
rect 1860 16584 1912 16590
rect 1860 16526 1912 16532
rect 1596 15910 1624 16526
rect 1964 16402 1992 16918
rect 2056 16454 2084 17614
rect 1872 16374 1992 16402
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 1584 15904 1636 15910
rect 1584 15846 1636 15852
rect 1412 15660 1532 15688
rect 1308 15360 1360 15366
rect 1308 15302 1360 15308
rect 1320 15026 1348 15302
rect 1308 15020 1360 15026
rect 1308 14962 1360 14968
rect 1124 14068 1176 14074
rect 1124 14010 1176 14016
rect 1136 13462 1164 14010
rect 1412 13954 1440 15660
rect 1596 15586 1624 15846
rect 1596 15558 1716 15586
rect 1688 15502 1716 15558
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1688 14822 1716 15438
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1320 13938 1440 13954
rect 1308 13932 1440 13938
rect 1360 13926 1440 13932
rect 1308 13874 1360 13880
rect 1124 13456 1176 13462
rect 1124 13398 1176 13404
rect 1308 13320 1360 13326
rect 1308 13262 1360 13268
rect 1320 12850 1348 13262
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 1032 12436 1084 12442
rect 1032 12378 1084 12384
rect 1216 12300 1268 12306
rect 1216 12242 1268 12248
rect 1228 12209 1256 12242
rect 1320 12238 1348 12786
rect 1308 12232 1360 12238
rect 1214 12200 1270 12209
rect 1308 12174 1360 12180
rect 1214 12135 1270 12144
rect 940 11688 992 11694
rect 940 11630 992 11636
rect 1216 11688 1268 11694
rect 1216 11630 1268 11636
rect 940 10124 992 10130
rect 940 10066 992 10072
rect 952 9586 980 10066
rect 940 9580 992 9586
rect 940 9522 992 9528
rect 1228 8974 1256 11630
rect 1320 11354 1348 12174
rect 1412 11558 1440 13926
rect 1504 13326 1532 14418
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1688 13326 1716 14350
rect 1780 13530 1808 14894
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1688 12646 1716 13262
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1688 12306 1716 12582
rect 1766 12336 1822 12345
rect 1676 12300 1728 12306
rect 1766 12271 1822 12280
rect 1676 12242 1728 12248
rect 1688 11778 1716 12242
rect 1780 12238 1808 12271
rect 1768 12232 1820 12238
rect 1768 12174 1820 12180
rect 1688 11750 1808 11778
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1308 11348 1360 11354
rect 1308 11290 1360 11296
rect 1320 10674 1348 11290
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 1320 10266 1348 10610
rect 1308 10260 1360 10266
rect 1308 10202 1360 10208
rect 1308 9172 1360 9178
rect 1308 9114 1360 9120
rect 1216 8968 1268 8974
rect 1216 8910 1268 8916
rect 1228 8634 1256 8910
rect 1216 8628 1268 8634
rect 1216 8570 1268 8576
rect 1320 8514 1348 9114
rect 1412 9042 1440 11494
rect 1596 11218 1624 11494
rect 1584 11212 1636 11218
rect 1584 11154 1636 11160
rect 1490 10160 1546 10169
rect 1490 10095 1546 10104
rect 1504 10062 1532 10095
rect 1492 10056 1544 10062
rect 1688 10033 1716 11630
rect 1780 11354 1808 11750
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1780 10470 1808 11290
rect 1872 10985 1900 16374
rect 2148 16017 2176 19246
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2332 16250 2360 18770
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2134 16008 2190 16017
rect 2134 15943 2190 15952
rect 2044 15496 2096 15502
rect 2042 15464 2044 15473
rect 2096 15464 2098 15473
rect 2042 15399 2098 15408
rect 2134 15056 2190 15065
rect 2134 14991 2136 15000
rect 2188 14991 2190 15000
rect 2136 14962 2188 14968
rect 2042 14512 2098 14521
rect 2042 14447 2098 14456
rect 2056 14414 2084 14447
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 1950 13424 2006 13433
rect 1950 13359 2006 13368
rect 1964 13326 1992 13359
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 1950 11248 2006 11257
rect 1950 11183 2006 11192
rect 1964 11150 1992 11183
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1858 10976 1914 10985
rect 1858 10911 1914 10920
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1780 10266 1808 10406
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1492 9998 1544 10004
rect 1674 10024 1730 10033
rect 1674 9959 1730 9968
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1228 8486 1348 8514
rect 1032 8424 1084 8430
rect 1032 8366 1084 8372
rect 1044 7886 1072 8366
rect 1124 7948 1176 7954
rect 1124 7890 1176 7896
rect 1032 7880 1084 7886
rect 1032 7822 1084 7828
rect 940 7744 992 7750
rect 940 7686 992 7692
rect 952 7546 980 7686
rect 940 7540 992 7546
rect 940 7482 992 7488
rect 1044 7342 1072 7822
rect 1032 7336 1084 7342
rect 1032 7278 1084 7284
rect 1044 6730 1072 7278
rect 1136 7177 1164 7890
rect 1122 7168 1178 7177
rect 1122 7103 1178 7112
rect 1032 6724 1084 6730
rect 1032 6666 1084 6672
rect 940 5704 992 5710
rect 940 5646 992 5652
rect 952 5370 980 5646
rect 940 5364 992 5370
rect 940 5306 992 5312
rect 848 4820 900 4826
rect 848 4762 900 4768
rect 756 3732 808 3738
rect 756 3674 808 3680
rect 952 3534 980 5306
rect 1032 4072 1084 4078
rect 1032 4014 1084 4020
rect 940 3528 992 3534
rect 940 3470 992 3476
rect 664 2644 716 2650
rect 664 2586 716 2592
rect 1044 2514 1072 4014
rect 1136 3670 1164 7103
rect 1124 3664 1176 3670
rect 1124 3606 1176 3612
rect 1228 3602 1256 8486
rect 1308 6112 1360 6118
rect 1308 6054 1360 6060
rect 1320 5710 1348 6054
rect 1308 5704 1360 5710
rect 1308 5646 1360 5652
rect 1320 5234 1348 5646
rect 1412 5409 1440 8978
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1596 8090 1624 8230
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1492 7880 1544 7886
rect 1490 7848 1492 7857
rect 1544 7848 1546 7857
rect 1490 7783 1546 7792
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1398 5400 1454 5409
rect 1398 5335 1454 5344
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 1320 4690 1348 5170
rect 1308 4684 1360 4690
rect 1308 4626 1360 4632
rect 1320 4146 1348 4626
rect 1504 4146 1532 7686
rect 1596 7206 1624 8026
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 7002 1624 7142
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1582 6352 1638 6361
rect 1582 6287 1638 6296
rect 1596 6254 1624 6287
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1596 5778 1624 6054
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1596 4690 1624 4966
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1308 4140 1360 4146
rect 1308 4082 1360 4088
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1216 3596 1268 3602
rect 1216 3538 1268 3544
rect 1320 3058 1348 4082
rect 1688 3466 1716 9454
rect 1780 9382 1808 10202
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1766 9072 1822 9081
rect 1766 9007 1768 9016
rect 1820 9007 1822 9016
rect 1768 8978 1820 8984
rect 1766 7304 1822 7313
rect 1766 7239 1822 7248
rect 1780 6798 1808 7239
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1780 5030 1808 6054
rect 1872 5914 1900 9998
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 3942 1808 4966
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1674 3088 1730 3097
rect 1308 3052 1360 3058
rect 1674 3023 1730 3032
rect 1308 2994 1360 3000
rect 1688 2990 1716 3023
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1780 2854 1808 3878
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 1400 2644 1452 2650
rect 1400 2586 1452 2592
rect 1032 2508 1084 2514
rect 1032 2450 1084 2456
rect 1412 1986 1440 2586
rect 1228 1958 1440 1986
rect 1674 2000 1730 2009
rect 1492 1964 1544 1970
rect 1228 1562 1256 1958
rect 1674 1935 1676 1944
rect 1492 1906 1544 1912
rect 1728 1935 1730 1944
rect 1676 1906 1728 1912
rect 1308 1896 1360 1902
rect 1308 1838 1360 1844
rect 1216 1556 1268 1562
rect 1216 1498 1268 1504
rect 1320 1358 1348 1838
rect 1308 1352 1360 1358
rect 1308 1294 1360 1300
rect 1320 1018 1348 1294
rect 1308 1012 1360 1018
rect 1308 954 1360 960
rect 1504 785 1532 1906
rect 1676 1760 1728 1766
rect 1676 1702 1728 1708
rect 1688 1358 1716 1702
rect 1780 1562 1808 2790
rect 1964 2650 1992 7822
rect 2056 6662 2084 13262
rect 2134 12880 2190 12889
rect 2134 12815 2136 12824
rect 2188 12815 2190 12824
rect 2136 12786 2188 12792
rect 2332 12481 2360 13874
rect 2424 13569 2452 17070
rect 2700 16153 2728 18226
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2686 16144 2742 16153
rect 2686 16079 2742 16088
rect 2792 15162 2820 17138
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 2504 15088 2556 15094
rect 2504 15030 2556 15036
rect 2516 14618 2544 15030
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 2596 14612 2648 14618
rect 2596 14554 2648 14560
rect 2608 14482 2636 14554
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2410 13560 2466 13569
rect 2410 13495 2466 13504
rect 2318 12472 2374 12481
rect 2136 12436 2188 12442
rect 2318 12407 2374 12416
rect 2136 12378 2188 12384
rect 2148 12238 2176 12378
rect 2226 12336 2282 12345
rect 2226 12271 2282 12280
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2136 12096 2188 12102
rect 2136 12038 2188 12044
rect 2148 11218 2176 12038
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2240 9178 2268 12271
rect 2608 9994 2636 13806
rect 2778 13288 2834 13297
rect 2778 13223 2834 13232
rect 2792 11898 2820 13223
rect 2884 12866 2912 21354
rect 3252 20924 3280 21422
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3884 21344 3936 21350
rect 3884 21286 3936 21292
rect 3620 21146 3648 21286
rect 3608 21140 3660 21146
rect 3608 21082 3660 21088
rect 3332 20936 3384 20942
rect 3252 20896 3332 20924
rect 3332 20878 3384 20884
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 2964 20800 3016 20806
rect 2962 20768 2964 20777
rect 3016 20768 3018 20777
rect 2962 20703 3018 20712
rect 3148 19916 3200 19922
rect 3148 19858 3200 19864
rect 3056 19372 3108 19378
rect 3056 19314 3108 19320
rect 3068 16794 3096 19314
rect 3160 18970 3188 19858
rect 3344 19854 3372 20878
rect 3620 20602 3648 20878
rect 3608 20596 3660 20602
rect 3608 20538 3660 20544
rect 3424 20392 3476 20398
rect 3424 20334 3476 20340
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 3344 19514 3372 19790
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 3344 18222 3372 19450
rect 3436 18358 3464 20334
rect 3700 20324 3752 20330
rect 3700 20266 3752 20272
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3620 19825 3648 19858
rect 3606 19816 3662 19825
rect 3606 19751 3662 19760
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 3424 18352 3476 18358
rect 3424 18294 3476 18300
rect 3332 18216 3384 18222
rect 3332 18158 3384 18164
rect 3148 18080 3200 18086
rect 3148 18022 3200 18028
rect 3160 17882 3188 18022
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3148 17740 3200 17746
rect 3148 17682 3200 17688
rect 3056 16788 3108 16794
rect 3056 16730 3108 16736
rect 3160 15706 3188 17682
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 3252 17338 3280 17478
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3068 14550 3096 15642
rect 3252 14958 3280 17070
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3528 15910 3556 16526
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3528 15502 3556 15846
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 3516 15088 3568 15094
rect 3516 15030 3568 15036
rect 3240 14952 3292 14958
rect 3240 14894 3292 14900
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3056 14544 3108 14550
rect 3056 14486 3108 14492
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3056 13864 3108 13870
rect 3054 13832 3056 13841
rect 3108 13832 3110 13841
rect 3054 13767 3110 13776
rect 3160 12986 3188 14350
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 2884 12838 3188 12866
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2976 10130 3004 11494
rect 3160 11098 3188 12838
rect 3252 12782 3280 13670
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3252 11529 3280 12582
rect 3436 11642 3464 14554
rect 3528 12968 3556 15030
rect 3620 14822 3648 19246
rect 3712 18222 3740 20266
rect 3896 19922 3924 21286
rect 4080 20058 4108 21422
rect 4193 20700 4501 20709
rect 4193 20698 4199 20700
rect 4255 20698 4279 20700
rect 4335 20698 4359 20700
rect 4415 20698 4439 20700
rect 4495 20698 4501 20700
rect 4255 20646 4257 20698
rect 4437 20646 4439 20698
rect 4193 20644 4199 20646
rect 4255 20644 4279 20646
rect 4335 20644 4359 20646
rect 4415 20644 4439 20646
rect 4495 20644 4501 20646
rect 4193 20635 4501 20644
rect 4712 20596 4764 20602
rect 4712 20538 4764 20544
rect 4528 20392 4580 20398
rect 4528 20334 4580 20340
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 3884 19916 3936 19922
rect 3884 19858 3936 19864
rect 3896 19378 3924 19858
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 3884 19236 3936 19242
rect 3884 19178 3936 19184
rect 3896 19145 3924 19178
rect 3882 19136 3938 19145
rect 3882 19071 3938 19080
rect 3896 18834 3924 19071
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3700 18216 3752 18222
rect 3700 18158 3752 18164
rect 3712 17678 3740 18158
rect 3804 17785 3832 18566
rect 4080 18426 4108 19790
rect 4193 19612 4501 19621
rect 4193 19610 4199 19612
rect 4255 19610 4279 19612
rect 4335 19610 4359 19612
rect 4415 19610 4439 19612
rect 4495 19610 4501 19612
rect 4255 19558 4257 19610
rect 4437 19558 4439 19610
rect 4193 19556 4199 19558
rect 4255 19556 4279 19558
rect 4335 19556 4359 19558
rect 4415 19556 4439 19558
rect 4495 19556 4501 19558
rect 4193 19547 4501 19556
rect 4540 19310 4568 20334
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4724 18902 4752 20538
rect 4816 19242 4844 21830
rect 5460 21486 5488 21898
rect 7576 21690 7604 22102
rect 7748 21956 7800 21962
rect 7748 21898 7800 21904
rect 7564 21684 7616 21690
rect 7564 21626 7616 21632
rect 5448 21480 5500 21486
rect 6184 21480 6236 21486
rect 5448 21422 5500 21428
rect 5906 21448 5962 21457
rect 5356 21412 5408 21418
rect 5356 21354 5408 21360
rect 4896 20392 4948 20398
rect 4896 20334 4948 20340
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 4712 18896 4764 18902
rect 4712 18838 4764 18844
rect 4193 18524 4501 18533
rect 4193 18522 4199 18524
rect 4255 18522 4279 18524
rect 4335 18522 4359 18524
rect 4415 18522 4439 18524
rect 4495 18522 4501 18524
rect 4255 18470 4257 18522
rect 4437 18470 4439 18522
rect 4193 18468 4199 18470
rect 4255 18468 4279 18470
rect 4335 18468 4359 18470
rect 4415 18468 4439 18470
rect 4495 18468 4501 18470
rect 4193 18459 4501 18468
rect 4618 18456 4674 18465
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4160 18420 4212 18426
rect 4674 18414 4844 18442
rect 4618 18391 4674 18400
rect 4160 18362 4212 18368
rect 4172 18306 4200 18362
rect 4080 18290 4200 18306
rect 4068 18284 4200 18290
rect 4120 18278 4200 18284
rect 4068 18226 4120 18232
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4528 18080 4580 18086
rect 4632 18057 4660 18158
rect 4528 18022 4580 18028
rect 4618 18048 4674 18057
rect 4540 17882 4568 18022
rect 4618 17983 4674 17992
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 3790 17776 3846 17785
rect 3790 17711 3846 17720
rect 3700 17672 3752 17678
rect 3700 17614 3752 17620
rect 3712 17270 3740 17614
rect 4193 17436 4501 17445
rect 4193 17434 4199 17436
rect 4255 17434 4279 17436
rect 4335 17434 4359 17436
rect 4415 17434 4439 17436
rect 4495 17434 4501 17436
rect 4255 17382 4257 17434
rect 4437 17382 4439 17434
rect 4193 17380 4199 17382
rect 4255 17380 4279 17382
rect 4335 17380 4359 17382
rect 4415 17380 4439 17382
rect 4495 17380 4501 17382
rect 4193 17371 4501 17380
rect 3700 17264 3752 17270
rect 3700 17206 3752 17212
rect 3712 16182 3740 17206
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 4080 16658 4108 17138
rect 4540 16998 4568 17818
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4712 16652 4764 16658
rect 4712 16594 4764 16600
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3976 16584 4028 16590
rect 4066 16552 4122 16561
rect 4028 16532 4066 16538
rect 3976 16526 4066 16532
rect 3792 16448 3844 16454
rect 3792 16390 3844 16396
rect 3804 16182 3832 16390
rect 3700 16176 3752 16182
rect 3700 16118 3752 16124
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 3896 15910 3924 16526
rect 3988 16510 4066 16526
rect 4066 16487 4122 16496
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 15502 3924 15846
rect 4080 15502 4108 16390
rect 4193 16348 4501 16357
rect 4193 16346 4199 16348
rect 4255 16346 4279 16348
rect 4335 16346 4359 16348
rect 4415 16346 4439 16348
rect 4495 16346 4501 16348
rect 4255 16294 4257 16346
rect 4437 16294 4439 16346
rect 4193 16292 4199 16294
rect 4255 16292 4279 16294
rect 4335 16292 4359 16294
rect 4415 16292 4439 16294
rect 4495 16292 4501 16294
rect 4193 16283 4501 16292
rect 4436 16040 4488 16046
rect 4436 15982 4488 15988
rect 4448 15910 4476 15982
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 4068 15496 4120 15502
rect 4068 15438 4120 15444
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 15026 3832 15302
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3896 14958 3924 15438
rect 4193 15260 4501 15269
rect 4193 15258 4199 15260
rect 4255 15258 4279 15260
rect 4335 15258 4359 15260
rect 4415 15258 4439 15260
rect 4495 15258 4501 15260
rect 4255 15206 4257 15258
rect 4437 15206 4439 15258
rect 4193 15204 4199 15206
rect 4255 15204 4279 15206
rect 4335 15204 4359 15206
rect 4415 15204 4439 15206
rect 4495 15204 4501 15206
rect 4193 15195 4501 15204
rect 4540 15042 4568 15506
rect 4448 15014 4568 15042
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 4448 14618 4476 15014
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4540 14618 4568 14894
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4632 14482 4660 14758
rect 4724 14482 4752 16594
rect 4436 14476 4488 14482
rect 4620 14476 4672 14482
rect 4488 14436 4568 14464
rect 4436 14418 4488 14424
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3804 14006 3832 14350
rect 4193 14172 4501 14181
rect 4193 14170 4199 14172
rect 4255 14170 4279 14172
rect 4335 14170 4359 14172
rect 4415 14170 4439 14172
rect 4495 14170 4501 14172
rect 4255 14118 4257 14170
rect 4437 14118 4439 14170
rect 4193 14116 4199 14118
rect 4255 14116 4279 14118
rect 4335 14116 4359 14118
rect 4415 14116 4439 14118
rect 4495 14116 4501 14118
rect 4193 14107 4501 14116
rect 3792 14000 3844 14006
rect 3792 13942 3844 13948
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3804 13190 3832 13806
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3896 13326 3924 13670
rect 3884 13320 3936 13326
rect 3936 13268 4016 13274
rect 3884 13262 4016 13268
rect 3896 13246 4016 13262
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3608 12980 3660 12986
rect 3528 12940 3608 12968
rect 3608 12922 3660 12928
rect 3620 12782 3648 12922
rect 3804 12782 3832 13126
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3516 12232 3568 12238
rect 3804 12220 3832 12718
rect 3988 12646 4016 13246
rect 4193 13084 4501 13093
rect 4193 13082 4199 13084
rect 4255 13082 4279 13084
rect 4335 13082 4359 13084
rect 4415 13082 4439 13084
rect 4495 13082 4501 13084
rect 4255 13030 4257 13082
rect 4437 13030 4439 13082
rect 4193 13028 4199 13030
rect 4255 13028 4279 13030
rect 4335 13028 4359 13030
rect 4415 13028 4439 13030
rect 4495 13028 4501 13030
rect 4193 13019 4501 13028
rect 3976 12640 4028 12646
rect 4028 12600 4108 12628
rect 3976 12582 4028 12588
rect 3568 12192 3832 12220
rect 3516 12174 3568 12180
rect 3528 11762 3556 12174
rect 3804 11880 3832 12192
rect 3884 12232 3936 12238
rect 4080 12220 4108 12600
rect 4540 12434 4568 14436
rect 4620 14418 4672 14424
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4816 14385 4844 18414
rect 4802 14376 4858 14385
rect 4712 14340 4764 14346
rect 4802 14311 4858 14320
rect 4712 14282 4764 14288
rect 4724 13938 4752 14282
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4632 12850 4660 13874
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4816 12434 4844 14214
rect 4540 12406 4660 12434
rect 3936 12192 4108 12220
rect 3884 12174 3936 12180
rect 3804 11852 4016 11880
rect 3700 11824 3752 11830
rect 3752 11784 3832 11812
rect 3700 11766 3752 11772
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3436 11614 3740 11642
rect 3424 11552 3476 11558
rect 3238 11520 3294 11529
rect 3424 11494 3476 11500
rect 3516 11552 3568 11558
rect 3516 11494 3568 11500
rect 3238 11455 3294 11464
rect 3436 11393 3464 11494
rect 3422 11384 3478 11393
rect 3422 11319 3478 11328
rect 3160 11070 3464 11098
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3056 10532 3108 10538
rect 3056 10474 3108 10480
rect 3068 10266 3096 10474
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 3068 9586 3096 9862
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 3160 9110 3188 10542
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3252 9518 3280 9998
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 3252 8974 3280 9454
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2148 7528 2176 8366
rect 2148 7500 2268 7528
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2148 7002 2176 7346
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 2148 5137 2176 6190
rect 2134 5128 2190 5137
rect 2134 5063 2190 5072
rect 2240 2774 2268 7500
rect 2318 6896 2374 6905
rect 2318 6831 2320 6840
rect 2372 6831 2374 6840
rect 2320 6802 2372 6808
rect 2424 6118 2452 8502
rect 2504 8424 2556 8430
rect 2502 8392 2504 8401
rect 2556 8392 2558 8401
rect 2502 8327 2558 8336
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2686 7440 2742 7449
rect 2608 7398 2686 7426
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2502 5672 2558 5681
rect 2502 5607 2558 5616
rect 2516 5370 2544 5607
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2608 5234 2636 7398
rect 2686 7375 2742 7384
rect 2686 6080 2742 6089
rect 2686 6015 2742 6024
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2332 4865 2360 5102
rect 2318 4856 2374 4865
rect 2318 4791 2374 4800
rect 2700 4146 2728 6015
rect 2792 4690 2820 8230
rect 2884 5642 2912 8570
rect 3054 8120 3110 8129
rect 3054 8055 3110 8064
rect 3068 7546 3096 8055
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2884 5234 2912 5578
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2870 4992 2926 5001
rect 2870 4927 2926 4936
rect 2884 4826 2912 4927
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2778 4040 2834 4049
rect 2778 3975 2834 3984
rect 2792 3942 2820 3975
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2976 3058 3004 7142
rect 3160 7002 3188 7686
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3252 7002 3280 7210
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 3146 6760 3202 6769
rect 3146 6695 3202 6704
rect 3160 5658 3188 6695
rect 3068 5630 3188 5658
rect 3344 5658 3372 10406
rect 3436 9353 3464 11070
rect 3528 9602 3556 11494
rect 3606 10704 3662 10713
rect 3606 10639 3662 10648
rect 3620 10606 3648 10639
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3620 9674 3648 10542
rect 3712 10305 3740 11614
rect 3698 10296 3754 10305
rect 3698 10231 3754 10240
rect 3804 10130 3832 11784
rect 3882 11520 3938 11529
rect 3882 11455 3938 11464
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 3896 9674 3924 11455
rect 3988 11150 4016 11852
rect 4080 11558 4108 12192
rect 4193 11996 4501 12005
rect 4193 11994 4199 11996
rect 4255 11994 4279 11996
rect 4335 11994 4359 11996
rect 4415 11994 4439 11996
rect 4495 11994 4501 11996
rect 4255 11942 4257 11994
rect 4437 11942 4439 11994
rect 4193 11940 4199 11942
rect 4255 11940 4279 11942
rect 4335 11940 4359 11942
rect 4415 11940 4439 11942
rect 4495 11940 4501 11942
rect 4193 11931 4501 11940
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4080 11286 4108 11494
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 3974 10568 4030 10577
rect 3974 10503 4030 10512
rect 3988 10470 4016 10503
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3974 10296 4030 10305
rect 4080 10266 4108 11222
rect 4172 10996 4200 11630
rect 4264 11218 4292 11698
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4540 11234 4568 11494
rect 4632 11370 4660 12406
rect 4724 12406 4844 12434
rect 4724 12306 4752 12406
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4802 11384 4858 11393
rect 4632 11342 4802 11370
rect 4802 11319 4858 11328
rect 4252 11212 4304 11218
rect 4540 11206 4660 11234
rect 4252 11154 4304 11160
rect 4632 11082 4660 11206
rect 4710 11112 4766 11121
rect 4620 11076 4672 11082
rect 4710 11047 4766 11056
rect 4620 11018 4672 11024
rect 4172 10968 4568 10996
rect 4193 10908 4501 10917
rect 4193 10906 4199 10908
rect 4255 10906 4279 10908
rect 4335 10906 4359 10908
rect 4415 10906 4439 10908
rect 4495 10906 4501 10908
rect 4255 10854 4257 10906
rect 4437 10854 4439 10906
rect 4193 10852 4199 10854
rect 4255 10852 4279 10854
rect 4335 10852 4359 10854
rect 4415 10852 4439 10854
rect 4495 10852 4501 10854
rect 4193 10843 4501 10852
rect 3974 10231 4030 10240
rect 4068 10260 4120 10266
rect 3620 9646 3740 9674
rect 3528 9574 3648 9602
rect 3620 9518 3648 9574
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3608 9376 3660 9382
rect 3422 9344 3478 9353
rect 3608 9318 3660 9324
rect 3422 9279 3478 9288
rect 3620 8974 3648 9318
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3528 7886 3556 8026
rect 3608 8016 3660 8022
rect 3608 7958 3660 7964
rect 3712 7970 3740 9646
rect 3804 9646 3924 9674
rect 3804 9042 3832 9646
rect 3988 9586 4016 10231
rect 4068 10202 4120 10208
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 4080 9382 4108 10202
rect 4193 9820 4501 9829
rect 4193 9818 4199 9820
rect 4255 9818 4279 9820
rect 4335 9818 4359 9820
rect 4415 9818 4439 9820
rect 4495 9818 4501 9820
rect 4255 9766 4257 9818
rect 4437 9766 4439 9818
rect 4193 9764 4199 9766
rect 4255 9764 4279 9766
rect 4335 9764 4359 9766
rect 4415 9764 4439 9766
rect 4495 9764 4501 9766
rect 4193 9755 4501 9764
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4344 9376 4396 9382
rect 4344 9318 4396 9324
rect 4434 9344 4490 9353
rect 4080 9178 4108 9318
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3884 8968 3936 8974
rect 3804 8916 3884 8922
rect 3804 8910 3936 8916
rect 3804 8894 3924 8910
rect 3804 8634 3832 8894
rect 3884 8832 3936 8838
rect 4356 8820 4384 9318
rect 4434 9279 4490 9288
rect 4448 8974 4476 9279
rect 4540 9217 4568 10968
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4526 9208 4582 9217
rect 4526 9143 4582 9152
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4356 8792 4568 8820
rect 3884 8774 3936 8780
rect 3896 8634 3924 8774
rect 4193 8732 4501 8741
rect 4193 8730 4199 8732
rect 4255 8730 4279 8732
rect 4335 8730 4359 8732
rect 4415 8730 4439 8732
rect 4495 8730 4501 8732
rect 4255 8678 4257 8730
rect 4437 8678 4439 8730
rect 4193 8676 4199 8678
rect 4255 8676 4279 8678
rect 4335 8676 4359 8678
rect 4415 8676 4439 8678
rect 4495 8676 4501 8678
rect 4193 8667 4501 8676
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3884 8628 3936 8634
rect 3884 8570 3936 8576
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 3804 8350 4016 8378
rect 3804 8294 3832 8350
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3516 7880 3568 7886
rect 3514 7848 3516 7857
rect 3620 7868 3648 7958
rect 3712 7942 3832 7970
rect 3700 7880 3752 7886
rect 3568 7848 3570 7857
rect 3620 7840 3700 7868
rect 3700 7822 3752 7828
rect 3514 7783 3570 7792
rect 3528 7546 3556 7783
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3528 6866 3556 7482
rect 3620 6934 3648 7482
rect 3712 7410 3740 7822
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3608 6928 3660 6934
rect 3608 6870 3660 6876
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3528 6322 3556 6802
rect 3712 6798 3740 7346
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3712 6322 3740 6734
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3528 5914 3556 6258
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3344 5630 3556 5658
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 3068 2774 3096 5630
rect 3332 5568 3384 5574
rect 3146 5536 3202 5545
rect 3332 5510 3384 5516
rect 3146 5471 3202 5480
rect 3160 4826 3188 5471
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3252 4146 3280 5170
rect 3344 4146 3372 5510
rect 3422 5264 3478 5273
rect 3422 5199 3478 5208
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3252 3670 3280 4082
rect 3436 4078 3464 5199
rect 3528 4554 3556 5630
rect 3804 4706 3832 7942
rect 3896 7886 3924 8230
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3988 6361 4016 8350
rect 4080 7546 4108 8434
rect 4160 7880 4212 7886
rect 4158 7848 4160 7857
rect 4212 7848 4214 7857
rect 4158 7783 4214 7792
rect 4193 7644 4501 7653
rect 4193 7642 4199 7644
rect 4255 7642 4279 7644
rect 4335 7642 4359 7644
rect 4415 7642 4439 7644
rect 4495 7642 4501 7644
rect 4255 7590 4257 7642
rect 4437 7590 4439 7642
rect 4193 7588 4199 7590
rect 4255 7588 4279 7590
rect 4335 7588 4359 7590
rect 4415 7588 4439 7590
rect 4495 7588 4501 7590
rect 4193 7579 4501 7588
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4158 6896 4214 6905
rect 4540 6882 4568 8792
rect 4214 6854 4568 6882
rect 4158 6831 4214 6840
rect 4172 6746 4200 6831
rect 4080 6718 4200 6746
rect 3974 6352 4030 6361
rect 4080 6338 4108 6718
rect 4193 6556 4501 6565
rect 4193 6554 4199 6556
rect 4255 6554 4279 6556
rect 4335 6554 4359 6556
rect 4415 6554 4439 6556
rect 4495 6554 4501 6556
rect 4255 6502 4257 6554
rect 4437 6502 4439 6554
rect 4193 6500 4199 6502
rect 4255 6500 4279 6502
rect 4335 6500 4359 6502
rect 4415 6500 4439 6502
rect 4495 6500 4501 6502
rect 4193 6491 4501 6500
rect 4632 6338 4660 9998
rect 4080 6310 4200 6338
rect 3974 6287 4030 6296
rect 3988 5778 4016 6287
rect 4172 5778 4200 6310
rect 4448 6310 4660 6338
rect 4448 5930 4476 6310
rect 4528 6112 4580 6118
rect 4580 6072 4660 6100
rect 4528 6054 4580 6060
rect 4448 5902 4568 5930
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 3896 5574 3924 5714
rect 3988 5574 4016 5714
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3620 4690 3832 4706
rect 3608 4684 3832 4690
rect 3660 4678 3832 4684
rect 3608 4626 3660 4632
rect 3516 4548 3568 4554
rect 3516 4490 3568 4496
rect 3424 4072 3476 4078
rect 3424 4014 3476 4020
rect 3330 3904 3386 3913
rect 3330 3839 3386 3848
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 3252 2990 3280 3606
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 2148 2746 2268 2774
rect 2976 2746 3096 2774
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 1858 2544 1914 2553
rect 1858 2479 1914 2488
rect 1952 2508 2004 2514
rect 1872 2446 1900 2479
rect 2056 2496 2084 2586
rect 2004 2468 2084 2496
rect 1952 2450 2004 2456
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 1768 1556 1820 1562
rect 1768 1498 1820 1504
rect 2148 1465 2176 2746
rect 2134 1456 2190 1465
rect 2134 1391 2190 1400
rect 1676 1352 1728 1358
rect 2044 1352 2096 1358
rect 1676 1294 1728 1300
rect 2042 1320 2044 1329
rect 2096 1320 2098 1329
rect 1688 1034 1716 1294
rect 2042 1255 2098 1264
rect 2504 1216 2556 1222
rect 2504 1158 2556 1164
rect 1688 1006 1808 1034
rect 1674 912 1730 921
rect 1584 876 1636 882
rect 1674 847 1676 856
rect 1584 818 1636 824
rect 1728 847 1730 856
rect 1676 818 1728 824
rect 1490 776 1546 785
rect 1490 711 1546 720
rect 1596 474 1624 818
rect 1780 678 1808 1006
rect 2516 950 2544 1158
rect 2976 1018 3004 2746
rect 3056 2576 3108 2582
rect 3056 2518 3108 2524
rect 3068 2310 3096 2518
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 3252 2038 3280 2246
rect 3344 2106 3372 3839
rect 3620 3670 3648 4626
rect 3608 3664 3660 3670
rect 3608 3606 3660 3612
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3332 2100 3384 2106
rect 3332 2042 3384 2048
rect 3240 2032 3292 2038
rect 3240 1974 3292 1980
rect 3424 1896 3476 1902
rect 3424 1838 3476 1844
rect 2964 1012 3016 1018
rect 2964 954 3016 960
rect 2504 944 2556 950
rect 2504 886 2556 892
rect 3436 746 3464 1838
rect 3528 1358 3556 2926
rect 3620 1902 3648 3606
rect 3896 2961 3924 5510
rect 4193 5468 4501 5477
rect 4193 5466 4199 5468
rect 4255 5466 4279 5468
rect 4335 5466 4359 5468
rect 4415 5466 4439 5468
rect 4495 5466 4501 5468
rect 4255 5414 4257 5466
rect 4437 5414 4439 5466
rect 4193 5412 4199 5414
rect 4255 5412 4279 5414
rect 4335 5412 4359 5414
rect 4415 5412 4439 5414
rect 4495 5412 4501 5414
rect 3974 5400 4030 5409
rect 4193 5403 4501 5412
rect 4540 5352 4568 5902
rect 3974 5335 4030 5344
rect 3988 5030 4016 5335
rect 4448 5324 4568 5352
rect 3976 5024 4028 5030
rect 4448 5001 4476 5324
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 3976 4966 4028 4972
rect 4434 4992 4490 5001
rect 3988 3942 4016 4966
rect 4434 4927 4490 4936
rect 4193 4380 4501 4389
rect 4193 4378 4199 4380
rect 4255 4378 4279 4380
rect 4335 4378 4359 4380
rect 4415 4378 4439 4380
rect 4495 4378 4501 4380
rect 4255 4326 4257 4378
rect 4437 4326 4439 4378
rect 4193 4324 4199 4326
rect 4255 4324 4279 4326
rect 4335 4324 4359 4326
rect 4415 4324 4439 4326
rect 4495 4324 4501 4326
rect 4193 4315 4501 4324
rect 3976 3936 4028 3942
rect 4028 3896 4108 3924
rect 3976 3878 4028 3884
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3882 2952 3938 2961
rect 3882 2887 3938 2896
rect 3988 2496 4016 3470
rect 4080 3176 4108 3896
rect 4540 3738 4568 5102
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4250 3632 4306 3641
rect 4250 3567 4252 3576
rect 4304 3567 4306 3576
rect 4252 3538 4304 3544
rect 4193 3292 4501 3301
rect 4193 3290 4199 3292
rect 4255 3290 4279 3292
rect 4335 3290 4359 3292
rect 4415 3290 4439 3292
rect 4495 3290 4501 3292
rect 4255 3238 4257 3290
rect 4437 3238 4439 3290
rect 4193 3236 4199 3238
rect 4255 3236 4279 3238
rect 4335 3236 4359 3238
rect 4415 3236 4439 3238
rect 4495 3236 4501 3238
rect 4193 3227 4501 3236
rect 4080 3148 4200 3176
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3896 2468 4016 2496
rect 3608 1896 3660 1902
rect 3608 1838 3660 1844
rect 3896 1562 3924 2468
rect 3974 2408 4030 2417
rect 3974 2343 4030 2352
rect 3988 1970 4016 2343
rect 3976 1964 4028 1970
rect 3976 1906 4028 1912
rect 3884 1556 3936 1562
rect 3884 1498 3936 1504
rect 3516 1352 3568 1358
rect 3516 1294 3568 1300
rect 3976 1352 4028 1358
rect 4080 1306 4108 2994
rect 4172 2854 4200 3148
rect 4632 3058 4660 6072
rect 4724 5642 4752 11047
rect 4908 10266 4936 20334
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 5080 18896 5132 18902
rect 5078 18864 5080 18873
rect 5132 18864 5134 18873
rect 5078 18799 5134 18808
rect 5080 17128 5132 17134
rect 5080 17070 5132 17076
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 5000 16658 5028 16934
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 4988 16040 5040 16046
rect 4988 15982 5040 15988
rect 5000 14618 5028 15982
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 5000 14074 5028 14418
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 4988 13252 5040 13258
rect 4988 13194 5040 13200
rect 5000 12209 5028 13194
rect 4986 12200 5042 12209
rect 4986 12135 5042 12144
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 5000 9674 5028 12135
rect 4908 9646 5028 9674
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4816 6254 4844 9318
rect 4908 6746 4936 9646
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5000 6866 5028 9522
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4908 6718 5028 6746
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4908 6390 4936 6598
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4896 5772 4948 5778
rect 5000 5760 5028 6718
rect 5092 5914 5120 17070
rect 5184 11694 5212 19790
rect 5368 19446 5396 21354
rect 5460 21010 5488 21422
rect 5724 21412 5776 21418
rect 5644 21372 5724 21400
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 5552 20890 5580 20946
rect 5460 20862 5580 20890
rect 5460 20369 5488 20862
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5446 20360 5502 20369
rect 5446 20295 5502 20304
rect 5460 19854 5488 20295
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 5460 19310 5488 19790
rect 5448 19304 5500 19310
rect 5448 19246 5500 19252
rect 5446 18728 5502 18737
rect 5446 18663 5502 18672
rect 5354 18184 5410 18193
rect 5354 18119 5356 18128
rect 5408 18119 5410 18128
rect 5356 18090 5408 18096
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 5276 13530 5304 17614
rect 5460 16969 5488 18663
rect 5552 18306 5580 20742
rect 5644 19514 5672 21372
rect 6184 21422 6236 21428
rect 7380 21480 7432 21486
rect 7380 21422 7432 21428
rect 5906 21383 5962 21392
rect 5724 21354 5776 21360
rect 5920 21350 5948 21383
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 6092 21344 6144 21350
rect 6092 21286 6144 21292
rect 5816 21140 5868 21146
rect 5816 21082 5868 21088
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5736 19514 5764 20334
rect 5828 20262 5856 21082
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5828 20058 5856 20198
rect 5816 20052 5868 20058
rect 5816 19994 5868 20000
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 5644 19417 5672 19450
rect 5630 19408 5686 19417
rect 5630 19343 5686 19352
rect 5736 19174 5764 19450
rect 5828 19174 5856 19994
rect 5908 19984 5960 19990
rect 5908 19926 5960 19932
rect 5920 19700 5948 19926
rect 6104 19700 6132 21286
rect 6196 20398 6224 21422
rect 7288 21412 7340 21418
rect 7288 21354 7340 21360
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 6472 20482 6500 21286
rect 6552 21140 6604 21146
rect 6552 21082 6604 21088
rect 6288 20466 6500 20482
rect 6276 20460 6500 20466
rect 6328 20454 6500 20460
rect 6276 20402 6328 20408
rect 6184 20392 6236 20398
rect 6184 20334 6236 20340
rect 6182 19952 6238 19961
rect 6182 19887 6238 19896
rect 5920 19672 6132 19700
rect 6000 19372 6052 19378
rect 6104 19360 6132 19672
rect 6052 19332 6132 19360
rect 6000 19314 6052 19320
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 5552 18278 5764 18306
rect 5632 18216 5684 18222
rect 5632 18158 5684 18164
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5446 16960 5502 16969
rect 5446 16895 5502 16904
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 5460 14618 5488 15914
rect 5552 15706 5580 17138
rect 5644 16726 5672 18158
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5630 16280 5686 16289
rect 5630 16215 5632 16224
rect 5684 16215 5686 16224
rect 5632 16186 5684 16192
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5368 13530 5396 14350
rect 5552 14113 5580 14758
rect 5736 14346 5764 18278
rect 5920 18222 5948 18770
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5828 16182 5856 17614
rect 5920 17202 5948 18158
rect 6012 17814 6040 18226
rect 6104 18086 6132 18770
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 6196 16697 6224 19887
rect 6460 19848 6512 19854
rect 6380 19808 6460 19836
rect 6274 19544 6330 19553
rect 6274 19479 6330 19488
rect 6182 16688 6238 16697
rect 6182 16623 6238 16632
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 6092 16040 6144 16046
rect 6144 16000 6224 16028
rect 6092 15982 6144 15988
rect 6196 15366 6224 16000
rect 6288 15609 6316 19479
rect 6380 17678 6408 19808
rect 6460 19790 6512 19796
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 6472 19009 6500 19246
rect 6458 19000 6514 19009
rect 6458 18935 6514 18944
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6472 18426 6500 18702
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 6564 17746 6592 21082
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6748 20777 6776 20878
rect 6734 20768 6790 20777
rect 6734 20703 6790 20712
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6656 19156 6684 20402
rect 6748 19334 6776 20402
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6932 19961 6960 20334
rect 7300 20262 7328 21354
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 6918 19952 6974 19961
rect 6918 19887 6974 19896
rect 6920 19440 6972 19446
rect 6918 19408 6920 19417
rect 6972 19408 6974 19417
rect 6918 19343 6974 19352
rect 6748 19306 6868 19334
rect 6736 19168 6788 19174
rect 6656 19128 6736 19156
rect 6736 19110 6788 19116
rect 6840 18970 6868 19306
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6736 18760 6788 18766
rect 6736 18702 6788 18708
rect 6748 18057 6776 18702
rect 6828 18080 6880 18086
rect 6734 18048 6790 18057
rect 6828 18022 6880 18028
rect 6734 17983 6790 17992
rect 6840 17882 6868 18022
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6472 17202 6500 17614
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6564 16794 6592 17138
rect 6840 16998 6868 17818
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6932 17338 6960 17614
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 7010 16960 7066 16969
rect 7010 16895 7066 16904
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6274 15600 6330 15609
rect 6274 15535 6330 15544
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6196 15201 6224 15302
rect 6182 15192 6238 15201
rect 6182 15127 6238 15136
rect 6092 15088 6144 15094
rect 6092 15030 6144 15036
rect 6104 14929 6132 15030
rect 6090 14920 6146 14929
rect 6090 14855 6146 14864
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 6092 14816 6144 14822
rect 6196 14804 6224 15127
rect 6288 15026 6316 15302
rect 6380 15162 6408 16526
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6472 15570 6500 16050
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6144 14776 6224 14804
rect 6092 14758 6144 14764
rect 5920 14482 5948 14758
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5724 14340 5776 14346
rect 5724 14282 5776 14288
rect 5538 14104 5594 14113
rect 5538 14039 5594 14048
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5184 11014 5212 11154
rect 5172 11008 5224 11014
rect 5368 10985 5396 12718
rect 5460 11762 5488 13126
rect 5552 12306 5580 14039
rect 5736 12986 5764 14282
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 5828 14074 5856 14214
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5552 11234 5580 12242
rect 5630 11384 5686 11393
rect 5630 11319 5686 11328
rect 5460 11206 5580 11234
rect 5172 10950 5224 10956
rect 5354 10976 5410 10985
rect 5354 10911 5410 10920
rect 5354 10704 5410 10713
rect 5354 10639 5356 10648
rect 5408 10639 5410 10648
rect 5356 10610 5408 10616
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5170 9888 5226 9897
rect 5170 9823 5226 9832
rect 5184 9654 5212 9823
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 5276 6497 5304 10542
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5368 9761 5396 10474
rect 5354 9752 5410 9761
rect 5354 9687 5410 9696
rect 5460 9602 5488 11206
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5552 10606 5580 11086
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5368 9574 5488 9602
rect 5368 9450 5396 9574
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5552 9058 5580 10542
rect 5460 9030 5580 9058
rect 5644 9042 5672 11319
rect 5632 9036 5684 9042
rect 5460 8430 5488 9030
rect 5632 8978 5684 8984
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5552 8294 5580 8910
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5460 7954 5488 8026
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5552 7449 5580 7686
rect 5538 7440 5594 7449
rect 5538 7375 5594 7384
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5262 6488 5318 6497
rect 5368 6458 5396 6598
rect 5460 6458 5488 6938
rect 5262 6423 5318 6432
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5644 6225 5672 8978
rect 5736 7342 5764 12922
rect 5828 12442 5856 13262
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5920 11762 5948 13806
rect 6012 12646 6040 14214
rect 6104 13870 6132 14758
rect 6380 14618 6408 14894
rect 6472 14822 6500 15506
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6288 14226 6316 14418
rect 6380 14346 6408 14418
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6366 14240 6422 14249
rect 6288 14198 6366 14226
rect 6366 14175 6422 14184
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6104 13326 6132 13466
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6104 12753 6132 13262
rect 6090 12744 6146 12753
rect 6090 12679 6146 12688
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 6012 12170 6040 12582
rect 6288 12442 6316 13398
rect 6380 13394 6408 14175
rect 6472 13734 6500 14758
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 6458 13560 6514 13569
rect 6458 13495 6514 13504
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6472 13161 6500 13495
rect 6458 13152 6514 13161
rect 6458 13087 6514 13096
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 6012 11694 6040 12106
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6012 11150 6040 11630
rect 6472 11558 6500 12582
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6472 11234 6500 11494
rect 6380 11218 6500 11234
rect 6368 11212 6500 11218
rect 6420 11206 6500 11212
rect 6368 11154 6420 11160
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 5814 10704 5870 10713
rect 5814 10639 5870 10648
rect 5828 9586 5856 10639
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6104 10130 6132 10542
rect 6092 10124 6144 10130
rect 6012 10084 6092 10112
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5814 9344 5870 9353
rect 5814 9279 5870 9288
rect 5828 9042 5856 9279
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5920 8498 5948 9862
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 6012 8294 6040 10084
rect 6092 10066 6144 10072
rect 6196 9674 6224 10542
rect 6104 9646 6224 9674
rect 6000 8288 6052 8294
rect 5814 8256 5870 8265
rect 6000 8230 6052 8236
rect 5814 8191 5870 8200
rect 5828 7546 5856 8191
rect 6000 7948 6052 7954
rect 5920 7908 6000 7936
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5814 7440 5870 7449
rect 5814 7375 5870 7384
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5828 6730 5856 7375
rect 5920 7342 5948 7908
rect 6000 7890 6052 7896
rect 6104 7585 6132 9646
rect 6184 9444 6236 9450
rect 6184 9386 6236 9392
rect 6196 9058 6224 9386
rect 6288 9178 6316 11086
rect 6380 10674 6408 11154
rect 6460 11144 6512 11150
rect 6564 11121 6592 16594
rect 7024 16590 7052 16895
rect 7012 16584 7064 16590
rect 6734 16552 6790 16561
rect 7012 16526 7064 16532
rect 6734 16487 6790 16496
rect 6748 15162 6776 16487
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 7116 14618 7144 15438
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6656 14278 6684 14418
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6656 13308 6684 14214
rect 7024 13326 7052 14350
rect 7208 14074 7236 16390
rect 7300 14929 7328 19246
rect 7392 16726 7420 21422
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7564 20392 7616 20398
rect 7562 20360 7564 20369
rect 7616 20360 7618 20369
rect 7562 20295 7618 20304
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7484 20058 7512 20198
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7562 19000 7618 19009
rect 7562 18935 7618 18944
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7380 16720 7432 16726
rect 7380 16662 7432 16668
rect 7484 16658 7512 17070
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7470 15464 7526 15473
rect 7470 15399 7526 15408
rect 7286 14920 7342 14929
rect 7286 14855 7342 14864
rect 7300 14618 7328 14855
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7196 13728 7248 13734
rect 7116 13688 7196 13716
rect 6736 13320 6788 13326
rect 6656 13280 6736 13308
rect 6736 13262 6788 13268
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6644 13184 6696 13190
rect 6696 13144 6776 13172
rect 6644 13126 6696 13132
rect 6748 12850 6776 13144
rect 6644 12844 6696 12850
rect 6644 12786 6696 12792
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6656 12628 6684 12786
rect 6656 12600 6776 12628
rect 6748 12102 6776 12600
rect 7024 12594 7052 13262
rect 7116 12866 7144 13688
rect 7196 13670 7248 13676
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7208 12986 7236 13262
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7116 12838 7236 12866
rect 7104 12640 7156 12646
rect 7024 12588 7104 12594
rect 7024 12582 7156 12588
rect 7024 12566 7144 12582
rect 7010 12472 7066 12481
rect 6828 12436 6880 12442
rect 7116 12442 7144 12566
rect 7010 12407 7066 12416
rect 7104 12436 7156 12442
rect 6828 12378 6880 12384
rect 6840 12238 6868 12378
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 7024 12102 7052 12407
rect 7104 12378 7156 12384
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 7102 12064 7158 12073
rect 7102 11999 7158 12008
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6826 11384 6882 11393
rect 6826 11319 6882 11328
rect 6840 11218 6868 11319
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6460 11086 6512 11092
rect 6550 11112 6606 11121
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6380 9586 6408 9998
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6380 9178 6408 9318
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6196 9030 6316 9058
rect 6288 8838 6316 9030
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6196 8498 6224 8774
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6090 7576 6146 7585
rect 6090 7511 6146 7520
rect 6000 7472 6052 7478
rect 5998 7440 6000 7449
rect 6052 7440 6054 7449
rect 5998 7375 6054 7384
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 6196 7256 6224 8230
rect 6380 8022 6408 8910
rect 6368 8016 6420 8022
rect 6368 7958 6420 7964
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6012 7228 6224 7256
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 6012 6338 6040 7228
rect 6182 7168 6238 7177
rect 6182 7103 6238 7112
rect 6196 6934 6224 7103
rect 6184 6928 6236 6934
rect 6184 6870 6236 6876
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 5828 6310 6040 6338
rect 5630 6216 5686 6225
rect 5630 6151 5632 6160
rect 5684 6151 5686 6160
rect 5632 6122 5684 6128
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5184 5914 5212 6054
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 4948 5732 5028 5760
rect 5540 5772 5592 5778
rect 4896 5714 4948 5720
rect 5540 5714 5592 5720
rect 5552 5681 5580 5714
rect 5538 5672 5594 5681
rect 4712 5636 4764 5642
rect 5538 5607 5594 5616
rect 4712 5578 4764 5584
rect 5172 5568 5224 5574
rect 5078 5536 5134 5545
rect 4908 5494 5078 5522
rect 4908 4622 4936 5494
rect 5172 5510 5224 5516
rect 5078 5471 5134 5480
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4896 4616 4948 4622
rect 4710 4584 4766 4593
rect 4896 4558 4948 4564
rect 4710 4519 4766 4528
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4540 2446 4568 2790
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4193 2204 4501 2213
rect 4193 2202 4199 2204
rect 4255 2202 4279 2204
rect 4335 2202 4359 2204
rect 4415 2202 4439 2204
rect 4495 2202 4501 2204
rect 4255 2150 4257 2202
rect 4437 2150 4439 2202
rect 4193 2148 4199 2150
rect 4255 2148 4279 2150
rect 4335 2148 4359 2150
rect 4415 2148 4439 2150
rect 4495 2148 4501 2150
rect 4193 2139 4501 2148
rect 4540 1562 4568 2382
rect 4528 1556 4580 1562
rect 4528 1498 4580 1504
rect 4724 1358 4752 4519
rect 5000 4146 5028 5306
rect 5184 5001 5212 5510
rect 5448 5024 5500 5030
rect 5170 4992 5226 5001
rect 5448 4966 5500 4972
rect 5170 4927 5226 4936
rect 5078 4720 5134 4729
rect 5460 4706 5488 4966
rect 5460 4678 5580 4706
rect 5078 4655 5134 4664
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4802 4040 4858 4049
rect 4802 3975 4858 3984
rect 4028 1300 4108 1306
rect 3976 1294 4108 1300
rect 4712 1352 4764 1358
rect 4712 1294 4764 1300
rect 3988 1278 4108 1294
rect 4193 1116 4501 1125
rect 4193 1114 4199 1116
rect 4255 1114 4279 1116
rect 4335 1114 4359 1116
rect 4415 1114 4439 1116
rect 4495 1114 4501 1116
rect 4255 1062 4257 1114
rect 4437 1062 4439 1114
rect 4193 1060 4199 1062
rect 4255 1060 4279 1062
rect 4335 1060 4359 1062
rect 4415 1060 4439 1062
rect 4495 1060 4501 1062
rect 4193 1051 4501 1060
rect 4816 1018 4844 3975
rect 5092 2514 5120 4655
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5276 3194 5304 4558
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 4988 2372 5040 2378
rect 4988 2314 5040 2320
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 4804 1012 4856 1018
rect 4804 954 4856 960
rect 4908 882 4936 2246
rect 4896 876 4948 882
rect 4896 818 4948 824
rect 4712 808 4764 814
rect 4712 750 4764 756
rect 3424 740 3476 746
rect 3424 682 3476 688
rect 1768 672 1820 678
rect 1768 614 1820 620
rect 2688 672 2740 678
rect 2688 614 2740 620
rect 1584 468 1636 474
rect 1584 410 1636 416
rect 2700 338 2728 614
rect 2688 332 2740 338
rect 2688 274 2740 280
rect 4724 66 4752 750
rect 4804 672 4856 678
rect 4896 672 4948 678
rect 4804 614 4856 620
rect 4894 640 4896 649
rect 4948 640 4950 649
rect 4816 241 4844 614
rect 4894 575 4950 584
rect 4802 232 4858 241
rect 5000 202 5028 2314
rect 5080 1216 5132 1222
rect 5080 1158 5132 1164
rect 5092 202 5120 1158
rect 5184 1018 5212 2926
rect 5264 2032 5316 2038
rect 5264 1974 5316 1980
rect 5172 1012 5224 1018
rect 5172 954 5224 960
rect 5276 814 5304 1974
rect 5368 814 5396 4150
rect 5552 4146 5580 4678
rect 5644 4282 5672 6122
rect 5828 4690 5856 6310
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5828 4486 5856 4626
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3738 5580 3878
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5828 3534 5856 4014
rect 5632 3528 5684 3534
rect 5630 3496 5632 3505
rect 5816 3528 5868 3534
rect 5684 3496 5686 3505
rect 5816 3470 5868 3476
rect 5630 3431 5686 3440
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5460 3126 5488 3334
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5552 2106 5580 2790
rect 5736 2650 5764 2790
rect 5828 2650 5856 3470
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5540 2100 5592 2106
rect 5540 2042 5592 2048
rect 5828 1902 5856 2586
rect 5920 1902 5948 6190
rect 6104 5846 6132 6802
rect 6092 5840 6144 5846
rect 6092 5782 6144 5788
rect 6196 5681 6224 6870
rect 6288 5914 6316 7346
rect 6380 5914 6408 7822
rect 6472 7002 6500 11086
rect 6550 11047 6606 11056
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6564 10198 6592 10950
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 6564 9353 6592 10134
rect 6644 10056 6696 10062
rect 6828 10056 6880 10062
rect 6696 10004 6776 10010
rect 6644 9998 6776 10004
rect 6828 9998 6880 10004
rect 6656 9982 6776 9998
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6656 9625 6684 9658
rect 6642 9616 6698 9625
rect 6642 9551 6698 9560
rect 6550 9344 6606 9353
rect 6550 9279 6606 9288
rect 6564 8294 6592 9279
rect 6656 9042 6684 9551
rect 6644 9036 6696 9042
rect 6748 9024 6776 9982
rect 6840 9722 6868 9998
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6932 9602 6960 11494
rect 7116 10690 7144 11999
rect 7024 10662 7144 10690
rect 7024 9897 7052 10662
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 7010 9888 7066 9897
rect 7010 9823 7066 9832
rect 7012 9716 7064 9722
rect 7116 9674 7144 10474
rect 7064 9664 7144 9674
rect 7012 9658 7144 9664
rect 7024 9646 7144 9658
rect 6840 9574 6960 9602
rect 6840 9518 6868 9574
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6748 8996 6868 9024
rect 6644 8978 6696 8984
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6550 7712 6606 7721
rect 6550 7647 6606 7656
rect 6564 7410 6592 7647
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6656 7342 6684 7822
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6472 6322 6500 6734
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6564 6118 6592 7142
rect 6656 6798 6684 7278
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6748 6322 6776 8842
rect 6840 8276 6868 8996
rect 6932 8634 6960 9454
rect 7116 9382 7144 9646
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7208 9178 7236 12838
rect 7300 11898 7328 14350
rect 7392 13530 7420 14350
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7484 13410 7512 15399
rect 7576 14414 7604 18935
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7392 13382 7512 13410
rect 7392 12617 7420 13382
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7484 12986 7512 13262
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7470 12744 7526 12753
rect 7470 12679 7526 12688
rect 7484 12646 7512 12679
rect 7472 12640 7524 12646
rect 7378 12608 7434 12617
rect 7472 12582 7524 12588
rect 7378 12543 7434 12552
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7576 11778 7604 13806
rect 7668 12209 7696 20742
rect 7654 12200 7710 12209
rect 7654 12135 7710 12144
rect 7392 11750 7604 11778
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7116 9058 7144 9114
rect 7012 9036 7064 9042
rect 7116 9030 7236 9058
rect 7012 8978 7064 8984
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 7024 8498 7052 8978
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7012 8288 7064 8294
rect 6840 8248 7012 8276
rect 7012 8230 7064 8236
rect 6918 7984 6974 7993
rect 7116 7954 7144 8774
rect 6918 7919 6974 7928
rect 7104 7948 7156 7954
rect 6932 7886 6960 7919
rect 7104 7890 7156 7896
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 7010 7848 7066 7857
rect 6840 7698 6868 7822
rect 7010 7783 7066 7792
rect 6840 7670 6960 7698
rect 6826 7576 6882 7585
rect 6826 7511 6828 7520
rect 6880 7511 6882 7520
rect 6828 7482 6880 7488
rect 6932 7206 6960 7670
rect 7024 7546 7052 7783
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7010 7440 7066 7449
rect 7010 7375 7066 7384
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6932 7002 6960 7142
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6918 6896 6974 6905
rect 6918 6831 6974 6840
rect 6932 6798 6960 6831
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6920 6248 6972 6254
rect 7024 6236 7052 7375
rect 7102 7032 7158 7041
rect 7102 6967 7158 6976
rect 6972 6208 7052 6236
rect 6920 6190 6972 6196
rect 6552 6112 6604 6118
rect 6736 6112 6788 6118
rect 6552 6054 6604 6060
rect 6734 6080 6736 6089
rect 6788 6080 6790 6089
rect 6734 6015 6790 6024
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6472 5778 6500 5850
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 6736 5704 6788 5710
rect 6182 5672 6238 5681
rect 6920 5704 6972 5710
rect 6736 5646 6788 5652
rect 6840 5664 6920 5692
rect 6182 5607 6238 5616
rect 6460 5636 6512 5642
rect 6196 4672 6224 5607
rect 6460 5578 6512 5584
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6288 4826 6316 5170
rect 6472 4865 6500 5578
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6458 4856 6514 4865
rect 6276 4820 6328 4826
rect 6458 4791 6514 4800
rect 6276 4762 6328 4768
rect 6104 4644 6224 4672
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6012 3942 6040 4558
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6012 3670 6040 3878
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 6012 2514 6040 2994
rect 6104 2582 6132 4644
rect 6460 4616 6512 4622
rect 6564 4604 6592 5306
rect 6512 4576 6592 4604
rect 6460 4558 6512 4564
rect 6184 3596 6236 3602
rect 6184 3538 6236 3544
rect 6092 2576 6144 2582
rect 6092 2518 6144 2524
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 5998 2408 6054 2417
rect 5998 2343 6000 2352
rect 6052 2343 6054 2352
rect 6000 2314 6052 2320
rect 6196 1970 6224 3538
rect 6472 2514 6500 4558
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6564 3602 6592 3674
rect 6656 3602 6684 5510
rect 6748 5273 6776 5646
rect 6840 5370 6868 5664
rect 6920 5646 6972 5652
rect 6920 5568 6972 5574
rect 6918 5536 6920 5545
rect 6972 5536 6974 5545
rect 6918 5471 6974 5480
rect 7024 5370 7052 5714
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6734 5264 6790 5273
rect 7024 5250 7052 5306
rect 6734 5199 6736 5208
rect 6788 5199 6790 5208
rect 6840 5222 7052 5250
rect 6736 5170 6788 5176
rect 6840 4282 6868 5222
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6932 4826 6960 4966
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6932 2854 6960 4762
rect 7116 4706 7144 6967
rect 7208 5386 7236 9030
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7300 8673 7328 8978
rect 7286 8664 7342 8673
rect 7286 8599 7342 8608
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7300 5778 7328 8434
rect 7392 5914 7420 11750
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7484 8974 7512 11154
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7576 9908 7604 10474
rect 7668 10130 7696 11086
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7656 9920 7708 9926
rect 7576 9880 7656 9908
rect 7656 9862 7708 9868
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7576 9217 7604 9386
rect 7562 9208 7618 9217
rect 7562 9143 7618 9152
rect 7576 9042 7604 9143
rect 7668 9042 7696 9862
rect 7760 9761 7788 21898
rect 8312 21542 8616 21570
rect 9140 21554 9168 22170
rect 15936 22160 15988 22166
rect 15936 22102 15988 22108
rect 10508 22092 10560 22098
rect 10508 22034 10560 22040
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 8312 21486 8340 21542
rect 8300 21480 8352 21486
rect 8300 21422 8352 21428
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 7988 21244 8296 21253
rect 7988 21242 7994 21244
rect 8050 21242 8074 21244
rect 8130 21242 8154 21244
rect 8210 21242 8234 21244
rect 8290 21242 8296 21244
rect 8050 21190 8052 21242
rect 8232 21190 8234 21242
rect 7988 21188 7994 21190
rect 8050 21188 8074 21190
rect 8130 21188 8154 21190
rect 8210 21188 8234 21190
rect 8290 21188 8296 21190
rect 7988 21179 8296 21188
rect 8404 21026 8432 21422
rect 8404 20998 8524 21026
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 7840 20800 7892 20806
rect 7840 20742 7892 20748
rect 7852 20369 7880 20742
rect 7838 20360 7894 20369
rect 7838 20295 7894 20304
rect 7988 20156 8296 20165
rect 7988 20154 7994 20156
rect 8050 20154 8074 20156
rect 8130 20154 8154 20156
rect 8210 20154 8234 20156
rect 8290 20154 8296 20156
rect 8050 20102 8052 20154
rect 8232 20102 8234 20154
rect 7988 20100 7994 20102
rect 8050 20100 8074 20102
rect 8130 20100 8154 20102
rect 8210 20100 8234 20102
rect 8290 20100 8296 20102
rect 7988 20091 8296 20100
rect 8404 19990 8432 20878
rect 8496 20806 8524 20998
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8392 19984 8444 19990
rect 8392 19926 8444 19932
rect 8496 19854 8524 20742
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8312 19514 8340 19654
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 7840 19236 7892 19242
rect 7840 19178 7892 19184
rect 7852 19145 7880 19178
rect 7838 19136 7894 19145
rect 7838 19071 7894 19080
rect 7852 18737 7880 19071
rect 7988 19068 8296 19077
rect 7988 19066 7994 19068
rect 8050 19066 8074 19068
rect 8130 19066 8154 19068
rect 8210 19066 8234 19068
rect 8290 19066 8296 19068
rect 8050 19014 8052 19066
rect 8232 19014 8234 19066
rect 7988 19012 7994 19014
rect 8050 19012 8074 19014
rect 8130 19012 8154 19014
rect 8210 19012 8234 19014
rect 8290 19012 8296 19014
rect 7988 19003 8296 19012
rect 7838 18728 7894 18737
rect 8404 18698 8432 19790
rect 8496 19242 8524 19790
rect 8588 19530 8616 21542
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 8680 21350 8708 21490
rect 9402 21448 9458 21457
rect 9402 21383 9458 21392
rect 8668 21344 8720 21350
rect 8720 21304 8800 21332
rect 8668 21286 8720 21292
rect 8772 21010 8800 21304
rect 8942 21040 8998 21049
rect 8760 21004 8812 21010
rect 8942 20975 8998 20984
rect 9128 21004 9180 21010
rect 8760 20946 8812 20952
rect 8956 20942 8984 20975
rect 9128 20946 9180 20952
rect 8668 20936 8720 20942
rect 8668 20878 8720 20884
rect 8944 20936 8996 20942
rect 8944 20878 8996 20884
rect 9036 20936 9088 20942
rect 9036 20878 9088 20884
rect 8680 19718 8708 20878
rect 9048 20788 9076 20878
rect 8772 20760 9076 20788
rect 8772 20398 8800 20760
rect 8942 20632 8998 20641
rect 9140 20602 9168 20946
rect 8942 20567 8998 20576
rect 9128 20596 9180 20602
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8850 20360 8906 20369
rect 8668 19712 8720 19718
rect 8772 19700 8800 20334
rect 8850 20295 8906 20304
rect 8864 19836 8892 20295
rect 8956 19938 8984 20567
rect 9128 20538 9180 20544
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 8956 19922 9076 19938
rect 8956 19916 9088 19922
rect 8956 19910 9036 19916
rect 9036 19858 9088 19864
rect 8944 19848 8996 19854
rect 8864 19808 8944 19836
rect 9140 19802 9168 20198
rect 8944 19790 8996 19796
rect 9048 19774 9168 19802
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 8772 19672 8984 19700
rect 8668 19654 8720 19660
rect 8588 19502 8892 19530
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8484 19236 8536 19242
rect 8484 19178 8536 19184
rect 8482 19136 8538 19145
rect 8482 19071 8538 19080
rect 8496 18766 8524 19071
rect 8588 18902 8616 19314
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8576 18896 8628 18902
rect 8576 18838 8628 18844
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 7838 18663 7894 18672
rect 8392 18692 8444 18698
rect 8392 18634 8444 18640
rect 8588 18601 8616 18702
rect 8574 18592 8630 18601
rect 8574 18527 8630 18536
rect 8208 18352 8260 18358
rect 8206 18320 8208 18329
rect 8260 18320 8262 18329
rect 8206 18255 8262 18264
rect 8482 18320 8538 18329
rect 8482 18255 8538 18264
rect 8392 18148 8444 18154
rect 8392 18090 8444 18096
rect 7988 17980 8296 17989
rect 7988 17978 7994 17980
rect 8050 17978 8074 17980
rect 8130 17978 8154 17980
rect 8210 17978 8234 17980
rect 8290 17978 8296 17980
rect 8050 17926 8052 17978
rect 8232 17926 8234 17978
rect 7988 17924 7994 17926
rect 8050 17924 8074 17926
rect 8130 17924 8154 17926
rect 8210 17924 8234 17926
rect 8290 17924 8296 17926
rect 7988 17915 8296 17924
rect 8404 17513 8432 18090
rect 8390 17504 8446 17513
rect 8390 17439 8446 17448
rect 8496 17338 8524 18255
rect 8576 18216 8628 18222
rect 8680 18204 8708 19246
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8628 18176 8708 18204
rect 8576 18158 8628 18164
rect 8680 17678 8708 18176
rect 8668 17672 8720 17678
rect 8772 17649 8800 18770
rect 8668 17614 8720 17620
rect 8758 17640 8814 17649
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8390 17232 8446 17241
rect 8680 17202 8708 17614
rect 8758 17575 8814 17584
rect 8390 17167 8392 17176
rect 8444 17167 8446 17176
rect 8668 17196 8720 17202
rect 8392 17138 8444 17144
rect 8668 17138 8720 17144
rect 8482 17096 8538 17105
rect 8482 17031 8538 17040
rect 7988 16892 8296 16901
rect 7988 16890 7994 16892
rect 8050 16890 8074 16892
rect 8130 16890 8154 16892
rect 8210 16890 8234 16892
rect 8290 16890 8296 16892
rect 8050 16838 8052 16890
rect 8232 16838 8234 16890
rect 7988 16836 7994 16838
rect 8050 16836 8074 16838
rect 8130 16836 8154 16838
rect 8210 16836 8234 16838
rect 8290 16836 8296 16838
rect 7988 16827 8296 16836
rect 7840 16720 7892 16726
rect 7840 16662 7892 16668
rect 7852 13025 7880 16662
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 8128 16250 8156 16526
rect 8496 16522 8524 17031
rect 8864 16674 8892 19502
rect 8956 19378 8984 19672
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8956 18601 8984 19314
rect 9048 19258 9076 19774
rect 9232 19417 9260 19790
rect 9218 19408 9274 19417
rect 9218 19343 9274 19352
rect 9416 19310 9444 21383
rect 9600 20806 9628 21490
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9404 19304 9456 19310
rect 9048 19230 9352 19258
rect 9404 19246 9456 19252
rect 9600 19258 9628 19450
rect 9678 19272 9734 19281
rect 9600 19230 9678 19258
rect 9048 18834 9076 19230
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9036 18828 9088 18834
rect 9036 18770 9088 18776
rect 8942 18592 8998 18601
rect 8942 18527 8998 18536
rect 8942 18320 8998 18329
rect 8998 18290 9076 18306
rect 8998 18284 9088 18290
rect 8998 18278 9036 18284
rect 8942 18255 8998 18264
rect 9036 18226 9088 18232
rect 8942 18184 8998 18193
rect 8942 18119 8998 18128
rect 8956 16810 8984 18119
rect 9036 18080 9088 18086
rect 9140 18068 9168 19110
rect 9324 18850 9352 19230
rect 9678 19207 9734 19216
rect 9678 19136 9734 19145
rect 9784 19122 9812 21422
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9734 19094 9812 19122
rect 9862 19136 9918 19145
rect 9678 19071 9734 19080
rect 9862 19071 9918 19080
rect 9324 18822 9536 18850
rect 9508 18766 9536 18822
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9416 18630 9444 18702
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 9088 18040 9168 18068
rect 9036 18022 9088 18028
rect 9036 17672 9088 17678
rect 9140 17660 9168 18040
rect 9088 17632 9168 17660
rect 9036 17614 9088 17620
rect 9048 17202 9076 17614
rect 9126 17504 9182 17513
rect 9126 17439 9182 17448
rect 9140 17202 9168 17439
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 8956 16782 9168 16810
rect 8668 16652 8720 16658
rect 8864 16646 9076 16674
rect 8668 16594 8720 16600
rect 8484 16516 8536 16522
rect 8484 16458 8536 16464
rect 8116 16244 8168 16250
rect 8496 16232 8524 16458
rect 8496 16204 8616 16232
rect 8116 16186 8168 16192
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 7988 15804 8296 15813
rect 7988 15802 7994 15804
rect 8050 15802 8074 15804
rect 8130 15802 8154 15804
rect 8210 15802 8234 15804
rect 8290 15802 8296 15804
rect 8050 15750 8052 15802
rect 8232 15750 8234 15802
rect 7988 15748 7994 15750
rect 8050 15748 8074 15750
rect 8130 15748 8154 15750
rect 8210 15748 8234 15750
rect 8290 15748 8296 15750
rect 7988 15739 8296 15748
rect 8298 15600 8354 15609
rect 8298 15535 8300 15544
rect 8352 15535 8354 15544
rect 8300 15506 8352 15512
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8220 15201 8248 15438
rect 8206 15192 8262 15201
rect 8206 15127 8262 15136
rect 8220 15026 8248 15127
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8496 14929 8524 16050
rect 8482 14920 8538 14929
rect 8482 14855 8538 14864
rect 7988 14716 8296 14725
rect 7988 14714 7994 14716
rect 8050 14714 8074 14716
rect 8130 14714 8154 14716
rect 8210 14714 8234 14716
rect 8290 14714 8296 14716
rect 8050 14662 8052 14714
rect 8232 14662 8234 14714
rect 7988 14660 7994 14662
rect 8050 14660 8074 14662
rect 8130 14660 8154 14662
rect 8210 14660 8234 14662
rect 8290 14660 8296 14662
rect 7988 14651 8296 14660
rect 8392 14340 8444 14346
rect 8392 14282 8444 14288
rect 7988 13628 8296 13637
rect 7988 13626 7994 13628
rect 8050 13626 8074 13628
rect 8130 13626 8154 13628
rect 8210 13626 8234 13628
rect 8290 13626 8296 13628
rect 8050 13574 8052 13626
rect 8232 13574 8234 13626
rect 7988 13572 7994 13574
rect 8050 13572 8074 13574
rect 8130 13572 8154 13574
rect 8210 13572 8234 13574
rect 8290 13572 8296 13574
rect 7988 13563 8296 13572
rect 8404 13258 8432 14282
rect 8588 14249 8616 16204
rect 8680 16046 8708 16594
rect 8944 16584 8996 16590
rect 9048 16561 9076 16646
rect 8944 16526 8996 16532
rect 9034 16552 9090 16561
rect 8956 16046 8984 16526
rect 9034 16487 9090 16496
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 8680 15570 8708 15982
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8956 15502 8984 15982
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8956 14822 8984 15438
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8956 14618 8984 14758
rect 9048 14618 9076 16487
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 9140 14498 9168 16782
rect 9218 16688 9274 16697
rect 9218 16623 9220 16632
rect 9272 16623 9274 16632
rect 9220 16594 9272 16600
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 9232 16114 9260 16390
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9324 15722 9352 18158
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9048 14470 9168 14498
rect 9232 15694 9352 15722
rect 8574 14240 8630 14249
rect 8574 14175 8630 14184
rect 8588 13682 8616 14175
rect 8944 13932 8996 13938
rect 8864 13892 8944 13920
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8588 13654 8708 13682
rect 8680 13530 8708 13654
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 7932 13184 7984 13190
rect 7930 13152 7932 13161
rect 7984 13152 7986 13161
rect 7930 13087 7986 13096
rect 7838 13016 7894 13025
rect 7838 12951 7894 12960
rect 7840 12912 7892 12918
rect 7840 12854 7892 12860
rect 7852 11762 7880 12854
rect 7988 12540 8296 12549
rect 7988 12538 7994 12540
rect 8050 12538 8074 12540
rect 8130 12538 8154 12540
rect 8210 12538 8234 12540
rect 8290 12538 8296 12540
rect 8050 12486 8052 12538
rect 8232 12486 8234 12538
rect 7988 12484 7994 12486
rect 8050 12484 8074 12486
rect 8130 12484 8154 12486
rect 8210 12484 8234 12486
rect 8290 12484 8296 12486
rect 7988 12475 8296 12484
rect 8588 12374 8616 13466
rect 8576 12368 8628 12374
rect 8576 12310 8628 12316
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11937 8524 12038
rect 8482 11928 8538 11937
rect 8482 11863 8538 11872
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 7852 11082 7880 11562
rect 7988 11452 8296 11461
rect 7988 11450 7994 11452
rect 8050 11450 8074 11452
rect 8130 11450 8154 11452
rect 8210 11450 8234 11452
rect 8290 11450 8296 11452
rect 8050 11398 8052 11450
rect 8232 11398 8234 11450
rect 7988 11396 7994 11398
rect 8050 11396 8074 11398
rect 8130 11396 8154 11398
rect 8210 11396 8234 11398
rect 8290 11396 8296 11398
rect 7988 11387 8296 11396
rect 8496 11354 8524 11562
rect 8666 11384 8722 11393
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8576 11348 8628 11354
rect 8666 11319 8722 11328
rect 8576 11290 8628 11296
rect 8404 11234 8432 11290
rect 8588 11234 8616 11290
rect 8404 11206 8616 11234
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7746 9752 7802 9761
rect 7746 9687 7802 9696
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7760 9178 7788 9318
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7852 9058 7880 10610
rect 8312 10538 8340 11086
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 7988 10364 8296 10373
rect 7988 10362 7994 10364
rect 8050 10362 8074 10364
rect 8130 10362 8154 10364
rect 8210 10362 8234 10364
rect 8290 10362 8296 10364
rect 8050 10310 8052 10362
rect 8232 10310 8234 10362
rect 7988 10308 7994 10310
rect 8050 10308 8074 10310
rect 8130 10308 8154 10310
rect 8210 10308 8234 10310
rect 8290 10308 8296 10310
rect 7988 10299 8296 10308
rect 8404 10146 8432 11206
rect 8482 10976 8538 10985
rect 8482 10911 8538 10920
rect 8496 10554 8524 10911
rect 8680 10606 8708 11319
rect 8772 11121 8800 13806
rect 8864 12782 8892 13892
rect 8944 13874 8996 13880
rect 8942 13696 8998 13705
rect 8942 13631 8998 13640
rect 8956 13530 8984 13631
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8852 12640 8904 12646
rect 8850 12608 8852 12617
rect 8904 12608 8906 12617
rect 8850 12543 8906 12552
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8864 11150 8892 12174
rect 9048 11762 9076 14470
rect 9126 14376 9182 14385
rect 9126 14311 9182 14320
rect 9140 13734 9168 14311
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9232 13530 9260 15694
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9324 14618 9352 15438
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9324 13938 9352 14418
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9324 13394 9352 13874
rect 9416 13530 9444 17614
rect 9600 17513 9628 18022
rect 9586 17504 9642 17513
rect 9586 17439 9642 17448
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 16590 9536 16934
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9494 16144 9550 16153
rect 9494 16079 9550 16088
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9220 13252 9272 13258
rect 9220 13194 9272 13200
rect 9232 12646 9260 13194
rect 9324 12986 9352 13330
rect 9508 13326 9536 16079
rect 9600 13530 9628 17138
rect 9692 16590 9720 19071
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9784 14906 9812 18362
rect 9876 17542 9904 19071
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9968 16794 9996 19178
rect 10152 17066 10180 21966
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 10416 21888 10468 21894
rect 10416 21830 10468 21836
rect 10232 21344 10284 21350
rect 10232 21286 10284 21292
rect 10244 21146 10272 21286
rect 10232 21140 10284 21146
rect 10232 21082 10284 21088
rect 10336 21010 10364 21830
rect 10428 21078 10456 21830
rect 10416 21072 10468 21078
rect 10416 21014 10468 21020
rect 10324 21004 10376 21010
rect 10324 20946 10376 20952
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10244 19514 10272 20402
rect 10520 20346 10548 22034
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 10428 20318 10548 20346
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 10428 18902 10456 20318
rect 10508 20256 10560 20262
rect 10508 20198 10560 20204
rect 10416 18896 10468 18902
rect 10416 18838 10468 18844
rect 10520 18850 10548 20198
rect 10612 19990 10640 21966
rect 11428 21956 11480 21962
rect 11428 21898 11480 21904
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 10874 20904 10930 20913
rect 10874 20839 10930 20848
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10600 19984 10652 19990
rect 10600 19926 10652 19932
rect 10704 19514 10732 20334
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10428 18737 10456 18838
rect 10520 18822 10640 18850
rect 10508 18760 10560 18766
rect 10414 18728 10470 18737
rect 10508 18702 10560 18708
rect 10414 18663 10470 18672
rect 10324 17740 10376 17746
rect 10324 17682 10376 17688
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10140 17060 10192 17066
rect 10140 17002 10192 17008
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9692 14618 9720 14894
rect 9784 14878 9904 14906
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9678 14104 9734 14113
rect 9784 14074 9812 14758
rect 9678 14039 9734 14048
rect 9772 14068 9824 14074
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9692 13394 9720 14039
rect 9772 14010 9824 14016
rect 9876 13802 9904 14878
rect 9968 14618 9996 16594
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10060 14618 10088 16526
rect 10138 15192 10194 15201
rect 10138 15127 10194 15136
rect 10152 15094 10180 15127
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 10244 15026 10272 17274
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10244 14482 10272 14962
rect 10336 14482 10364 17682
rect 10520 17338 10548 18702
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10428 16289 10456 16390
rect 10414 16280 10470 16289
rect 10414 16215 10470 16224
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10428 15706 10456 15846
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10520 15366 10548 16186
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10428 15065 10456 15302
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 10414 15056 10470 15065
rect 10414 14991 10470 15000
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9680 13388 9732 13394
rect 9864 13388 9916 13394
rect 9680 13330 9732 13336
rect 9784 13348 9864 13376
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9680 13184 9732 13190
rect 9678 13152 9680 13161
rect 9732 13152 9734 13161
rect 9678 13087 9734 13096
rect 9784 13002 9812 13348
rect 9864 13330 9916 13336
rect 9968 13240 9996 14418
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9508 12974 9812 13002
rect 9876 13212 9996 13240
rect 9508 12918 9536 12974
rect 9496 12912 9548 12918
rect 9496 12854 9548 12860
rect 9772 12844 9824 12850
rect 9680 12826 9732 12832
rect 9588 12776 9640 12782
rect 9494 12744 9550 12753
rect 9772 12786 9824 12792
rect 9680 12768 9732 12774
rect 9588 12718 9640 12724
rect 9494 12679 9550 12688
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9324 12306 9352 12582
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8852 11144 8904 11150
rect 8758 11112 8814 11121
rect 8852 11086 8904 11092
rect 8758 11047 8814 11056
rect 8864 10674 8892 11086
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8668 10600 8720 10606
rect 8496 10526 8616 10554
rect 8720 10560 8800 10588
rect 8668 10542 8720 10548
rect 8588 10441 8616 10526
rect 8574 10432 8630 10441
rect 8574 10367 8630 10376
rect 8404 10118 8524 10146
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 7988 9276 8296 9285
rect 7988 9274 7994 9276
rect 8050 9274 8074 9276
rect 8130 9274 8154 9276
rect 8210 9274 8234 9276
rect 8290 9274 8296 9276
rect 8050 9222 8052 9274
rect 8232 9222 8234 9274
rect 7988 9220 7994 9222
rect 8050 9220 8074 9222
rect 8130 9220 8154 9222
rect 8210 9220 8234 9222
rect 8290 9220 8296 9222
rect 7988 9211 8296 9220
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7656 9036 7708 9042
rect 7852 9030 8156 9058
rect 7656 8978 7708 8984
rect 8128 8974 8156 9030
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7656 8900 7708 8906
rect 7656 8842 7708 8848
rect 7562 8392 7618 8401
rect 7562 8327 7618 8336
rect 7576 7478 7604 8327
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7668 7290 7696 8842
rect 8404 8634 8432 9998
rect 8496 9518 8524 10118
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7760 7410 7788 8502
rect 8588 8294 8616 10367
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8680 9586 8708 9998
rect 8772 9908 8800 10560
rect 8956 10062 8984 11562
rect 9324 11558 9352 12038
rect 9508 11762 9536 12679
rect 9600 12102 9628 12718
rect 9692 12322 9720 12768
rect 9784 12442 9812 12786
rect 9876 12696 9904 13212
rect 9876 12668 9996 12696
rect 9862 12608 9918 12617
rect 9862 12543 9918 12552
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9770 12336 9826 12345
rect 9692 12294 9770 12322
rect 9770 12271 9826 12280
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9876 11762 9904 12543
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9968 11642 9996 12668
rect 9876 11614 9996 11642
rect 9312 11552 9364 11558
rect 9876 11529 9904 11614
rect 9956 11552 10008 11558
rect 9312 11494 9364 11500
rect 9862 11520 9918 11529
rect 9036 11144 9088 11150
rect 9034 11112 9036 11121
rect 9088 11112 9090 11121
rect 9034 11047 9090 11056
rect 9324 10606 9352 11494
rect 9956 11494 10008 11500
rect 9862 11455 9918 11464
rect 9496 11144 9548 11150
rect 9416 11092 9496 11098
rect 9416 11086 9548 11092
rect 9416 11070 9536 11086
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9048 10266 9076 10542
rect 9220 10464 9272 10470
rect 9218 10432 9220 10441
rect 9272 10432 9274 10441
rect 9218 10367 9274 10376
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 9312 10260 9364 10266
rect 9416 10248 9444 11070
rect 9876 11014 9904 11455
rect 9968 11121 9996 11494
rect 9954 11112 10010 11121
rect 9954 11047 10010 11056
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9586 10840 9642 10849
rect 9586 10775 9642 10784
rect 9600 10724 9628 10775
rect 9600 10696 9720 10724
rect 9692 10266 9720 10696
rect 9968 10674 9996 11047
rect 10060 10674 10088 14214
rect 10152 14074 10180 14282
rect 10244 14278 10272 14418
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10152 11898 10180 13874
rect 10336 13705 10364 14418
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10322 13696 10378 13705
rect 10428 13682 10456 14214
rect 10520 14074 10548 15098
rect 10612 15094 10640 18822
rect 10796 17814 10824 20742
rect 10888 20534 10916 20839
rect 10876 20528 10928 20534
rect 10876 20470 10928 20476
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 10888 18902 10916 20334
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10980 18612 11008 21286
rect 11072 20330 11100 21490
rect 11440 21486 11468 21898
rect 12530 21856 12586 21865
rect 11783 21788 12091 21797
rect 12530 21791 12586 21800
rect 11783 21786 11789 21788
rect 11845 21786 11869 21788
rect 11925 21786 11949 21788
rect 12005 21786 12029 21788
rect 12085 21786 12091 21788
rect 11845 21734 11847 21786
rect 12027 21734 12029 21786
rect 11783 21732 11789 21734
rect 11845 21732 11869 21734
rect 11925 21732 11949 21734
rect 12005 21732 12029 21734
rect 12085 21732 12091 21734
rect 11783 21723 12091 21732
rect 12544 21690 12572 21791
rect 11704 21684 11756 21690
rect 11704 21626 11756 21632
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 11428 21480 11480 21486
rect 11428 21422 11480 21428
rect 11256 21298 11284 21422
rect 11612 21344 11664 21350
rect 11256 21270 11376 21298
rect 11612 21286 11664 21292
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 10888 18584 11008 18612
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10692 15972 10744 15978
rect 10692 15914 10744 15920
rect 10600 15088 10652 15094
rect 10600 15030 10652 15036
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10612 13938 10640 14214
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10704 13802 10732 15914
rect 10796 15881 10824 17002
rect 10888 16794 10916 18584
rect 11072 18426 11100 19314
rect 11164 19174 11192 20878
rect 11244 20392 11296 20398
rect 11348 20346 11376 21270
rect 11428 20936 11480 20942
rect 11428 20878 11480 20884
rect 11440 20806 11468 20878
rect 11428 20800 11480 20806
rect 11428 20742 11480 20748
rect 11426 20496 11482 20505
rect 11426 20431 11482 20440
rect 11296 20340 11376 20346
rect 11244 20334 11376 20340
rect 11256 20318 11376 20334
rect 11348 19922 11376 20318
rect 11336 19916 11388 19922
rect 11336 19858 11388 19864
rect 11242 19816 11298 19825
rect 11242 19751 11298 19760
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11164 18766 11192 19110
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 11256 18306 11284 19751
rect 11348 18834 11376 19858
rect 11440 19174 11468 20431
rect 11624 20262 11652 21286
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11164 18278 11284 18306
rect 10968 18216 11020 18222
rect 10966 18184 10968 18193
rect 11020 18184 11022 18193
rect 10966 18119 11022 18128
rect 10966 18048 11022 18057
rect 10966 17983 11022 17992
rect 10980 17542 11008 17983
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10980 16454 11008 17070
rect 11072 16998 11100 18226
rect 11164 18154 11192 18278
rect 11244 18216 11296 18222
rect 11244 18158 11296 18164
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 11058 16688 11114 16697
rect 11058 16623 11114 16632
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 11072 16114 11100 16623
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 10782 15872 10838 15881
rect 10782 15807 10838 15816
rect 10796 14482 10824 15807
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10428 13654 10732 13682
rect 10322 13631 10378 13640
rect 10230 13560 10286 13569
rect 10230 13495 10286 13504
rect 10244 13394 10272 13495
rect 10336 13394 10364 13631
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10244 11762 10272 13126
rect 10322 13016 10378 13025
rect 10322 12951 10378 12960
rect 10428 12968 10456 13126
rect 10336 12170 10364 12951
rect 10428 12940 10548 12968
rect 10520 12850 10548 12940
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 10612 11218 10640 13126
rect 10704 12220 10732 13654
rect 10796 13394 10824 14418
rect 10888 14346 10916 14894
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 10876 14340 10928 14346
rect 10876 14282 10928 14288
rect 10980 13870 11008 14486
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10782 13152 10838 13161
rect 10782 13087 10838 13096
rect 10796 12782 10824 13087
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10784 12232 10836 12238
rect 10704 12192 10784 12220
rect 10784 12174 10836 12180
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11898 10732 12038
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9864 10464 9916 10470
rect 9784 10424 9864 10452
rect 9364 10220 9444 10248
rect 9680 10260 9732 10266
rect 9312 10202 9364 10208
rect 9680 10202 9732 10208
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 9048 9926 9076 10202
rect 9218 10160 9274 10169
rect 9218 10095 9274 10104
rect 9036 9920 9088 9926
rect 8772 9880 8984 9908
rect 8956 9722 8984 9880
rect 9036 9862 9088 9868
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8680 8673 8708 9318
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8666 8664 8722 8673
rect 8666 8599 8722 8608
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7668 7262 7788 7290
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7470 6488 7526 6497
rect 7470 6423 7526 6432
rect 7484 6322 7512 6423
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7576 5778 7604 7142
rect 7656 6248 7708 6254
rect 7654 6216 7656 6225
rect 7708 6216 7710 6225
rect 7654 6151 7710 6160
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7656 5772 7708 5778
rect 7760 5760 7788 7262
rect 7708 5732 7788 5760
rect 7656 5714 7708 5720
rect 7576 5681 7604 5714
rect 7562 5672 7618 5681
rect 7562 5607 7618 5616
rect 7380 5568 7432 5574
rect 7432 5516 7604 5522
rect 7380 5510 7604 5516
rect 7392 5494 7604 5510
rect 7208 5358 7420 5386
rect 7024 4678 7144 4706
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6932 2650 6960 2790
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 6472 2378 6500 2450
rect 6460 2372 6512 2378
rect 6460 2314 6512 2320
rect 6184 1964 6236 1970
rect 6184 1906 6236 1912
rect 6368 1964 6420 1970
rect 6368 1906 6420 1912
rect 5724 1896 5776 1902
rect 5724 1838 5776 1844
rect 5816 1896 5868 1902
rect 5816 1838 5868 1844
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 5736 1222 5764 1838
rect 5724 1216 5776 1222
rect 5724 1158 5776 1164
rect 5920 814 5948 1838
rect 6380 1290 6408 1906
rect 6472 1358 6500 2314
rect 6840 1426 6868 2450
rect 6932 1562 6960 2586
rect 6920 1556 6972 1562
rect 6920 1498 6972 1504
rect 6828 1420 6880 1426
rect 6828 1362 6880 1368
rect 7024 1358 7052 4678
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7116 3738 7144 4558
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7116 2514 7144 3538
rect 7208 2650 7236 4558
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7300 3602 7328 4422
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7286 3224 7342 3233
rect 7286 3159 7288 3168
rect 7340 3159 7342 3168
rect 7288 3130 7340 3136
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7392 2122 7420 5358
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7484 2446 7512 5170
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7208 2094 7420 2122
rect 7208 1358 7236 2094
rect 7576 1986 7604 5494
rect 7668 4078 7696 5714
rect 7852 5574 7880 8230
rect 7988 8188 8296 8197
rect 7988 8186 7994 8188
rect 8050 8186 8074 8188
rect 8130 8186 8154 8188
rect 8210 8186 8234 8188
rect 8290 8186 8296 8188
rect 8050 8134 8052 8186
rect 8232 8134 8234 8186
rect 7988 8132 7994 8134
rect 8050 8132 8074 8134
rect 8130 8132 8154 8134
rect 8210 8132 8234 8134
rect 8290 8132 8296 8134
rect 7988 8123 8296 8132
rect 8404 8090 8432 8230
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8588 7274 8616 8230
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 7988 7100 8296 7109
rect 7988 7098 7994 7100
rect 8050 7098 8074 7100
rect 8130 7098 8154 7100
rect 8210 7098 8234 7100
rect 8290 7098 8296 7100
rect 8050 7046 8052 7098
rect 8232 7046 8234 7098
rect 7988 7044 7994 7046
rect 8050 7044 8074 7046
rect 8130 7044 8154 7046
rect 8210 7044 8234 7046
rect 8290 7044 8296 7046
rect 7988 7035 8296 7044
rect 8496 6730 8524 7142
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 7944 6390 7972 6598
rect 8312 6458 8340 6598
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8680 6390 8708 8599
rect 8760 8560 8812 8566
rect 8760 8502 8812 8508
rect 8772 6866 8800 8502
rect 8864 8294 8892 8774
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 8668 6384 8720 6390
rect 8668 6326 8720 6332
rect 8484 6180 8536 6186
rect 8484 6122 8536 6128
rect 7988 6012 8296 6021
rect 7988 6010 7994 6012
rect 8050 6010 8074 6012
rect 8130 6010 8154 6012
rect 8210 6010 8234 6012
rect 8290 6010 8296 6012
rect 8050 5958 8052 6010
rect 8232 5958 8234 6010
rect 7988 5956 7994 5958
rect 8050 5956 8074 5958
rect 8130 5956 8154 5958
rect 8210 5956 8234 5958
rect 8290 5956 8296 5958
rect 7988 5947 8296 5956
rect 8496 5914 8524 6122
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7944 5234 7972 5714
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 8036 5098 8064 5646
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7852 4826 7880 4966
rect 7988 4924 8296 4933
rect 7988 4922 7994 4924
rect 8050 4922 8074 4924
rect 8130 4922 8154 4924
rect 8210 4922 8234 4924
rect 8290 4922 8296 4924
rect 8050 4870 8052 4922
rect 8232 4870 8234 4922
rect 7988 4868 7994 4870
rect 8050 4868 8074 4870
rect 8130 4868 8154 4870
rect 8210 4868 8234 4870
rect 8290 4868 8296 4870
rect 7988 4859 8296 4868
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 8404 4146 8432 5646
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8496 4826 8524 5170
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 8496 4010 8524 4762
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 7988 3836 8296 3845
rect 7988 3834 7994 3836
rect 8050 3834 8074 3836
rect 8130 3834 8154 3836
rect 8210 3834 8234 3836
rect 8290 3834 8296 3836
rect 8050 3782 8052 3834
rect 8232 3782 8234 3834
rect 7988 3780 7994 3782
rect 8050 3780 8074 3782
rect 8130 3780 8154 3782
rect 8210 3780 8234 3782
rect 8290 3780 8296 3782
rect 7988 3771 8296 3780
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8128 3194 8156 3538
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7760 2446 7788 2994
rect 7988 2748 8296 2757
rect 7988 2746 7994 2748
rect 8050 2746 8074 2748
rect 8130 2746 8154 2748
rect 8210 2746 8234 2748
rect 8290 2746 8296 2748
rect 8050 2694 8052 2746
rect 8232 2694 8234 2746
rect 7988 2692 7994 2694
rect 8050 2692 8074 2694
rect 8130 2692 8154 2694
rect 8210 2692 8234 2694
rect 8290 2692 8296 2694
rect 7988 2683 8296 2692
rect 8404 2650 8432 3470
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 7748 2440 7800 2446
rect 7852 2417 7880 2450
rect 8208 2440 8260 2446
rect 7748 2382 7800 2388
rect 7838 2408 7894 2417
rect 8208 2382 8260 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 7838 2343 7894 2352
rect 8220 2106 8248 2382
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 7300 1970 7604 1986
rect 7288 1964 7604 1970
rect 7340 1958 7604 1964
rect 7288 1906 7340 1912
rect 8312 1902 8340 2382
rect 8300 1896 8352 1902
rect 8300 1838 8352 1844
rect 8404 1737 8432 2586
rect 8390 1728 8446 1737
rect 7988 1660 8296 1669
rect 8390 1663 8446 1672
rect 7988 1658 7994 1660
rect 8050 1658 8074 1660
rect 8130 1658 8154 1660
rect 8210 1658 8234 1660
rect 8290 1658 8296 1660
rect 8050 1606 8052 1658
rect 8232 1606 8234 1658
rect 7988 1604 7994 1606
rect 8050 1604 8074 1606
rect 8130 1604 8154 1606
rect 8210 1604 8234 1606
rect 8290 1604 8296 1606
rect 7988 1595 8296 1604
rect 6460 1352 6512 1358
rect 6460 1294 6512 1300
rect 7012 1352 7064 1358
rect 7012 1294 7064 1300
rect 7196 1352 7248 1358
rect 7196 1294 7248 1300
rect 6368 1284 6420 1290
rect 6368 1226 6420 1232
rect 7564 1216 7616 1222
rect 6090 1184 6146 1193
rect 7564 1158 7616 1164
rect 6090 1119 6146 1128
rect 6104 950 6132 1119
rect 7576 1018 7604 1158
rect 7564 1012 7616 1018
rect 7564 954 7616 960
rect 6092 944 6144 950
rect 6092 886 6144 892
rect 6644 876 6696 882
rect 6644 818 6696 824
rect 5264 808 5316 814
rect 5264 750 5316 756
rect 5356 808 5408 814
rect 5356 750 5408 756
rect 5908 808 5960 814
rect 5908 750 5960 756
rect 6184 808 6236 814
rect 6184 750 6236 756
rect 5816 672 5868 678
rect 5816 614 5868 620
rect 6000 672 6052 678
rect 6196 649 6224 750
rect 6460 672 6512 678
rect 6000 614 6052 620
rect 6182 640 6238 649
rect 5828 474 5856 614
rect 5816 468 5868 474
rect 5816 410 5868 416
rect 4802 167 4858 176
rect 4988 196 5040 202
rect 4988 138 5040 144
rect 5080 196 5132 202
rect 5080 138 5132 144
rect 6012 66 6040 614
rect 6656 660 6684 818
rect 8496 796 8524 3946
rect 8588 3942 8616 5646
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8588 2514 8616 2994
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8680 1902 8708 6326
rect 8864 5778 8892 8230
rect 8956 6202 8984 9658
rect 9036 9444 9088 9450
rect 9088 9404 9168 9432
rect 9036 9386 9088 9392
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9048 8430 9076 8910
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 9140 8294 9168 9404
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 9048 7342 9076 7890
rect 9128 7880 9180 7886
rect 9126 7848 9128 7857
rect 9180 7848 9182 7857
rect 9126 7783 9182 7792
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 6866 9076 7278
rect 9128 7268 9180 7274
rect 9128 7210 9180 7216
rect 9140 7177 9168 7210
rect 9126 7168 9182 7177
rect 9126 7103 9182 7112
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9048 6322 9076 6802
rect 9126 6760 9182 6769
rect 9126 6695 9182 6704
rect 9140 6458 9168 6695
rect 9232 6458 9260 10095
rect 9324 9586 9352 10202
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 9600 9926 9628 9998
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9324 9042 9352 9522
rect 9508 9178 9536 9522
rect 9784 9518 9812 10424
rect 9864 10406 9916 10412
rect 10612 10130 10640 10950
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10704 9722 10732 10542
rect 10796 10062 10824 12174
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9692 9178 9720 9454
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9784 9058 9812 9454
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9692 9030 9812 9058
rect 10414 9072 10470 9081
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9508 8430 9536 8774
rect 9692 8446 9720 9030
rect 10414 9007 10470 9016
rect 10598 9072 10654 9081
rect 10598 9007 10600 9016
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9680 8440 9732 8446
rect 9496 8424 9548 8430
rect 9784 8430 9812 8910
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9876 8498 9904 8774
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9680 8382 9732 8388
rect 9772 8424 9824 8430
rect 9496 8366 9548 8372
rect 9772 8366 9824 8372
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9324 6746 9352 8298
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9416 7886 9444 8230
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9508 7426 9536 8026
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9416 7410 9536 7426
rect 9404 7404 9536 7410
rect 9456 7398 9536 7404
rect 9404 7346 9456 7352
rect 9508 7002 9536 7398
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9324 6718 9444 6746
rect 9416 6662 9444 6718
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9324 6322 9352 6598
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 8956 6174 9352 6202
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 8772 5098 8800 5306
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8772 4282 8800 5034
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 8864 4622 8892 4966
rect 9048 4622 9076 4966
rect 9232 4826 9260 5306
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8864 4146 8892 4558
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8864 3534 8892 4082
rect 9048 4078 9076 4558
rect 9324 4298 9352 6174
rect 9416 6118 9444 6598
rect 9508 6118 9536 6938
rect 9692 6458 9720 7482
rect 9968 7177 9996 8230
rect 10428 8022 10456 9007
rect 10652 9007 10654 9016
rect 10692 9036 10744 9042
rect 10600 8978 10652 8984
rect 10692 8978 10744 8984
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 10506 7576 10562 7585
rect 10506 7511 10562 7520
rect 9954 7168 10010 7177
rect 9954 7103 10010 7112
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9416 5930 9444 6054
rect 9416 5902 9720 5930
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9416 4690 9444 5578
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9600 5166 9628 5510
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9324 4270 9536 4298
rect 9324 4078 9352 4270
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9416 4078 9444 4150
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9048 3534 9076 4014
rect 9232 3738 9260 4014
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9324 3602 9352 3878
rect 9508 3602 9536 4270
rect 9692 4026 9720 5902
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9784 5234 9812 5510
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9600 3998 9720 4026
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8864 3126 8892 3470
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 8864 2922 8892 3062
rect 9048 2938 9076 3470
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9232 3097 9260 3334
rect 9218 3088 9274 3097
rect 9218 3023 9274 3032
rect 9600 2938 9628 3998
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9692 3058 9720 3878
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 8852 2916 8904 2922
rect 9048 2910 9444 2938
rect 9600 2910 9720 2938
rect 8852 2858 8904 2864
rect 8864 2310 8892 2858
rect 9416 2854 9444 2910
rect 9312 2848 9364 2854
rect 9312 2790 9364 2796
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 8864 1970 8892 2246
rect 8852 1964 8904 1970
rect 8852 1906 8904 1912
rect 8668 1896 8720 1902
rect 8668 1838 8720 1844
rect 8668 1760 8720 1766
rect 8668 1702 8720 1708
rect 8760 1760 8812 1766
rect 8760 1702 8812 1708
rect 8680 1601 8708 1702
rect 8666 1592 8722 1601
rect 8666 1527 8722 1536
rect 8772 1426 8800 1702
rect 8760 1420 8812 1426
rect 8760 1362 8812 1368
rect 8576 808 8628 814
rect 8496 768 8576 796
rect 8576 750 8628 756
rect 8760 740 8812 746
rect 8864 728 8892 1906
rect 8944 1760 8996 1766
rect 8944 1702 8996 1708
rect 8956 1562 8984 1702
rect 8944 1556 8996 1562
rect 8944 1498 8996 1504
rect 9128 1352 9180 1358
rect 9128 1294 9180 1300
rect 9140 1018 9168 1294
rect 9324 1018 9352 2790
rect 9416 1766 9444 2790
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9404 1760 9456 1766
rect 9404 1702 9456 1708
rect 9128 1012 9180 1018
rect 9128 954 9180 960
rect 9312 1012 9364 1018
rect 9312 954 9364 960
rect 8812 700 8892 728
rect 8760 682 8812 688
rect 9416 678 9444 1702
rect 9508 1426 9536 2450
rect 9692 2446 9720 2910
rect 9784 2650 9812 3470
rect 9876 3194 9904 3878
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9968 2530 9996 7103
rect 10520 7002 10548 7511
rect 10612 7206 10640 8978
rect 10704 8294 10732 8978
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10888 8090 10916 13806
rect 11072 13394 11100 16050
rect 11164 14958 11192 18090
rect 11256 17678 11284 18158
rect 11336 18080 11388 18086
rect 11388 18040 11468 18068
rect 11336 18022 11388 18028
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11256 17134 11284 17614
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 11256 16046 11284 17070
rect 11336 16720 11388 16726
rect 11336 16662 11388 16668
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11256 15434 11284 15982
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11256 14958 11284 15370
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11164 13530 11192 14894
rect 11256 14482 11284 14894
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11256 13870 11284 14418
rect 11348 14113 11376 16662
rect 11334 14104 11390 14113
rect 11334 14039 11390 14048
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11244 13728 11296 13734
rect 11296 13688 11376 13716
rect 11244 13670 11296 13676
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 11242 13016 11298 13025
rect 11242 12951 11298 12960
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11058 12200 11114 12209
rect 11058 12135 11114 12144
rect 11072 12102 11100 12135
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10980 10674 11008 12038
rect 11164 11694 11192 12786
rect 11256 12442 11284 12951
rect 11348 12918 11376 13688
rect 11440 13530 11468 18040
rect 11532 17338 11560 18158
rect 11612 18080 11664 18086
rect 11612 18022 11664 18028
rect 11624 17746 11652 18022
rect 11716 17762 11744 21626
rect 15580 21622 15608 21966
rect 15568 21616 15620 21622
rect 14002 21584 14058 21593
rect 15568 21558 15620 21564
rect 14002 21519 14058 21528
rect 13820 21412 13872 21418
rect 13820 21354 13872 21360
rect 12348 21344 12400 21350
rect 12348 21286 12400 21292
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 11783 20700 12091 20709
rect 11783 20698 11789 20700
rect 11845 20698 11869 20700
rect 11925 20698 11949 20700
rect 12005 20698 12029 20700
rect 12085 20698 12091 20700
rect 11845 20646 11847 20698
rect 12027 20646 12029 20698
rect 11783 20644 11789 20646
rect 11845 20644 11869 20646
rect 11925 20644 11949 20646
rect 12005 20644 12029 20646
rect 12085 20644 12091 20646
rect 11783 20635 12091 20644
rect 12072 20392 12124 20398
rect 12072 20334 12124 20340
rect 12084 19990 12112 20334
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 11980 19848 12032 19854
rect 12360 19836 12388 21286
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12440 19848 12492 19854
rect 12032 19808 12296 19836
rect 11980 19790 12032 19796
rect 11783 19612 12091 19621
rect 11783 19610 11789 19612
rect 11845 19610 11869 19612
rect 11925 19610 11949 19612
rect 12005 19610 12029 19612
rect 12085 19610 12091 19612
rect 11845 19558 11847 19610
rect 12027 19558 12029 19610
rect 11783 19556 11789 19558
rect 11845 19556 11869 19558
rect 11925 19556 11949 19558
rect 12005 19556 12029 19558
rect 12085 19556 12091 19558
rect 11783 19547 12091 19556
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 11992 18970 12020 19246
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 11794 18728 11850 18737
rect 11794 18663 11796 18672
rect 11848 18663 11850 18672
rect 11796 18634 11848 18640
rect 11783 18524 12091 18533
rect 11783 18522 11789 18524
rect 11845 18522 11869 18524
rect 11925 18522 11949 18524
rect 12005 18522 12029 18524
rect 12085 18522 12091 18524
rect 11845 18470 11847 18522
rect 12027 18470 12029 18522
rect 11783 18468 11789 18470
rect 11845 18468 11869 18470
rect 11925 18468 11949 18470
rect 12005 18468 12029 18470
rect 12085 18468 12091 18470
rect 11783 18459 12091 18468
rect 12072 18080 12124 18086
rect 12176 18068 12204 19110
rect 12268 18136 12296 19808
rect 12360 19808 12440 19836
rect 12360 18970 12388 19808
rect 12440 19790 12492 19796
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12544 18834 12572 19110
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12346 18728 12402 18737
rect 12402 18686 12480 18714
rect 12346 18663 12402 18672
rect 12268 18108 12388 18136
rect 12124 18040 12204 18068
rect 12072 18022 12124 18028
rect 12254 17912 12310 17921
rect 12072 17876 12124 17882
rect 12254 17847 12256 17856
rect 12072 17818 12124 17824
rect 12308 17847 12310 17856
rect 12256 17818 12308 17824
rect 11612 17740 11664 17746
rect 11716 17734 11928 17762
rect 11612 17682 11664 17688
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11624 16998 11652 17682
rect 11900 17678 11928 17734
rect 12084 17678 12112 17818
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 11783 17436 12091 17445
rect 11783 17434 11789 17436
rect 11845 17434 11869 17436
rect 11925 17434 11949 17436
rect 12005 17434 12029 17436
rect 12085 17434 12091 17436
rect 11845 17382 11847 17434
rect 12027 17382 12029 17434
rect 11783 17380 11789 17382
rect 11845 17380 11869 17382
rect 11925 17380 11949 17382
rect 12005 17380 12029 17382
rect 12085 17380 12091 17382
rect 11783 17371 12091 17380
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11624 16114 11652 16934
rect 11716 16833 11744 17274
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11702 16824 11758 16833
rect 11702 16759 11758 16768
rect 11808 16697 11836 17138
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 11886 16824 11942 16833
rect 11886 16759 11888 16768
rect 11940 16759 11942 16768
rect 11888 16730 11940 16736
rect 11794 16688 11850 16697
rect 11992 16658 12020 17070
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 12084 16658 12112 16934
rect 12360 16658 12388 18108
rect 12452 16726 12480 18686
rect 12636 18630 12664 20946
rect 12716 20800 12768 20806
rect 12716 20742 12768 20748
rect 12728 19854 12756 20742
rect 13004 20602 13032 21286
rect 13176 20800 13228 20806
rect 13176 20742 13228 20748
rect 12992 20596 13044 20602
rect 12992 20538 13044 20544
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 13096 20058 13124 20198
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12636 17320 12664 18566
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12544 17292 12664 17320
rect 12440 16720 12492 16726
rect 12440 16662 12492 16668
rect 11794 16623 11850 16632
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16153 11744 16526
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 11783 16348 12091 16357
rect 11783 16346 11789 16348
rect 11845 16346 11869 16348
rect 11925 16346 11949 16348
rect 12005 16346 12029 16348
rect 12085 16346 12091 16348
rect 11845 16294 11847 16346
rect 12027 16294 12029 16346
rect 11783 16292 11789 16294
rect 11845 16292 11869 16294
rect 11925 16292 11949 16294
rect 12005 16292 12029 16294
rect 12085 16292 12091 16294
rect 11783 16283 12091 16292
rect 11702 16144 11758 16153
rect 11612 16108 11664 16114
rect 11702 16079 11758 16088
rect 11612 16050 11664 16056
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11532 15706 11560 15846
rect 11624 15706 11652 16050
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11624 15026 11652 15642
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 11783 15260 12091 15269
rect 11783 15258 11789 15260
rect 11845 15258 11869 15260
rect 11925 15258 11949 15260
rect 12005 15258 12029 15260
rect 12085 15258 12091 15260
rect 11845 15206 11847 15258
rect 12027 15206 12029 15258
rect 11783 15204 11789 15206
rect 11845 15204 11869 15206
rect 11925 15204 11949 15206
rect 12005 15204 12029 15206
rect 12085 15204 12091 15206
rect 11783 15195 12091 15204
rect 11900 15116 12112 15144
rect 11900 15026 11928 15116
rect 12084 15026 12112 15116
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11980 15018 12032 15024
rect 11520 14544 11572 14550
rect 11624 14498 11652 14962
rect 11980 14960 12032 14966
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 11992 14618 12020 14960
rect 11980 14612 12032 14618
rect 12360 14600 12388 15438
rect 11980 14554 12032 14560
rect 12176 14572 12388 14600
rect 11572 14492 11652 14498
rect 11520 14486 11652 14492
rect 11532 14470 11652 14486
rect 11624 13938 11652 14470
rect 11796 14408 11848 14414
rect 11794 14376 11796 14385
rect 11848 14376 11850 14385
rect 11794 14311 11850 14320
rect 11783 14172 12091 14181
rect 11783 14170 11789 14172
rect 11845 14170 11869 14172
rect 11925 14170 11949 14172
rect 12005 14170 12029 14172
rect 12085 14170 12091 14172
rect 11845 14118 11847 14170
rect 12027 14118 12029 14170
rect 11783 14116 11789 14118
rect 11845 14116 11869 14118
rect 11925 14116 11949 14118
rect 12005 14116 12029 14118
rect 12085 14116 12091 14118
rect 11783 14107 12091 14116
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11900 13530 11928 13670
rect 12176 13530 12204 14572
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11440 12986 11468 13330
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11348 12646 11376 12718
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11058 11384 11114 11393
rect 11440 11354 11468 12922
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11532 12345 11560 12786
rect 11518 12336 11574 12345
rect 11624 12322 11652 13398
rect 12268 13190 12296 14350
rect 12256 13184 12308 13190
rect 12452 13138 12480 16390
rect 12544 14113 12572 17292
rect 12728 17082 12756 18022
rect 12820 17882 12848 19790
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13004 18834 13032 19110
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 13188 18154 13216 20742
rect 13726 20632 13782 20641
rect 13726 20567 13782 20576
rect 13740 19718 13768 20567
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13268 19304 13320 19310
rect 13268 19246 13320 19252
rect 13358 19272 13414 19281
rect 13176 18148 13228 18154
rect 13176 18090 13228 18096
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 12728 17054 12848 17082
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12728 14278 12756 16934
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12530 14104 12586 14113
rect 12530 14039 12586 14048
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12256 13126 12308 13132
rect 12360 13110 12480 13138
rect 11783 13084 12091 13093
rect 11783 13082 11789 13084
rect 11845 13082 11869 13084
rect 11925 13082 11949 13084
rect 12005 13082 12029 13084
rect 12085 13082 12091 13084
rect 11845 13030 11847 13082
rect 12027 13030 12029 13082
rect 11783 13028 11789 13030
rect 11845 13028 11869 13030
rect 11925 13028 11949 13030
rect 12005 13028 12029 13030
rect 12085 13028 12091 13030
rect 11783 13019 12091 13028
rect 12360 13025 12388 13110
rect 12346 13016 12402 13025
rect 12346 12951 12402 12960
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 11716 12442 11744 12718
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11624 12294 11744 12322
rect 11518 12271 11520 12280
rect 11572 12271 11574 12280
rect 11520 12242 11572 12248
rect 11610 12064 11666 12073
rect 11610 11999 11666 12008
rect 11624 11830 11652 11999
rect 11612 11824 11664 11830
rect 11518 11792 11574 11801
rect 11612 11766 11664 11772
rect 11518 11727 11574 11736
rect 11532 11354 11560 11727
rect 11716 11626 11744 12294
rect 11783 11996 12091 12005
rect 11783 11994 11789 11996
rect 11845 11994 11869 11996
rect 11925 11994 11949 11996
rect 12005 11994 12029 11996
rect 12085 11994 12091 11996
rect 11845 11942 11847 11994
rect 12027 11942 12029 11994
rect 11783 11940 11789 11942
rect 11845 11940 11869 11942
rect 11925 11940 11949 11942
rect 12005 11940 12029 11942
rect 12085 11940 12091 11942
rect 11783 11931 12091 11940
rect 12176 11937 12204 12718
rect 12162 11928 12218 11937
rect 12162 11863 12218 11872
rect 12176 11830 12204 11863
rect 12164 11824 12216 11830
rect 12164 11766 12216 11772
rect 12360 11744 12388 12951
rect 12544 12832 12572 13466
rect 12716 13320 12768 13326
rect 12716 13262 12768 13268
rect 12452 12804 12572 12832
rect 12624 12844 12676 12850
rect 12452 12306 12480 12804
rect 12624 12786 12676 12792
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12544 12345 12572 12650
rect 12530 12336 12586 12345
rect 12440 12300 12492 12306
rect 12530 12271 12586 12280
rect 12440 12242 12492 12248
rect 12544 11830 12572 12271
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12268 11716 12388 11744
rect 11704 11620 11756 11626
rect 11704 11562 11756 11568
rect 12164 11552 12216 11558
rect 12070 11520 12126 11529
rect 12164 11494 12216 11500
rect 12070 11455 12126 11464
rect 11058 11319 11114 11328
rect 11428 11348 11480 11354
rect 11072 11218 11100 11319
rect 11428 11290 11480 11296
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11060 11212 11112 11218
rect 11440 11200 11468 11290
rect 12084 11286 12112 11455
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 11520 11212 11572 11218
rect 11440 11172 11520 11200
rect 11060 11154 11112 11160
rect 11520 11154 11572 11160
rect 12176 11150 12204 11494
rect 12268 11200 12296 11716
rect 12346 11656 12402 11665
rect 12346 11591 12402 11600
rect 12360 11558 12388 11591
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12268 11172 12388 11200
rect 12164 11144 12216 11150
rect 11532 11082 11836 11098
rect 12164 11086 12216 11092
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11520 11076 11848 11082
rect 11572 11070 11796 11076
rect 11520 11018 11572 11024
rect 11796 11018 11848 11024
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 11164 10062 11192 10474
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 9586 11100 9862
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11164 9518 11192 9998
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11164 9042 11192 9454
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11150 8936 11206 8945
rect 11150 8871 11152 8880
rect 11204 8871 11206 8880
rect 11152 8842 11204 8848
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 11058 7304 11114 7313
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10152 5914 10180 6054
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10612 5846 10640 7142
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10060 4146 10088 5646
rect 10508 5568 10560 5574
rect 10704 5545 10732 6938
rect 10980 6866 11008 7278
rect 11058 7239 11114 7248
rect 11072 7206 11100 7239
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11164 6984 11192 8842
rect 11256 8498 11284 11018
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11348 8430 11376 11018
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11716 10742 11744 10950
rect 11783 10908 12091 10917
rect 11783 10906 11789 10908
rect 11845 10906 11869 10908
rect 11925 10906 11949 10908
rect 12005 10906 12029 10908
rect 12085 10906 12091 10908
rect 11845 10854 11847 10906
rect 12027 10854 12029 10906
rect 11783 10852 11789 10854
rect 11845 10852 11869 10854
rect 11925 10852 11949 10854
rect 12005 10852 12029 10854
rect 12085 10852 12091 10854
rect 11783 10843 12091 10852
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11532 10062 11560 10610
rect 11992 10470 12020 10678
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11532 9518 11560 9998
rect 11624 9722 11652 9998
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11532 9178 11560 9454
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11716 9058 11744 9998
rect 11783 9820 12091 9829
rect 11783 9818 11789 9820
rect 11845 9818 11869 9820
rect 11925 9818 11949 9820
rect 12005 9818 12029 9820
rect 12085 9818 12091 9820
rect 11845 9766 11847 9818
rect 12027 9766 12029 9818
rect 11783 9764 11789 9766
rect 11845 9764 11869 9766
rect 11925 9764 11949 9766
rect 12005 9764 12029 9766
rect 12085 9764 12091 9766
rect 11783 9755 12091 9764
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 11624 9030 11744 9058
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11256 7410 11284 7822
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 11348 6984 11376 8366
rect 11072 6956 11192 6984
rect 11256 6956 11376 6984
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 11072 6474 11100 6956
rect 11256 6882 11284 6956
rect 11164 6866 11284 6882
rect 11152 6860 11284 6866
rect 11204 6854 11284 6860
rect 11152 6802 11204 6808
rect 11072 6446 11192 6474
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11072 5846 11100 6326
rect 11164 5846 11192 6446
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 10968 5636 11020 5642
rect 10968 5578 11020 5584
rect 10508 5510 10560 5516
rect 10690 5536 10746 5545
rect 10520 4146 10548 5510
rect 10690 5471 10746 5480
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10980 3738 11008 5578
rect 11072 5166 11100 5646
rect 11164 5370 11192 5782
rect 11256 5642 11284 6854
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11348 6338 11376 6802
rect 11440 6458 11468 8570
rect 11532 8498 11560 8910
rect 11624 8838 11652 9030
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11716 8634 11744 8910
rect 11783 8732 12091 8741
rect 11783 8730 11789 8732
rect 11845 8730 11869 8732
rect 11925 8730 11949 8732
rect 12005 8730 12029 8732
rect 12085 8730 12091 8732
rect 11845 8678 11847 8730
rect 12027 8678 12029 8730
rect 11783 8676 11789 8678
rect 11845 8676 11869 8678
rect 11925 8676 11949 8678
rect 12005 8676 12029 8678
rect 12085 8676 12091 8678
rect 11783 8667 12091 8676
rect 12176 8634 12204 9454
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12268 8514 12296 11018
rect 12360 10470 12388 11172
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 12176 8486 12296 8514
rect 12176 8362 12204 8486
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 11518 8256 11574 8265
rect 11518 8191 11574 8200
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11426 6352 11482 6361
rect 11348 6310 11426 6338
rect 11348 5681 11376 6310
rect 11426 6287 11482 6296
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11334 5672 11390 5681
rect 11244 5636 11296 5642
rect 11334 5607 11390 5616
rect 11244 5578 11296 5584
rect 11336 5568 11388 5574
rect 11336 5510 11388 5516
rect 11152 5364 11204 5370
rect 11204 5324 11284 5352
rect 11152 5306 11204 5312
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 11072 4486 11100 5102
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9784 2502 9996 2530
rect 9784 2446 9812 2502
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9588 1964 9640 1970
rect 9588 1906 9640 1912
rect 9496 1420 9548 1426
rect 9496 1362 9548 1368
rect 9600 1193 9628 1906
rect 9586 1184 9642 1193
rect 9586 1119 9642 1128
rect 6512 632 6684 660
rect 9404 672 9456 678
rect 6460 614 6512 620
rect 9404 614 9456 620
rect 6182 575 6238 584
rect 7988 572 8296 581
rect 7988 570 7994 572
rect 8050 570 8074 572
rect 8130 570 8154 572
rect 8210 570 8234 572
rect 8290 570 8296 572
rect 8050 518 8052 570
rect 8232 518 8234 570
rect 7988 516 7994 518
rect 8050 516 8074 518
rect 8130 516 8154 518
rect 8210 516 8234 518
rect 8290 516 8296 518
rect 7988 507 8296 516
rect 9128 400 9180 406
rect 9128 342 9180 348
rect 9140 134 9168 342
rect 9128 128 9180 134
rect 9128 70 9180 76
rect 9784 66 9812 2382
rect 10060 2378 10088 2586
rect 10520 2514 10548 3674
rect 11072 3466 11100 4422
rect 11256 4146 11284 5324
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11150 3904 11206 3913
rect 11150 3839 11206 3848
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 10612 2553 10640 2586
rect 10598 2544 10654 2553
rect 10508 2508 10560 2514
rect 10598 2479 10654 2488
rect 10508 2450 10560 2456
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 10520 1494 10548 2450
rect 10888 2106 10916 2586
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 10784 1896 10836 1902
rect 10784 1838 10836 1844
rect 10508 1488 10560 1494
rect 10508 1430 10560 1436
rect 10796 1222 10824 1838
rect 10876 1760 10928 1766
rect 10876 1702 10928 1708
rect 10888 1562 10916 1702
rect 10980 1562 11008 3130
rect 11072 2990 11100 3402
rect 11164 3233 11192 3839
rect 11150 3224 11206 3233
rect 11150 3159 11206 3168
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11072 2514 11100 2926
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11072 1902 11100 2450
rect 11164 2258 11192 3159
rect 11256 2360 11284 4082
rect 11348 2990 11376 5510
rect 11440 4826 11468 5714
rect 11532 5642 11560 8191
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 11624 6934 11652 7958
rect 11716 7002 11744 8026
rect 12268 7750 12296 8298
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 11783 7644 12091 7653
rect 11783 7642 11789 7644
rect 11845 7642 11869 7644
rect 11925 7642 11949 7644
rect 12005 7642 12029 7644
rect 12085 7642 12091 7644
rect 11845 7590 11847 7642
rect 12027 7590 12029 7642
rect 11783 7588 11789 7590
rect 11845 7588 11869 7590
rect 11925 7588 11949 7590
rect 12005 7588 12029 7590
rect 12085 7588 12091 7590
rect 11783 7579 12091 7588
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11612 6928 11664 6934
rect 11612 6870 11664 6876
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11716 6118 11744 6802
rect 11900 6662 11928 7278
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12084 7002 12112 7142
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12268 6866 12296 7686
rect 12360 7410 12388 9862
rect 12452 9081 12480 11018
rect 12532 11008 12584 11014
rect 12636 10996 12664 12786
rect 12728 12238 12756 13262
rect 12820 12986 12848 17054
rect 12912 16794 12940 17614
rect 13004 17542 13032 18022
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 12990 16960 13046 16969
rect 12990 16895 13046 16904
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 13004 16658 13032 16895
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 13096 15910 13124 17478
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13188 13682 13216 18090
rect 13280 17746 13308 19246
rect 13358 19207 13414 19216
rect 13372 18426 13400 19207
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13268 17740 13320 17746
rect 13320 17700 13400 17728
rect 13268 17682 13320 17688
rect 13268 17264 13320 17270
rect 13266 17232 13268 17241
rect 13320 17232 13322 17241
rect 13266 17167 13322 17176
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 13280 16658 13308 16934
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13372 16538 13400 17700
rect 12912 13654 13216 13682
rect 13280 16510 13400 16538
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12728 11898 12756 12174
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12728 11150 12756 11834
rect 12820 11354 12848 12378
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12584 10968 12664 10996
rect 12532 10950 12584 10956
rect 12728 10742 12756 11086
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12820 9110 12848 10474
rect 12912 10010 12940 13654
rect 12990 13560 13046 13569
rect 13280 13530 13308 16510
rect 13360 16448 13412 16454
rect 13358 16416 13360 16425
rect 13412 16416 13414 16425
rect 13358 16351 13414 16360
rect 13464 16250 13492 19450
rect 13832 18970 13860 21354
rect 14016 20602 14044 21519
rect 14186 21448 14242 21457
rect 15948 21418 15976 22102
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 16132 21486 16160 22034
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 14186 21383 14242 21392
rect 15936 21412 15988 21418
rect 14200 21350 14228 21383
rect 15936 21354 15988 21360
rect 14188 21344 14240 21350
rect 14188 21286 14240 21292
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 15384 21140 15436 21146
rect 15488 21128 15516 21286
rect 15578 21244 15886 21253
rect 15578 21242 15584 21244
rect 15640 21242 15664 21244
rect 15720 21242 15744 21244
rect 15800 21242 15824 21244
rect 15880 21242 15886 21244
rect 15640 21190 15642 21242
rect 15822 21190 15824 21242
rect 15578 21188 15584 21190
rect 15640 21188 15664 21190
rect 15720 21188 15744 21190
rect 15800 21188 15824 21190
rect 15880 21188 15886 21190
rect 15578 21179 15886 21188
rect 15660 21140 15712 21146
rect 15488 21100 15660 21128
rect 15384 21082 15436 21088
rect 15660 21082 15712 21088
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14004 20324 14056 20330
rect 14004 20266 14056 20272
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13544 18352 13596 18358
rect 13544 18294 13596 18300
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13556 16114 13584 18294
rect 13924 18222 13952 19654
rect 14016 19514 14044 20266
rect 14200 19922 14228 20402
rect 14476 20262 14504 21082
rect 14844 21026 14872 21082
rect 15106 21040 15162 21049
rect 14844 20998 15106 21026
rect 14844 20330 14872 20998
rect 15106 20975 15162 20984
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 14200 19378 14228 19858
rect 14476 19417 14504 20198
rect 14462 19408 14518 19417
rect 14188 19372 14240 19378
rect 14844 19378 14872 20266
rect 15396 20262 15424 21082
rect 16120 21004 16172 21010
rect 16120 20946 16172 20952
rect 16132 20330 16160 20946
rect 16120 20324 16172 20330
rect 16120 20266 16172 20272
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15396 19922 15424 20198
rect 15578 20156 15886 20165
rect 15578 20154 15584 20156
rect 15640 20154 15664 20156
rect 15720 20154 15744 20156
rect 15800 20154 15824 20156
rect 15880 20154 15886 20156
rect 15640 20102 15642 20154
rect 15822 20102 15824 20154
rect 15578 20100 15584 20102
rect 15640 20100 15664 20102
rect 15720 20100 15744 20102
rect 15800 20100 15824 20102
rect 15880 20100 15886 20102
rect 15578 20091 15886 20100
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15856 19378 15884 19654
rect 14462 19343 14518 19352
rect 14832 19372 14884 19378
rect 14188 19314 14240 19320
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13832 17678 13860 18158
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14292 17882 14320 18022
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13648 17105 13676 17478
rect 13634 17096 13690 17105
rect 13634 17031 13690 17040
rect 13832 16590 13860 17614
rect 14004 17128 14056 17134
rect 14096 17128 14148 17134
rect 14004 17070 14056 17076
rect 14094 17096 14096 17105
rect 14148 17096 14150 17105
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13634 16280 13690 16289
rect 13634 16215 13690 16224
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13648 15994 13676 16215
rect 13832 16046 13860 16526
rect 13556 15978 13676 15994
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13544 15972 13676 15978
rect 13596 15966 13676 15972
rect 13544 15914 13596 15920
rect 13556 15745 13584 15914
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13542 15736 13598 15745
rect 13452 15700 13504 15706
rect 13542 15671 13598 15680
rect 13452 15642 13504 15648
rect 13464 15609 13492 15642
rect 13450 15600 13506 15609
rect 13450 15535 13506 15544
rect 13740 15162 13768 15846
rect 13832 15502 13860 15982
rect 13924 15881 13952 15982
rect 14016 15978 14044 17070
rect 14094 17031 14150 17040
rect 14188 16584 14240 16590
rect 14292 16572 14320 17818
rect 14476 17270 14504 19343
rect 14832 19314 14884 19320
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 14554 18864 14610 18873
rect 14554 18799 14556 18808
rect 14608 18799 14610 18808
rect 14556 18770 14608 18776
rect 14464 17264 14516 17270
rect 14464 17206 14516 17212
rect 14648 17060 14700 17066
rect 14844 17048 14872 19314
rect 15948 19310 15976 19790
rect 16132 19514 16160 20266
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 15936 19304 15988 19310
rect 15106 19272 15162 19281
rect 15162 19230 15240 19258
rect 15936 19246 15988 19252
rect 15106 19207 15162 19216
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 15028 18170 15056 18226
rect 15028 18142 15148 18170
rect 15120 18086 15148 18142
rect 15108 18080 15160 18086
rect 15108 18022 15160 18028
rect 15212 17338 15240 19230
rect 15578 19068 15886 19077
rect 15578 19066 15584 19068
rect 15640 19066 15664 19068
rect 15720 19066 15744 19068
rect 15800 19066 15824 19068
rect 15880 19066 15886 19068
rect 15640 19014 15642 19066
rect 15822 19014 15824 19066
rect 15578 19012 15584 19014
rect 15640 19012 15664 19014
rect 15720 19012 15744 19014
rect 15800 19012 15824 19014
rect 15880 19012 15886 19014
rect 15578 19003 15886 19012
rect 15948 18834 15976 19246
rect 16028 19168 16080 19174
rect 16028 19110 16080 19116
rect 16040 18970 16068 19110
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15856 18290 15884 18702
rect 15384 18284 15436 18290
rect 15384 18226 15436 18232
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 14700 17020 14872 17048
rect 14924 17060 14976 17066
rect 14648 17002 14700 17008
rect 14924 17002 14976 17008
rect 14554 16960 14610 16969
rect 14660 16946 14688 17002
rect 14610 16918 14688 16946
rect 14554 16895 14610 16904
rect 14240 16544 14320 16572
rect 14936 16561 14964 17002
rect 15028 16590 15056 17070
rect 15200 17060 15252 17066
rect 15200 17002 15252 17008
rect 15106 16824 15162 16833
rect 15212 16794 15240 17002
rect 15106 16759 15162 16768
rect 15200 16788 15252 16794
rect 15016 16584 15068 16590
rect 14922 16552 14978 16561
rect 14188 16526 14240 16532
rect 14004 15972 14056 15978
rect 14004 15914 14056 15920
rect 13910 15872 13966 15881
rect 13910 15807 13966 15816
rect 14200 15570 14228 16526
rect 15016 16526 15068 16532
rect 14922 16487 14978 16496
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 15120 16402 15148 16759
rect 15200 16730 15252 16736
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14476 15502 14504 16390
rect 15120 16374 15240 16402
rect 15212 16130 15240 16374
rect 15304 16250 15332 18158
rect 15396 17882 15424 18226
rect 15578 17980 15886 17989
rect 15578 17978 15584 17980
rect 15640 17978 15664 17980
rect 15720 17978 15744 17980
rect 15800 17978 15824 17980
rect 15880 17978 15886 17980
rect 15640 17926 15642 17978
rect 15822 17926 15824 17978
rect 15578 17924 15584 17926
rect 15640 17924 15664 17926
rect 15720 17924 15744 17926
rect 15800 17924 15824 17926
rect 15880 17924 15886 17926
rect 15578 17915 15886 17924
rect 16132 17882 16160 19450
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 15568 17808 15620 17814
rect 15568 17750 15620 17756
rect 16026 17776 16082 17785
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15384 17264 15436 17270
rect 15384 17206 15436 17212
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15212 16102 15332 16130
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14832 15904 14884 15910
rect 14832 15846 14884 15852
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13450 14920 13506 14929
rect 13450 14855 13506 14864
rect 13464 14618 13492 14855
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13648 14074 13676 14758
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13740 13705 13768 15098
rect 13832 14958 13860 15438
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13832 14822 13860 14894
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13832 14414 13860 14758
rect 13820 14408 13872 14414
rect 14464 14408 14516 14414
rect 13820 14350 13872 14356
rect 14278 14376 14334 14385
rect 14462 14376 14464 14385
rect 14556 14408 14608 14414
rect 14516 14376 14518 14385
rect 14334 14334 14412 14362
rect 14278 14311 14334 14320
rect 14188 14272 14240 14278
rect 14094 14240 14150 14249
rect 14188 14214 14240 14220
rect 14094 14175 14150 14184
rect 14108 13870 14136 14175
rect 14200 13870 14228 14214
rect 14278 13968 14334 13977
rect 14278 13903 14334 13912
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 13358 13696 13414 13705
rect 13358 13631 13414 13640
rect 13726 13696 13782 13705
rect 13726 13631 13782 13640
rect 12990 13495 13046 13504
rect 13268 13524 13320 13530
rect 13004 12782 13032 13495
rect 13268 13466 13320 13472
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13188 12782 13216 13262
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13004 11830 13032 12718
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 12992 11824 13044 11830
rect 12992 11766 13044 11772
rect 13096 11218 13124 12582
rect 13188 12306 13216 12582
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13280 12102 13308 13262
rect 13372 12782 13400 13631
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13452 12912 13504 12918
rect 13452 12854 13504 12860
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13174 11928 13230 11937
rect 13174 11863 13230 11872
rect 13268 11892 13320 11898
rect 13188 11694 13216 11863
rect 13268 11834 13320 11840
rect 13280 11694 13308 11834
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13176 11552 13228 11558
rect 13174 11520 13176 11529
rect 13268 11552 13320 11558
rect 13228 11520 13230 11529
rect 13268 11494 13320 11500
rect 13174 11455 13230 11464
rect 13280 11354 13308 11494
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13372 11218 13400 12718
rect 13464 12238 13492 12854
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13176 11144 13228 11150
rect 13004 11092 13176 11098
rect 13004 11086 13228 11092
rect 13004 11070 13216 11086
rect 13004 10305 13032 11070
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 12990 10296 13046 10305
rect 12990 10231 13046 10240
rect 13096 10130 13124 10474
rect 13464 10198 13492 11766
rect 13556 11694 13584 12718
rect 13648 12646 13676 13262
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13648 12442 13676 12582
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13832 11898 13860 13806
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13924 11393 13952 12786
rect 14292 12442 14320 13903
rect 14384 13274 14412 14334
rect 14556 14350 14608 14356
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14462 14311 14518 14320
rect 14568 13530 14596 14350
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14660 13410 14688 14350
rect 14568 13382 14688 13410
rect 14384 13246 14504 13274
rect 14476 13190 14504 13246
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14280 12436 14332 12442
rect 14384 12434 14412 13126
rect 14568 12753 14596 13382
rect 14648 12776 14700 12782
rect 14554 12744 14610 12753
rect 14648 12718 14700 12724
rect 14554 12679 14610 12688
rect 14384 12406 14504 12434
rect 14280 12378 14332 12384
rect 14278 12336 14334 12345
rect 14004 12300 14056 12306
rect 14278 12271 14334 12280
rect 14004 12242 14056 12248
rect 13910 11384 13966 11393
rect 13910 11319 13966 11328
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 10266 13584 10406
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 12912 9982 13124 10010
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12808 9104 12860 9110
rect 12438 9072 12494 9081
rect 12494 9030 12572 9058
rect 12808 9046 12860 9052
rect 12438 9007 12494 9016
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11783 6556 12091 6565
rect 11783 6554 11789 6556
rect 11845 6554 11869 6556
rect 11925 6554 11949 6556
rect 12005 6554 12029 6556
rect 12085 6554 12091 6556
rect 11845 6502 11847 6554
rect 12027 6502 12029 6554
rect 11783 6500 11789 6502
rect 11845 6500 11869 6502
rect 11925 6500 11949 6502
rect 12005 6500 12029 6502
rect 12085 6500 12091 6502
rect 11783 6491 12091 6500
rect 12544 6254 12572 9030
rect 12820 8945 12848 9046
rect 12806 8936 12862 8945
rect 12806 8871 12862 8880
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12728 7886 12756 8774
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12820 7954 12848 8230
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12808 7472 12860 7478
rect 12808 7414 12860 7420
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12636 6322 12664 7142
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12256 6248 12308 6254
rect 12532 6248 12584 6254
rect 12308 6196 12480 6202
rect 12256 6190 12480 6196
rect 12532 6190 12584 6196
rect 12268 6174 12480 6190
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 11796 5704 11848 5710
rect 11716 5664 11796 5692
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 11716 5030 11744 5664
rect 11796 5646 11848 5652
rect 11783 5468 12091 5477
rect 11783 5466 11789 5468
rect 11845 5466 11869 5468
rect 11925 5466 11949 5468
rect 12005 5466 12029 5468
rect 12085 5466 12091 5468
rect 11845 5414 11847 5466
rect 12027 5414 12029 5466
rect 11783 5412 11789 5414
rect 11845 5412 11869 5414
rect 11925 5412 11949 5414
rect 12005 5412 12029 5414
rect 12085 5412 12091 5414
rect 11783 5403 12091 5412
rect 12176 5234 12204 6054
rect 12254 5808 12310 5817
rect 12254 5743 12310 5752
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 4826 11744 4966
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11716 3618 11744 4762
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 11783 4380 12091 4389
rect 11783 4378 11789 4380
rect 11845 4378 11869 4380
rect 11925 4378 11949 4380
rect 12005 4378 12029 4380
rect 12085 4378 12091 4380
rect 11845 4326 11847 4378
rect 12027 4326 12029 4378
rect 11783 4324 11789 4326
rect 11845 4324 11869 4326
rect 11925 4324 11949 4326
rect 12005 4324 12029 4326
rect 12085 4324 12091 4326
rect 11783 4315 12091 4324
rect 12176 4282 12204 4558
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12072 3936 12124 3942
rect 12268 3913 12296 5743
rect 12360 4690 12388 6054
rect 12452 5914 12480 6174
rect 12728 6118 12756 7278
rect 12820 6866 12848 7414
rect 12912 6866 12940 8502
rect 13004 6866 13032 9318
rect 13096 7478 13124 9982
rect 13464 9674 13492 10134
rect 13740 9994 13768 10950
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13464 9646 13676 9674
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 7546 13492 7686
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13084 7472 13136 7478
rect 13084 7414 13136 7420
rect 13648 6866 13676 9646
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 9178 13768 9318
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13740 8634 13768 8910
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13832 8430 13860 10678
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13924 10130 13952 10542
rect 14016 10538 14044 12242
rect 14292 12238 14320 12271
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14096 11688 14148 11694
rect 14096 11630 14148 11636
rect 14108 11529 14136 11630
rect 14094 11520 14150 11529
rect 14094 11455 14150 11464
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14004 10532 14056 10538
rect 14056 10492 14136 10520
rect 14004 10474 14056 10480
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13924 9518 13952 10066
rect 14002 10024 14058 10033
rect 14002 9959 14058 9968
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13924 8974 13952 9454
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13832 7410 13860 7822
rect 14016 7546 14044 9959
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 14108 7426 14136 10492
rect 14200 8498 14228 11290
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14292 10266 14320 10610
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14292 9382 14320 10202
rect 14476 10010 14504 12406
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14568 10674 14596 12038
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14660 10470 14688 12718
rect 14752 11150 14780 15846
rect 14844 15570 14872 15846
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 14844 14822 14872 15506
rect 15106 14920 15162 14929
rect 15106 14855 15162 14864
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14844 14618 14872 14758
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14844 13734 14872 14554
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14844 13530 14872 13670
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14936 13394 14964 14554
rect 15120 13938 15148 14855
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15198 13832 15254 13841
rect 15198 13767 15254 13776
rect 15108 13524 15160 13530
rect 15028 13484 15108 13512
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14752 10674 14780 10950
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14648 10464 14700 10470
rect 14648 10406 14700 10412
rect 14384 9982 14504 10010
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14384 9586 14412 9982
rect 14568 9926 14596 9998
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14292 9058 14320 9318
rect 14292 9042 14412 9058
rect 14292 9036 14424 9042
rect 14292 9030 14372 9036
rect 14372 8978 14424 8984
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14292 8498 14320 8774
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14384 8430 14412 8978
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14372 7744 14424 7750
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13924 7398 14136 7426
rect 14200 7704 14372 7732
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13648 6186 13676 6802
rect 13832 6730 13860 7142
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13832 6322 13860 6666
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 13924 6186 13952 7398
rect 14200 7290 14228 7704
rect 14372 7686 14424 7692
rect 14568 7546 14596 7822
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14108 7262 14228 7290
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12438 5808 12494 5817
rect 12636 5778 12664 6054
rect 13648 5914 13676 6122
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 12438 5743 12494 5752
rect 12624 5772 12676 5778
rect 12452 5710 12480 5743
rect 12624 5714 12676 5720
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13450 5400 13506 5409
rect 13450 5335 13506 5344
rect 13266 5264 13322 5273
rect 13266 5199 13322 5208
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12544 4282 12572 4558
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12072 3878 12124 3884
rect 12254 3904 12310 3913
rect 12084 3738 12112 3878
rect 12254 3839 12310 3848
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 11532 3590 11836 3618
rect 11532 3534 11560 3590
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11716 2854 11744 3590
rect 11808 3534 11836 3590
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 11783 3292 12091 3301
rect 11783 3290 11789 3292
rect 11845 3290 11869 3292
rect 11925 3290 11949 3292
rect 12005 3290 12029 3292
rect 12085 3290 12091 3292
rect 11845 3238 11847 3290
rect 12027 3238 12029 3290
rect 11783 3236 11789 3238
rect 11845 3236 11869 3238
rect 11925 3236 11949 3238
rect 12005 3236 12029 3238
rect 12085 3236 12091 3238
rect 11783 3227 12091 3236
rect 12254 3088 12310 3097
rect 12254 3023 12310 3032
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 11256 2332 11376 2360
rect 11164 2230 11284 2258
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 11060 1896 11112 1902
rect 11060 1838 11112 1844
rect 10876 1556 10928 1562
rect 10876 1498 10928 1504
rect 10968 1556 11020 1562
rect 10968 1498 11020 1504
rect 11060 1556 11112 1562
rect 11060 1498 11112 1504
rect 11072 1465 11100 1498
rect 11058 1456 11114 1465
rect 11058 1391 11114 1400
rect 10784 1216 10836 1222
rect 10784 1158 10836 1164
rect 11164 1034 11192 2042
rect 11072 1018 11192 1034
rect 11060 1012 11192 1018
rect 11112 1006 11192 1012
rect 11060 954 11112 960
rect 11256 882 11284 2230
rect 11348 1426 11376 2332
rect 11532 1902 11560 2518
rect 11716 2446 11744 2790
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 11520 1896 11572 1902
rect 11520 1838 11572 1844
rect 11716 1766 11744 2382
rect 11783 2204 12091 2213
rect 11783 2202 11789 2204
rect 11845 2202 11869 2204
rect 11925 2202 11949 2204
rect 12005 2202 12029 2204
rect 12085 2202 12091 2204
rect 11845 2150 11847 2202
rect 12027 2150 12029 2202
rect 11783 2148 11789 2150
rect 11845 2148 11869 2150
rect 11925 2148 11949 2150
rect 12005 2148 12029 2150
rect 12085 2148 12091 2150
rect 11783 2139 12091 2148
rect 12176 2106 12204 2382
rect 12164 2100 12216 2106
rect 12164 2042 12216 2048
rect 11888 1896 11940 1902
rect 11808 1844 11888 1850
rect 11808 1838 11940 1844
rect 11808 1822 11928 1838
rect 11704 1760 11756 1766
rect 11426 1728 11482 1737
rect 11704 1702 11756 1708
rect 11426 1663 11482 1672
rect 11440 1465 11468 1663
rect 11426 1456 11482 1465
rect 11336 1420 11388 1426
rect 11426 1391 11482 1400
rect 11612 1420 11664 1426
rect 11336 1362 11388 1368
rect 11612 1362 11664 1368
rect 11244 876 11296 882
rect 11244 818 11296 824
rect 11348 814 11376 1362
rect 11624 1306 11652 1362
rect 11808 1306 11836 1822
rect 11888 1760 11940 1766
rect 11888 1702 11940 1708
rect 11900 1358 11928 1702
rect 11440 1290 11652 1306
rect 11428 1284 11652 1290
rect 11480 1278 11652 1284
rect 11716 1278 11836 1306
rect 11888 1352 11940 1358
rect 11888 1294 11940 1300
rect 12164 1352 12216 1358
rect 12164 1294 12216 1300
rect 11428 1226 11480 1232
rect 11336 808 11388 814
rect 11336 750 11388 756
rect 11612 672 11664 678
rect 11610 640 11612 649
rect 11664 640 11666 649
rect 11610 575 11666 584
rect 11716 474 11744 1278
rect 11783 1116 12091 1125
rect 11783 1114 11789 1116
rect 11845 1114 11869 1116
rect 11925 1114 11949 1116
rect 12005 1114 12029 1116
rect 12085 1114 12091 1116
rect 11845 1062 11847 1114
rect 12027 1062 12029 1114
rect 11783 1060 11789 1062
rect 11845 1060 11869 1062
rect 11925 1060 11949 1062
rect 12005 1060 12029 1062
rect 12085 1060 12091 1062
rect 11783 1051 12091 1060
rect 11980 1012 12032 1018
rect 11980 954 12032 960
rect 11796 876 11848 882
rect 11796 818 11848 824
rect 11704 468 11756 474
rect 11704 410 11756 416
rect 11808 134 11836 818
rect 11992 814 12020 954
rect 11980 808 12032 814
rect 11980 750 12032 756
rect 11992 241 12020 750
rect 12176 377 12204 1294
rect 12268 678 12296 3023
rect 12360 1970 12388 3470
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 12348 1964 12400 1970
rect 12348 1906 12400 1912
rect 12348 1216 12400 1222
rect 12348 1158 12400 1164
rect 12360 882 12388 1158
rect 13188 1018 13216 2042
rect 13280 1018 13308 5199
rect 13464 5166 13492 5335
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13728 5160 13780 5166
rect 13832 5148 13860 5646
rect 13780 5120 13860 5148
rect 13728 5102 13780 5108
rect 13832 4622 13860 5120
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 13464 4010 13492 4422
rect 13832 4078 13860 4558
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 13636 4072 13688 4078
rect 13634 4040 13636 4049
rect 13820 4072 13872 4078
rect 13688 4040 13690 4049
rect 13452 4004 13504 4010
rect 13820 4014 13872 4020
rect 13634 3975 13690 3984
rect 13452 3946 13504 3952
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13556 3534 13584 3878
rect 13832 3534 13860 4014
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 13924 3670 13952 3946
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13648 1766 13676 2926
rect 13728 2440 13780 2446
rect 13832 2428 13860 3470
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13780 2400 13860 2428
rect 13728 2382 13780 2388
rect 13740 1902 13768 2382
rect 13728 1896 13780 1902
rect 13728 1838 13780 1844
rect 13636 1760 13688 1766
rect 13636 1702 13688 1708
rect 13360 1216 13412 1222
rect 13360 1158 13412 1164
rect 13176 1012 13228 1018
rect 13176 954 13228 960
rect 13268 1012 13320 1018
rect 13268 954 13320 960
rect 12348 876 12400 882
rect 12348 818 12400 824
rect 12256 672 12308 678
rect 12256 614 12308 620
rect 12162 368 12218 377
rect 12162 303 12218 312
rect 13372 270 13400 1158
rect 13648 814 13676 1702
rect 13740 1358 13768 1838
rect 13820 1556 13872 1562
rect 13924 1544 13952 2790
rect 14016 2650 14044 4082
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14016 1902 14044 2586
rect 14004 1896 14056 1902
rect 14004 1838 14056 1844
rect 14016 1562 14044 1838
rect 13872 1516 13952 1544
rect 14004 1556 14056 1562
rect 13820 1498 13872 1504
rect 14004 1498 14056 1504
rect 13818 1456 13874 1465
rect 13818 1391 13874 1400
rect 13728 1352 13780 1358
rect 13728 1294 13780 1300
rect 13636 808 13688 814
rect 13636 750 13688 756
rect 13832 678 13860 1391
rect 14108 882 14136 7262
rect 14476 7002 14504 7278
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14660 6866 14688 9318
rect 14844 9042 14872 11018
rect 14936 9042 14964 11494
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14936 8090 14964 8230
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14752 7410 14780 7822
rect 14830 7576 14886 7585
rect 14830 7511 14886 7520
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14200 5234 14228 5646
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14200 4826 14228 5170
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14200 4146 14228 4762
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14200 3738 14228 4082
rect 14292 3942 14320 6258
rect 14384 5778 14412 6326
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14476 4690 14504 6394
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14568 5234 14596 6054
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14464 4684 14516 4690
rect 14464 4626 14516 4632
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14372 4072 14424 4078
rect 14476 4049 14504 4082
rect 14372 4014 14424 4020
rect 14462 4040 14518 4049
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14292 3194 14320 3470
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14384 3074 14412 4014
rect 14462 3975 14518 3984
rect 14292 3046 14412 3074
rect 14292 2990 14320 3046
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14384 2514 14412 2926
rect 14462 2544 14518 2553
rect 14372 2508 14424 2514
rect 14462 2479 14518 2488
rect 14372 2450 14424 2456
rect 14476 2446 14504 2479
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14200 1970 14228 2246
rect 14188 1964 14240 1970
rect 14188 1906 14240 1912
rect 14462 1592 14518 1601
rect 14462 1527 14518 1536
rect 14476 1358 14504 1527
rect 14464 1352 14516 1358
rect 14464 1294 14516 1300
rect 14096 876 14148 882
rect 14096 818 14148 824
rect 14568 814 14596 4218
rect 14660 4078 14688 6802
rect 14752 6254 14780 7346
rect 14844 7274 14872 7511
rect 14936 7410 14964 8026
rect 15028 7750 15056 13484
rect 15108 13466 15160 13472
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15120 12782 15148 13262
rect 15212 12850 15240 13767
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15304 12730 15332 16102
rect 15396 15502 15424 17206
rect 15488 16794 15516 17478
rect 15580 16998 15608 17750
rect 16026 17711 16082 17720
rect 16120 17740 16172 17746
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15578 16892 15886 16901
rect 15578 16890 15584 16892
rect 15640 16890 15664 16892
rect 15720 16890 15744 16892
rect 15800 16890 15824 16892
rect 15880 16890 15886 16892
rect 15640 16838 15642 16890
rect 15822 16838 15824 16890
rect 15578 16836 15584 16838
rect 15640 16836 15664 16838
rect 15720 16836 15744 16838
rect 15800 16836 15824 16838
rect 15880 16836 15886 16838
rect 15578 16827 15886 16836
rect 15948 16794 15976 17070
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 15934 16688 15990 16697
rect 15568 16652 15620 16658
rect 15934 16623 15990 16632
rect 15568 16594 15620 16600
rect 15474 16280 15530 16289
rect 15474 16215 15476 16224
rect 15528 16215 15530 16224
rect 15476 16186 15528 16192
rect 15580 16130 15608 16594
rect 15488 16102 15608 16130
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15488 15348 15516 16102
rect 15578 15804 15886 15813
rect 15578 15802 15584 15804
rect 15640 15802 15664 15804
rect 15720 15802 15744 15804
rect 15800 15802 15824 15804
rect 15880 15802 15886 15804
rect 15640 15750 15642 15802
rect 15822 15750 15824 15802
rect 15578 15748 15584 15750
rect 15640 15748 15664 15750
rect 15720 15748 15744 15750
rect 15800 15748 15824 15750
rect 15880 15748 15886 15750
rect 15578 15739 15886 15748
rect 15948 15638 15976 16623
rect 16040 16522 16068 17711
rect 16120 17682 16172 17688
rect 16132 16726 16160 17682
rect 16120 16720 16172 16726
rect 16120 16662 16172 16668
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 15936 15632 15988 15638
rect 15936 15574 15988 15580
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 15396 15320 15516 15348
rect 15568 15360 15620 15366
rect 15396 14414 15424 15320
rect 15568 15302 15620 15308
rect 15580 14906 15608 15302
rect 15488 14878 15608 14906
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15382 13696 15438 13705
rect 15382 13631 15438 13640
rect 15396 13462 15424 13631
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15488 13002 15516 14878
rect 15578 14716 15886 14725
rect 15578 14714 15584 14716
rect 15640 14714 15664 14716
rect 15720 14714 15744 14716
rect 15800 14714 15824 14716
rect 15880 14714 15886 14716
rect 15640 14662 15642 14714
rect 15822 14662 15824 14714
rect 15578 14660 15584 14662
rect 15640 14660 15664 14662
rect 15720 14660 15744 14662
rect 15800 14660 15824 14662
rect 15880 14660 15886 14662
rect 15578 14651 15886 14660
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 15578 13628 15886 13637
rect 15578 13626 15584 13628
rect 15640 13626 15664 13628
rect 15720 13626 15744 13628
rect 15800 13626 15824 13628
rect 15880 13626 15886 13628
rect 15640 13574 15642 13626
rect 15822 13574 15824 13626
rect 15578 13572 15584 13574
rect 15640 13572 15664 13574
rect 15720 13572 15744 13574
rect 15800 13572 15824 13574
rect 15880 13572 15886 13574
rect 15578 13563 15886 13572
rect 15752 13184 15804 13190
rect 15948 13172 15976 13738
rect 16040 13394 16068 15438
rect 16028 13388 16080 13394
rect 16132 13376 16160 15982
rect 16224 13802 16252 22222
rect 16764 22228 16816 22234
rect 16764 22170 16816 22176
rect 16856 22228 16908 22234
rect 16856 22170 16908 22176
rect 16670 21448 16726 21457
rect 16670 21383 16726 21392
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16592 21049 16620 21082
rect 16578 21040 16634 21049
rect 16684 21010 16712 21383
rect 16578 20975 16634 20984
rect 16672 21004 16724 21010
rect 16672 20946 16724 20952
rect 16684 20398 16712 20946
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 16684 19417 16712 20334
rect 16670 19408 16726 19417
rect 16670 19343 16726 19352
rect 16302 19272 16358 19281
rect 16302 19207 16358 19216
rect 16486 19272 16542 19281
rect 16542 19230 16620 19258
rect 16486 19207 16542 19216
rect 16316 19174 16344 19207
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16302 18184 16358 18193
rect 16358 18142 16436 18170
rect 16302 18119 16358 18128
rect 16408 17320 16436 18142
rect 16592 17882 16620 19230
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16684 17762 16712 19343
rect 16592 17746 16712 17762
rect 16580 17740 16712 17746
rect 16632 17734 16712 17740
rect 16580 17682 16632 17688
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16408 17292 16620 17320
rect 16486 17232 16542 17241
rect 16486 17167 16542 17176
rect 16500 17066 16528 17167
rect 16488 17060 16540 17066
rect 16488 17002 16540 17008
rect 16302 16824 16358 16833
rect 16302 16759 16358 16768
rect 16316 16658 16344 16759
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16396 16516 16448 16522
rect 16396 16458 16448 16464
rect 16304 16176 16356 16182
rect 16302 16144 16304 16153
rect 16356 16144 16358 16153
rect 16302 16079 16358 16088
rect 16408 15366 16436 16458
rect 16592 15994 16620 17292
rect 16684 16794 16712 17614
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16684 16250 16712 16458
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16776 16130 16804 22170
rect 16868 21690 16896 22170
rect 18696 22092 18748 22098
rect 18696 22034 18748 22040
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 16856 21684 16908 21690
rect 16856 21626 16908 21632
rect 16868 21486 16896 21626
rect 17130 21584 17186 21593
rect 17130 21519 17186 21528
rect 16856 21480 16908 21486
rect 16856 21422 16908 21428
rect 17144 21146 17172 21519
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17512 21010 17540 21830
rect 18510 21448 18566 21457
rect 18510 21383 18512 21392
rect 18564 21383 18566 21392
rect 18512 21354 18564 21360
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18616 21146 18644 21286
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 17880 21049 17908 21082
rect 17866 21040 17922 21049
rect 17500 21004 17552 21010
rect 17500 20946 17552 20952
rect 17788 20998 17866 21026
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 17512 20058 17540 20198
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 17236 19310 17264 19790
rect 17788 19378 17816 20998
rect 17866 20975 17922 20984
rect 18708 20505 18736 22034
rect 18892 21690 18920 22238
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 24124 22092 24176 22098
rect 24124 22034 24176 22040
rect 18880 21684 18932 21690
rect 18880 21626 18932 21632
rect 19260 21486 19288 22034
rect 19708 21888 19760 21894
rect 19708 21830 19760 21836
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 23388 21888 23440 21894
rect 23388 21830 23440 21836
rect 19373 21788 19681 21797
rect 19373 21786 19379 21788
rect 19435 21786 19459 21788
rect 19515 21786 19539 21788
rect 19595 21786 19619 21788
rect 19675 21786 19681 21788
rect 19435 21734 19437 21786
rect 19617 21734 19619 21786
rect 19373 21732 19379 21734
rect 19435 21732 19459 21734
rect 19515 21732 19539 21734
rect 19595 21732 19619 21734
rect 19675 21732 19681 21734
rect 19373 21723 19681 21732
rect 19720 21486 19748 21830
rect 19248 21480 19300 21486
rect 19248 21422 19300 21428
rect 19708 21480 19760 21486
rect 19708 21422 19760 21428
rect 19260 21146 19288 21422
rect 19248 21140 19300 21146
rect 19248 21082 19300 21088
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19373 20700 19681 20709
rect 19373 20698 19379 20700
rect 19435 20698 19459 20700
rect 19515 20698 19539 20700
rect 19595 20698 19619 20700
rect 19675 20698 19681 20700
rect 19435 20646 19437 20698
rect 19617 20646 19619 20698
rect 19373 20644 19379 20646
rect 19435 20644 19459 20646
rect 19515 20644 19539 20646
rect 19595 20644 19619 20646
rect 19675 20644 19681 20646
rect 19373 20635 19681 20644
rect 18694 20496 18750 20505
rect 19720 20466 19748 20878
rect 18694 20431 18696 20440
rect 18748 20431 18750 20440
rect 19708 20460 19760 20466
rect 18696 20402 18748 20408
rect 19708 20402 19760 20408
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 18880 20392 18932 20398
rect 18880 20334 18932 20340
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17880 19854 17908 20198
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17776 19372 17828 19378
rect 17682 19348 17738 19357
rect 17224 19304 17276 19310
rect 17776 19314 17828 19320
rect 17682 19283 17684 19292
rect 17224 19246 17276 19252
rect 17736 19283 17738 19292
rect 17684 19246 17736 19252
rect 17236 18834 17264 19246
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 17052 18057 17080 18226
rect 17038 18048 17094 18057
rect 17038 17983 17094 17992
rect 17788 17882 17816 19314
rect 17972 18970 18000 19858
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 18064 18222 18092 20334
rect 18892 20058 18920 20334
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18156 18834 18184 19654
rect 18248 19378 18276 19790
rect 19156 19712 19208 19718
rect 19156 19654 19208 19660
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18892 18290 18920 18634
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 19076 18290 19104 18566
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17052 17134 17080 17614
rect 17040 17128 17092 17134
rect 16854 17096 16910 17105
rect 17040 17070 17092 17076
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 16854 17031 16910 17040
rect 16868 16658 16896 17031
rect 17052 16658 17080 17070
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 17144 16250 17172 17070
rect 17512 16998 17540 17614
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 16776 16102 17080 16130
rect 16948 16040 17000 16046
rect 16592 15966 16712 15994
rect 16948 15982 17000 15988
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 16592 15706 16620 15846
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16408 15065 16436 15302
rect 16394 15056 16450 15065
rect 16592 15026 16620 15302
rect 16394 14991 16450 15000
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16408 14074 16436 14758
rect 16592 14278 16620 14962
rect 16684 14482 16712 15966
rect 16960 15706 16988 15982
rect 17052 15706 17080 16102
rect 17130 16008 17186 16017
rect 17130 15943 17186 15952
rect 17144 15910 17172 15943
rect 17236 15910 17264 16594
rect 17512 16590 17540 16934
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 17040 15700 17092 15706
rect 17040 15642 17092 15648
rect 17236 15502 17264 15846
rect 17512 15570 17540 16526
rect 17604 16454 17632 17478
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17696 16046 17724 16390
rect 17880 16250 17908 17614
rect 18788 17128 18840 17134
rect 18892 17116 18920 18226
rect 18970 17640 19026 17649
rect 19026 17598 19104 17626
rect 18970 17575 19026 17584
rect 18840 17088 18920 17116
rect 18788 17070 18840 17076
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17592 16040 17644 16046
rect 17592 15982 17644 15988
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17604 15706 17632 15982
rect 17868 15972 17920 15978
rect 17868 15914 17920 15920
rect 17592 15700 17644 15706
rect 17592 15642 17644 15648
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 16764 15496 16816 15502
rect 17224 15496 17276 15502
rect 16764 15438 16816 15444
rect 16854 15464 16910 15473
rect 16776 14822 16804 15438
rect 17224 15438 17276 15444
rect 16854 15399 16856 15408
rect 16908 15399 16910 15408
rect 16856 15370 16908 15376
rect 17880 15094 17908 15914
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16776 14482 16804 14758
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16592 13938 16620 14214
rect 16684 13977 16712 14418
rect 16670 13968 16726 13977
rect 16580 13932 16632 13938
rect 16776 13938 16804 14418
rect 16670 13903 16726 13912
rect 16764 13932 16816 13938
rect 16580 13874 16632 13880
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16132 13348 16252 13376
rect 16028 13330 16080 13336
rect 16224 13240 16252 13348
rect 16304 13320 16356 13326
rect 16580 13320 16632 13326
rect 16356 13280 16436 13308
rect 16304 13262 16356 13268
rect 15804 13144 15976 13172
rect 16132 13212 16252 13240
rect 15752 13126 15804 13132
rect 15488 12974 15976 13002
rect 15200 12708 15252 12714
rect 15304 12702 15424 12730
rect 15200 12650 15252 12656
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 15120 11354 15148 12582
rect 15212 12434 15240 12650
rect 15396 12434 15424 12702
rect 15578 12540 15886 12549
rect 15578 12538 15584 12540
rect 15640 12538 15664 12540
rect 15720 12538 15744 12540
rect 15800 12538 15824 12540
rect 15880 12538 15886 12540
rect 15640 12486 15642 12538
rect 15822 12486 15824 12538
rect 15578 12484 15584 12486
rect 15640 12484 15664 12486
rect 15720 12484 15744 12486
rect 15800 12484 15824 12486
rect 15880 12484 15886 12486
rect 15578 12475 15886 12484
rect 15212 12406 15332 12434
rect 15396 12406 15516 12434
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14832 7268 14884 7274
rect 14832 7210 14884 7216
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14936 6118 14964 7346
rect 15120 6322 15148 8774
rect 15212 6866 15240 11154
rect 15304 10577 15332 12406
rect 15488 11014 15516 12406
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15580 11801 15608 12038
rect 15948 11898 15976 12974
rect 16132 12442 16160 13212
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 15566 11792 15622 11801
rect 15566 11727 15622 11736
rect 15578 11452 15886 11461
rect 15578 11450 15584 11452
rect 15640 11450 15664 11452
rect 15720 11450 15744 11452
rect 15800 11450 15824 11452
rect 15880 11450 15886 11452
rect 15640 11398 15642 11450
rect 15822 11398 15824 11450
rect 15578 11396 15584 11398
rect 15640 11396 15664 11398
rect 15720 11396 15744 11398
rect 15800 11396 15824 11398
rect 15880 11396 15886 11398
rect 15578 11387 15886 11396
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15488 10810 15516 10950
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15290 10568 15346 10577
rect 15290 10503 15346 10512
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15304 8090 15332 10406
rect 15578 10364 15886 10373
rect 15578 10362 15584 10364
rect 15640 10362 15664 10364
rect 15720 10362 15744 10364
rect 15800 10362 15824 10364
rect 15880 10362 15886 10364
rect 15640 10310 15642 10362
rect 15822 10310 15824 10362
rect 15578 10308 15584 10310
rect 15640 10308 15664 10310
rect 15720 10308 15744 10310
rect 15800 10308 15824 10310
rect 15880 10308 15886 10310
rect 15578 10299 15886 10308
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15396 7410 15424 9318
rect 15578 9276 15886 9285
rect 15578 9274 15584 9276
rect 15640 9274 15664 9276
rect 15720 9274 15744 9276
rect 15800 9274 15824 9276
rect 15880 9274 15886 9276
rect 15640 9222 15642 9274
rect 15822 9222 15824 9274
rect 15578 9220 15584 9222
rect 15640 9220 15664 9222
rect 15720 9220 15744 9222
rect 15800 9220 15824 9222
rect 15880 9220 15886 9222
rect 15578 9211 15886 9220
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 15578 8188 15886 8197
rect 15578 8186 15584 8188
rect 15640 8186 15664 8188
rect 15720 8186 15744 8188
rect 15800 8186 15824 8188
rect 15880 8186 15886 8188
rect 15640 8134 15642 8186
rect 15822 8134 15824 8186
rect 15578 8132 15584 8134
rect 15640 8132 15664 8134
rect 15720 8132 15744 8134
rect 15800 8132 15824 8134
rect 15880 8132 15886 8134
rect 15578 8123 15886 8132
rect 15948 7954 15976 8366
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 15658 7848 15714 7857
rect 15658 7783 15660 7792
rect 15712 7783 15714 7792
rect 15660 7754 15712 7760
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15396 6322 15424 7142
rect 15488 7002 15516 7346
rect 15578 7100 15886 7109
rect 15578 7098 15584 7100
rect 15640 7098 15664 7100
rect 15720 7098 15744 7100
rect 15800 7098 15824 7100
rect 15880 7098 15886 7100
rect 15640 7046 15642 7098
rect 15822 7046 15824 7098
rect 15578 7044 15584 7046
rect 15640 7044 15664 7046
rect 15720 7044 15744 7046
rect 15800 7044 15824 7046
rect 15880 7044 15886 7046
rect 15578 7035 15886 7044
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 15290 5128 15346 5137
rect 15290 5063 15346 5072
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 15106 3088 15162 3097
rect 15106 3023 15108 3032
rect 15160 3023 15162 3032
rect 15108 2994 15160 3000
rect 15016 2848 15068 2854
rect 15200 2848 15252 2854
rect 15016 2790 15068 2796
rect 15120 2796 15200 2802
rect 15120 2790 15252 2796
rect 14280 808 14332 814
rect 14280 750 14332 756
rect 14556 808 14608 814
rect 14556 750 14608 756
rect 13820 672 13872 678
rect 13820 614 13872 620
rect 14292 474 14320 750
rect 15028 678 15056 2790
rect 15120 2774 15240 2790
rect 15016 672 15068 678
rect 15016 614 15068 620
rect 14280 468 14332 474
rect 14280 410 14332 416
rect 13360 264 13412 270
rect 11978 232 12034 241
rect 13360 206 13412 212
rect 15120 202 15148 2774
rect 15304 1018 15332 5063
rect 15292 1012 15344 1018
rect 15292 954 15344 960
rect 15488 950 15516 6598
rect 15578 6012 15886 6021
rect 15578 6010 15584 6012
rect 15640 6010 15664 6012
rect 15720 6010 15744 6012
rect 15800 6010 15824 6012
rect 15880 6010 15886 6012
rect 15640 5958 15642 6010
rect 15822 5958 15824 6010
rect 15578 5956 15584 5958
rect 15640 5956 15664 5958
rect 15720 5956 15744 5958
rect 15800 5956 15824 5958
rect 15880 5956 15886 5958
rect 15578 5947 15886 5956
rect 16040 5914 16068 9454
rect 16224 6769 16252 12922
rect 16408 12850 16436 13280
rect 16578 13288 16580 13297
rect 16632 13288 16634 13297
rect 16578 13223 16634 13232
rect 16684 13002 16712 13903
rect 16764 13874 16816 13880
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16500 12974 16712 13002
rect 16762 13016 16818 13025
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16302 12744 16358 12753
rect 16302 12679 16358 12688
rect 16316 11286 16344 12679
rect 16500 12288 16528 12974
rect 16868 12986 16896 13262
rect 17972 12986 18000 15438
rect 18064 15162 18092 16526
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18616 15570 18644 15982
rect 18972 15904 19024 15910
rect 18972 15846 19024 15852
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 18326 15056 18382 15065
rect 18326 14991 18382 15000
rect 18340 14618 18368 14991
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18708 14278 18736 14894
rect 18984 14890 19012 15846
rect 19076 15450 19104 17598
rect 19168 17202 19196 19654
rect 19373 19612 19681 19621
rect 19373 19610 19379 19612
rect 19435 19610 19459 19612
rect 19515 19610 19539 19612
rect 19595 19610 19619 19612
rect 19675 19610 19681 19612
rect 19435 19558 19437 19610
rect 19617 19558 19619 19610
rect 19373 19556 19379 19558
rect 19435 19556 19459 19558
rect 19515 19556 19539 19558
rect 19595 19556 19619 19558
rect 19675 19556 19681 19558
rect 19373 19547 19681 19556
rect 19996 19334 20024 20402
rect 20640 19922 20668 21830
rect 23400 21690 23428 21830
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 21456 21480 21508 21486
rect 21456 21422 21508 21428
rect 21364 21344 21416 21350
rect 21364 21286 21416 21292
rect 21376 21146 21404 21286
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20732 20534 20760 20946
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 20720 20528 20772 20534
rect 20720 20470 20772 20476
rect 21284 20398 21312 20878
rect 21364 20528 21416 20534
rect 21364 20470 21416 20476
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 21376 20262 21404 20470
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 20996 19984 21048 19990
rect 20994 19952 20996 19961
rect 21048 19952 21050 19961
rect 20628 19916 20680 19922
rect 20628 19858 20680 19864
rect 20904 19916 20956 19922
rect 20994 19887 21050 19896
rect 20904 19858 20956 19864
rect 19904 19306 20024 19334
rect 19904 18834 19932 19306
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 19892 18828 19944 18834
rect 19892 18770 19944 18776
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 19373 18524 19681 18533
rect 19373 18522 19379 18524
rect 19435 18522 19459 18524
rect 19515 18522 19539 18524
rect 19595 18522 19619 18524
rect 19675 18522 19681 18524
rect 19435 18470 19437 18522
rect 19617 18470 19619 18522
rect 19373 18468 19379 18470
rect 19435 18468 19459 18470
rect 19515 18468 19539 18470
rect 19595 18468 19619 18470
rect 19675 18468 19681 18470
rect 19373 18459 19681 18468
rect 19720 18358 19748 18702
rect 20088 18426 20116 19110
rect 20456 18834 20484 19246
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20456 18698 20484 18770
rect 20444 18692 20496 18698
rect 20444 18634 20496 18640
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 19708 18352 19760 18358
rect 19708 18294 19760 18300
rect 19340 18080 19392 18086
rect 19246 18048 19302 18057
rect 19340 18022 19392 18028
rect 19246 17983 19302 17992
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 19260 16538 19288 17983
rect 19352 17746 19380 18022
rect 19340 17740 19392 17746
rect 19340 17682 19392 17688
rect 20456 17678 20484 18634
rect 20548 18426 20576 19246
rect 20640 18970 20668 19858
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20536 18420 20588 18426
rect 20536 18362 20588 18368
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 19982 17504 20038 17513
rect 19373 17436 19681 17445
rect 19982 17439 20038 17448
rect 19373 17434 19379 17436
rect 19435 17434 19459 17436
rect 19515 17434 19539 17436
rect 19595 17434 19619 17436
rect 19675 17434 19681 17436
rect 19435 17382 19437 17434
rect 19617 17382 19619 17434
rect 19373 17380 19379 17382
rect 19435 17380 19459 17382
rect 19515 17380 19539 17382
rect 19595 17380 19619 17382
rect 19675 17380 19681 17382
rect 19373 17371 19681 17380
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19338 16552 19394 16561
rect 19260 16510 19338 16538
rect 19260 16232 19288 16510
rect 19338 16487 19394 16496
rect 19373 16348 19681 16357
rect 19373 16346 19379 16348
rect 19435 16346 19459 16348
rect 19515 16346 19539 16348
rect 19595 16346 19619 16348
rect 19675 16346 19681 16348
rect 19435 16294 19437 16346
rect 19617 16294 19619 16346
rect 19373 16292 19379 16294
rect 19435 16292 19459 16294
rect 19515 16292 19539 16294
rect 19595 16292 19619 16294
rect 19675 16292 19681 16294
rect 19373 16283 19681 16292
rect 19904 16250 19932 16934
rect 19892 16244 19944 16250
rect 19260 16204 19380 16232
rect 19076 15422 19196 15450
rect 19064 15360 19116 15366
rect 19064 15302 19116 15308
rect 19076 14929 19104 15302
rect 19062 14920 19118 14929
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18972 14884 19024 14890
rect 19062 14855 19118 14864
rect 18972 14826 19024 14832
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 16762 12951 16818 12960
rect 16856 12980 16908 12986
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16408 12260 16528 12288
rect 16408 11354 16436 12260
rect 16684 12186 16712 12786
rect 16776 12782 16804 12951
rect 16856 12922 16908 12928
rect 17960 12980 18012 12986
rect 17960 12922 18012 12928
rect 18616 12850 18644 13262
rect 18708 13190 18736 14214
rect 18892 14006 18920 14826
rect 19062 14784 19118 14793
rect 19062 14719 19118 14728
rect 18970 14376 19026 14385
rect 18970 14311 18972 14320
rect 19024 14311 19026 14320
rect 18972 14282 19024 14288
rect 18970 14104 19026 14113
rect 19076 14090 19104 14719
rect 19026 14062 19104 14090
rect 18970 14039 19026 14048
rect 18880 14000 18932 14006
rect 18880 13942 18932 13948
rect 18984 13870 19012 14039
rect 19168 14006 19196 15422
rect 19352 15348 19380 16204
rect 19892 16186 19944 16192
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19536 15638 19564 15846
rect 19614 15736 19670 15745
rect 19614 15671 19670 15680
rect 19524 15632 19576 15638
rect 19524 15574 19576 15580
rect 19432 15496 19484 15502
rect 19628 15484 19656 15671
rect 19706 15600 19762 15609
rect 19706 15535 19708 15544
rect 19760 15535 19762 15544
rect 19800 15564 19852 15570
rect 19708 15506 19760 15512
rect 19800 15506 19852 15512
rect 19484 15456 19656 15484
rect 19812 15450 19840 15506
rect 19432 15438 19484 15444
rect 19720 15422 19840 15450
rect 19720 15366 19748 15422
rect 19311 15320 19380 15348
rect 19708 15360 19760 15366
rect 19311 15144 19339 15320
rect 19708 15302 19760 15308
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19373 15260 19681 15269
rect 19373 15258 19379 15260
rect 19435 15258 19459 15260
rect 19515 15258 19539 15260
rect 19595 15258 19619 15260
rect 19675 15258 19681 15260
rect 19435 15206 19437 15258
rect 19617 15206 19619 15258
rect 19373 15204 19379 15206
rect 19435 15204 19459 15206
rect 19515 15204 19539 15206
rect 19595 15204 19619 15206
rect 19675 15204 19681 15206
rect 19373 15195 19681 15204
rect 19311 15116 19380 15144
rect 19352 14362 19380 15116
rect 19812 15026 19840 15302
rect 19904 15026 19932 16186
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19260 14334 19380 14362
rect 19156 14000 19208 14006
rect 19156 13942 19208 13948
rect 19260 13954 19288 14334
rect 19373 14172 19681 14181
rect 19373 14170 19379 14172
rect 19435 14170 19459 14172
rect 19515 14170 19539 14172
rect 19595 14170 19619 14172
rect 19675 14170 19681 14172
rect 19435 14118 19437 14170
rect 19617 14118 19619 14170
rect 19373 14116 19379 14118
rect 19435 14116 19459 14118
rect 19515 14116 19539 14118
rect 19595 14116 19619 14118
rect 19675 14116 19681 14118
rect 19373 14107 19681 14116
rect 18972 13864 19024 13870
rect 18892 13812 18972 13818
rect 18892 13806 19024 13812
rect 19168 13818 19196 13942
rect 19260 13938 19472 13954
rect 19260 13932 19484 13938
rect 19260 13926 19432 13932
rect 19432 13874 19484 13880
rect 18892 13790 19012 13806
rect 19168 13790 19288 13818
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 16500 12158 16712 12186
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16408 9586 16436 10542
rect 16500 10169 16528 12158
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16684 11354 16712 12038
rect 16776 11558 16804 12038
rect 17236 11558 17264 12378
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17512 12102 17540 12174
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16776 11150 16804 11494
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16578 10704 16634 10713
rect 16578 10639 16580 10648
rect 16632 10639 16634 10648
rect 16580 10610 16632 10616
rect 16486 10160 16542 10169
rect 16868 10130 16896 11222
rect 17236 11150 17264 11494
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 16486 10095 16542 10104
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16500 9178 16528 9862
rect 16578 9616 16634 9625
rect 16578 9551 16580 9560
rect 16632 9551 16634 9560
rect 16580 9522 16632 9528
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16316 8634 16344 8774
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16316 7449 16344 8570
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16408 8090 16436 8230
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16394 7984 16450 7993
rect 16394 7919 16450 7928
rect 16408 7886 16436 7919
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16302 7440 16358 7449
rect 16302 7375 16358 7384
rect 16500 7274 16528 9114
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16488 7268 16540 7274
rect 16488 7210 16540 7216
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16304 6792 16356 6798
rect 16210 6760 16266 6769
rect 16304 6734 16356 6740
rect 16210 6695 16266 6704
rect 16028 5908 16080 5914
rect 16028 5850 16080 5856
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 15844 5160 15896 5166
rect 16040 5148 16068 5646
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 15896 5120 16068 5148
rect 15844 5102 15896 5108
rect 15578 4924 15886 4933
rect 15578 4922 15584 4924
rect 15640 4922 15664 4924
rect 15720 4922 15744 4924
rect 15800 4922 15824 4924
rect 15880 4922 15886 4924
rect 15640 4870 15642 4922
rect 15822 4870 15824 4922
rect 15578 4868 15584 4870
rect 15640 4868 15664 4870
rect 15720 4868 15744 4870
rect 15800 4868 15824 4870
rect 15880 4868 15886 4870
rect 15578 4859 15886 4868
rect 16040 4604 16068 5120
rect 16132 4758 16160 5170
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 16120 4616 16172 4622
rect 16040 4576 16120 4604
rect 16120 4558 16172 4564
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 15578 3836 15886 3845
rect 15578 3834 15584 3836
rect 15640 3834 15664 3836
rect 15720 3834 15744 3836
rect 15800 3834 15824 3836
rect 15880 3834 15886 3836
rect 15640 3782 15642 3834
rect 15822 3782 15824 3834
rect 15578 3780 15584 3782
rect 15640 3780 15664 3782
rect 15720 3780 15744 3782
rect 15800 3780 15824 3782
rect 15880 3780 15886 3782
rect 15578 3771 15886 3780
rect 16040 3058 16068 3878
rect 16132 3534 16160 4558
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16224 3738 16252 4014
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 16132 2990 16160 3470
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 15578 2748 15886 2757
rect 15578 2746 15584 2748
rect 15640 2746 15664 2748
rect 15720 2746 15744 2748
rect 15800 2746 15824 2748
rect 15880 2746 15886 2748
rect 15640 2694 15642 2746
rect 15822 2694 15824 2746
rect 15578 2692 15584 2694
rect 15640 2692 15664 2694
rect 15720 2692 15744 2694
rect 15800 2692 15824 2694
rect 15880 2692 15886 2694
rect 15578 2683 15886 2692
rect 16132 2514 16160 2926
rect 16120 2508 16172 2514
rect 16120 2450 16172 2456
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 15936 2304 15988 2310
rect 15936 2246 15988 2252
rect 15578 1660 15886 1669
rect 15578 1658 15584 1660
rect 15640 1658 15664 1660
rect 15720 1658 15744 1660
rect 15800 1658 15824 1660
rect 15880 1658 15886 1660
rect 15640 1606 15642 1658
rect 15822 1606 15824 1658
rect 15578 1604 15584 1606
rect 15640 1604 15664 1606
rect 15720 1604 15744 1606
rect 15800 1604 15824 1606
rect 15880 1604 15886 1606
rect 15578 1595 15886 1604
rect 15948 1426 15976 2246
rect 16040 1562 16068 2382
rect 16132 1902 16160 2450
rect 16120 1896 16172 1902
rect 16120 1838 16172 1844
rect 16028 1556 16080 1562
rect 16028 1498 16080 1504
rect 16132 1426 16160 1838
rect 15936 1420 15988 1426
rect 15936 1362 15988 1368
rect 16120 1420 16172 1426
rect 16120 1362 16172 1368
rect 16224 1018 16252 2450
rect 16212 1012 16264 1018
rect 16212 954 16264 960
rect 15384 944 15436 950
rect 15384 886 15436 892
rect 15476 944 15528 950
rect 15476 886 15528 892
rect 15396 649 15424 886
rect 16316 814 16344 6734
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16408 6322 16436 6598
rect 16500 6458 16528 6802
rect 16592 6746 16620 8366
rect 16684 7993 16712 9998
rect 16868 9042 16896 10066
rect 16960 9518 16988 10542
rect 17144 10305 17172 10542
rect 17236 10470 17264 11086
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17130 10296 17186 10305
rect 17130 10231 17186 10240
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17144 9722 17172 10066
rect 17236 10062 17264 10406
rect 17224 10056 17276 10062
rect 17224 9998 17276 10004
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 17420 9518 17448 9998
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 17408 9512 17460 9518
rect 17604 9489 17632 12582
rect 17972 12306 18000 12582
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 18064 12186 18092 12242
rect 17972 12158 18092 12186
rect 17972 11898 18000 12158
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17408 9454 17460 9460
rect 17590 9480 17646 9489
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16670 7984 16726 7993
rect 16670 7919 16726 7928
rect 16670 7848 16726 7857
rect 16670 7783 16726 7792
rect 16684 7478 16712 7783
rect 16672 7472 16724 7478
rect 16672 7414 16724 7420
rect 16592 6730 16712 6746
rect 16592 6724 16724 6730
rect 16592 6718 16672 6724
rect 16672 6666 16724 6672
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16592 6338 16620 6598
rect 16670 6488 16726 6497
rect 16670 6423 16672 6432
rect 16724 6423 16726 6432
rect 16672 6394 16724 6400
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16500 6310 16620 6338
rect 16500 5914 16528 6310
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16408 4622 16436 5510
rect 16592 5030 16620 5850
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16684 5370 16712 5646
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16592 4826 16620 4966
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16394 4176 16450 4185
rect 16394 4111 16450 4120
rect 16408 4078 16436 4111
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16592 3738 16620 4762
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16500 3398 16528 3674
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16408 3058 16436 3334
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16592 2854 16620 3674
rect 16684 3602 16712 3878
rect 16672 3596 16724 3602
rect 16672 3538 16724 3544
rect 16580 2848 16632 2854
rect 16776 2825 16804 8774
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16868 7002 16896 7822
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 16960 6798 16988 9454
rect 17420 9042 17448 9454
rect 17590 9415 17646 9424
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 17328 7585 17356 8978
rect 17314 7576 17370 7585
rect 17314 7511 17370 7520
rect 17224 7200 17276 7206
rect 17222 7168 17224 7177
rect 17276 7168 17278 7177
rect 17222 7103 17278 7112
rect 16948 6792 17000 6798
rect 16868 6740 16948 6746
rect 16868 6734 17000 6740
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 16868 6718 16988 6734
rect 16868 6458 16896 6718
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16868 3369 16896 6394
rect 16948 6180 17000 6186
rect 16948 6122 17000 6128
rect 17132 6180 17184 6186
rect 17132 6122 17184 6128
rect 16960 5778 16988 6122
rect 17144 5914 17172 6122
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16946 5400 17002 5409
rect 16946 5335 16948 5344
rect 17000 5335 17002 5344
rect 16948 5306 17000 5312
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16854 3360 16910 3369
rect 16854 3295 16910 3304
rect 16960 3194 16988 4082
rect 17236 3942 17264 6734
rect 17328 6254 17356 7511
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17420 6361 17448 7278
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17512 7041 17540 7142
rect 17498 7032 17554 7041
rect 17498 6967 17554 6976
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17406 6352 17462 6361
rect 17406 6287 17462 6296
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 17328 5166 17356 6190
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17420 5234 17448 6054
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17512 4282 17540 6734
rect 17696 6458 17724 6734
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17696 4690 17724 6054
rect 17788 5137 17816 9522
rect 17880 9450 17908 10202
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 17880 9178 17908 9386
rect 18156 9382 18184 12718
rect 18616 12458 18644 12786
rect 18616 12430 18736 12458
rect 18800 12442 18828 13262
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 10266 18460 12038
rect 18708 11694 18736 12430
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18892 12374 18920 13790
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 18708 10606 18736 11630
rect 18984 11354 19012 12922
rect 19064 12776 19116 12782
rect 19168 12730 19196 13466
rect 19116 12724 19196 12730
rect 19064 12718 19196 12724
rect 19076 12702 19196 12718
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19076 11694 19104 12038
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19168 11558 19196 12702
rect 19260 12170 19288 13790
rect 19720 13410 19748 14894
rect 19904 14657 19932 14962
rect 19996 14890 20024 17439
rect 20640 16658 20668 18770
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20732 17678 20760 18158
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20732 17134 20760 17614
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20718 16144 20774 16153
rect 20824 16114 20852 18226
rect 20916 16658 20944 19858
rect 21284 19825 21312 19994
rect 21468 19922 21496 21422
rect 21732 20800 21784 20806
rect 21732 20742 21784 20748
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21560 19922 21588 20334
rect 21364 19916 21416 19922
rect 21364 19858 21416 19864
rect 21456 19916 21508 19922
rect 21456 19858 21508 19864
rect 21548 19916 21600 19922
rect 21548 19858 21600 19864
rect 21270 19816 21326 19825
rect 21270 19751 21326 19760
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21284 18766 21312 19654
rect 21376 19530 21404 19858
rect 21468 19700 21496 19858
rect 21548 19712 21600 19718
rect 21468 19672 21548 19700
rect 21548 19654 21600 19660
rect 21376 19502 21588 19530
rect 21560 19446 21588 19502
rect 21548 19440 21600 19446
rect 21548 19382 21600 19388
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21548 18760 21600 18766
rect 21548 18702 21600 18708
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20718 16079 20774 16088
rect 20812 16108 20864 16114
rect 20732 15706 20760 16079
rect 20812 16050 20864 16056
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20534 15192 20590 15201
rect 20534 15127 20590 15136
rect 20548 15026 20576 15127
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 19984 14884 20036 14890
rect 19984 14826 20036 14832
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 19890 14648 19946 14657
rect 19890 14583 19946 14592
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19812 14006 19840 14214
rect 19800 14000 19852 14006
rect 19800 13942 19852 13948
rect 19904 13870 19932 14583
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 20180 14385 20208 14418
rect 20166 14376 20222 14385
rect 20166 14311 20222 14320
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19720 13382 19840 13410
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19373 13084 19681 13093
rect 19373 13082 19379 13084
rect 19435 13082 19459 13084
rect 19515 13082 19539 13084
rect 19595 13082 19619 13084
rect 19675 13082 19681 13084
rect 19435 13030 19437 13082
rect 19617 13030 19619 13082
rect 19373 13028 19379 13030
rect 19435 13028 19459 13030
rect 19515 13028 19539 13030
rect 19595 13028 19619 13030
rect 19675 13028 19681 13030
rect 19373 13019 19681 13028
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19248 12164 19300 12170
rect 19248 12106 19300 12112
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 19168 11286 19196 11494
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19260 11132 19288 12106
rect 19444 12102 19472 12718
rect 19536 12330 19564 12718
rect 19720 12442 19748 13262
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19524 12324 19576 12330
rect 19812 12306 19840 13382
rect 20180 13326 20208 14311
rect 20272 13734 20300 14758
rect 20640 14618 20668 14962
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20732 14482 20760 14962
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20548 14249 20576 14418
rect 20626 14376 20682 14385
rect 20626 14311 20682 14320
rect 20534 14240 20590 14249
rect 20534 14175 20590 14184
rect 20640 13938 20668 14311
rect 20628 13932 20680 13938
rect 20628 13874 20680 13880
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 20168 13320 20220 13326
rect 20168 13262 20220 13268
rect 20626 13288 20682 13297
rect 20180 12306 20208 13262
rect 20626 13223 20682 13232
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 20364 12986 20392 13126
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 20640 12306 20668 13223
rect 20732 12782 20760 14418
rect 21008 14278 21036 18566
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 21086 17776 21142 17785
rect 21086 17711 21142 17720
rect 21100 16726 21128 17711
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20996 14272 21048 14278
rect 20996 14214 21048 14220
rect 20824 13870 20852 14214
rect 21192 13938 21220 18362
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21468 17678 21496 18022
rect 21456 17672 21508 17678
rect 21270 17640 21326 17649
rect 21456 17614 21508 17620
rect 21270 17575 21326 17584
rect 21284 17202 21312 17575
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21468 16998 21496 17614
rect 21560 17338 21588 18702
rect 21744 18426 21772 20742
rect 21916 20596 21968 20602
rect 21916 20538 21968 20544
rect 21824 20052 21876 20058
rect 21824 19994 21876 20000
rect 21836 19961 21864 19994
rect 21928 19990 21956 20538
rect 22112 20330 22140 21490
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 22296 21146 22324 21422
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 22284 21140 22336 21146
rect 22284 21082 22336 21088
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22100 20324 22152 20330
rect 22100 20266 22152 20272
rect 21916 19984 21968 19990
rect 21822 19952 21878 19961
rect 21916 19926 21968 19932
rect 22204 19922 22232 20742
rect 21822 19887 21878 19896
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22006 18456 22062 18465
rect 21732 18420 21784 18426
rect 21732 18362 21784 18368
rect 21928 18414 22006 18442
rect 21928 18170 21956 18414
rect 22006 18391 22062 18400
rect 22664 18290 22692 19654
rect 23032 19310 23060 21286
rect 23168 21244 23476 21253
rect 23168 21242 23174 21244
rect 23230 21242 23254 21244
rect 23310 21242 23334 21244
rect 23390 21242 23414 21244
rect 23470 21242 23476 21244
rect 23230 21190 23232 21242
rect 23412 21190 23414 21242
rect 23168 21188 23174 21190
rect 23230 21188 23254 21190
rect 23310 21188 23334 21190
rect 23390 21188 23414 21190
rect 23470 21188 23476 21190
rect 23168 21179 23476 21188
rect 23388 21140 23440 21146
rect 23388 21082 23440 21088
rect 23112 21004 23164 21010
rect 23112 20946 23164 20952
rect 23124 20330 23152 20946
rect 23400 20398 23428 21082
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23112 20324 23164 20330
rect 23112 20266 23164 20272
rect 23168 20156 23476 20165
rect 23168 20154 23174 20156
rect 23230 20154 23254 20156
rect 23310 20154 23334 20156
rect 23390 20154 23414 20156
rect 23470 20154 23476 20156
rect 23230 20102 23232 20154
rect 23412 20102 23414 20154
rect 23168 20100 23174 20102
rect 23230 20100 23254 20102
rect 23310 20100 23334 20102
rect 23390 20100 23414 20102
rect 23470 20100 23476 20102
rect 23168 20091 23476 20100
rect 23480 19780 23532 19786
rect 23480 19722 23532 19728
rect 23492 19514 23520 19722
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23480 19508 23532 19514
rect 23480 19450 23532 19456
rect 23584 19378 23612 19654
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 23020 19304 23072 19310
rect 23020 19246 23072 19252
rect 23570 19272 23626 19281
rect 22836 19236 22888 19242
rect 23570 19207 23572 19216
rect 22836 19178 22888 19184
rect 23624 19207 23626 19216
rect 23572 19178 23624 19184
rect 22848 18970 22876 19178
rect 23168 19068 23476 19077
rect 23168 19066 23174 19068
rect 23230 19066 23254 19068
rect 23310 19066 23334 19068
rect 23390 19066 23414 19068
rect 23470 19066 23476 19068
rect 23230 19014 23232 19066
rect 23412 19014 23414 19066
rect 23168 19012 23174 19014
rect 23230 19012 23254 19014
rect 23310 19012 23334 19014
rect 23390 19012 23414 19014
rect 23470 19012 23476 19014
rect 23168 19003 23476 19012
rect 23676 18970 23704 21422
rect 23848 20596 23900 20602
rect 23848 20538 23900 20544
rect 23756 20324 23808 20330
rect 23756 20266 23808 20272
rect 23768 19990 23796 20266
rect 23756 19984 23808 19990
rect 23756 19926 23808 19932
rect 23860 19825 23888 20538
rect 23952 20058 23980 21490
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 23846 19816 23902 19825
rect 23846 19751 23902 19760
rect 22836 18964 22888 18970
rect 22836 18906 22888 18912
rect 23664 18964 23716 18970
rect 23664 18906 23716 18912
rect 23860 18408 23888 19751
rect 24136 19242 24164 22034
rect 24228 21622 24256 22238
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 24216 21616 24268 21622
rect 24216 21558 24268 21564
rect 24400 21548 24452 21554
rect 24400 21490 24452 21496
rect 24412 20505 24440 21490
rect 24398 20496 24454 20505
rect 24398 20431 24454 20440
rect 24214 20224 24270 20233
rect 24214 20159 24270 20168
rect 24228 19242 24256 20159
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 24412 19514 24440 19790
rect 24400 19508 24452 19514
rect 24400 19450 24452 19456
rect 24504 19310 24532 21626
rect 24492 19304 24544 19310
rect 24492 19246 24544 19252
rect 24124 19236 24176 19242
rect 24124 19178 24176 19184
rect 24216 19236 24268 19242
rect 24216 19178 24268 19184
rect 24492 19168 24544 19174
rect 24596 19122 24624 21830
rect 25056 21486 25084 22238
rect 27620 22228 27672 22234
rect 27620 22170 27672 22176
rect 25872 22160 25924 22166
rect 25872 22102 25924 22108
rect 25688 21548 25740 21554
rect 25688 21490 25740 21496
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 25044 21480 25096 21486
rect 25044 21422 25096 21428
rect 24872 21298 24900 21422
rect 24780 21270 24900 21298
rect 25320 21344 25372 21350
rect 25320 21286 25372 21292
rect 24780 21146 24808 21270
rect 25134 21176 25190 21185
rect 24768 21140 24820 21146
rect 25332 21146 25360 21286
rect 25134 21111 25190 21120
rect 25320 21140 25372 21146
rect 24768 21082 24820 21088
rect 25148 21078 25176 21111
rect 25320 21082 25372 21088
rect 25136 21072 25188 21078
rect 25136 21014 25188 21020
rect 25148 20398 25176 21014
rect 25596 21004 25648 21010
rect 25596 20946 25648 20952
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 24768 20256 24820 20262
rect 24768 20198 24820 20204
rect 24674 20088 24730 20097
rect 24674 20023 24730 20032
rect 24544 19116 24624 19122
rect 24492 19110 24624 19116
rect 24504 19094 24624 19110
rect 24122 18864 24178 18873
rect 24122 18799 24178 18808
rect 24228 18834 24440 18850
rect 24228 18828 24452 18834
rect 24228 18822 24400 18828
rect 24136 18766 24164 18799
rect 24124 18760 24176 18766
rect 24124 18702 24176 18708
rect 24228 18612 24256 18822
rect 24400 18770 24452 18776
rect 24308 18760 24360 18766
rect 24504 18714 24532 19094
rect 24582 19000 24638 19009
rect 24582 18935 24638 18944
rect 24360 18708 24532 18714
rect 24308 18702 24532 18708
rect 24320 18686 24532 18702
rect 24228 18584 24348 18612
rect 23860 18380 24256 18408
rect 23846 18320 23902 18329
rect 22652 18284 22704 18290
rect 23846 18255 23902 18264
rect 22652 18226 22704 18232
rect 22928 18216 22980 18222
rect 21744 18142 21956 18170
rect 22926 18184 22928 18193
rect 23664 18216 23716 18222
rect 22980 18184 22982 18193
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 21548 17332 21600 17338
rect 21548 17274 21600 17280
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21468 16590 21496 16934
rect 21652 16697 21680 17818
rect 21638 16688 21694 16697
rect 21638 16623 21694 16632
rect 21272 16584 21324 16590
rect 21272 16526 21324 16532
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21284 15502 21312 16526
rect 21468 15978 21496 16526
rect 21456 15972 21508 15978
rect 21456 15914 21508 15920
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21284 14657 21312 15438
rect 21270 14648 21326 14657
rect 21270 14583 21326 14592
rect 21284 14414 21312 14583
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21376 14006 21404 15506
rect 21468 15502 21496 15914
rect 21744 15745 21772 18142
rect 23664 18158 23716 18164
rect 22926 18119 22982 18128
rect 21824 18080 21876 18086
rect 21824 18022 21876 18028
rect 22558 18048 22614 18057
rect 21836 17134 21864 18022
rect 22558 17983 22614 17992
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 21928 17377 21956 17614
rect 22008 17536 22060 17542
rect 22008 17478 22060 17484
rect 22282 17504 22338 17513
rect 21914 17368 21970 17377
rect 21914 17303 21970 17312
rect 22020 17134 22048 17478
rect 22282 17439 22338 17448
rect 22466 17504 22522 17513
rect 22466 17439 22522 17448
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 21824 17128 21876 17134
rect 21824 17070 21876 17076
rect 22008 17128 22060 17134
rect 22008 17070 22060 17076
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 22008 16992 22060 16998
rect 22112 16946 22140 17274
rect 22296 17202 22324 17439
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22480 17105 22508 17439
rect 22466 17096 22522 17105
rect 22466 17031 22522 17040
rect 22060 16940 22140 16946
rect 22008 16934 22140 16940
rect 22468 16992 22520 16998
rect 22468 16934 22520 16940
rect 21836 16590 21864 16934
rect 22020 16918 22140 16934
rect 22480 16794 22508 16934
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 21824 16584 21876 16590
rect 21824 16526 21876 16532
rect 21916 16584 21968 16590
rect 21916 16526 21968 16532
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 21822 16416 21878 16425
rect 21822 16351 21878 16360
rect 21836 16114 21864 16351
rect 21824 16108 21876 16114
rect 21824 16050 21876 16056
rect 21928 15910 21956 16526
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 21916 15904 21968 15910
rect 21916 15846 21968 15852
rect 21730 15736 21786 15745
rect 21730 15671 21786 15680
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21468 14822 21496 15438
rect 21744 14906 21772 15671
rect 21916 15496 21968 15502
rect 21916 15438 21968 15444
rect 21928 15162 21956 15438
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 22020 14929 22048 16050
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22006 14920 22062 14929
rect 21744 14878 21864 14906
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 21468 14414 21496 14758
rect 21744 14618 21772 14758
rect 21732 14612 21784 14618
rect 21732 14554 21784 14560
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 21836 13938 21864 14878
rect 22006 14855 22062 14864
rect 22100 14476 22152 14482
rect 22100 14418 22152 14424
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 19524 12266 19576 12272
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 20168 12300 20220 12306
rect 20628 12300 20680 12306
rect 20168 12242 20220 12248
rect 20548 12260 20628 12288
rect 20548 12170 20576 12260
rect 20628 12242 20680 12248
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19373 11996 19681 12005
rect 19373 11994 19379 11996
rect 19435 11994 19459 11996
rect 19515 11994 19539 11996
rect 19595 11994 19619 11996
rect 19675 11994 19681 11996
rect 19435 11942 19437 11994
rect 19617 11942 19619 11994
rect 19373 11940 19379 11942
rect 19435 11940 19459 11942
rect 19515 11940 19539 11942
rect 19595 11940 19619 11942
rect 19675 11940 19681 11942
rect 19373 11931 19681 11940
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19168 11104 19288 11132
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 19076 10606 19104 10950
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17972 7834 18000 9318
rect 18144 8968 18196 8974
rect 18524 8945 18552 10474
rect 18708 10112 18736 10542
rect 18788 10124 18840 10130
rect 18708 10084 18788 10112
rect 18788 10066 18840 10072
rect 19168 9926 19196 11104
rect 19373 10908 19681 10917
rect 19373 10906 19379 10908
rect 19435 10906 19459 10908
rect 19515 10906 19539 10908
rect 19595 10906 19619 10908
rect 19675 10906 19681 10908
rect 19435 10854 19437 10906
rect 19617 10854 19619 10906
rect 19373 10852 19379 10854
rect 19435 10852 19459 10854
rect 19515 10852 19539 10854
rect 19595 10852 19619 10854
rect 19675 10852 19681 10854
rect 19373 10843 19681 10852
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19156 9920 19208 9926
rect 19156 9862 19208 9868
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18144 8910 18196 8916
rect 18510 8936 18566 8945
rect 18156 8634 18184 8910
rect 18510 8871 18566 8880
rect 18800 8838 18828 9386
rect 19064 8900 19116 8906
rect 19064 8842 19116 8848
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 19076 8430 19104 8842
rect 19260 8634 19288 9998
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19373 9820 19681 9829
rect 19373 9818 19379 9820
rect 19435 9818 19459 9820
rect 19515 9818 19539 9820
rect 19595 9818 19619 9820
rect 19675 9818 19681 9820
rect 19435 9766 19437 9818
rect 19617 9766 19619 9818
rect 19373 9764 19379 9766
rect 19435 9764 19459 9766
rect 19515 9764 19539 9766
rect 19595 9764 19619 9766
rect 19675 9764 19681 9766
rect 19373 9755 19681 9764
rect 19720 9518 19748 9862
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19708 9512 19760 9518
rect 19708 9454 19760 9460
rect 19352 9178 19380 9454
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19812 9110 19840 11834
rect 20824 11762 20852 12650
rect 21008 12646 21036 13670
rect 22112 13326 22140 14418
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 21640 12776 21692 12782
rect 21640 12718 21692 12724
rect 20996 12640 21048 12646
rect 20996 12582 21048 12588
rect 21008 12434 21036 12582
rect 21008 12406 21128 12434
rect 21100 12306 21128 12406
rect 21284 12306 21312 12718
rect 21652 12442 21680 12718
rect 21732 12640 21784 12646
rect 21732 12582 21784 12588
rect 21744 12442 21772 12582
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 21284 11694 21312 12242
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21468 11762 21496 12038
rect 21744 11898 21772 12174
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21928 11558 21956 12378
rect 22296 11665 22324 15982
rect 22388 12102 22416 16526
rect 22466 15464 22522 15473
rect 22466 15399 22522 15408
rect 22480 15094 22508 15399
rect 22468 15088 22520 15094
rect 22468 15030 22520 15036
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22480 12442 22508 13262
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22572 12209 22600 17983
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22650 16824 22706 16833
rect 22650 16759 22652 16768
rect 22704 16759 22706 16768
rect 22652 16730 22704 16736
rect 22756 16250 22784 17478
rect 22940 16454 22968 18119
rect 23018 18048 23074 18057
rect 23018 17983 23074 17992
rect 23032 17882 23060 17983
rect 23168 17980 23476 17989
rect 23168 17978 23174 17980
rect 23230 17978 23254 17980
rect 23310 17978 23334 17980
rect 23390 17978 23414 17980
rect 23470 17978 23476 17980
rect 23230 17926 23232 17978
rect 23412 17926 23414 17978
rect 23168 17924 23174 17926
rect 23230 17924 23254 17926
rect 23310 17924 23334 17926
rect 23390 17924 23414 17926
rect 23470 17924 23476 17926
rect 23168 17915 23476 17924
rect 23020 17876 23072 17882
rect 23020 17818 23072 17824
rect 23676 17746 23704 18158
rect 23664 17740 23716 17746
rect 23664 17682 23716 17688
rect 23756 17740 23808 17746
rect 23756 17682 23808 17688
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 23032 16590 23060 17138
rect 23584 16998 23612 17614
rect 23676 17270 23704 17682
rect 23664 17264 23716 17270
rect 23664 17206 23716 17212
rect 23768 17202 23796 17682
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23664 17128 23716 17134
rect 23860 17105 23888 18255
rect 23938 18184 23994 18193
rect 23938 18119 23994 18128
rect 23664 17070 23716 17076
rect 23846 17096 23902 17105
rect 23572 16992 23624 16998
rect 23572 16934 23624 16940
rect 23168 16892 23476 16901
rect 23168 16890 23174 16892
rect 23230 16890 23254 16892
rect 23310 16890 23334 16892
rect 23390 16890 23414 16892
rect 23470 16890 23476 16892
rect 23230 16838 23232 16890
rect 23412 16838 23414 16890
rect 23168 16836 23174 16838
rect 23230 16836 23254 16838
rect 23310 16836 23334 16838
rect 23390 16836 23414 16838
rect 23470 16836 23476 16838
rect 23168 16827 23476 16836
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 23480 16584 23532 16590
rect 23584 16572 23612 16934
rect 23676 16697 23704 17070
rect 23846 17031 23902 17040
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 23860 16794 23888 16934
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23662 16688 23718 16697
rect 23662 16623 23718 16632
rect 23532 16544 23612 16572
rect 23664 16584 23716 16590
rect 23480 16526 23532 16532
rect 23664 16526 23716 16532
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 23020 16448 23072 16454
rect 23020 16390 23072 16396
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 22928 16244 22980 16250
rect 22928 16186 22980 16192
rect 22650 16144 22706 16153
rect 22650 16079 22706 16088
rect 22664 15910 22692 16079
rect 22834 16008 22890 16017
rect 22834 15943 22890 15952
rect 22652 15904 22704 15910
rect 22652 15846 22704 15852
rect 22848 15706 22876 15943
rect 22836 15700 22888 15706
rect 22836 15642 22888 15648
rect 22940 15314 22968 16186
rect 23032 15706 23060 16390
rect 23492 16046 23520 16526
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 23168 15804 23476 15813
rect 23168 15802 23174 15804
rect 23230 15802 23254 15804
rect 23310 15802 23334 15804
rect 23390 15802 23414 15804
rect 23470 15802 23476 15804
rect 23230 15750 23232 15802
rect 23412 15750 23414 15802
rect 23168 15748 23174 15750
rect 23230 15748 23254 15750
rect 23310 15748 23334 15750
rect 23390 15748 23414 15750
rect 23470 15748 23476 15750
rect 23168 15739 23476 15748
rect 23020 15700 23072 15706
rect 23020 15642 23072 15648
rect 23676 15450 23704 16526
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 23756 15972 23808 15978
rect 23756 15914 23808 15920
rect 23768 15570 23796 15914
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23860 15502 23888 15982
rect 23584 15422 23704 15450
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 22940 15286 23060 15314
rect 23032 15042 23060 15286
rect 23584 15094 23612 15422
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23754 15328 23810 15337
rect 23676 15201 23704 15302
rect 23754 15263 23810 15272
rect 23662 15192 23718 15201
rect 23662 15127 23718 15136
rect 22836 15020 22888 15026
rect 22836 14962 22888 14968
rect 22940 15014 23060 15042
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 23768 15026 23796 15263
rect 23756 15020 23808 15026
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22664 14618 22692 14758
rect 22652 14612 22704 14618
rect 22652 14554 22704 14560
rect 22848 14482 22876 14962
rect 22836 14476 22888 14482
rect 22836 14418 22888 14424
rect 22940 14414 22968 15014
rect 23756 14962 23808 14968
rect 23860 14958 23888 15438
rect 23204 14952 23256 14958
rect 23848 14952 23900 14958
rect 23256 14912 23612 14940
rect 23204 14894 23256 14900
rect 23020 14884 23072 14890
rect 23020 14826 23072 14832
rect 22928 14408 22980 14414
rect 22928 14350 22980 14356
rect 22652 13320 22704 13326
rect 22652 13262 22704 13268
rect 22664 12986 22692 13262
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22928 12844 22980 12850
rect 22928 12786 22980 12792
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22756 12374 22784 12582
rect 22744 12368 22796 12374
rect 22744 12310 22796 12316
rect 22558 12200 22614 12209
rect 22558 12135 22614 12144
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 22940 11898 22968 12786
rect 23032 12782 23060 14826
rect 23168 14716 23476 14725
rect 23168 14714 23174 14716
rect 23230 14714 23254 14716
rect 23310 14714 23334 14716
rect 23390 14714 23414 14716
rect 23470 14714 23476 14716
rect 23230 14662 23232 14714
rect 23412 14662 23414 14714
rect 23168 14660 23174 14662
rect 23230 14660 23254 14662
rect 23310 14660 23334 14662
rect 23390 14660 23414 14662
rect 23470 14660 23476 14662
rect 23168 14651 23476 14660
rect 23584 14657 23612 14912
rect 23848 14894 23900 14900
rect 23846 14784 23902 14793
rect 23768 14742 23846 14770
rect 23570 14648 23626 14657
rect 23570 14583 23626 14592
rect 23664 14612 23716 14618
rect 23296 14272 23348 14278
rect 23584 14249 23612 14583
rect 23768 14600 23796 14742
rect 23846 14719 23902 14728
rect 23716 14572 23796 14600
rect 23664 14554 23716 14560
rect 23768 14482 23796 14572
rect 23848 14612 23900 14618
rect 23848 14554 23900 14560
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 23756 14476 23808 14482
rect 23756 14418 23808 14424
rect 23296 14214 23348 14220
rect 23570 14240 23626 14249
rect 23308 14074 23336 14214
rect 23570 14175 23626 14184
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 23168 13628 23476 13637
rect 23168 13626 23174 13628
rect 23230 13626 23254 13628
rect 23310 13626 23334 13628
rect 23390 13626 23414 13628
rect 23470 13626 23476 13628
rect 23230 13574 23232 13626
rect 23412 13574 23414 13626
rect 23168 13572 23174 13574
rect 23230 13572 23254 13574
rect 23310 13572 23334 13574
rect 23390 13572 23414 13574
rect 23470 13572 23476 13574
rect 23168 13563 23476 13572
rect 23584 12986 23612 14175
rect 23676 13870 23704 14418
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23664 13388 23716 13394
rect 23664 13330 23716 13336
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23676 12782 23704 13330
rect 23020 12776 23072 12782
rect 23020 12718 23072 12724
rect 23480 12776 23532 12782
rect 23664 12776 23716 12782
rect 23532 12736 23612 12764
rect 23480 12718 23532 12724
rect 23168 12540 23476 12549
rect 23168 12538 23174 12540
rect 23230 12538 23254 12540
rect 23310 12538 23334 12540
rect 23390 12538 23414 12540
rect 23470 12538 23476 12540
rect 23230 12486 23232 12538
rect 23412 12486 23414 12538
rect 23168 12484 23174 12486
rect 23230 12484 23254 12486
rect 23310 12484 23334 12486
rect 23390 12484 23414 12486
rect 23470 12484 23476 12486
rect 23168 12475 23476 12484
rect 23296 12096 23348 12102
rect 23296 12038 23348 12044
rect 23308 11898 23336 12038
rect 22928 11892 22980 11898
rect 22928 11834 22980 11840
rect 23296 11892 23348 11898
rect 23296 11834 23348 11840
rect 23308 11694 23336 11834
rect 22928 11688 22980 11694
rect 22282 11656 22338 11665
rect 22928 11630 22980 11636
rect 23296 11688 23348 11694
rect 23296 11630 23348 11636
rect 22282 11591 22338 11600
rect 21916 11552 21968 11558
rect 21916 11494 21968 11500
rect 22376 11552 22428 11558
rect 22376 11494 22428 11500
rect 22560 11552 22612 11558
rect 22560 11494 22612 11500
rect 22388 11354 22416 11494
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 22008 11348 22060 11354
rect 22008 11290 22060 11296
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 20364 10266 20392 11290
rect 21364 11280 21416 11286
rect 21416 11240 21496 11268
rect 21364 11222 21416 11228
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 20536 10600 20588 10606
rect 20588 10548 20760 10554
rect 20536 10542 20760 10548
rect 20548 10526 20760 10542
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20444 10192 20496 10198
rect 20442 10160 20444 10169
rect 20496 10160 20498 10169
rect 19892 10124 19944 10130
rect 20442 10095 20498 10104
rect 20628 10124 20680 10130
rect 19892 10066 19944 10072
rect 20628 10066 20680 10072
rect 19800 9104 19852 9110
rect 19800 9046 19852 9052
rect 19708 8832 19760 8838
rect 19708 8774 19760 8780
rect 19373 8732 19681 8741
rect 19373 8730 19379 8732
rect 19435 8730 19459 8732
rect 19515 8730 19539 8732
rect 19595 8730 19619 8732
rect 19675 8730 19681 8732
rect 19435 8678 19437 8730
rect 19617 8678 19619 8730
rect 19373 8676 19379 8678
rect 19435 8676 19459 8678
rect 19515 8676 19539 8678
rect 19595 8676 19619 8678
rect 19675 8676 19681 8678
rect 19373 8667 19681 8676
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 18328 8288 18380 8294
rect 18328 8230 18380 8236
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 17880 7806 18000 7834
rect 17880 7342 17908 7806
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17868 7336 17920 7342
rect 17972 7313 18000 7686
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 18064 7342 18092 7414
rect 18156 7342 18184 8026
rect 18236 7472 18288 7478
rect 18340 7426 18368 8230
rect 18708 7750 18736 8366
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19168 7886 19196 8230
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18880 7744 18932 7750
rect 18880 7686 18932 7692
rect 18288 7420 18368 7426
rect 18236 7414 18368 7420
rect 18248 7398 18368 7414
rect 18340 7342 18368 7398
rect 18708 7342 18736 7686
rect 18892 7410 18920 7686
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18052 7336 18104 7342
rect 17868 7278 17920 7284
rect 17958 7304 18014 7313
rect 18052 7278 18104 7284
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18696 7336 18748 7342
rect 18984 7313 19012 7822
rect 19076 7546 19104 7822
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 19064 7404 19116 7410
rect 19168 7392 19196 7822
rect 19444 7750 19472 8366
rect 19720 7993 19748 8774
rect 19904 8090 19932 10066
rect 20640 9110 20668 10066
rect 20732 9722 20760 10526
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20824 9586 20852 11086
rect 20996 10124 21048 10130
rect 20996 10066 21048 10072
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20628 9104 20680 9110
rect 20628 9046 20680 9052
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20180 8090 20208 8910
rect 19892 8084 19944 8090
rect 20168 8084 20220 8090
rect 19944 8044 20024 8072
rect 19892 8026 19944 8032
rect 19706 7984 19762 7993
rect 19706 7919 19762 7928
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19373 7644 19681 7653
rect 19373 7642 19379 7644
rect 19435 7642 19459 7644
rect 19515 7642 19539 7644
rect 19595 7642 19619 7644
rect 19675 7642 19681 7644
rect 19435 7590 19437 7642
rect 19617 7590 19619 7642
rect 19373 7588 19379 7590
rect 19435 7588 19459 7590
rect 19515 7588 19539 7590
rect 19595 7588 19619 7590
rect 19675 7588 19681 7590
rect 19373 7579 19681 7588
rect 19116 7364 19288 7392
rect 19064 7346 19116 7352
rect 18696 7278 18748 7284
rect 18970 7304 19026 7313
rect 17958 7239 18014 7248
rect 17960 6860 18012 6866
rect 18156 6848 18184 7278
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18248 7002 18276 7142
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18012 6820 18184 6848
rect 17960 6802 18012 6808
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17972 6254 18000 6394
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 17960 6112 18012 6118
rect 17960 6054 18012 6060
rect 17972 5914 18000 6054
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 18156 5234 18184 5510
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18248 5166 18276 5510
rect 18236 5160 18288 5166
rect 17774 5128 17830 5137
rect 18236 5102 18288 5108
rect 17774 5063 17830 5072
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17972 4826 18000 5034
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 17684 4684 17736 4690
rect 17684 4626 17736 4632
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17500 4276 17552 4282
rect 17500 4218 17552 4224
rect 17880 4146 17908 4422
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16580 2790 16632 2796
rect 16762 2816 16818 2825
rect 16592 2650 16620 2790
rect 16762 2751 16818 2760
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16592 1766 16620 2586
rect 16776 2106 16804 2751
rect 16764 2100 16816 2106
rect 16764 2042 16816 2048
rect 16580 1760 16632 1766
rect 16580 1702 16632 1708
rect 16592 1562 16620 1702
rect 16580 1556 16632 1562
rect 16580 1498 16632 1504
rect 16856 876 16908 882
rect 16856 818 16908 824
rect 16304 808 16356 814
rect 16304 750 16356 756
rect 16488 808 16540 814
rect 16488 750 16540 756
rect 15382 640 15438 649
rect 15382 575 15438 584
rect 15578 572 15886 581
rect 15578 570 15584 572
rect 15640 570 15664 572
rect 15720 570 15744 572
rect 15800 570 15824 572
rect 15880 570 15886 572
rect 15640 518 15642 570
rect 15822 518 15824 570
rect 15578 516 15584 518
rect 15640 516 15664 518
rect 15720 516 15744 518
rect 15800 516 15824 518
rect 15880 516 15886 518
rect 15578 507 15886 516
rect 16500 202 16528 750
rect 16868 474 16896 818
rect 16856 468 16908 474
rect 16856 410 16908 416
rect 17052 338 17080 3878
rect 17866 3632 17922 3641
rect 17866 3567 17922 3576
rect 17880 1873 17908 3567
rect 17958 2408 18014 2417
rect 17958 2343 18014 2352
rect 17972 2106 18000 2343
rect 17960 2100 18012 2106
rect 17960 2042 18012 2048
rect 18340 2038 18368 7278
rect 18970 7239 19026 7248
rect 19260 7206 19288 7364
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 19154 6896 19210 6905
rect 19154 6831 19210 6840
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18800 6361 18828 6598
rect 18786 6352 18842 6361
rect 18786 6287 18842 6296
rect 18880 6112 18932 6118
rect 18880 6054 18932 6060
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18696 5704 18748 5710
rect 18696 5646 18748 5652
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18524 5166 18552 5646
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18524 4622 18552 5102
rect 18708 5030 18736 5646
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18696 4820 18748 4826
rect 18800 4808 18828 5646
rect 18748 4780 18828 4808
rect 18696 4762 18748 4768
rect 18892 4690 18920 6054
rect 18984 5166 19012 6734
rect 19064 6248 19116 6254
rect 19168 6236 19196 6831
rect 19260 6440 19288 7142
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19352 6662 19380 6802
rect 19996 6746 20024 8044
rect 20168 8026 20220 8032
rect 19996 6718 20208 6746
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 19373 6556 19681 6565
rect 19373 6554 19379 6556
rect 19435 6554 19459 6556
rect 19515 6554 19539 6556
rect 19595 6554 19619 6556
rect 19675 6554 19681 6556
rect 19435 6502 19437 6554
rect 19617 6502 19619 6554
rect 19373 6500 19379 6502
rect 19435 6500 19459 6502
rect 19515 6500 19539 6502
rect 19595 6500 19619 6502
rect 19675 6500 19681 6502
rect 19373 6491 19681 6500
rect 19892 6452 19944 6458
rect 19260 6412 19380 6440
rect 19352 6322 19380 6412
rect 19892 6394 19944 6400
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19248 6248 19300 6254
rect 19168 6208 19248 6236
rect 19064 6190 19116 6196
rect 19248 6190 19300 6196
rect 19076 5914 19104 6190
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 19260 5574 19288 6190
rect 19524 6180 19576 6186
rect 19524 6122 19576 6128
rect 19536 5778 19564 6122
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19248 5568 19300 5574
rect 19248 5510 19300 5516
rect 18972 5160 19024 5166
rect 18972 5102 19024 5108
rect 18972 5024 19024 5030
rect 18972 4966 19024 4972
rect 18984 4826 19012 4966
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18524 4282 18552 4558
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18524 3534 18552 4218
rect 18984 3738 19012 4762
rect 19062 3768 19118 3777
rect 18972 3732 19024 3738
rect 19062 3703 19118 3712
rect 18972 3674 19024 3680
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18524 2990 18552 3470
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 18694 2952 18750 2961
rect 18524 2446 18552 2926
rect 18694 2887 18750 2896
rect 18512 2440 18564 2446
rect 18564 2400 18644 2428
rect 18512 2382 18564 2388
rect 18328 2032 18380 2038
rect 18328 1974 18380 1980
rect 18616 1970 18644 2400
rect 18604 1964 18656 1970
rect 18604 1906 18656 1912
rect 18236 1896 18288 1902
rect 17866 1864 17922 1873
rect 18236 1838 18288 1844
rect 17866 1799 17922 1808
rect 18144 1828 18196 1834
rect 18144 1770 18196 1776
rect 17960 1760 18012 1766
rect 17960 1702 18012 1708
rect 17972 1358 18000 1702
rect 18156 1562 18184 1770
rect 18144 1556 18196 1562
rect 18144 1498 18196 1504
rect 18248 1494 18276 1838
rect 18236 1488 18288 1494
rect 18236 1430 18288 1436
rect 18616 1358 18644 1906
rect 17960 1352 18012 1358
rect 17960 1294 18012 1300
rect 18604 1352 18656 1358
rect 18604 1294 18656 1300
rect 18708 1018 18736 2887
rect 18984 2854 19012 3674
rect 18972 2848 19024 2854
rect 18972 2790 19024 2796
rect 18984 2650 19012 2790
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 18788 2440 18840 2446
rect 18786 2408 18788 2417
rect 18840 2408 18842 2417
rect 18786 2343 18842 2352
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 18800 1358 18828 2246
rect 18984 1766 19012 2586
rect 18972 1760 19024 1766
rect 18972 1702 19024 1708
rect 18984 1562 19012 1702
rect 18972 1556 19024 1562
rect 18972 1498 19024 1504
rect 18788 1352 18840 1358
rect 18788 1294 18840 1300
rect 18696 1012 18748 1018
rect 18696 954 18748 960
rect 19076 814 19104 3703
rect 19260 3534 19288 5510
rect 19373 5468 19681 5477
rect 19373 5466 19379 5468
rect 19435 5466 19459 5468
rect 19515 5466 19539 5468
rect 19595 5466 19619 5468
rect 19675 5466 19681 5468
rect 19435 5414 19437 5466
rect 19617 5414 19619 5466
rect 19373 5412 19379 5414
rect 19435 5412 19459 5414
rect 19515 5412 19539 5414
rect 19595 5412 19619 5414
rect 19675 5412 19681 5414
rect 19373 5403 19681 5412
rect 19720 5166 19748 6326
rect 19904 6254 19932 6394
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 19996 5574 20024 6190
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19708 5160 19760 5166
rect 19708 5102 19760 5108
rect 19800 4684 19852 4690
rect 19720 4644 19800 4672
rect 19373 4380 19681 4389
rect 19373 4378 19379 4380
rect 19435 4378 19459 4380
rect 19515 4378 19539 4380
rect 19595 4378 19619 4380
rect 19675 4378 19681 4380
rect 19435 4326 19437 4378
rect 19617 4326 19619 4378
rect 19373 4324 19379 4326
rect 19435 4324 19459 4326
rect 19515 4324 19539 4326
rect 19595 4324 19619 4326
rect 19675 4324 19681 4326
rect 19373 4315 19681 4324
rect 19616 4072 19668 4078
rect 19720 4060 19748 4644
rect 19800 4626 19852 4632
rect 19800 4548 19852 4554
rect 19800 4490 19852 4496
rect 19812 4078 19840 4490
rect 19996 4078 20024 5510
rect 20088 4593 20116 6598
rect 20074 4584 20130 4593
rect 20074 4519 20130 4528
rect 19668 4032 19748 4060
rect 19800 4072 19852 4078
rect 19616 4014 19668 4020
rect 19800 4014 19852 4020
rect 19984 4072 20036 4078
rect 19984 4014 20036 4020
rect 19340 3936 19392 3942
rect 19340 3878 19392 3884
rect 19352 3602 19380 3878
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19524 3392 19576 3398
rect 19628 3380 19656 4014
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19576 3352 19656 3380
rect 19524 3334 19576 3340
rect 19373 3292 19681 3301
rect 19373 3290 19379 3292
rect 19435 3290 19459 3292
rect 19515 3290 19539 3292
rect 19595 3290 19619 3292
rect 19675 3290 19681 3292
rect 19435 3238 19437 3290
rect 19617 3238 19619 3290
rect 19373 3236 19379 3238
rect 19435 3236 19459 3238
rect 19515 3236 19539 3238
rect 19595 3236 19619 3238
rect 19675 3236 19681 3238
rect 19373 3227 19681 3236
rect 19720 2990 19748 3878
rect 19996 3466 20024 4014
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 19260 1850 19288 2382
rect 20180 2310 20208 6718
rect 20456 6338 20484 8978
rect 20732 7478 20760 9522
rect 20812 9444 20864 9450
rect 20812 9386 20864 9392
rect 20824 8974 20852 9386
rect 20916 9042 20944 9862
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20902 8528 20958 8537
rect 20902 8463 20958 8472
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 20272 6322 20484 6338
rect 20260 6316 20484 6322
rect 20312 6310 20484 6316
rect 20260 6258 20312 6264
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 20364 5914 20392 6190
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20456 5710 20484 6310
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20548 4758 20576 6802
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20640 6225 20668 6734
rect 20720 6248 20772 6254
rect 20626 6216 20682 6225
rect 20720 6190 20772 6196
rect 20626 6151 20682 6160
rect 20732 5914 20760 6190
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20916 5778 20944 8463
rect 21008 8022 21036 10066
rect 21100 9722 21128 11086
rect 21364 10804 21416 10810
rect 21468 10792 21496 11240
rect 22020 11150 22048 11290
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 21416 10764 21496 10792
rect 21364 10746 21416 10752
rect 21180 10600 21232 10606
rect 21180 10542 21232 10548
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 21192 10062 21220 10542
rect 21270 10160 21326 10169
rect 21270 10095 21272 10104
rect 21324 10095 21326 10104
rect 21272 10066 21324 10072
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21376 9722 21404 10542
rect 21468 10062 21496 10764
rect 21560 10470 21588 11086
rect 22572 10606 22600 11494
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22284 10532 22336 10538
rect 22284 10474 22336 10480
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21560 9926 21588 10406
rect 21928 10130 21956 10406
rect 22296 10266 22324 10474
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22388 10130 22416 10406
rect 21916 10124 21968 10130
rect 21916 10066 21968 10072
rect 22376 10124 22428 10130
rect 22376 10066 22428 10072
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21100 9489 21128 9658
rect 21640 9512 21692 9518
rect 21086 9480 21142 9489
rect 21916 9512 21968 9518
rect 21640 9454 21692 9460
rect 21836 9472 21916 9500
rect 21086 9415 21142 9424
rect 21100 9110 21128 9415
rect 21652 9178 21680 9454
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21088 9104 21140 9110
rect 21088 9046 21140 9052
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21192 8430 21220 8842
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21362 8392 21418 8401
rect 20996 8016 21048 8022
rect 21048 7976 21128 8004
rect 20996 7958 21048 7964
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20732 5234 20760 5510
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 20536 4752 20588 4758
rect 20536 4694 20588 4700
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 20364 4146 20392 4422
rect 20824 4146 20852 5510
rect 21008 5166 21036 6054
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 20902 4720 20958 4729
rect 20902 4655 20904 4664
rect 20956 4655 20958 4664
rect 20904 4626 20956 4632
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20626 4040 20682 4049
rect 20626 3975 20682 3984
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 20168 2304 20220 2310
rect 20168 2246 20220 2252
rect 19373 2204 19681 2213
rect 19373 2202 19379 2204
rect 19435 2202 19459 2204
rect 19515 2202 19539 2204
rect 19595 2202 19619 2204
rect 19675 2202 19681 2204
rect 19435 2150 19437 2202
rect 19617 2150 19619 2202
rect 19373 2148 19379 2150
rect 19435 2148 19459 2150
rect 19515 2148 19539 2150
rect 19595 2148 19619 2150
rect 19675 2148 19681 2150
rect 19373 2139 19681 2148
rect 19260 1822 19380 1850
rect 19352 1766 19380 1822
rect 19340 1760 19392 1766
rect 19340 1702 19392 1708
rect 20180 1494 20208 2246
rect 20548 2145 20576 2450
rect 20534 2136 20590 2145
rect 20534 2071 20590 2080
rect 20444 1896 20496 1902
rect 20444 1838 20496 1844
rect 20168 1488 20220 1494
rect 20168 1430 20220 1436
rect 20074 1184 20130 1193
rect 19373 1116 19681 1125
rect 20074 1119 20130 1128
rect 19373 1114 19379 1116
rect 19435 1114 19459 1116
rect 19515 1114 19539 1116
rect 19595 1114 19619 1116
rect 19675 1114 19681 1116
rect 19435 1062 19437 1114
rect 19617 1062 19619 1114
rect 19373 1060 19379 1062
rect 19435 1060 19459 1062
rect 19515 1060 19539 1062
rect 19595 1060 19619 1062
rect 19675 1060 19681 1062
rect 19373 1051 19681 1060
rect 20088 1018 20116 1119
rect 19340 1012 19392 1018
rect 19340 954 19392 960
rect 20076 1012 20128 1018
rect 20076 954 20128 960
rect 19352 814 19380 954
rect 17132 808 17184 814
rect 19064 808 19116 814
rect 17132 750 17184 756
rect 18234 776 18290 785
rect 17144 474 17172 750
rect 19064 750 19116 756
rect 19340 808 19392 814
rect 19340 750 19392 756
rect 18234 711 18290 720
rect 18248 678 18276 711
rect 17960 672 18012 678
rect 17960 614 18012 620
rect 18236 672 18288 678
rect 18236 614 18288 620
rect 18328 672 18380 678
rect 18328 614 18380 620
rect 17132 468 17184 474
rect 17132 410 17184 416
rect 17972 338 18000 614
rect 17040 332 17092 338
rect 17040 274 17092 280
rect 17960 332 18012 338
rect 17960 274 18012 280
rect 11978 167 12034 176
rect 15108 196 15160 202
rect 15108 138 15160 144
rect 16488 196 16540 202
rect 16488 138 16540 144
rect 18340 134 18368 614
rect 19352 270 19380 750
rect 20456 746 20484 1838
rect 20640 814 20668 3975
rect 21008 3942 21036 5102
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 21008 3738 21036 3878
rect 20996 3732 21048 3738
rect 20996 3674 21048 3680
rect 21008 3602 21036 3674
rect 20996 3596 21048 3602
rect 20996 3538 21048 3544
rect 20904 3460 20956 3466
rect 20904 3402 20956 3408
rect 20916 2990 20944 3402
rect 21100 3380 21128 7976
rect 21192 7868 21220 8366
rect 21362 8327 21418 8336
rect 21376 8294 21404 8327
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21468 7886 21496 8230
rect 21272 7880 21324 7886
rect 21192 7840 21272 7868
rect 21192 7410 21220 7840
rect 21272 7822 21324 7828
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 21192 6866 21220 7346
rect 21364 7200 21416 7206
rect 21468 7188 21496 7822
rect 21416 7160 21496 7188
rect 21364 7142 21416 7148
rect 21468 7002 21496 7160
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21456 6996 21508 7002
rect 21456 6938 21508 6944
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 21284 4690 21312 6938
rect 21560 6798 21588 8570
rect 21836 8430 21864 9472
rect 21916 9454 21968 9460
rect 22008 9376 22060 9382
rect 22008 9318 22060 9324
rect 22020 9178 22048 9318
rect 22664 9178 22692 11154
rect 22940 11150 22968 11630
rect 23168 11452 23476 11461
rect 23168 11450 23174 11452
rect 23230 11450 23254 11452
rect 23310 11450 23334 11452
rect 23390 11450 23414 11452
rect 23470 11450 23476 11452
rect 23230 11398 23232 11450
rect 23412 11398 23414 11450
rect 23168 11396 23174 11398
rect 23230 11396 23254 11398
rect 23310 11396 23334 11398
rect 23390 11396 23414 11398
rect 23470 11396 23476 11398
rect 23168 11387 23476 11396
rect 23020 11280 23072 11286
rect 23020 11222 23072 11228
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 23032 10810 23060 11222
rect 23020 10804 23072 10810
rect 23020 10746 23072 10752
rect 23168 10364 23476 10373
rect 23168 10362 23174 10364
rect 23230 10362 23254 10364
rect 23310 10362 23334 10364
rect 23390 10362 23414 10364
rect 23470 10362 23476 10364
rect 23230 10310 23232 10362
rect 23412 10310 23414 10362
rect 23168 10308 23174 10310
rect 23230 10308 23254 10310
rect 23310 10308 23334 10310
rect 23390 10308 23414 10310
rect 23470 10308 23476 10310
rect 23168 10299 23476 10308
rect 23584 9674 23612 12736
rect 23664 12718 23716 12724
rect 23676 12238 23704 12718
rect 23768 12714 23796 14418
rect 23860 14074 23888 14554
rect 23952 14346 23980 18119
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 24044 14618 24072 18022
rect 24228 17270 24256 18380
rect 24124 17264 24176 17270
rect 24124 17206 24176 17212
rect 24216 17264 24268 17270
rect 24216 17206 24268 17212
rect 24136 16289 24164 17206
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 24122 16280 24178 16289
rect 24122 16215 24178 16224
rect 24228 16114 24256 16730
rect 24320 16153 24348 18584
rect 24398 18592 24454 18601
rect 24398 18527 24454 18536
rect 24412 18154 24440 18527
rect 24504 18290 24532 18686
rect 24596 18358 24624 18935
rect 24584 18352 24636 18358
rect 24584 18294 24636 18300
rect 24492 18284 24544 18290
rect 24492 18226 24544 18232
rect 24400 18148 24452 18154
rect 24400 18090 24452 18096
rect 24596 18034 24624 18294
rect 24412 18006 24624 18034
rect 24412 16561 24440 18006
rect 24584 17876 24636 17882
rect 24584 17818 24636 17824
rect 24492 17672 24544 17678
rect 24492 17614 24544 17620
rect 24504 17202 24532 17614
rect 24492 17196 24544 17202
rect 24492 17138 24544 17144
rect 24504 16794 24532 17138
rect 24492 16788 24544 16794
rect 24492 16730 24544 16736
rect 24398 16552 24454 16561
rect 24398 16487 24454 16496
rect 24306 16144 24362 16153
rect 24216 16108 24268 16114
rect 24306 16079 24362 16088
rect 24400 16108 24452 16114
rect 24216 16050 24268 16056
rect 24400 16050 24452 16056
rect 24228 15706 24256 16050
rect 24216 15700 24268 15706
rect 24136 15660 24216 15688
rect 24136 15008 24164 15660
rect 24216 15642 24268 15648
rect 24216 15496 24268 15502
rect 24412 15473 24440 16050
rect 24492 16040 24544 16046
rect 24492 15982 24544 15988
rect 24504 15706 24532 15982
rect 24492 15700 24544 15706
rect 24492 15642 24544 15648
rect 24216 15438 24268 15444
rect 24398 15464 24454 15473
rect 24228 15162 24256 15438
rect 24398 15399 24454 15408
rect 24216 15156 24268 15162
rect 24216 15098 24268 15104
rect 24216 15020 24268 15026
rect 24136 14980 24216 15008
rect 24216 14962 24268 14968
rect 24596 14906 24624 17818
rect 24688 17678 24716 20023
rect 24780 18630 24808 20198
rect 25148 20058 25176 20334
rect 25608 20233 25636 20946
rect 25700 20262 25728 21490
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25792 20602 25820 21286
rect 25780 20596 25832 20602
rect 25780 20538 25832 20544
rect 25688 20256 25740 20262
rect 25594 20224 25650 20233
rect 25688 20198 25740 20204
rect 25594 20159 25650 20168
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 25148 19230 25636 19258
rect 25148 19174 25176 19230
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 25504 19168 25556 19174
rect 25504 19110 25556 19116
rect 24860 18760 24912 18766
rect 24860 18702 24912 18708
rect 24872 18630 24900 18702
rect 24768 18624 24820 18630
rect 24768 18566 24820 18572
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 24860 18216 24912 18222
rect 24912 18164 24992 18170
rect 24860 18158 24992 18164
rect 24768 18148 24820 18154
rect 24872 18142 24992 18158
rect 24768 18090 24820 18096
rect 24780 17882 24808 18090
rect 24858 18048 24914 18057
rect 24858 17983 24914 17992
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 24872 17678 24900 17983
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 24688 16425 24716 17206
rect 24860 17128 24912 17134
rect 24964 17116 24992 18142
rect 25056 17678 25084 18226
rect 25044 17672 25096 17678
rect 25044 17614 25096 17620
rect 24912 17088 24992 17116
rect 24860 17070 24912 17076
rect 24964 16726 24992 17088
rect 24952 16720 25004 16726
rect 24952 16662 25004 16668
rect 24674 16416 24730 16425
rect 24674 16351 24730 16360
rect 24688 15881 24716 16351
rect 24858 16008 24914 16017
rect 25148 15994 25176 19110
rect 25228 18964 25280 18970
rect 25228 18906 25280 18912
rect 25320 18964 25372 18970
rect 25320 18906 25372 18912
rect 25240 18766 25268 18906
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 25240 17202 25268 18022
rect 25332 17202 25360 18906
rect 25516 18714 25544 19110
rect 25608 18902 25636 19230
rect 25596 18896 25648 18902
rect 25596 18838 25648 18844
rect 25686 18864 25742 18873
rect 25686 18799 25742 18808
rect 25516 18698 25636 18714
rect 25516 18692 25648 18698
rect 25516 18686 25596 18692
rect 25516 18222 25544 18686
rect 25596 18634 25648 18640
rect 25504 18216 25556 18222
rect 25504 18158 25556 18164
rect 25504 17536 25556 17542
rect 25504 17478 25556 17484
rect 25516 17202 25544 17478
rect 25594 17368 25650 17377
rect 25594 17303 25650 17312
rect 25228 17196 25280 17202
rect 25228 17138 25280 17144
rect 25320 17196 25372 17202
rect 25320 17138 25372 17144
rect 25504 17196 25556 17202
rect 25504 17138 25556 17144
rect 25240 16726 25268 17138
rect 25608 16998 25636 17303
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25228 16720 25280 16726
rect 25228 16662 25280 16668
rect 25700 16590 25728 18799
rect 25884 18714 25912 22102
rect 25964 21888 26016 21894
rect 25964 21830 26016 21836
rect 25976 21690 26004 21830
rect 26963 21788 27271 21797
rect 26963 21786 26969 21788
rect 27025 21786 27049 21788
rect 27105 21786 27129 21788
rect 27185 21786 27209 21788
rect 27265 21786 27271 21788
rect 27025 21734 27027 21786
rect 27207 21734 27209 21786
rect 26963 21732 26969 21734
rect 27025 21732 27049 21734
rect 27105 21732 27129 21734
rect 27185 21732 27209 21734
rect 27265 21732 27271 21734
rect 26963 21723 27271 21732
rect 25964 21684 26016 21690
rect 25964 21626 26016 21632
rect 26792 21548 26844 21554
rect 26792 21490 26844 21496
rect 26332 21480 26384 21486
rect 26332 21422 26384 21428
rect 26056 21072 26108 21078
rect 26056 21014 26108 21020
rect 26068 20641 26096 21014
rect 26148 21004 26200 21010
rect 26148 20946 26200 20952
rect 26054 20632 26110 20641
rect 26054 20567 26110 20576
rect 25964 19848 26016 19854
rect 25964 19790 26016 19796
rect 25976 18834 26004 19790
rect 26056 19168 26108 19174
rect 26056 19110 26108 19116
rect 25964 18828 26016 18834
rect 25964 18770 26016 18776
rect 25792 18686 25912 18714
rect 25688 16584 25740 16590
rect 25688 16526 25740 16532
rect 24914 15966 25176 15994
rect 24858 15943 24914 15952
rect 24674 15872 24730 15881
rect 24674 15807 24730 15816
rect 25502 15600 25558 15609
rect 24676 15564 24728 15570
rect 25502 15535 25558 15544
rect 24676 15506 24728 15512
rect 24688 15065 24716 15506
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24674 15056 24730 15065
rect 24674 14991 24730 15000
rect 24596 14878 24808 14906
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 24032 14408 24084 14414
rect 24032 14350 24084 14356
rect 23940 14340 23992 14346
rect 23940 14282 23992 14288
rect 24044 14074 24072 14350
rect 24228 14113 24256 14758
rect 24400 14612 24452 14618
rect 24400 14554 24452 14560
rect 24214 14104 24270 14113
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 24032 14068 24084 14074
rect 24084 14028 24164 14056
rect 24214 14039 24270 14048
rect 24032 14010 24084 14016
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23860 13705 23888 13874
rect 23938 13832 23994 13841
rect 23938 13767 23994 13776
rect 23846 13696 23902 13705
rect 23846 13631 23902 13640
rect 23848 12980 23900 12986
rect 23848 12922 23900 12928
rect 23756 12708 23808 12714
rect 23756 12650 23808 12656
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23860 11694 23888 12922
rect 23952 12753 23980 13767
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 23938 12744 23994 12753
rect 23938 12679 23994 12688
rect 24044 12628 24072 13466
rect 24136 13326 24164 14028
rect 24412 13938 24440 14554
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24124 13320 24176 13326
rect 24124 13262 24176 13268
rect 24124 13184 24176 13190
rect 24308 13184 24360 13190
rect 24176 13132 24256 13138
rect 24124 13126 24256 13132
rect 24308 13126 24360 13132
rect 24136 13110 24256 13126
rect 24124 12640 24176 12646
rect 24044 12600 24124 12628
rect 24124 12582 24176 12588
rect 24136 12442 24164 12582
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24228 12306 24256 13110
rect 24216 12300 24268 12306
rect 24216 12242 24268 12248
rect 24216 12096 24268 12102
rect 24216 12038 24268 12044
rect 23940 11892 23992 11898
rect 23992 11852 24072 11880
rect 23940 11834 23992 11840
rect 23848 11688 23900 11694
rect 23676 11648 23848 11676
rect 23676 10538 23704 11648
rect 23848 11630 23900 11636
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 23952 11558 23980 11630
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 24044 11150 24072 11852
rect 24228 11694 24256 12038
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 24320 11257 24348 13126
rect 24504 12986 24532 14350
rect 24676 14272 24728 14278
rect 24676 14214 24728 14220
rect 24688 13938 24716 14214
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24492 12980 24544 12986
rect 24492 12922 24544 12928
rect 24596 12442 24624 13874
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24584 12436 24636 12442
rect 24584 12378 24636 12384
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24306 11248 24362 11257
rect 24306 11183 24362 11192
rect 23848 11144 23900 11150
rect 23846 11112 23848 11121
rect 23940 11144 23992 11150
rect 23900 11112 23902 11121
rect 23940 11086 23992 11092
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 23846 11047 23902 11056
rect 23756 11008 23808 11014
rect 23756 10950 23808 10956
rect 23768 10674 23796 10950
rect 23756 10668 23808 10674
rect 23756 10610 23808 10616
rect 23664 10532 23716 10538
rect 23664 10474 23716 10480
rect 23756 10532 23808 10538
rect 23756 10474 23808 10480
rect 23768 10169 23796 10474
rect 23952 10266 23980 11086
rect 23940 10260 23992 10266
rect 23940 10202 23992 10208
rect 23754 10160 23810 10169
rect 23754 10095 23810 10104
rect 23584 9646 23704 9674
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22020 9081 22048 9114
rect 22006 9072 22062 9081
rect 22006 9007 22062 9016
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22466 8800 22522 8809
rect 22466 8735 22522 8744
rect 21824 8424 21876 8430
rect 22284 8424 22336 8430
rect 21824 8366 21876 8372
rect 22282 8392 22284 8401
rect 22336 8392 22338 8401
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21456 6112 21508 6118
rect 21456 6054 21508 6060
rect 21468 5778 21496 6054
rect 21560 5817 21588 6734
rect 21652 6458 21680 7278
rect 21836 6497 21864 8366
rect 22282 8327 22338 8336
rect 22480 8090 22508 8735
rect 22664 8090 22692 8910
rect 22468 8084 22520 8090
rect 22468 8026 22520 8032
rect 22652 8084 22704 8090
rect 22652 8026 22704 8032
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 21928 6866 21956 7142
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 21822 6488 21878 6497
rect 21640 6452 21692 6458
rect 22572 6458 22600 6734
rect 21822 6423 21878 6432
rect 22560 6452 22612 6458
rect 21640 6394 21692 6400
rect 21546 5808 21602 5817
rect 21456 5772 21508 5778
rect 21836 5778 21864 6423
rect 22560 6394 22612 6400
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22572 5778 22600 6054
rect 21546 5743 21602 5752
rect 21824 5772 21876 5778
rect 21456 5714 21508 5720
rect 21824 5714 21876 5720
rect 22560 5772 22612 5778
rect 22560 5714 22612 5720
rect 21916 5704 21968 5710
rect 21916 5646 21968 5652
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 21456 5636 21508 5642
rect 21456 5578 21508 5584
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21376 4486 21404 5306
rect 21468 5234 21496 5578
rect 21548 5364 21600 5370
rect 21548 5306 21600 5312
rect 21456 5228 21508 5234
rect 21456 5170 21508 5176
rect 21456 4684 21508 4690
rect 21456 4626 21508 4632
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21008 3352 21128 3380
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 20916 2650 20944 2926
rect 20904 2644 20956 2650
rect 20904 2586 20956 2592
rect 20720 2100 20772 2106
rect 20720 2042 20772 2048
rect 21008 2088 21036 3352
rect 21284 2990 21312 4422
rect 21272 2984 21324 2990
rect 21272 2926 21324 2932
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21364 2508 21416 2514
rect 21468 2496 21496 4626
rect 21560 4282 21588 5306
rect 21928 5166 21956 5646
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 21640 4752 21692 4758
rect 21640 4694 21692 4700
rect 21652 4282 21680 4694
rect 21928 4690 21956 5102
rect 21916 4684 21968 4690
rect 21916 4626 21968 4632
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 21824 4480 21876 4486
rect 22020 4457 22048 4558
rect 21824 4422 21876 4428
rect 22006 4448 22062 4457
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21548 3732 21600 3738
rect 21548 3674 21600 3680
rect 21560 2854 21588 3674
rect 21836 3602 21864 4422
rect 22006 4383 22062 4392
rect 22204 4214 22232 4558
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22192 4208 22244 4214
rect 22296 4185 22324 4422
rect 22192 4150 22244 4156
rect 22282 4176 22338 4185
rect 22388 4146 22416 5646
rect 22560 5568 22612 5574
rect 22664 5545 22692 7822
rect 22756 7546 22784 9522
rect 23572 9376 23624 9382
rect 23572 9318 23624 9324
rect 23168 9276 23476 9285
rect 23168 9274 23174 9276
rect 23230 9274 23254 9276
rect 23310 9274 23334 9276
rect 23390 9274 23414 9276
rect 23470 9274 23476 9276
rect 23230 9222 23232 9274
rect 23412 9222 23414 9274
rect 23168 9220 23174 9222
rect 23230 9220 23254 9222
rect 23310 9220 23334 9222
rect 23390 9220 23414 9222
rect 23470 9220 23476 9222
rect 23168 9211 23476 9220
rect 23584 9178 23612 9318
rect 23572 9172 23624 9178
rect 23572 9114 23624 9120
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23492 8498 23520 8774
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23168 8188 23476 8197
rect 23168 8186 23174 8188
rect 23230 8186 23254 8188
rect 23310 8186 23334 8188
rect 23390 8186 23414 8188
rect 23470 8186 23476 8188
rect 23230 8134 23232 8186
rect 23412 8134 23414 8186
rect 23168 8132 23174 8134
rect 23230 8132 23254 8134
rect 23310 8132 23334 8134
rect 23390 8132 23414 8134
rect 23470 8132 23476 8134
rect 23168 8123 23476 8132
rect 23584 8090 23612 8230
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 22836 7880 22888 7886
rect 22836 7822 22888 7828
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 22848 7750 22876 7822
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 23216 7274 23244 7822
rect 23204 7268 23256 7274
rect 23204 7210 23256 7216
rect 23572 7268 23624 7274
rect 23572 7210 23624 7216
rect 23168 7100 23476 7109
rect 23168 7098 23174 7100
rect 23230 7098 23254 7100
rect 23310 7098 23334 7100
rect 23390 7098 23414 7100
rect 23470 7098 23476 7100
rect 23230 7046 23232 7098
rect 23412 7046 23414 7098
rect 23168 7044 23174 7046
rect 23230 7044 23254 7046
rect 23310 7044 23334 7046
rect 23390 7044 23414 7046
rect 23470 7044 23476 7046
rect 23168 7035 23476 7044
rect 23584 6798 23612 7210
rect 23676 7154 23704 9646
rect 23940 9376 23992 9382
rect 23940 9318 23992 9324
rect 23756 9172 23808 9178
rect 23756 9114 23808 9120
rect 23768 9081 23796 9114
rect 23754 9072 23810 9081
rect 23754 9007 23810 9016
rect 23768 8362 23796 9007
rect 23952 8430 23980 9318
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 23940 8424 23992 8430
rect 23940 8366 23992 8372
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23860 7342 23888 8366
rect 24044 8242 24072 11086
rect 24412 10674 24440 11698
rect 24688 11558 24716 12582
rect 24780 11801 24808 14878
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24872 13705 24900 14418
rect 24964 13938 24992 15098
rect 25042 14104 25098 14113
rect 25042 14039 25098 14048
rect 24952 13932 25004 13938
rect 24952 13874 25004 13880
rect 24858 13696 24914 13705
rect 24858 13631 24914 13640
rect 24872 12782 24900 13631
rect 24964 12850 24992 13874
rect 25056 13326 25084 14039
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 24952 12844 25004 12850
rect 24952 12786 25004 12792
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 25516 12102 25544 15535
rect 25688 14816 25740 14822
rect 25688 14758 25740 14764
rect 25700 14385 25728 14758
rect 25686 14376 25742 14385
rect 25686 14311 25742 14320
rect 25504 12096 25556 12102
rect 25504 12038 25556 12044
rect 24766 11792 24822 11801
rect 24766 11727 24822 11736
rect 25320 11688 25372 11694
rect 25320 11630 25372 11636
rect 24676 11552 24728 11558
rect 24676 11494 24728 11500
rect 25332 11354 25360 11630
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25596 11212 25648 11218
rect 25596 11154 25648 11160
rect 24400 10668 24452 10674
rect 24400 10610 24452 10616
rect 25320 10668 25372 10674
rect 25320 10610 25372 10616
rect 25332 10470 25360 10610
rect 25320 10464 25372 10470
rect 25320 10406 25372 10412
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24124 10056 24176 10062
rect 24124 9998 24176 10004
rect 24136 9518 24164 9998
rect 24124 9512 24176 9518
rect 24122 9480 24124 9489
rect 24176 9480 24178 9489
rect 24122 9415 24178 9424
rect 24136 9178 24164 9415
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 24228 8537 24256 10202
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 24872 9722 24900 9998
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24860 9716 24912 9722
rect 24860 9658 24912 9664
rect 24492 9648 24544 9654
rect 24492 9590 24544 9596
rect 24308 9512 24360 9518
rect 24308 9454 24360 9460
rect 24214 8528 24270 8537
rect 24214 8463 24270 8472
rect 23952 8214 24072 8242
rect 24216 8288 24268 8294
rect 24216 8230 24268 8236
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 23676 7126 23888 7154
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23216 6458 23244 6734
rect 23204 6452 23256 6458
rect 23204 6394 23256 6400
rect 22836 6384 22888 6390
rect 22836 6326 22888 6332
rect 22848 6254 22876 6326
rect 22836 6248 22888 6254
rect 22836 6190 22888 6196
rect 22744 6112 22796 6118
rect 22744 6054 22796 6060
rect 23756 6112 23808 6118
rect 23756 6054 23808 6060
rect 22756 5574 22784 6054
rect 23168 6012 23476 6021
rect 23168 6010 23174 6012
rect 23230 6010 23254 6012
rect 23310 6010 23334 6012
rect 23390 6010 23414 6012
rect 23470 6010 23476 6012
rect 23230 5958 23232 6010
rect 23412 5958 23414 6010
rect 23168 5956 23174 5958
rect 23230 5956 23254 5958
rect 23310 5956 23334 5958
rect 23390 5956 23414 5958
rect 23470 5956 23476 5958
rect 23168 5947 23476 5956
rect 22928 5908 22980 5914
rect 22928 5850 22980 5856
rect 23388 5908 23440 5914
rect 23388 5850 23440 5856
rect 22744 5568 22796 5574
rect 22560 5510 22612 5516
rect 22650 5536 22706 5545
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 22480 4690 22508 4966
rect 22572 4690 22600 5510
rect 22744 5510 22796 5516
rect 22650 5471 22706 5480
rect 22940 5030 22968 5850
rect 23400 5273 23428 5850
rect 23572 5704 23624 5710
rect 23570 5672 23572 5681
rect 23624 5672 23626 5681
rect 23570 5607 23626 5616
rect 23386 5264 23442 5273
rect 23386 5199 23442 5208
rect 23662 5264 23718 5273
rect 23768 5234 23796 6054
rect 23662 5199 23718 5208
rect 23756 5228 23808 5234
rect 23676 5098 23704 5199
rect 23756 5170 23808 5176
rect 23664 5092 23716 5098
rect 23664 5034 23716 5040
rect 23756 5092 23808 5098
rect 23756 5034 23808 5040
rect 22928 5024 22980 5030
rect 22928 4966 22980 4972
rect 22468 4684 22520 4690
rect 22468 4626 22520 4632
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 22834 4448 22890 4457
rect 22834 4383 22890 4392
rect 22848 4214 22876 4383
rect 22836 4208 22888 4214
rect 22836 4150 22888 4156
rect 22282 4111 22338 4120
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 22940 4078 22968 4966
rect 23168 4924 23476 4933
rect 23168 4922 23174 4924
rect 23230 4922 23254 4924
rect 23310 4922 23334 4924
rect 23390 4922 23414 4924
rect 23470 4922 23476 4924
rect 23230 4870 23232 4922
rect 23412 4870 23414 4922
rect 23168 4868 23174 4870
rect 23230 4868 23254 4870
rect 23310 4868 23334 4870
rect 23390 4868 23414 4870
rect 23470 4868 23476 4870
rect 23168 4859 23476 4868
rect 23572 4276 23624 4282
rect 23572 4218 23624 4224
rect 22652 4072 22704 4078
rect 22652 4014 22704 4020
rect 22928 4072 22980 4078
rect 22928 4014 22980 4020
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 22664 2990 22692 4014
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22848 3738 22876 3878
rect 22940 3738 22968 4014
rect 23168 3836 23476 3845
rect 23168 3834 23174 3836
rect 23230 3834 23254 3836
rect 23310 3834 23334 3836
rect 23390 3834 23414 3836
rect 23470 3834 23476 3836
rect 23230 3782 23232 3834
rect 23412 3782 23414 3834
rect 23168 3780 23174 3782
rect 23230 3780 23254 3782
rect 23310 3780 23334 3782
rect 23390 3780 23414 3782
rect 23470 3780 23476 3782
rect 23168 3771 23476 3780
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 22928 3732 22980 3738
rect 22928 3674 22980 3680
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 22742 3088 22798 3097
rect 23308 3058 23336 3334
rect 22742 3023 22798 3032
rect 23296 3052 23348 3058
rect 22652 2984 22704 2990
rect 22652 2926 22704 2932
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 21560 2650 21588 2790
rect 21548 2644 21600 2650
rect 21548 2586 21600 2592
rect 21416 2468 21496 2496
rect 21364 2450 21416 2456
rect 21088 2100 21140 2106
rect 21008 2060 21088 2088
rect 20732 814 20760 2042
rect 20812 1760 20864 1766
rect 20812 1702 20864 1708
rect 20824 1426 20852 1702
rect 21008 1562 21036 2060
rect 21088 2042 21140 2048
rect 21192 1902 21220 2450
rect 21180 1896 21232 1902
rect 21180 1838 21232 1844
rect 20996 1556 21048 1562
rect 20996 1498 21048 1504
rect 21008 1426 21036 1498
rect 21192 1426 21220 1838
rect 20812 1420 20864 1426
rect 20812 1362 20864 1368
rect 20996 1420 21048 1426
rect 20996 1362 21048 1368
rect 21180 1420 21232 1426
rect 21180 1362 21232 1368
rect 21376 882 21404 2450
rect 21456 2304 21508 2310
rect 21456 2246 21508 2252
rect 21468 1970 21496 2246
rect 21456 1964 21508 1970
rect 21456 1906 21508 1912
rect 21560 1766 21588 2586
rect 22008 2440 22060 2446
rect 22060 2400 22416 2428
rect 22008 2382 22060 2388
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 21548 1760 21600 1766
rect 21548 1702 21600 1708
rect 21560 1562 21588 1702
rect 21548 1556 21600 1562
rect 21548 1498 21600 1504
rect 21916 1352 21968 1358
rect 21916 1294 21968 1300
rect 21928 882 21956 1294
rect 22204 882 22232 2246
rect 22388 2106 22416 2400
rect 22376 2100 22428 2106
rect 22376 2042 22428 2048
rect 22652 1896 22704 1902
rect 22652 1838 22704 1844
rect 22664 1465 22692 1838
rect 22650 1456 22706 1465
rect 22650 1391 22706 1400
rect 22756 1018 22784 3023
rect 23296 2994 23348 3000
rect 23168 2748 23476 2757
rect 23168 2746 23174 2748
rect 23230 2746 23254 2748
rect 23310 2746 23334 2748
rect 23390 2746 23414 2748
rect 23470 2746 23476 2748
rect 23230 2694 23232 2746
rect 23412 2694 23414 2746
rect 23168 2692 23174 2694
rect 23230 2692 23254 2694
rect 23310 2692 23334 2694
rect 23390 2692 23414 2694
rect 23470 2692 23476 2694
rect 23168 2683 23476 2692
rect 22928 2372 22980 2378
rect 22928 2314 22980 2320
rect 22836 1760 22888 1766
rect 22836 1702 22888 1708
rect 22848 1358 22876 1702
rect 22836 1352 22888 1358
rect 22836 1294 22888 1300
rect 22652 1012 22704 1018
rect 22652 954 22704 960
rect 22744 1012 22796 1018
rect 22744 954 22796 960
rect 21364 876 21416 882
rect 21364 818 21416 824
rect 21916 876 21968 882
rect 21916 818 21968 824
rect 22192 876 22244 882
rect 22192 818 22244 824
rect 22664 814 22692 954
rect 22940 882 22968 2314
rect 23584 2258 23612 4218
rect 23768 4162 23796 5034
rect 23860 4978 23888 7126
rect 23952 5098 23980 8214
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 24044 6934 24072 7346
rect 24228 7206 24256 8230
rect 24216 7200 24268 7206
rect 24216 7142 24268 7148
rect 24032 6928 24084 6934
rect 24032 6870 24084 6876
rect 24320 6390 24348 9454
rect 24400 9376 24452 9382
rect 24400 9318 24452 9324
rect 24412 7410 24440 9318
rect 24504 9042 24532 9590
rect 24964 9518 24992 9862
rect 24952 9512 25004 9518
rect 24952 9454 25004 9460
rect 24584 9444 24636 9450
rect 24584 9386 24636 9392
rect 24492 9036 24544 9042
rect 24492 8978 24544 8984
rect 24596 8838 24624 9386
rect 24964 8906 24992 9454
rect 24952 8900 25004 8906
rect 24952 8842 25004 8848
rect 24584 8832 24636 8838
rect 24584 8774 24636 8780
rect 25056 7546 25084 9998
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25240 9178 25268 9454
rect 25228 9172 25280 9178
rect 25228 9114 25280 9120
rect 25320 8968 25372 8974
rect 25320 8910 25372 8916
rect 25228 8288 25280 8294
rect 25228 8230 25280 8236
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 24688 7206 24716 7482
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 24964 7002 24992 7346
rect 25044 7336 25096 7342
rect 25044 7278 25096 7284
rect 25056 7041 25084 7278
rect 25042 7032 25098 7041
rect 24860 6996 24912 7002
rect 24860 6938 24912 6944
rect 24952 6996 25004 7002
rect 25042 6967 25098 6976
rect 24952 6938 25004 6944
rect 24492 6656 24544 6662
rect 24492 6598 24544 6604
rect 24398 6488 24454 6497
rect 24398 6423 24454 6432
rect 24412 6390 24440 6423
rect 24308 6384 24360 6390
rect 24308 6326 24360 6332
rect 24400 6384 24452 6390
rect 24400 6326 24452 6332
rect 24504 6322 24532 6598
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 24044 5234 24072 6258
rect 24872 6118 24900 6938
rect 25044 6316 25096 6322
rect 25044 6258 25096 6264
rect 24492 6112 24544 6118
rect 24492 6054 24544 6060
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24860 6112 24912 6118
rect 24860 6054 24912 6060
rect 24400 5772 24452 5778
rect 24400 5714 24452 5720
rect 24124 5636 24176 5642
rect 24124 5578 24176 5584
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 23940 5092 23992 5098
rect 23940 5034 23992 5040
rect 23860 4950 23980 4978
rect 23676 4134 23796 4162
rect 23676 2514 23704 4134
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 23768 2990 23796 3470
rect 23860 3126 23888 3470
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 23756 2984 23808 2990
rect 23756 2926 23808 2932
rect 23664 2508 23716 2514
rect 23664 2450 23716 2456
rect 23492 2230 23612 2258
rect 23662 2272 23718 2281
rect 23492 2106 23520 2230
rect 23662 2207 23718 2216
rect 23480 2100 23532 2106
rect 23480 2042 23532 2048
rect 23676 2038 23704 2207
rect 23664 2032 23716 2038
rect 23664 1974 23716 1980
rect 23480 1964 23532 1970
rect 23480 1906 23532 1912
rect 23492 1850 23520 1906
rect 23768 1902 23796 2926
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 23860 2582 23888 2790
rect 23848 2576 23900 2582
rect 23848 2518 23900 2524
rect 23952 2514 23980 4950
rect 24032 4616 24084 4622
rect 24136 4570 24164 5578
rect 24412 4622 24440 5714
rect 24504 4672 24532 6054
rect 24780 5778 24808 6054
rect 24768 5772 24820 5778
rect 24768 5714 24820 5720
rect 24676 5704 24728 5710
rect 24674 5672 24676 5681
rect 24728 5672 24730 5681
rect 24674 5607 24730 5616
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24688 5234 24716 5306
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 24584 4684 24636 4690
rect 24504 4644 24584 4672
rect 24584 4626 24636 4632
rect 24084 4564 24164 4570
rect 24032 4558 24164 4564
rect 24400 4616 24452 4622
rect 24400 4558 24452 4564
rect 24044 4542 24164 4558
rect 24136 4468 24164 4542
rect 24136 4440 24256 4468
rect 24228 4282 24256 4440
rect 24216 4276 24268 4282
rect 24216 4218 24268 4224
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 23848 2304 23900 2310
rect 23848 2246 23900 2252
rect 23756 1896 23808 1902
rect 23020 1828 23072 1834
rect 23492 1822 23704 1850
rect 23756 1838 23808 1844
rect 23020 1770 23072 1776
rect 23032 1562 23060 1770
rect 23572 1760 23624 1766
rect 23572 1702 23624 1708
rect 23168 1660 23476 1669
rect 23168 1658 23174 1660
rect 23230 1658 23254 1660
rect 23310 1658 23334 1660
rect 23390 1658 23414 1660
rect 23470 1658 23476 1660
rect 23230 1606 23232 1658
rect 23412 1606 23414 1658
rect 23168 1604 23174 1606
rect 23230 1604 23254 1606
rect 23310 1604 23334 1606
rect 23390 1604 23414 1606
rect 23470 1604 23476 1606
rect 23168 1595 23476 1604
rect 23020 1556 23072 1562
rect 23020 1498 23072 1504
rect 23480 1352 23532 1358
rect 23584 1340 23612 1702
rect 23532 1312 23612 1340
rect 23480 1294 23532 1300
rect 23676 950 23704 1822
rect 23756 1760 23808 1766
rect 23756 1702 23808 1708
rect 23768 1562 23796 1702
rect 23860 1562 23888 2246
rect 23940 1760 23992 1766
rect 23940 1702 23992 1708
rect 23756 1556 23808 1562
rect 23756 1498 23808 1504
rect 23848 1556 23900 1562
rect 23848 1498 23900 1504
rect 23756 1420 23808 1426
rect 23952 1408 23980 1702
rect 23808 1380 23980 1408
rect 23756 1362 23808 1368
rect 23664 944 23716 950
rect 23664 886 23716 892
rect 22928 876 22980 882
rect 22928 818 22980 824
rect 20628 808 20680 814
rect 20628 750 20680 756
rect 20720 808 20772 814
rect 21456 808 21508 814
rect 20720 750 20772 756
rect 21454 776 21456 785
rect 22652 808 22704 814
rect 21508 776 21510 785
rect 20444 740 20496 746
rect 22652 750 22704 756
rect 21454 711 21510 720
rect 20444 682 20496 688
rect 23768 678 23796 1362
rect 24044 950 24072 3878
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 24136 2854 24164 3674
rect 24124 2848 24176 2854
rect 24124 2790 24176 2796
rect 24136 1766 24164 2790
rect 24228 2514 24256 4218
rect 24412 4026 24440 4558
rect 24582 4448 24638 4457
rect 24582 4383 24638 4392
rect 24412 3998 24532 4026
rect 24504 3942 24532 3998
rect 24400 3936 24452 3942
rect 24400 3878 24452 3884
rect 24492 3936 24544 3942
rect 24492 3878 24544 3884
rect 24412 3058 24440 3878
rect 24504 3602 24532 3878
rect 24596 3738 24624 4383
rect 24780 4146 24808 5306
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 24858 4720 24914 4729
rect 24858 4655 24860 4664
rect 24912 4655 24914 4664
rect 24860 4626 24912 4632
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 24688 4026 24716 4082
rect 24964 4026 24992 4966
rect 24688 3998 24992 4026
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 24492 3596 24544 3602
rect 24492 3538 24544 3544
rect 24400 3052 24452 3058
rect 24400 2994 24452 3000
rect 24216 2508 24268 2514
rect 24216 2450 24268 2456
rect 24124 1760 24176 1766
rect 24124 1702 24176 1708
rect 24124 1556 24176 1562
rect 24124 1498 24176 1504
rect 24136 1426 24164 1498
rect 24124 1420 24176 1426
rect 24124 1362 24176 1368
rect 24032 944 24084 950
rect 24032 886 24084 892
rect 23940 808 23992 814
rect 23938 776 23940 785
rect 24124 808 24176 814
rect 23992 776 23994 785
rect 24228 796 24256 2450
rect 24504 2446 24532 3538
rect 24676 2848 24728 2854
rect 24676 2790 24728 2796
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 24306 2136 24362 2145
rect 24306 2071 24362 2080
rect 24320 1562 24348 2071
rect 24308 1556 24360 1562
rect 24308 1498 24360 1504
rect 24306 1456 24362 1465
rect 24306 1391 24308 1400
rect 24360 1391 24362 1400
rect 24308 1362 24360 1368
rect 24176 768 24256 796
rect 24124 750 24176 756
rect 23938 711 23994 720
rect 23756 672 23808 678
rect 23756 614 23808 620
rect 23940 672 23992 678
rect 23940 614 23992 620
rect 23168 572 23476 581
rect 23168 570 23174 572
rect 23230 570 23254 572
rect 23310 570 23334 572
rect 23390 570 23414 572
rect 23470 570 23476 572
rect 23230 518 23232 570
rect 23412 518 23414 570
rect 23168 516 23174 518
rect 23230 516 23254 518
rect 23310 516 23334 518
rect 23390 516 23414 518
rect 23470 516 23476 518
rect 23168 507 23476 516
rect 23952 338 23980 614
rect 23940 332 23992 338
rect 23940 274 23992 280
rect 19340 264 19392 270
rect 19340 206 19392 212
rect 24136 202 24164 750
rect 24504 678 24532 2382
rect 24688 882 24716 2790
rect 25056 2774 25084 6258
rect 25240 4078 25268 8230
rect 25332 8090 25360 8910
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25320 8084 25372 8090
rect 25320 8026 25372 8032
rect 25424 4622 25452 8570
rect 25608 7834 25636 11154
rect 25792 10130 25820 18686
rect 26068 18630 26096 19110
rect 25872 18624 25924 18630
rect 25872 18566 25924 18572
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 26056 18624 26108 18630
rect 26056 18566 26108 18572
rect 25884 16250 25912 18566
rect 25976 18290 26004 18566
rect 25964 18284 26016 18290
rect 25964 18226 26016 18232
rect 25964 16516 26016 16522
rect 25964 16458 26016 16464
rect 25872 16244 25924 16250
rect 25872 16186 25924 16192
rect 25870 16144 25926 16153
rect 25976 16114 26004 16458
rect 25870 16079 25872 16088
rect 25924 16079 25926 16088
rect 25964 16108 26016 16114
rect 25872 16050 25924 16056
rect 25964 16050 26016 16056
rect 25976 15978 26004 16050
rect 25964 15972 26016 15978
rect 25964 15914 26016 15920
rect 25976 15570 26004 15914
rect 25872 15564 25924 15570
rect 25872 15506 25924 15512
rect 25964 15564 26016 15570
rect 25964 15506 26016 15512
rect 25884 14074 25912 15506
rect 25976 15026 26004 15506
rect 26054 15464 26110 15473
rect 26054 15399 26110 15408
rect 26068 15094 26096 15399
rect 26056 15088 26108 15094
rect 26056 15030 26108 15036
rect 25964 15020 26016 15026
rect 25964 14962 26016 14968
rect 26056 14816 26108 14822
rect 26056 14758 26108 14764
rect 26068 14618 26096 14758
rect 26056 14612 26108 14618
rect 26056 14554 26108 14560
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 26160 12434 26188 20946
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 26252 19922 26280 20878
rect 26344 20262 26372 21422
rect 26700 20460 26752 20466
rect 26700 20402 26752 20408
rect 26332 20256 26384 20262
rect 26332 20198 26384 20204
rect 26240 19916 26292 19922
rect 26240 19858 26292 19864
rect 26252 18766 26280 19858
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 26252 18290 26280 18702
rect 26240 18284 26292 18290
rect 26240 18226 26292 18232
rect 26344 18034 26372 20198
rect 26424 19780 26476 19786
rect 26424 19722 26476 19728
rect 26252 18006 26372 18034
rect 26252 16538 26280 18006
rect 26436 17678 26464 19722
rect 26516 19508 26568 19514
rect 26516 19450 26568 19456
rect 26528 19242 26556 19450
rect 26712 19378 26740 20402
rect 26700 19372 26752 19378
rect 26700 19314 26752 19320
rect 26516 19236 26568 19242
rect 26516 19178 26568 19184
rect 26528 19009 26556 19178
rect 26608 19168 26660 19174
rect 26608 19110 26660 19116
rect 26514 19000 26570 19009
rect 26514 18935 26570 18944
rect 26516 18828 26568 18834
rect 26516 18770 26568 18776
rect 26528 18290 26556 18770
rect 26516 18284 26568 18290
rect 26516 18226 26568 18232
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 26424 17536 26476 17542
rect 26424 17478 26476 17484
rect 26436 17134 26464 17478
rect 26620 17377 26648 19110
rect 26712 18873 26740 19314
rect 26698 18864 26754 18873
rect 26698 18799 26754 18808
rect 26700 18080 26752 18086
rect 26700 18022 26752 18028
rect 26712 17649 26740 18022
rect 26698 17640 26754 17649
rect 26698 17575 26754 17584
rect 26606 17368 26662 17377
rect 26606 17303 26662 17312
rect 26424 17128 26476 17134
rect 26424 17070 26476 17076
rect 26252 16510 26556 16538
rect 26332 16040 26384 16046
rect 26238 16008 26294 16017
rect 26332 15982 26384 15988
rect 26238 15943 26294 15952
rect 26252 15638 26280 15943
rect 26240 15632 26292 15638
rect 26240 15574 26292 15580
rect 26252 15337 26280 15574
rect 26238 15328 26294 15337
rect 26238 15263 26294 15272
rect 26344 14074 26372 15982
rect 26528 15892 26556 16510
rect 26436 15864 26556 15892
rect 26436 14482 26464 15864
rect 26514 15192 26570 15201
rect 26514 15127 26570 15136
rect 26528 14498 26556 15127
rect 26620 15026 26648 17303
rect 26700 16448 26752 16454
rect 26700 16390 26752 16396
rect 26712 15910 26740 16390
rect 26700 15904 26752 15910
rect 26700 15846 26752 15852
rect 26712 15570 26740 15846
rect 26804 15586 26832 21490
rect 27632 21486 27660 22170
rect 28724 22092 28776 22098
rect 28724 22034 28776 22040
rect 27804 21888 27856 21894
rect 27804 21830 27856 21836
rect 27816 21690 27844 21830
rect 27804 21684 27856 21690
rect 27804 21626 27856 21632
rect 27344 21480 27396 21486
rect 27344 21422 27396 21428
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 28356 21480 28408 21486
rect 28356 21422 28408 21428
rect 26976 21004 27028 21010
rect 26976 20946 27028 20952
rect 26988 20890 27016 20946
rect 26896 20862 27016 20890
rect 26896 20466 26924 20862
rect 26963 20700 27271 20709
rect 26963 20698 26969 20700
rect 27025 20698 27049 20700
rect 27105 20698 27129 20700
rect 27185 20698 27209 20700
rect 27265 20698 27271 20700
rect 27025 20646 27027 20698
rect 27207 20646 27209 20698
rect 26963 20644 26969 20646
rect 27025 20644 27049 20646
rect 27105 20644 27129 20646
rect 27185 20644 27209 20646
rect 27265 20644 27271 20646
rect 26963 20635 27271 20644
rect 26884 20460 26936 20466
rect 26884 20402 26936 20408
rect 26896 19394 26924 20402
rect 27356 20058 27384 21422
rect 27436 20936 27488 20942
rect 27436 20878 27488 20884
rect 27528 20936 27580 20942
rect 27528 20878 27580 20884
rect 27344 20052 27396 20058
rect 27344 19994 27396 20000
rect 26963 19612 27271 19621
rect 26963 19610 26969 19612
rect 27025 19610 27049 19612
rect 27105 19610 27129 19612
rect 27185 19610 27209 19612
rect 27265 19610 27271 19612
rect 27025 19558 27027 19610
rect 27207 19558 27209 19610
rect 26963 19556 26969 19558
rect 27025 19556 27049 19558
rect 27105 19556 27129 19558
rect 27185 19556 27209 19558
rect 27265 19556 27271 19558
rect 26963 19547 27271 19556
rect 26896 19366 27108 19394
rect 27080 19334 27108 19366
rect 27344 19372 27396 19378
rect 27080 19310 27200 19334
rect 27344 19314 27396 19320
rect 27068 19306 27200 19310
rect 27068 19304 27120 19306
rect 27068 19246 27120 19252
rect 27172 18873 27200 19306
rect 27158 18864 27214 18873
rect 27158 18799 27214 18808
rect 26963 18524 27271 18533
rect 26963 18522 26969 18524
rect 27025 18522 27049 18524
rect 27105 18522 27129 18524
rect 27185 18522 27209 18524
rect 27265 18522 27271 18524
rect 27025 18470 27027 18522
rect 27207 18470 27209 18522
rect 26963 18468 26969 18470
rect 27025 18468 27049 18470
rect 27105 18468 27129 18470
rect 27185 18468 27209 18470
rect 27265 18468 27271 18470
rect 26963 18459 27271 18468
rect 26884 18420 26936 18426
rect 26884 18362 26936 18368
rect 26896 16674 26924 18362
rect 27068 18352 27120 18358
rect 27068 18294 27120 18300
rect 27080 18222 27108 18294
rect 27068 18216 27120 18222
rect 27068 18158 27120 18164
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 27172 17785 27200 18158
rect 27158 17776 27214 17785
rect 27356 17762 27384 19314
rect 27448 17882 27476 20878
rect 27540 20602 27568 20878
rect 28264 20800 28316 20806
rect 28264 20742 28316 20748
rect 27528 20596 27580 20602
rect 27528 20538 27580 20544
rect 28172 20596 28224 20602
rect 28172 20538 28224 20544
rect 27528 20256 27580 20262
rect 27528 20198 27580 20204
rect 27436 17876 27488 17882
rect 27436 17818 27488 17824
rect 27356 17734 27476 17762
rect 27158 17711 27214 17720
rect 27344 17672 27396 17678
rect 27344 17614 27396 17620
rect 26963 17436 27271 17445
rect 26963 17434 26969 17436
rect 27025 17434 27049 17436
rect 27105 17434 27129 17436
rect 27185 17434 27209 17436
rect 27265 17434 27271 17436
rect 27025 17382 27027 17434
rect 27207 17382 27209 17434
rect 26963 17380 26969 17382
rect 27025 17380 27049 17382
rect 27105 17380 27129 17382
rect 27185 17380 27209 17382
rect 27265 17380 27271 17382
rect 26963 17371 27271 17380
rect 26896 16646 27016 16674
rect 26988 16590 27016 16646
rect 26976 16584 27028 16590
rect 26976 16526 27028 16532
rect 26963 16348 27271 16357
rect 26963 16346 26969 16348
rect 27025 16346 27049 16348
rect 27105 16346 27129 16348
rect 27185 16346 27209 16348
rect 27265 16346 27271 16348
rect 27025 16294 27027 16346
rect 27207 16294 27209 16346
rect 26963 16292 26969 16294
rect 27025 16292 27049 16294
rect 27105 16292 27129 16294
rect 27185 16292 27209 16294
rect 27265 16292 27271 16294
rect 26963 16283 27271 16292
rect 26804 15570 27016 15586
rect 26700 15564 26752 15570
rect 26804 15564 27028 15570
rect 26804 15558 26976 15564
rect 26700 15506 26752 15512
rect 26976 15506 27028 15512
rect 26608 15020 26660 15026
rect 26608 14962 26660 14968
rect 26712 14822 26740 15506
rect 26884 15496 26936 15502
rect 26884 15438 26936 15444
rect 26700 14816 26752 14822
rect 26700 14758 26752 14764
rect 26792 14816 26844 14822
rect 26792 14758 26844 14764
rect 26804 14634 26832 14758
rect 26712 14606 26832 14634
rect 26424 14476 26476 14482
rect 26528 14470 26648 14498
rect 26424 14418 26476 14424
rect 26516 14272 26568 14278
rect 26516 14214 26568 14220
rect 26332 14068 26384 14074
rect 26332 14010 26384 14016
rect 26528 12782 26556 14214
rect 26620 13802 26648 14470
rect 26712 13938 26740 14606
rect 26792 14544 26844 14550
rect 26792 14486 26844 14492
rect 26700 13932 26752 13938
rect 26700 13874 26752 13880
rect 26608 13796 26660 13802
rect 26608 13738 26660 13744
rect 26620 13433 26648 13738
rect 26606 13424 26662 13433
rect 26606 13359 26662 13368
rect 26608 13320 26660 13326
rect 26712 13308 26740 13874
rect 26804 13870 26832 14486
rect 26792 13864 26844 13870
rect 26792 13806 26844 13812
rect 26804 13394 26832 13806
rect 26896 13530 26924 15438
rect 26963 15260 27271 15269
rect 26963 15258 26969 15260
rect 27025 15258 27049 15260
rect 27105 15258 27129 15260
rect 27185 15258 27209 15260
rect 27265 15258 27271 15260
rect 27025 15206 27027 15258
rect 27207 15206 27209 15258
rect 26963 15204 26969 15206
rect 27025 15204 27049 15206
rect 27105 15204 27129 15206
rect 27185 15204 27209 15206
rect 27265 15204 27271 15206
rect 26963 15195 27271 15204
rect 27066 14648 27122 14657
rect 27356 14618 27384 17614
rect 27066 14583 27122 14592
rect 27344 14612 27396 14618
rect 27080 14482 27108 14583
rect 27344 14554 27396 14560
rect 27068 14476 27120 14482
rect 27068 14418 27120 14424
rect 27344 14272 27396 14278
rect 27344 14214 27396 14220
rect 26963 14172 27271 14181
rect 26963 14170 26969 14172
rect 27025 14170 27049 14172
rect 27105 14170 27129 14172
rect 27185 14170 27209 14172
rect 27265 14170 27271 14172
rect 27025 14118 27027 14170
rect 27207 14118 27209 14170
rect 26963 14116 26969 14118
rect 27025 14116 27049 14118
rect 27105 14116 27129 14118
rect 27185 14116 27209 14118
rect 27265 14116 27271 14118
rect 26963 14107 27271 14116
rect 26884 13524 26936 13530
rect 26884 13466 26936 13472
rect 26792 13388 26844 13394
rect 26792 13330 26844 13336
rect 27356 13326 27384 14214
rect 27448 14074 27476 17734
rect 27540 16658 27568 20198
rect 27896 19984 27948 19990
rect 27896 19926 27948 19932
rect 27712 19168 27764 19174
rect 27712 19110 27764 19116
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27632 18222 27660 18702
rect 27620 18216 27672 18222
rect 27620 18158 27672 18164
rect 27528 16652 27580 16658
rect 27528 16594 27580 16600
rect 27724 16182 27752 19110
rect 27804 16652 27856 16658
rect 27804 16594 27856 16600
rect 27712 16176 27764 16182
rect 27712 16118 27764 16124
rect 27712 15972 27764 15978
rect 27712 15914 27764 15920
rect 27528 15904 27580 15910
rect 27528 15846 27580 15852
rect 27540 15162 27568 15846
rect 27528 15156 27580 15162
rect 27528 15098 27580 15104
rect 27618 14920 27674 14929
rect 27618 14855 27674 14864
rect 27528 14816 27580 14822
rect 27528 14758 27580 14764
rect 27540 14550 27568 14758
rect 27528 14544 27580 14550
rect 27528 14486 27580 14492
rect 27436 14068 27488 14074
rect 27436 14010 27488 14016
rect 27632 13530 27660 14855
rect 27724 14278 27752 15914
rect 27816 15162 27844 16594
rect 27908 15994 27936 19926
rect 28078 18864 28134 18873
rect 28078 18799 28134 18808
rect 27988 16992 28040 16998
rect 27988 16934 28040 16940
rect 28000 16794 28028 16934
rect 27988 16788 28040 16794
rect 27988 16730 28040 16736
rect 28092 16454 28120 18799
rect 28080 16448 28132 16454
rect 28080 16390 28132 16396
rect 27908 15966 28028 15994
rect 27896 15904 27948 15910
rect 27896 15846 27948 15852
rect 27908 15473 27936 15846
rect 27894 15464 27950 15473
rect 27894 15399 27950 15408
rect 28000 15314 28028 15966
rect 28078 15872 28134 15881
rect 28078 15807 28134 15816
rect 27908 15286 28028 15314
rect 27804 15156 27856 15162
rect 27804 15098 27856 15104
rect 27802 14648 27858 14657
rect 27802 14583 27858 14592
rect 27712 14272 27764 14278
rect 27712 14214 27764 14220
rect 27724 13734 27752 14214
rect 27712 13728 27764 13734
rect 27712 13670 27764 13676
rect 27620 13524 27672 13530
rect 27620 13466 27672 13472
rect 26660 13280 26740 13308
rect 26884 13320 26936 13326
rect 26608 13262 26660 13268
rect 26884 13262 26936 13268
rect 27344 13320 27396 13326
rect 27344 13262 27396 13268
rect 26608 12844 26660 12850
rect 26608 12786 26660 12792
rect 26516 12776 26568 12782
rect 26516 12718 26568 12724
rect 26068 12406 26188 12434
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 25872 11008 25924 11014
rect 25872 10950 25924 10956
rect 25780 10124 25832 10130
rect 25780 10066 25832 10072
rect 25688 9512 25740 9518
rect 25688 9454 25740 9460
rect 25700 9178 25728 9454
rect 25688 9172 25740 9178
rect 25688 9114 25740 9120
rect 25516 7806 25636 7834
rect 25412 4616 25464 4622
rect 25412 4558 25464 4564
rect 25228 4072 25280 4078
rect 25228 4014 25280 4020
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 25148 3641 25176 3878
rect 25134 3632 25190 3641
rect 25516 3602 25544 7806
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25700 6866 25728 7686
rect 25884 7342 25912 10950
rect 25976 10810 26004 11698
rect 25964 10804 26016 10810
rect 25964 10746 26016 10752
rect 26068 10062 26096 12406
rect 26424 12368 26476 12374
rect 26424 12310 26476 12316
rect 26436 11694 26464 12310
rect 26528 12306 26556 12718
rect 26516 12300 26568 12306
rect 26516 12242 26568 12248
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 26436 11354 26464 11630
rect 26424 11348 26476 11354
rect 26424 11290 26476 11296
rect 26148 11212 26200 11218
rect 26148 11154 26200 11160
rect 26332 11212 26384 11218
rect 26332 11154 26384 11160
rect 26160 10810 26188 11154
rect 26344 11082 26372 11154
rect 26436 11121 26464 11290
rect 26422 11112 26478 11121
rect 26332 11076 26384 11082
rect 26422 11047 26478 11056
rect 26332 11018 26384 11024
rect 26240 11008 26292 11014
rect 26240 10950 26292 10956
rect 26148 10804 26200 10810
rect 26148 10746 26200 10752
rect 26252 10606 26280 10950
rect 26240 10600 26292 10606
rect 26240 10542 26292 10548
rect 26148 10464 26200 10470
rect 26148 10406 26200 10412
rect 26160 10266 26188 10406
rect 26148 10260 26200 10266
rect 26148 10202 26200 10208
rect 26252 10062 26280 10542
rect 26332 10464 26384 10470
rect 26332 10406 26384 10412
rect 26344 10198 26372 10406
rect 26332 10192 26384 10198
rect 26332 10134 26384 10140
rect 26056 10056 26108 10062
rect 26056 9998 26108 10004
rect 26240 10056 26292 10062
rect 26240 9998 26292 10004
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 25976 8974 26004 9454
rect 26056 9036 26108 9042
rect 26056 8978 26108 8984
rect 25964 8968 26016 8974
rect 25964 8910 26016 8916
rect 25976 8430 26004 8910
rect 26068 8838 26096 8978
rect 26056 8832 26108 8838
rect 26056 8774 26108 8780
rect 26252 8498 26280 9998
rect 26332 9512 26384 9518
rect 26332 9454 26384 9460
rect 26240 8492 26292 8498
rect 26240 8434 26292 8440
rect 25964 8424 26016 8430
rect 25964 8366 26016 8372
rect 26344 7954 26372 9454
rect 26436 7954 26464 11047
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 26528 10266 26556 10610
rect 26516 10260 26568 10266
rect 26516 10202 26568 10208
rect 26528 8498 26556 10202
rect 26516 8492 26568 8498
rect 26516 8434 26568 8440
rect 26514 8392 26570 8401
rect 26514 8327 26570 8336
rect 26528 8106 26556 8327
rect 26620 8294 26648 12786
rect 26792 12640 26844 12646
rect 26792 12582 26844 12588
rect 26804 12442 26832 12582
rect 26792 12436 26844 12442
rect 26792 12378 26844 12384
rect 26896 12322 26924 13262
rect 26963 13084 27271 13093
rect 26963 13082 26969 13084
rect 27025 13082 27049 13084
rect 27105 13082 27129 13084
rect 27185 13082 27209 13084
rect 27265 13082 27271 13084
rect 27025 13030 27027 13082
rect 27207 13030 27209 13082
rect 26963 13028 26969 13030
rect 27025 13028 27049 13030
rect 27105 13028 27129 13030
rect 27185 13028 27209 13030
rect 27265 13028 27271 13030
rect 26963 13019 27271 13028
rect 27816 12646 27844 14583
rect 27804 12640 27856 12646
rect 26804 12294 26924 12322
rect 27724 12600 27804 12628
rect 26804 11898 26832 12294
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 26896 11898 26924 12174
rect 26963 11996 27271 12005
rect 26963 11994 26969 11996
rect 27025 11994 27049 11996
rect 27105 11994 27129 11996
rect 27185 11994 27209 11996
rect 27265 11994 27271 11996
rect 27025 11942 27027 11994
rect 27207 11942 27209 11994
rect 26963 11940 26969 11942
rect 27025 11940 27049 11942
rect 27105 11940 27129 11942
rect 27185 11940 27209 11942
rect 27265 11940 27271 11942
rect 26963 11931 27271 11940
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26884 11892 26936 11898
rect 26884 11834 26936 11840
rect 27160 11688 27212 11694
rect 27160 11630 27212 11636
rect 26700 11552 26752 11558
rect 26700 11494 26752 11500
rect 26712 11286 26740 11494
rect 27172 11354 27200 11630
rect 27724 11354 27752 12600
rect 27804 12582 27856 12588
rect 27804 12232 27856 12238
rect 27804 12174 27856 12180
rect 27816 11354 27844 12174
rect 27908 11354 27936 15286
rect 27988 14884 28040 14890
rect 27988 14826 28040 14832
rect 28000 13297 28028 14826
rect 28092 13852 28120 15807
rect 28184 15144 28212 20538
rect 28276 16658 28304 20742
rect 28368 20602 28396 21422
rect 28736 21350 28764 22034
rect 30288 22024 30340 22030
rect 30288 21966 30340 21972
rect 29092 21480 29144 21486
rect 29092 21422 29144 21428
rect 29276 21480 29328 21486
rect 29328 21440 29500 21468
rect 29276 21422 29328 21428
rect 28724 21344 28776 21350
rect 28724 21286 28776 21292
rect 28540 20800 28592 20806
rect 28540 20742 28592 20748
rect 28356 20596 28408 20602
rect 28356 20538 28408 20544
rect 28552 20097 28580 20742
rect 28538 20088 28594 20097
rect 28538 20023 28594 20032
rect 28354 19952 28410 19961
rect 28354 19887 28356 19896
rect 28408 19887 28410 19896
rect 28356 19858 28408 19864
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28460 18834 28488 19790
rect 28540 19168 28592 19174
rect 28540 19110 28592 19116
rect 28552 18970 28580 19110
rect 28540 18964 28592 18970
rect 28540 18906 28592 18912
rect 28448 18828 28500 18834
rect 28500 18788 28580 18816
rect 28448 18770 28500 18776
rect 28356 18624 28408 18630
rect 28356 18566 28408 18572
rect 28368 17270 28396 18566
rect 28448 18080 28500 18086
rect 28448 18022 28500 18028
rect 28356 17264 28408 17270
rect 28354 17232 28356 17241
rect 28408 17232 28410 17241
rect 28460 17202 28488 18022
rect 28552 17678 28580 18788
rect 28736 17762 28764 21286
rect 29000 20936 29052 20942
rect 29000 20878 29052 20884
rect 28908 20528 28960 20534
rect 28908 20470 28960 20476
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28828 18970 28856 19790
rect 28920 19378 28948 20470
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 28816 18964 28868 18970
rect 28816 18906 28868 18912
rect 28828 17882 28856 18906
rect 28908 18760 28960 18766
rect 28908 18702 28960 18708
rect 28816 17876 28868 17882
rect 28816 17818 28868 17824
rect 28736 17734 28856 17762
rect 28540 17672 28592 17678
rect 28540 17614 28592 17620
rect 28354 17167 28410 17176
rect 28448 17196 28500 17202
rect 28448 17138 28500 17144
rect 28264 16652 28316 16658
rect 28264 16594 28316 16600
rect 28448 16176 28500 16182
rect 28448 16118 28500 16124
rect 28184 15116 28396 15144
rect 28172 15020 28224 15026
rect 28172 14962 28224 14968
rect 28184 14006 28212 14962
rect 28172 14000 28224 14006
rect 28172 13942 28224 13948
rect 28092 13824 28212 13852
rect 27986 13288 28042 13297
rect 27986 13223 28042 13232
rect 28080 12300 28132 12306
rect 28080 12242 28132 12248
rect 27160 11348 27212 11354
rect 27160 11290 27212 11296
rect 27712 11348 27764 11354
rect 27712 11290 27764 11296
rect 27804 11348 27856 11354
rect 27804 11290 27856 11296
rect 27896 11348 27948 11354
rect 27896 11290 27948 11296
rect 26700 11280 26752 11286
rect 26700 11222 26752 11228
rect 26608 8288 26660 8294
rect 26608 8230 26660 8236
rect 26528 8078 26648 8106
rect 26712 8090 26740 11222
rect 28092 11150 28120 12242
rect 28080 11144 28132 11150
rect 28080 11086 28132 11092
rect 26963 10908 27271 10917
rect 26963 10906 26969 10908
rect 27025 10906 27049 10908
rect 27105 10906 27129 10908
rect 27185 10906 27209 10908
rect 27265 10906 27271 10908
rect 27025 10854 27027 10906
rect 27207 10854 27209 10906
rect 26963 10852 26969 10854
rect 27025 10852 27049 10854
rect 27105 10852 27129 10854
rect 27185 10852 27209 10854
rect 27265 10852 27271 10854
rect 26963 10843 27271 10852
rect 28184 10810 28212 13824
rect 28264 13728 28316 13734
rect 28264 13670 28316 13676
rect 28276 12442 28304 13670
rect 28368 13394 28396 15116
rect 28460 13682 28488 16118
rect 28552 15026 28580 17614
rect 28724 17060 28776 17066
rect 28724 17002 28776 17008
rect 28632 16992 28684 16998
rect 28632 16934 28684 16940
rect 28644 16590 28672 16934
rect 28632 16584 28684 16590
rect 28632 16526 28684 16532
rect 28630 16144 28686 16153
rect 28630 16079 28686 16088
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28538 13832 28594 13841
rect 28538 13767 28540 13776
rect 28592 13767 28594 13776
rect 28540 13738 28592 13744
rect 28644 13734 28672 16079
rect 28736 15570 28764 17002
rect 28724 15564 28776 15570
rect 28724 15506 28776 15512
rect 28828 15502 28856 17734
rect 28816 15496 28868 15502
rect 28816 15438 28868 15444
rect 28816 15360 28868 15366
rect 28816 15302 28868 15308
rect 28724 14952 28776 14958
rect 28724 14894 28776 14900
rect 28736 14793 28764 14894
rect 28828 14890 28856 15302
rect 28816 14884 28868 14890
rect 28816 14826 28868 14832
rect 28722 14784 28778 14793
rect 28722 14719 28778 14728
rect 28722 14648 28778 14657
rect 28722 14583 28724 14592
rect 28776 14583 28778 14592
rect 28724 14554 28776 14560
rect 28724 14408 28776 14414
rect 28724 14350 28776 14356
rect 28816 14408 28868 14414
rect 28816 14350 28868 14356
rect 28632 13728 28684 13734
rect 28460 13654 28580 13682
rect 28632 13670 28684 13676
rect 28356 13388 28408 13394
rect 28356 13330 28408 13336
rect 28448 12776 28500 12782
rect 28448 12718 28500 12724
rect 28264 12436 28316 12442
rect 28264 12378 28316 12384
rect 28460 11898 28488 12718
rect 28552 12220 28580 13654
rect 28632 12232 28684 12238
rect 28552 12192 28632 12220
rect 28632 12174 28684 12180
rect 28448 11892 28500 11898
rect 28448 11834 28500 11840
rect 28172 10804 28224 10810
rect 28172 10746 28224 10752
rect 28448 10736 28500 10742
rect 28448 10678 28500 10684
rect 27988 10600 28040 10606
rect 27988 10542 28040 10548
rect 27804 10532 27856 10538
rect 27804 10474 27856 10480
rect 26884 10056 26936 10062
rect 26884 9998 26936 10004
rect 27620 10056 27672 10062
rect 27620 9998 27672 10004
rect 26896 9722 26924 9998
rect 26963 9820 27271 9829
rect 26963 9818 26969 9820
rect 27025 9818 27049 9820
rect 27105 9818 27129 9820
rect 27185 9818 27209 9820
rect 27265 9818 27271 9820
rect 27025 9766 27027 9818
rect 27207 9766 27209 9818
rect 26963 9764 26969 9766
rect 27025 9764 27049 9766
rect 27105 9764 27129 9766
rect 27185 9764 27209 9766
rect 27265 9764 27271 9766
rect 26963 9755 27271 9764
rect 27632 9722 27660 9998
rect 26884 9716 26936 9722
rect 26884 9658 26936 9664
rect 27620 9716 27672 9722
rect 27620 9658 27672 9664
rect 27252 9580 27304 9586
rect 27252 9522 27304 9528
rect 26792 9444 26844 9450
rect 26792 9386 26844 9392
rect 26804 8945 26832 9386
rect 27264 9382 27292 9522
rect 27816 9450 27844 10474
rect 28000 9722 28028 10542
rect 28356 10532 28408 10538
rect 28356 10474 28408 10480
rect 28172 9920 28224 9926
rect 28172 9862 28224 9868
rect 27988 9716 28040 9722
rect 27988 9658 28040 9664
rect 27804 9444 27856 9450
rect 27804 9386 27856 9392
rect 27252 9376 27304 9382
rect 27252 9318 27304 9324
rect 27988 9376 28040 9382
rect 27988 9318 28040 9324
rect 28080 9376 28132 9382
rect 28080 9318 28132 9324
rect 26884 8968 26936 8974
rect 26790 8936 26846 8945
rect 26884 8910 26936 8916
rect 26790 8871 26846 8880
rect 26792 8832 26844 8838
rect 26792 8774 26844 8780
rect 26332 7948 26384 7954
rect 26252 7908 26332 7936
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 25964 7744 26016 7750
rect 25964 7686 26016 7692
rect 25872 7336 25924 7342
rect 25778 7304 25834 7313
rect 25872 7278 25924 7284
rect 25778 7239 25834 7248
rect 25688 6860 25740 6866
rect 25688 6802 25740 6808
rect 25596 6248 25648 6254
rect 25596 6190 25648 6196
rect 25608 5846 25636 6190
rect 25596 5840 25648 5846
rect 25596 5782 25648 5788
rect 25134 3567 25190 3576
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 25320 3392 25372 3398
rect 25320 3334 25372 3340
rect 25056 2746 25176 2774
rect 24860 1760 24912 1766
rect 24860 1702 24912 1708
rect 24676 876 24728 882
rect 24676 818 24728 824
rect 24492 672 24544 678
rect 24492 614 24544 620
rect 24872 406 24900 1702
rect 25148 1358 25176 2746
rect 25332 2514 25360 3334
rect 25516 3126 25544 3538
rect 25792 3466 25820 7239
rect 25872 6724 25924 6730
rect 25872 6666 25924 6672
rect 25884 5710 25912 6666
rect 25976 6322 26004 7686
rect 26068 6390 26096 7822
rect 26252 6798 26280 7908
rect 26332 7890 26384 7896
rect 26424 7948 26476 7954
rect 26424 7890 26476 7896
rect 26436 7410 26464 7890
rect 26424 7404 26476 7410
rect 26424 7346 26476 7352
rect 26332 7268 26384 7274
rect 26332 7210 26384 7216
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26056 6384 26108 6390
rect 26056 6326 26108 6332
rect 26238 6352 26294 6361
rect 25964 6316 26016 6322
rect 26238 6287 26240 6296
rect 25964 6258 26016 6264
rect 26292 6287 26294 6296
rect 26240 6258 26292 6264
rect 26344 6118 26372 7210
rect 26424 6860 26476 6866
rect 26424 6802 26476 6808
rect 26436 6662 26464 6802
rect 26424 6656 26476 6662
rect 26424 6598 26476 6604
rect 26516 6656 26568 6662
rect 26516 6598 26568 6604
rect 26436 6254 26464 6598
rect 26424 6248 26476 6254
rect 26424 6190 26476 6196
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 26436 5778 26464 6190
rect 26424 5772 26476 5778
rect 26424 5714 26476 5720
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 26240 5636 26292 5642
rect 26240 5578 26292 5584
rect 26148 5568 26200 5574
rect 25870 5536 25926 5545
rect 26148 5510 26200 5516
rect 25870 5471 25926 5480
rect 25780 3460 25832 3466
rect 25780 3402 25832 3408
rect 25884 3126 25912 5471
rect 26056 4480 26108 4486
rect 26056 4422 26108 4428
rect 26068 4146 26096 4422
rect 26056 4140 26108 4146
rect 26056 4082 26108 4088
rect 26056 3936 26108 3942
rect 26056 3878 26108 3884
rect 25964 3188 26016 3194
rect 25964 3130 26016 3136
rect 25504 3120 25556 3126
rect 25504 3062 25556 3068
rect 25872 3120 25924 3126
rect 25872 3062 25924 3068
rect 25976 2650 26004 3130
rect 25964 2644 26016 2650
rect 25964 2586 26016 2592
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 26068 2038 26096 3878
rect 26160 3058 26188 5510
rect 26252 5166 26280 5578
rect 26330 5536 26386 5545
rect 26330 5471 26386 5480
rect 26344 5234 26372 5471
rect 26332 5228 26384 5234
rect 26332 5170 26384 5176
rect 26436 5166 26464 5714
rect 26240 5160 26292 5166
rect 26240 5102 26292 5108
rect 26424 5160 26476 5166
rect 26424 5102 26476 5108
rect 26528 5098 26556 6598
rect 26620 5658 26648 8078
rect 26700 8084 26752 8090
rect 26700 8026 26752 8032
rect 26712 7546 26740 8026
rect 26804 7954 26832 8774
rect 26896 8634 26924 8910
rect 28000 8838 28028 9318
rect 27988 8832 28040 8838
rect 27988 8774 28040 8780
rect 26963 8732 27271 8741
rect 26963 8730 26969 8732
rect 27025 8730 27049 8732
rect 27105 8730 27129 8732
rect 27185 8730 27209 8732
rect 27265 8730 27271 8732
rect 27025 8678 27027 8730
rect 27207 8678 27209 8730
rect 26963 8676 26969 8678
rect 27025 8676 27049 8678
rect 27105 8676 27129 8678
rect 27185 8676 27209 8678
rect 27265 8676 27271 8678
rect 26963 8667 27271 8676
rect 26884 8628 26936 8634
rect 26884 8570 26936 8576
rect 28092 8430 28120 9318
rect 26976 8424 27028 8430
rect 26976 8366 27028 8372
rect 28080 8424 28132 8430
rect 28080 8366 28132 8372
rect 26792 7948 26844 7954
rect 26792 7890 26844 7896
rect 26884 7948 26936 7954
rect 26988 7936 27016 8366
rect 27988 8356 28040 8362
rect 27988 8298 28040 8304
rect 27068 8288 27120 8294
rect 27068 8230 27120 8236
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 27080 7954 27108 8230
rect 26936 7908 27016 7936
rect 27068 7948 27120 7954
rect 26884 7890 26936 7896
rect 27068 7890 27120 7896
rect 27528 7948 27580 7954
rect 27528 7890 27580 7896
rect 26792 7744 26844 7750
rect 26792 7686 26844 7692
rect 26700 7540 26752 7546
rect 26700 7482 26752 7488
rect 26700 6792 26752 6798
rect 26700 6734 26752 6740
rect 26712 5760 26740 6734
rect 26804 6254 26832 7686
rect 26896 6662 26924 7890
rect 26963 7644 27271 7653
rect 26963 7642 26969 7644
rect 27025 7642 27049 7644
rect 27105 7642 27129 7644
rect 27185 7642 27209 7644
rect 27265 7642 27271 7644
rect 27025 7590 27027 7642
rect 27207 7590 27209 7642
rect 26963 7588 26969 7590
rect 27025 7588 27049 7590
rect 27105 7588 27129 7590
rect 27185 7588 27209 7590
rect 27265 7588 27271 7590
rect 26963 7579 27271 7588
rect 26884 6656 26936 6662
rect 26884 6598 26936 6604
rect 27344 6656 27396 6662
rect 27344 6598 27396 6604
rect 26963 6556 27271 6565
rect 26963 6554 26969 6556
rect 27025 6554 27049 6556
rect 27105 6554 27129 6556
rect 27185 6554 27209 6556
rect 27265 6554 27271 6556
rect 27025 6502 27027 6554
rect 27207 6502 27209 6554
rect 26963 6500 26969 6502
rect 27025 6500 27049 6502
rect 27105 6500 27129 6502
rect 27185 6500 27209 6502
rect 27265 6500 27271 6502
rect 26963 6491 27271 6500
rect 27252 6316 27304 6322
rect 27252 6258 27304 6264
rect 26792 6248 26844 6254
rect 26792 6190 26844 6196
rect 27264 5778 27292 6258
rect 26792 5772 26844 5778
rect 26712 5732 26792 5760
rect 26792 5714 26844 5720
rect 27252 5772 27304 5778
rect 27252 5714 27304 5720
rect 26620 5630 26740 5658
rect 26608 5568 26660 5574
rect 26608 5510 26660 5516
rect 26516 5092 26568 5098
rect 26516 5034 26568 5040
rect 26240 4072 26292 4078
rect 26240 4014 26292 4020
rect 26148 3052 26200 3058
rect 26148 2994 26200 3000
rect 26252 2990 26280 4014
rect 26528 3738 26556 5034
rect 26516 3732 26568 3738
rect 26516 3674 26568 3680
rect 26424 3392 26476 3398
rect 26424 3334 26476 3340
rect 26240 2984 26292 2990
rect 26240 2926 26292 2932
rect 26252 2582 26280 2926
rect 26240 2576 26292 2582
rect 26240 2518 26292 2524
rect 26056 2032 26108 2038
rect 26056 1974 26108 1980
rect 26252 1970 26280 2518
rect 26436 2446 26464 3334
rect 26620 2990 26648 5510
rect 26712 4758 26740 5630
rect 26792 5636 26844 5642
rect 26792 5578 26844 5584
rect 26700 4752 26752 4758
rect 26700 4694 26752 4700
rect 26804 4146 26832 5578
rect 26884 5568 26936 5574
rect 26884 5510 26936 5516
rect 26792 4140 26844 4146
rect 26792 4082 26844 4088
rect 26700 3936 26752 3942
rect 26700 3878 26752 3884
rect 26712 3738 26740 3878
rect 26700 3732 26752 3738
rect 26700 3674 26752 3680
rect 26608 2984 26660 2990
rect 26608 2926 26660 2932
rect 26712 2854 26740 3674
rect 26700 2848 26752 2854
rect 26620 2796 26700 2802
rect 26620 2790 26752 2796
rect 26620 2774 26740 2790
rect 26424 2440 26476 2446
rect 26424 2382 26476 2388
rect 26422 2272 26478 2281
rect 26478 2230 26556 2258
rect 26422 2207 26478 2216
rect 26240 1964 26292 1970
rect 26240 1906 26292 1912
rect 26056 1896 26108 1902
rect 26056 1838 26108 1844
rect 26424 1896 26476 1902
rect 26528 1884 26556 2230
rect 26476 1856 26556 1884
rect 26424 1838 26476 1844
rect 25962 1456 26018 1465
rect 25962 1391 25964 1400
rect 26016 1391 26018 1400
rect 25964 1362 26016 1368
rect 25136 1352 25188 1358
rect 25136 1294 25188 1300
rect 25320 1216 25372 1222
rect 25320 1158 25372 1164
rect 25688 1216 25740 1222
rect 25688 1158 25740 1164
rect 24860 400 24912 406
rect 25332 377 25360 1158
rect 25700 474 25728 1158
rect 25778 776 25834 785
rect 25976 762 26004 1362
rect 26068 1018 26096 1838
rect 26332 1760 26384 1766
rect 26332 1702 26384 1708
rect 26240 1488 26292 1494
rect 26240 1430 26292 1436
rect 26056 1012 26108 1018
rect 26056 954 26108 960
rect 26252 921 26280 1430
rect 26344 1193 26372 1702
rect 26528 1426 26556 1856
rect 26620 1766 26648 2774
rect 26896 1986 26924 5510
rect 26963 5468 27271 5477
rect 26963 5466 26969 5468
rect 27025 5466 27049 5468
rect 27105 5466 27129 5468
rect 27185 5466 27209 5468
rect 27265 5466 27271 5468
rect 27025 5414 27027 5466
rect 27207 5414 27209 5466
rect 26963 5412 26969 5414
rect 27025 5412 27049 5414
rect 27105 5412 27129 5414
rect 27185 5412 27209 5414
rect 27265 5412 27271 5414
rect 26963 5403 27271 5412
rect 27356 5273 27384 6598
rect 27540 6322 27568 7890
rect 27712 7880 27764 7886
rect 27712 7822 27764 7828
rect 27724 6866 27752 7822
rect 27816 7410 27844 8230
rect 28000 7954 28028 8298
rect 28080 8084 28132 8090
rect 28080 8026 28132 8032
rect 27988 7948 28040 7954
rect 27988 7890 28040 7896
rect 27804 7404 27856 7410
rect 27804 7346 27856 7352
rect 27712 6860 27764 6866
rect 27712 6802 27764 6808
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 28000 6202 28028 7890
rect 28092 7002 28120 8026
rect 28184 7886 28212 9862
rect 28264 8832 28316 8838
rect 28264 8774 28316 8780
rect 28276 8634 28304 8774
rect 28264 8628 28316 8634
rect 28264 8570 28316 8576
rect 28172 7880 28224 7886
rect 28172 7822 28224 7828
rect 28264 7744 28316 7750
rect 28264 7686 28316 7692
rect 28080 6996 28132 7002
rect 28080 6938 28132 6944
rect 27816 6174 28028 6202
rect 27620 5908 27672 5914
rect 27620 5850 27672 5856
rect 27632 5817 27660 5850
rect 27618 5808 27674 5817
rect 27618 5743 27674 5752
rect 27528 5704 27580 5710
rect 27528 5646 27580 5652
rect 27342 5264 27398 5273
rect 27342 5199 27398 5208
rect 26963 4380 27271 4389
rect 26963 4378 26969 4380
rect 27025 4378 27049 4380
rect 27105 4378 27129 4380
rect 27185 4378 27209 4380
rect 27265 4378 27271 4380
rect 27025 4326 27027 4378
rect 27207 4326 27209 4378
rect 26963 4324 26969 4326
rect 27025 4324 27049 4326
rect 27105 4324 27129 4326
rect 27185 4324 27209 4326
rect 27265 4324 27271 4326
rect 26963 4315 27271 4324
rect 26963 3292 27271 3301
rect 26963 3290 26969 3292
rect 27025 3290 27049 3292
rect 27105 3290 27129 3292
rect 27185 3290 27209 3292
rect 27265 3290 27271 3292
rect 27025 3238 27027 3290
rect 27207 3238 27209 3290
rect 26963 3236 26969 3238
rect 27025 3236 27049 3238
rect 27105 3236 27129 3238
rect 27185 3236 27209 3238
rect 27265 3236 27271 3238
rect 26963 3227 27271 3236
rect 27068 3052 27120 3058
rect 27068 2994 27120 3000
rect 27080 2961 27108 2994
rect 27066 2952 27122 2961
rect 27066 2887 27122 2896
rect 27356 2514 27384 5199
rect 27540 4690 27568 5646
rect 27528 4684 27580 4690
rect 27528 4626 27580 4632
rect 27816 4622 27844 6174
rect 27896 6112 27948 6118
rect 27896 6054 27948 6060
rect 27908 5710 27936 6054
rect 27896 5704 27948 5710
rect 27896 5646 27948 5652
rect 27908 5030 27936 5646
rect 28172 5568 28224 5574
rect 28172 5510 28224 5516
rect 27896 5024 27948 5030
rect 27896 4966 27948 4972
rect 27908 4826 27936 4966
rect 27896 4820 27948 4826
rect 27896 4762 27948 4768
rect 27896 4684 27948 4690
rect 27896 4626 27948 4632
rect 27436 4616 27488 4622
rect 27804 4616 27856 4622
rect 27436 4558 27488 4564
rect 27618 4584 27674 4593
rect 27448 2990 27476 4558
rect 27804 4558 27856 4564
rect 27618 4519 27674 4528
rect 27632 3670 27660 4519
rect 27710 4176 27766 4185
rect 27710 4111 27766 4120
rect 27620 3664 27672 3670
rect 27620 3606 27672 3612
rect 27436 2984 27488 2990
rect 27436 2926 27488 2932
rect 27620 2848 27672 2854
rect 27620 2790 27672 2796
rect 27344 2508 27396 2514
rect 27344 2450 27396 2456
rect 27528 2508 27580 2514
rect 27528 2450 27580 2456
rect 26963 2204 27271 2213
rect 26963 2202 26969 2204
rect 27025 2202 27049 2204
rect 27105 2202 27129 2204
rect 27185 2202 27209 2204
rect 27265 2202 27271 2204
rect 27025 2150 27027 2202
rect 27207 2150 27209 2202
rect 26963 2148 26969 2150
rect 27025 2148 27049 2150
rect 27105 2148 27129 2150
rect 27185 2148 27209 2150
rect 27265 2148 27271 2150
rect 26963 2139 27271 2148
rect 26896 1970 27016 1986
rect 26896 1964 27028 1970
rect 26896 1958 26976 1964
rect 26976 1906 27028 1912
rect 26608 1760 26660 1766
rect 26608 1702 26660 1708
rect 26976 1760 27028 1766
rect 26976 1702 27028 1708
rect 26884 1556 26936 1562
rect 26884 1498 26936 1504
rect 26516 1420 26568 1426
rect 26516 1362 26568 1368
rect 26896 1329 26924 1498
rect 26988 1465 27016 1702
rect 26974 1456 27030 1465
rect 27356 1426 27384 2450
rect 27434 2000 27490 2009
rect 27434 1935 27490 1944
rect 27448 1562 27476 1935
rect 27540 1766 27568 2450
rect 27528 1760 27580 1766
rect 27528 1702 27580 1708
rect 27436 1556 27488 1562
rect 27436 1498 27488 1504
rect 26974 1391 26976 1400
rect 27028 1391 27030 1400
rect 27344 1420 27396 1426
rect 26976 1362 27028 1368
rect 27344 1362 27396 1368
rect 26882 1320 26938 1329
rect 26882 1255 26938 1264
rect 26330 1184 26386 1193
rect 26330 1119 26386 1128
rect 26963 1116 27271 1125
rect 26963 1114 26969 1116
rect 27025 1114 27049 1116
rect 27105 1114 27129 1116
rect 27185 1114 27209 1116
rect 27265 1114 27271 1116
rect 27025 1062 27027 1114
rect 27207 1062 27209 1114
rect 26963 1060 26969 1062
rect 27025 1060 27049 1062
rect 27105 1060 27129 1062
rect 27185 1060 27209 1062
rect 27265 1060 27271 1062
rect 26963 1051 27271 1060
rect 26238 912 26294 921
rect 26238 847 26294 856
rect 27356 814 27384 1362
rect 27632 882 27660 2790
rect 27724 2650 27752 4111
rect 27804 3664 27856 3670
rect 27804 3606 27856 3612
rect 27712 2644 27764 2650
rect 27712 2586 27764 2592
rect 27712 1760 27764 1766
rect 27712 1702 27764 1708
rect 27724 1358 27752 1702
rect 27816 1562 27844 3606
rect 27908 3602 27936 4626
rect 28080 3936 28132 3942
rect 28080 3878 28132 3884
rect 27896 3596 27948 3602
rect 27948 3556 28028 3584
rect 27896 3538 27948 3544
rect 27894 3496 27950 3505
rect 27894 3431 27950 3440
rect 27908 2378 27936 3431
rect 28000 2514 28028 3556
rect 27988 2508 28040 2514
rect 27988 2450 28040 2456
rect 27896 2372 27948 2378
rect 27896 2314 27948 2320
rect 27804 1556 27856 1562
rect 27804 1498 27856 1504
rect 27712 1352 27764 1358
rect 27712 1294 27764 1300
rect 27620 876 27672 882
rect 27620 818 27672 824
rect 25834 734 26004 762
rect 27344 808 27396 814
rect 27344 750 27396 756
rect 25778 711 25834 720
rect 27816 678 27844 1498
rect 28092 1358 28120 3878
rect 28184 1358 28212 5510
rect 28276 4622 28304 7686
rect 28368 6866 28396 10474
rect 28460 7954 28488 10678
rect 28540 10464 28592 10470
rect 28540 10406 28592 10412
rect 28552 9518 28580 10406
rect 28644 10130 28672 12174
rect 28632 10124 28684 10130
rect 28632 10066 28684 10072
rect 28540 9512 28592 9518
rect 28540 9454 28592 9460
rect 28540 8288 28592 8294
rect 28540 8230 28592 8236
rect 28448 7948 28500 7954
rect 28448 7890 28500 7896
rect 28448 7200 28500 7206
rect 28448 7142 28500 7148
rect 28356 6860 28408 6866
rect 28356 6802 28408 6808
rect 28460 5302 28488 7142
rect 28552 5778 28580 8230
rect 28736 7546 28764 14350
rect 28828 11898 28856 14350
rect 28920 12986 28948 18702
rect 29012 17882 29040 20878
rect 29104 20330 29132 21422
rect 29472 20534 29500 21440
rect 29828 21412 29880 21418
rect 29828 21354 29880 21360
rect 29920 21412 29972 21418
rect 29920 21354 29972 21360
rect 29736 21344 29788 21350
rect 29736 21286 29788 21292
rect 29460 20528 29512 20534
rect 29460 20470 29512 20476
rect 29472 20398 29500 20470
rect 29276 20392 29328 20398
rect 29276 20334 29328 20340
rect 29460 20392 29512 20398
rect 29460 20334 29512 20340
rect 29092 20324 29144 20330
rect 29092 20266 29144 20272
rect 29104 19394 29132 20266
rect 29104 19366 29224 19394
rect 29092 19236 29144 19242
rect 29092 19178 29144 19184
rect 29000 17876 29052 17882
rect 29000 17818 29052 17824
rect 29104 16425 29132 19178
rect 29196 18850 29224 19366
rect 29288 18970 29316 20334
rect 29460 20256 29512 20262
rect 29460 20198 29512 20204
rect 29552 20256 29604 20262
rect 29552 20198 29604 20204
rect 29276 18964 29328 18970
rect 29276 18906 29328 18912
rect 29196 18834 29316 18850
rect 29196 18828 29328 18834
rect 29196 18822 29276 18828
rect 29276 18770 29328 18776
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29196 16561 29224 18702
rect 29368 18148 29420 18154
rect 29368 18090 29420 18096
rect 29276 17536 29328 17542
rect 29276 17478 29328 17484
rect 29288 16998 29316 17478
rect 29276 16992 29328 16998
rect 29276 16934 29328 16940
rect 29288 16833 29316 16934
rect 29274 16824 29330 16833
rect 29380 16794 29408 18090
rect 29274 16759 29330 16768
rect 29368 16788 29420 16794
rect 29368 16730 29420 16736
rect 29182 16552 29238 16561
rect 29182 16487 29238 16496
rect 29090 16416 29146 16425
rect 29090 16351 29146 16360
rect 28998 16280 29054 16289
rect 28998 16215 29000 16224
rect 29052 16215 29054 16224
rect 29000 16186 29052 16192
rect 29366 16144 29422 16153
rect 29362 16088 29366 16130
rect 29362 16079 29422 16088
rect 29092 16040 29144 16046
rect 29092 15982 29144 15988
rect 29184 16040 29236 16046
rect 29362 15994 29390 16079
rect 29236 15988 29390 15994
rect 29184 15982 29390 15988
rect 29000 15972 29052 15978
rect 29000 15914 29052 15920
rect 29012 15570 29040 15914
rect 29104 15745 29132 15982
rect 29196 15966 29390 15982
rect 29368 15904 29420 15910
rect 29368 15846 29420 15852
rect 29090 15736 29146 15745
rect 29090 15671 29146 15680
rect 29000 15564 29052 15570
rect 29000 15506 29052 15512
rect 29104 14113 29132 15671
rect 29380 15586 29408 15846
rect 29196 15558 29408 15586
rect 29090 14104 29146 14113
rect 29090 14039 29146 14048
rect 29000 14000 29052 14006
rect 28998 13968 29000 13977
rect 29052 13968 29054 13977
rect 28998 13903 29054 13912
rect 29196 13870 29224 15558
rect 29368 15496 29420 15502
rect 29368 15438 29420 15444
rect 29276 14816 29328 14822
rect 29276 14758 29328 14764
rect 29288 14006 29316 14758
rect 29276 14000 29328 14006
rect 29276 13942 29328 13948
rect 29380 13870 29408 15438
rect 29000 13864 29052 13870
rect 29000 13806 29052 13812
rect 29184 13864 29236 13870
rect 29276 13864 29328 13870
rect 29184 13806 29236 13812
rect 29274 13832 29276 13841
rect 29368 13864 29420 13870
rect 29328 13832 29330 13841
rect 28908 12980 28960 12986
rect 28908 12922 28960 12928
rect 29012 12889 29040 13806
rect 29368 13806 29420 13812
rect 29274 13767 29330 13776
rect 29366 13696 29422 13705
rect 29366 13631 29422 13640
rect 29274 13560 29330 13569
rect 29274 13495 29276 13504
rect 29328 13495 29330 13504
rect 29276 13466 29328 13472
rect 29274 13424 29330 13433
rect 29274 13359 29330 13368
rect 29090 13016 29146 13025
rect 29090 12951 29092 12960
rect 29144 12951 29146 12960
rect 29092 12922 29144 12928
rect 28998 12880 29054 12889
rect 29288 12866 29316 13359
rect 28998 12815 29054 12824
rect 29104 12838 29316 12866
rect 29000 12640 29052 12646
rect 29000 12582 29052 12588
rect 28906 12336 28962 12345
rect 28906 12271 28908 12280
rect 28960 12271 28962 12280
rect 28908 12242 28960 12248
rect 29012 12186 29040 12582
rect 28920 12158 29040 12186
rect 28816 11892 28868 11898
rect 28816 11834 28868 11840
rect 28920 11762 28948 12158
rect 29104 12050 29132 12838
rect 29184 12776 29236 12782
rect 29184 12718 29236 12724
rect 29274 12744 29330 12753
rect 29012 12022 29132 12050
rect 28908 11756 28960 11762
rect 28908 11698 28960 11704
rect 28816 11552 28868 11558
rect 28816 11494 28868 11500
rect 28828 10606 28856 11494
rect 28816 10600 28868 10606
rect 28816 10542 28868 10548
rect 29012 9178 29040 12022
rect 29196 11914 29224 12718
rect 29274 12679 29276 12688
rect 29328 12679 29330 12688
rect 29276 12650 29328 12656
rect 29274 12472 29330 12481
rect 29274 12407 29330 12416
rect 29104 11886 29224 11914
rect 29104 11694 29132 11886
rect 29288 11762 29316 12407
rect 29184 11756 29236 11762
rect 29184 11698 29236 11704
rect 29276 11756 29328 11762
rect 29276 11698 29328 11704
rect 29092 11688 29144 11694
rect 29092 11630 29144 11636
rect 29196 11642 29224 11698
rect 29196 11614 29316 11642
rect 29092 11552 29144 11558
rect 29092 11494 29144 11500
rect 29104 10606 29132 11494
rect 29184 10736 29236 10742
rect 29184 10678 29236 10684
rect 29092 10600 29144 10606
rect 29092 10542 29144 10548
rect 29000 9172 29052 9178
rect 29000 9114 29052 9120
rect 28816 7744 28868 7750
rect 28816 7686 28868 7692
rect 28724 7540 28776 7546
rect 28724 7482 28776 7488
rect 28630 6216 28686 6225
rect 28630 6151 28686 6160
rect 28644 6118 28672 6151
rect 28632 6112 28684 6118
rect 28632 6054 28684 6060
rect 28540 5772 28592 5778
rect 28540 5714 28592 5720
rect 28448 5296 28500 5302
rect 28448 5238 28500 5244
rect 28722 5128 28778 5137
rect 28722 5063 28778 5072
rect 28356 4820 28408 4826
rect 28356 4762 28408 4768
rect 28264 4616 28316 4622
rect 28264 4558 28316 4564
rect 28264 3528 28316 3534
rect 28368 3516 28396 4762
rect 28538 4040 28594 4049
rect 28538 3975 28594 3984
rect 28552 3534 28580 3975
rect 28316 3488 28396 3516
rect 28540 3528 28592 3534
rect 28264 3470 28316 3476
rect 28540 3470 28592 3476
rect 28276 2514 28304 3470
rect 28264 2508 28316 2514
rect 28264 2450 28316 2456
rect 28736 2106 28764 5063
rect 28828 3534 28856 7686
rect 28908 7472 28960 7478
rect 28908 7414 28960 7420
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 28920 2514 28948 7414
rect 29000 7200 29052 7206
rect 29000 7142 29052 7148
rect 29012 5234 29040 7142
rect 29104 6662 29132 10542
rect 29196 9586 29224 10678
rect 29288 10538 29316 11614
rect 29276 10532 29328 10538
rect 29276 10474 29328 10480
rect 29184 9580 29236 9586
rect 29184 9522 29236 9528
rect 29092 6656 29144 6662
rect 29092 6598 29144 6604
rect 29196 5302 29224 9522
rect 29380 9178 29408 13631
rect 29472 12986 29500 20198
rect 29564 19417 29592 20198
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29550 19408 29606 19417
rect 29550 19343 29606 19352
rect 29552 19236 29604 19242
rect 29552 19178 29604 19184
rect 29564 18358 29592 19178
rect 29552 18352 29604 18358
rect 29552 18294 29604 18300
rect 29564 17270 29592 18294
rect 29552 17264 29604 17270
rect 29552 17206 29604 17212
rect 29564 17105 29592 17206
rect 29550 17096 29606 17105
rect 29550 17031 29606 17040
rect 29552 16992 29604 16998
rect 29552 16934 29604 16940
rect 29564 14958 29592 16934
rect 29552 14952 29604 14958
rect 29552 14894 29604 14900
rect 29564 13190 29592 14894
rect 29552 13184 29604 13190
rect 29552 13126 29604 13132
rect 29656 12986 29684 19790
rect 29748 18737 29776 21286
rect 29840 21026 29868 21354
rect 29932 21146 29960 21354
rect 29920 21140 29972 21146
rect 29920 21082 29972 21088
rect 29840 20998 29960 21026
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 29734 18728 29790 18737
rect 29734 18663 29790 18672
rect 29736 17672 29788 17678
rect 29736 17614 29788 17620
rect 29748 15638 29776 17614
rect 29736 15632 29788 15638
rect 29736 15574 29788 15580
rect 29736 14884 29788 14890
rect 29736 14826 29788 14832
rect 29460 12980 29512 12986
rect 29460 12922 29512 12928
rect 29644 12980 29696 12986
rect 29644 12922 29696 12928
rect 29460 11688 29512 11694
rect 29460 11630 29512 11636
rect 29472 11558 29500 11630
rect 29460 11552 29512 11558
rect 29460 11494 29512 11500
rect 29644 11552 29696 11558
rect 29644 11494 29696 11500
rect 29656 11286 29684 11494
rect 29644 11280 29696 11286
rect 29644 11222 29696 11228
rect 29552 11144 29604 11150
rect 29552 11086 29604 11092
rect 29460 11008 29512 11014
rect 29460 10950 29512 10956
rect 29368 9172 29420 9178
rect 29368 9114 29420 9120
rect 29472 8430 29500 10950
rect 29460 8424 29512 8430
rect 29460 8366 29512 8372
rect 29276 8288 29328 8294
rect 29276 8230 29328 8236
rect 29288 7342 29316 8230
rect 29564 8090 29592 11086
rect 29748 10810 29776 14826
rect 29840 12986 29868 20878
rect 29932 20398 29960 20998
rect 29920 20392 29972 20398
rect 29920 20334 29972 20340
rect 29932 19310 29960 20334
rect 30104 20324 30156 20330
rect 30104 20266 30156 20272
rect 30116 19514 30144 20266
rect 30104 19508 30156 19514
rect 30104 19450 30156 19456
rect 29920 19304 29972 19310
rect 29920 19246 29972 19252
rect 29932 18154 29960 19246
rect 30012 19168 30064 19174
rect 30012 19110 30064 19116
rect 30104 19168 30156 19174
rect 30104 19110 30156 19116
rect 30024 18834 30052 19110
rect 30012 18828 30064 18834
rect 30012 18770 30064 18776
rect 29920 18148 29972 18154
rect 29920 18090 29972 18096
rect 29932 17898 29960 18090
rect 30024 18068 30052 18770
rect 30116 18329 30144 19110
rect 30102 18320 30158 18329
rect 30102 18255 30158 18264
rect 30104 18080 30156 18086
rect 30024 18040 30104 18068
rect 30104 18022 30156 18028
rect 30196 18080 30248 18086
rect 30196 18022 30248 18028
rect 29932 17870 30052 17898
rect 29920 17672 29972 17678
rect 29920 17614 29972 17620
rect 29932 14618 29960 17614
rect 30024 17066 30052 17870
rect 30116 17542 30144 18022
rect 30104 17536 30156 17542
rect 30104 17478 30156 17484
rect 30012 17060 30064 17066
rect 30012 17002 30064 17008
rect 30024 16182 30052 17002
rect 30102 16688 30158 16697
rect 30102 16623 30104 16632
rect 30156 16623 30158 16632
rect 30104 16594 30156 16600
rect 30104 16448 30156 16454
rect 30104 16390 30156 16396
rect 30208 16402 30236 18022
rect 30300 16726 30328 21966
rect 30564 21616 30616 21622
rect 30564 21558 30616 21564
rect 30380 18080 30432 18086
rect 30378 18048 30380 18057
rect 30432 18048 30434 18057
rect 30378 17983 30434 17992
rect 30380 16992 30432 16998
rect 30380 16934 30432 16940
rect 30288 16720 30340 16726
rect 30288 16662 30340 16668
rect 30012 16176 30064 16182
rect 30012 16118 30064 16124
rect 30012 16040 30064 16046
rect 30012 15982 30064 15988
rect 30024 15881 30052 15982
rect 30116 15978 30144 16390
rect 30208 16374 30328 16402
rect 30194 16280 30250 16289
rect 30194 16215 30250 16224
rect 30104 15972 30156 15978
rect 30104 15914 30156 15920
rect 30010 15872 30066 15881
rect 30010 15807 30066 15816
rect 30012 15360 30064 15366
rect 30012 15302 30064 15308
rect 29920 14612 29972 14618
rect 29920 14554 29972 14560
rect 29918 14512 29974 14521
rect 29918 14447 29920 14456
rect 29972 14447 29974 14456
rect 29920 14418 29972 14424
rect 29920 14340 29972 14346
rect 29920 14282 29972 14288
rect 29828 12980 29880 12986
rect 29828 12922 29880 12928
rect 29932 12782 29960 14282
rect 30024 13394 30052 15302
rect 30104 15156 30156 15162
rect 30104 15098 30156 15104
rect 30012 13388 30064 13394
rect 30012 13330 30064 13336
rect 29920 12776 29972 12782
rect 30012 12776 30064 12782
rect 29920 12718 29972 12724
rect 30010 12744 30012 12753
rect 30064 12744 30066 12753
rect 29932 12374 29960 12718
rect 30010 12679 30066 12688
rect 29920 12368 29972 12374
rect 29840 12316 29920 12322
rect 29840 12310 29972 12316
rect 29840 12294 29960 12310
rect 29840 11694 29868 12294
rect 29918 12200 29974 12209
rect 29918 12135 29974 12144
rect 29932 11694 29960 12135
rect 29828 11688 29880 11694
rect 29828 11630 29880 11636
rect 29920 11688 29972 11694
rect 29920 11630 29972 11636
rect 30116 10810 30144 15098
rect 30208 12442 30236 16215
rect 30300 15502 30328 16374
rect 30288 15496 30340 15502
rect 30288 15438 30340 15444
rect 30288 14000 30340 14006
rect 30288 13942 30340 13948
rect 30300 13841 30328 13942
rect 30392 13938 30420 16934
rect 30472 16652 30524 16658
rect 30472 16594 30524 16600
rect 30484 14226 30512 16594
rect 30576 14482 30604 21558
rect 31116 21480 31168 21486
rect 31116 21422 31168 21428
rect 30758 21244 31066 21253
rect 30758 21242 30764 21244
rect 30820 21242 30844 21244
rect 30900 21242 30924 21244
rect 30980 21242 31004 21244
rect 31060 21242 31066 21244
rect 30820 21190 30822 21242
rect 31002 21190 31004 21242
rect 30758 21188 30764 21190
rect 30820 21188 30844 21190
rect 30900 21188 30924 21190
rect 30980 21188 31004 21190
rect 31060 21188 31066 21190
rect 30758 21179 31066 21188
rect 30758 20156 31066 20165
rect 30758 20154 30764 20156
rect 30820 20154 30844 20156
rect 30900 20154 30924 20156
rect 30980 20154 31004 20156
rect 31060 20154 31066 20156
rect 30820 20102 30822 20154
rect 31002 20102 31004 20154
rect 30758 20100 30764 20102
rect 30820 20100 30844 20102
rect 30900 20100 30924 20102
rect 30980 20100 31004 20102
rect 31060 20100 31066 20102
rect 30758 20091 31066 20100
rect 30656 19168 30708 19174
rect 30656 19110 30708 19116
rect 30668 18193 30696 19110
rect 30758 19068 31066 19077
rect 30758 19066 30764 19068
rect 30820 19066 30844 19068
rect 30900 19066 30924 19068
rect 30980 19066 31004 19068
rect 31060 19066 31066 19068
rect 30820 19014 30822 19066
rect 31002 19014 31004 19066
rect 30758 19012 30764 19014
rect 30820 19012 30844 19014
rect 30900 19012 30924 19014
rect 30980 19012 31004 19014
rect 31060 19012 31066 19014
rect 30758 19003 31066 19012
rect 30654 18184 30710 18193
rect 30654 18119 30710 18128
rect 30668 18086 30696 18119
rect 30656 18080 30708 18086
rect 30656 18022 30708 18028
rect 30668 15502 30696 18022
rect 30758 17980 31066 17989
rect 30758 17978 30764 17980
rect 30820 17978 30844 17980
rect 30900 17978 30924 17980
rect 30980 17978 31004 17980
rect 31060 17978 31066 17980
rect 30820 17926 30822 17978
rect 31002 17926 31004 17978
rect 30758 17924 30764 17926
rect 30820 17924 30844 17926
rect 30900 17924 30924 17926
rect 30980 17924 31004 17926
rect 31060 17924 31066 17926
rect 30758 17915 31066 17924
rect 30758 16892 31066 16901
rect 30758 16890 30764 16892
rect 30820 16890 30844 16892
rect 30900 16890 30924 16892
rect 30980 16890 31004 16892
rect 31060 16890 31066 16892
rect 30820 16838 30822 16890
rect 31002 16838 31004 16890
rect 30758 16836 30764 16838
rect 30820 16836 30844 16838
rect 30900 16836 30924 16838
rect 30980 16836 31004 16838
rect 31060 16836 31066 16838
rect 30758 16827 31066 16836
rect 31128 16017 31156 21422
rect 31114 16008 31170 16017
rect 31114 15943 31170 15952
rect 30758 15804 31066 15813
rect 30758 15802 30764 15804
rect 30820 15802 30844 15804
rect 30900 15802 30924 15804
rect 30980 15802 31004 15804
rect 31060 15802 31066 15804
rect 30820 15750 30822 15802
rect 31002 15750 31004 15802
rect 30758 15748 30764 15750
rect 30820 15748 30844 15750
rect 30900 15748 30924 15750
rect 30980 15748 31004 15750
rect 31060 15748 31066 15750
rect 30758 15739 31066 15748
rect 30656 15496 30708 15502
rect 30656 15438 30708 15444
rect 30564 14476 30616 14482
rect 30564 14418 30616 14424
rect 30564 14272 30616 14278
rect 30484 14220 30564 14226
rect 30484 14214 30616 14220
rect 30484 14198 30604 14214
rect 30484 14074 30512 14198
rect 30472 14068 30524 14074
rect 30472 14010 30524 14016
rect 30380 13932 30432 13938
rect 30380 13874 30432 13880
rect 30286 13832 30342 13841
rect 30286 13767 30342 13776
rect 30286 13696 30342 13705
rect 30286 13631 30342 13640
rect 30300 13530 30328 13631
rect 30392 13546 30420 13874
rect 30564 13728 30616 13734
rect 30564 13670 30616 13676
rect 30288 13524 30340 13530
rect 30392 13518 30512 13546
rect 30288 13466 30340 13472
rect 30484 13462 30512 13518
rect 30472 13456 30524 13462
rect 30472 13398 30524 13404
rect 30288 13184 30340 13190
rect 30288 13126 30340 13132
rect 30196 12436 30248 12442
rect 30196 12378 30248 12384
rect 30300 11898 30328 13126
rect 30288 11892 30340 11898
rect 30484 11880 30512 13398
rect 30576 12782 30604 13670
rect 30564 12776 30616 12782
rect 30564 12718 30616 12724
rect 30668 12714 30696 15438
rect 31116 14816 31168 14822
rect 31116 14758 31168 14764
rect 30758 14716 31066 14725
rect 30758 14714 30764 14716
rect 30820 14714 30844 14716
rect 30900 14714 30924 14716
rect 30980 14714 31004 14716
rect 31060 14714 31066 14716
rect 30820 14662 30822 14714
rect 31002 14662 31004 14714
rect 30758 14660 30764 14662
rect 30820 14660 30844 14662
rect 30900 14660 30924 14662
rect 30980 14660 31004 14662
rect 31060 14660 31066 14662
rect 30758 14651 31066 14660
rect 31128 14482 31156 14758
rect 31116 14476 31168 14482
rect 31116 14418 31168 14424
rect 30758 13628 31066 13637
rect 30758 13626 30764 13628
rect 30820 13626 30844 13628
rect 30900 13626 30924 13628
rect 30980 13626 31004 13628
rect 31060 13626 31066 13628
rect 30820 13574 30822 13626
rect 31002 13574 31004 13626
rect 30758 13572 30764 13574
rect 30820 13572 30844 13574
rect 30900 13572 30924 13574
rect 30980 13572 31004 13574
rect 31060 13572 31066 13574
rect 30758 13563 31066 13572
rect 30656 12708 30708 12714
rect 30656 12650 30708 12656
rect 30758 12540 31066 12549
rect 30758 12538 30764 12540
rect 30820 12538 30844 12540
rect 30900 12538 30924 12540
rect 30980 12538 31004 12540
rect 31060 12538 31066 12540
rect 30820 12486 30822 12538
rect 31002 12486 31004 12538
rect 30758 12484 30764 12486
rect 30820 12484 30844 12486
rect 30900 12484 30924 12486
rect 30980 12484 31004 12486
rect 31060 12484 31066 12486
rect 30758 12475 31066 12484
rect 30484 11852 30696 11880
rect 30288 11834 30340 11840
rect 30380 11824 30432 11830
rect 30286 11792 30342 11801
rect 30380 11766 30432 11772
rect 30286 11727 30342 11736
rect 30300 11218 30328 11727
rect 30392 11665 30420 11766
rect 30472 11756 30524 11762
rect 30472 11698 30524 11704
rect 30378 11656 30434 11665
rect 30378 11591 30434 11600
rect 30484 11354 30512 11698
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 30472 11348 30524 11354
rect 30472 11290 30524 11296
rect 30288 11212 30340 11218
rect 30288 11154 30340 11160
rect 29644 10804 29696 10810
rect 29644 10746 29696 10752
rect 29736 10804 29788 10810
rect 29736 10746 29788 10752
rect 30104 10804 30156 10810
rect 30104 10746 30156 10752
rect 29656 10130 29684 10746
rect 30104 10668 30156 10674
rect 30104 10610 30156 10616
rect 29828 10464 29880 10470
rect 29828 10406 29880 10412
rect 29920 10464 29972 10470
rect 29920 10406 29972 10412
rect 29644 10124 29696 10130
rect 29644 10066 29696 10072
rect 29736 8288 29788 8294
rect 29736 8230 29788 8236
rect 29552 8084 29604 8090
rect 29552 8026 29604 8032
rect 29644 7948 29696 7954
rect 29644 7890 29696 7896
rect 29276 7336 29328 7342
rect 29276 7278 29328 7284
rect 29184 5296 29236 5302
rect 29184 5238 29236 5244
rect 29000 5228 29052 5234
rect 29000 5170 29052 5176
rect 29000 5024 29052 5030
rect 29052 4984 29132 5012
rect 29000 4966 29052 4972
rect 29000 4684 29052 4690
rect 29000 4626 29052 4632
rect 28908 2508 28960 2514
rect 28908 2450 28960 2456
rect 28724 2100 28776 2106
rect 28724 2042 28776 2048
rect 29012 1562 29040 4626
rect 29000 1556 29052 1562
rect 29000 1498 29052 1504
rect 28080 1352 28132 1358
rect 28080 1294 28132 1300
rect 28172 1352 28224 1358
rect 28172 1294 28224 1300
rect 28172 1216 28224 1222
rect 28172 1158 28224 1164
rect 28184 950 28212 1158
rect 28172 944 28224 950
rect 28172 886 28224 892
rect 29104 814 29132 4984
rect 29288 1970 29316 7278
rect 29552 7200 29604 7206
rect 29552 7142 29604 7148
rect 29564 1970 29592 7142
rect 29656 2310 29684 7890
rect 29748 7274 29776 8230
rect 29736 7268 29788 7274
rect 29736 7210 29788 7216
rect 29840 6866 29868 10406
rect 29932 7410 29960 10406
rect 30012 9920 30064 9926
rect 30012 9862 30064 9868
rect 30024 9042 30052 9862
rect 30012 9036 30064 9042
rect 30012 8978 30064 8984
rect 30116 8922 30144 10610
rect 30024 8894 30144 8922
rect 30024 8362 30052 8894
rect 30012 8356 30064 8362
rect 30012 8298 30064 8304
rect 29920 7404 29972 7410
rect 29920 7346 29972 7352
rect 30024 7290 30052 8298
rect 30104 8288 30156 8294
rect 30104 8230 30156 8236
rect 30116 7954 30144 8230
rect 30104 7948 30156 7954
rect 30104 7890 30156 7896
rect 29932 7262 30052 7290
rect 29828 6860 29880 6866
rect 29828 6802 29880 6808
rect 29644 2304 29696 2310
rect 29644 2246 29696 2252
rect 29276 1964 29328 1970
rect 29276 1906 29328 1912
rect 29552 1964 29604 1970
rect 29552 1906 29604 1912
rect 29182 1864 29238 1873
rect 29182 1799 29238 1808
rect 29196 1766 29224 1799
rect 29184 1760 29236 1766
rect 29184 1702 29236 1708
rect 29932 1018 29960 7262
rect 30576 6254 30604 11630
rect 30668 11014 30696 11852
rect 31128 11762 31156 14418
rect 31220 13190 31248 22238
rect 31298 18728 31354 18737
rect 31298 18663 31354 18672
rect 31312 13433 31340 18663
rect 31390 16008 31446 16017
rect 31390 15943 31446 15952
rect 31298 13424 31354 13433
rect 31298 13359 31354 13368
rect 31208 13184 31260 13190
rect 31208 13126 31260 13132
rect 31208 12844 31260 12850
rect 31208 12786 31260 12792
rect 31116 11756 31168 11762
rect 31116 11698 31168 11704
rect 30758 11452 31066 11461
rect 30758 11450 30764 11452
rect 30820 11450 30844 11452
rect 30900 11450 30924 11452
rect 30980 11450 31004 11452
rect 31060 11450 31066 11452
rect 30820 11398 30822 11450
rect 31002 11398 31004 11450
rect 30758 11396 30764 11398
rect 30820 11396 30844 11398
rect 30900 11396 30924 11398
rect 30980 11396 31004 11398
rect 31060 11396 31066 11398
rect 30758 11387 31066 11396
rect 30656 11008 30708 11014
rect 30656 10950 30708 10956
rect 30758 10364 31066 10373
rect 30758 10362 30764 10364
rect 30820 10362 30844 10364
rect 30900 10362 30924 10364
rect 30980 10362 31004 10364
rect 31060 10362 31066 10364
rect 30820 10310 30822 10362
rect 31002 10310 31004 10362
rect 30758 10308 30764 10310
rect 30820 10308 30844 10310
rect 30900 10308 30924 10310
rect 30980 10308 31004 10310
rect 31060 10308 31066 10310
rect 30758 10299 31066 10308
rect 30758 9276 31066 9285
rect 30758 9274 30764 9276
rect 30820 9274 30844 9276
rect 30900 9274 30924 9276
rect 30980 9274 31004 9276
rect 31060 9274 31066 9276
rect 30820 9222 30822 9274
rect 31002 9222 31004 9274
rect 30758 9220 30764 9222
rect 30820 9220 30844 9222
rect 30900 9220 30924 9222
rect 30980 9220 31004 9222
rect 31060 9220 31066 9222
rect 30758 9211 31066 9220
rect 30758 8188 31066 8197
rect 30758 8186 30764 8188
rect 30820 8186 30844 8188
rect 30900 8186 30924 8188
rect 30980 8186 31004 8188
rect 31060 8186 31066 8188
rect 30820 8134 30822 8186
rect 31002 8134 31004 8186
rect 30758 8132 30764 8134
rect 30820 8132 30844 8134
rect 30900 8132 30924 8134
rect 30980 8132 31004 8134
rect 31060 8132 31066 8134
rect 30758 8123 31066 8132
rect 30758 7100 31066 7109
rect 30758 7098 30764 7100
rect 30820 7098 30844 7100
rect 30900 7098 30924 7100
rect 30980 7098 31004 7100
rect 31060 7098 31066 7100
rect 30820 7046 30822 7098
rect 31002 7046 31004 7098
rect 30758 7044 30764 7046
rect 30820 7044 30844 7046
rect 30900 7044 30924 7046
rect 30980 7044 31004 7046
rect 31060 7044 31066 7046
rect 30758 7035 31066 7044
rect 31220 6662 31248 12786
rect 31404 8430 31432 15943
rect 31392 8424 31444 8430
rect 31392 8366 31444 8372
rect 31208 6656 31260 6662
rect 31208 6598 31260 6604
rect 30564 6248 30616 6254
rect 30564 6190 30616 6196
rect 30758 6012 31066 6021
rect 30758 6010 30764 6012
rect 30820 6010 30844 6012
rect 30900 6010 30924 6012
rect 30980 6010 31004 6012
rect 31060 6010 31066 6012
rect 30820 5958 30822 6010
rect 31002 5958 31004 6010
rect 30758 5956 30764 5958
rect 30820 5956 30844 5958
rect 30900 5956 30924 5958
rect 30980 5956 31004 5958
rect 31060 5956 31066 5958
rect 30758 5947 31066 5956
rect 30758 4924 31066 4933
rect 30758 4922 30764 4924
rect 30820 4922 30844 4924
rect 30900 4922 30924 4924
rect 30980 4922 31004 4924
rect 31060 4922 31066 4924
rect 30820 4870 30822 4922
rect 31002 4870 31004 4922
rect 30758 4868 30764 4870
rect 30820 4868 30844 4870
rect 30900 4868 30924 4870
rect 30980 4868 31004 4870
rect 31060 4868 31066 4870
rect 30758 4859 31066 4868
rect 30758 3836 31066 3845
rect 30758 3834 30764 3836
rect 30820 3834 30844 3836
rect 30900 3834 30924 3836
rect 30980 3834 31004 3836
rect 31060 3834 31066 3836
rect 30820 3782 30822 3834
rect 31002 3782 31004 3834
rect 30758 3780 30764 3782
rect 30820 3780 30844 3782
rect 30900 3780 30924 3782
rect 30980 3780 31004 3782
rect 31060 3780 31066 3782
rect 30758 3771 31066 3780
rect 30012 3188 30064 3194
rect 30012 3130 30064 3136
rect 30024 2650 30052 3130
rect 30758 2748 31066 2757
rect 30758 2746 30764 2748
rect 30820 2746 30844 2748
rect 30900 2746 30924 2748
rect 30980 2746 31004 2748
rect 31060 2746 31066 2748
rect 30820 2694 30822 2746
rect 31002 2694 31004 2746
rect 30758 2692 30764 2694
rect 30820 2692 30844 2694
rect 30900 2692 30924 2694
rect 30980 2692 31004 2694
rect 31060 2692 31066 2694
rect 30758 2683 31066 2692
rect 30012 2644 30064 2650
rect 30012 2586 30064 2592
rect 30758 1660 31066 1669
rect 30758 1658 30764 1660
rect 30820 1658 30844 1660
rect 30900 1658 30924 1660
rect 30980 1658 31004 1660
rect 31060 1658 31066 1660
rect 30820 1606 30822 1658
rect 31002 1606 31004 1658
rect 30758 1604 30764 1606
rect 30820 1604 30844 1606
rect 30900 1604 30924 1606
rect 30980 1604 31004 1606
rect 31060 1604 31066 1606
rect 30758 1595 31066 1604
rect 29920 1012 29972 1018
rect 29920 954 29972 960
rect 29092 808 29144 814
rect 29092 750 29144 756
rect 27804 672 27856 678
rect 27804 614 27856 620
rect 30758 572 31066 581
rect 30758 570 30764 572
rect 30820 570 30844 572
rect 30900 570 30924 572
rect 30980 570 31004 572
rect 31060 570 31066 572
rect 30820 518 30822 570
rect 31002 518 31004 570
rect 30758 516 30764 518
rect 30820 516 30844 518
rect 30900 516 30924 518
rect 30980 516 31004 518
rect 31060 516 31066 518
rect 30758 507 31066 516
rect 25688 468 25740 474
rect 25688 410 25740 416
rect 24860 342 24912 348
rect 25318 368 25374 377
rect 25318 303 25374 312
rect 24124 196 24176 202
rect 24124 138 24176 144
rect 11796 128 11848 134
rect 11796 70 11848 76
rect 18328 128 18380 134
rect 18328 70 18380 76
rect 4712 60 4764 66
rect 4712 2 4764 8
rect 6000 60 6052 66
rect 6000 2 6052 8
rect 9772 60 9824 66
rect 9772 2 9824 8
<< via2 >>
rect 10966 22244 10968 22264
rect 10968 22244 11020 22264
rect 11020 22244 11022 22264
rect 10966 22208 11022 22244
rect 4199 21786 4255 21788
rect 4279 21786 4335 21788
rect 4359 21786 4415 21788
rect 4439 21786 4495 21788
rect 4199 21734 4245 21786
rect 4245 21734 4255 21786
rect 4279 21734 4309 21786
rect 4309 21734 4321 21786
rect 4321 21734 4335 21786
rect 4359 21734 4373 21786
rect 4373 21734 4385 21786
rect 4385 21734 4415 21786
rect 4439 21734 4449 21786
rect 4449 21734 4495 21786
rect 4199 21732 4255 21734
rect 4279 21732 4335 21734
rect 4359 21732 4415 21734
rect 4439 21732 4495 21734
rect 1674 21004 1730 21040
rect 1674 20984 1676 21004
rect 1676 20984 1728 21004
rect 1728 20984 1730 21004
rect 1674 20460 1730 20496
rect 1674 20440 1676 20460
rect 1676 20440 1728 20460
rect 1728 20440 1730 20460
rect 1398 18672 1454 18728
rect 1306 18128 1362 18184
rect 1674 19352 1730 19408
rect 1766 16768 1822 16824
rect 1214 12144 1270 12200
rect 1766 12280 1822 12336
rect 1490 10104 1546 10160
rect 2134 15952 2190 16008
rect 2042 15444 2044 15464
rect 2044 15444 2096 15464
rect 2096 15444 2098 15464
rect 2042 15408 2098 15444
rect 2134 15020 2190 15056
rect 2134 15000 2136 15020
rect 2136 15000 2188 15020
rect 2188 15000 2190 15020
rect 2042 14456 2098 14512
rect 1950 13368 2006 13424
rect 1950 11192 2006 11248
rect 1858 10920 1914 10976
rect 1674 9968 1730 10024
rect 1122 7112 1178 7168
rect 1490 7828 1492 7848
rect 1492 7828 1544 7848
rect 1544 7828 1546 7848
rect 1490 7792 1546 7828
rect 1398 5344 1454 5400
rect 1582 6296 1638 6352
rect 1766 9036 1822 9072
rect 1766 9016 1768 9036
rect 1768 9016 1820 9036
rect 1820 9016 1822 9036
rect 1766 7248 1822 7304
rect 1674 3032 1730 3088
rect 1674 1964 1730 2000
rect 1674 1944 1676 1964
rect 1676 1944 1728 1964
rect 1728 1944 1730 1964
rect 2134 12844 2190 12880
rect 2134 12824 2136 12844
rect 2136 12824 2188 12844
rect 2188 12824 2190 12844
rect 2686 16088 2742 16144
rect 2410 13504 2466 13560
rect 2318 12416 2374 12472
rect 2226 12280 2282 12336
rect 2778 13232 2834 13288
rect 2962 20748 2964 20768
rect 2964 20748 3016 20768
rect 3016 20748 3018 20768
rect 2962 20712 3018 20748
rect 3606 19760 3662 19816
rect 3054 13812 3056 13832
rect 3056 13812 3108 13832
rect 3108 13812 3110 13832
rect 3054 13776 3110 13812
rect 4199 20698 4255 20700
rect 4279 20698 4335 20700
rect 4359 20698 4415 20700
rect 4439 20698 4495 20700
rect 4199 20646 4245 20698
rect 4245 20646 4255 20698
rect 4279 20646 4309 20698
rect 4309 20646 4321 20698
rect 4321 20646 4335 20698
rect 4359 20646 4373 20698
rect 4373 20646 4385 20698
rect 4385 20646 4415 20698
rect 4439 20646 4449 20698
rect 4449 20646 4495 20698
rect 4199 20644 4255 20646
rect 4279 20644 4335 20646
rect 4359 20644 4415 20646
rect 4439 20644 4495 20646
rect 3882 19080 3938 19136
rect 4199 19610 4255 19612
rect 4279 19610 4335 19612
rect 4359 19610 4415 19612
rect 4439 19610 4495 19612
rect 4199 19558 4245 19610
rect 4245 19558 4255 19610
rect 4279 19558 4309 19610
rect 4309 19558 4321 19610
rect 4321 19558 4335 19610
rect 4359 19558 4373 19610
rect 4373 19558 4385 19610
rect 4385 19558 4415 19610
rect 4439 19558 4449 19610
rect 4449 19558 4495 19610
rect 4199 19556 4255 19558
rect 4279 19556 4335 19558
rect 4359 19556 4415 19558
rect 4439 19556 4495 19558
rect 4199 18522 4255 18524
rect 4279 18522 4335 18524
rect 4359 18522 4415 18524
rect 4439 18522 4495 18524
rect 4199 18470 4245 18522
rect 4245 18470 4255 18522
rect 4279 18470 4309 18522
rect 4309 18470 4321 18522
rect 4321 18470 4335 18522
rect 4359 18470 4373 18522
rect 4373 18470 4385 18522
rect 4385 18470 4415 18522
rect 4439 18470 4449 18522
rect 4449 18470 4495 18522
rect 4199 18468 4255 18470
rect 4279 18468 4335 18470
rect 4359 18468 4415 18470
rect 4439 18468 4495 18470
rect 4618 18400 4674 18456
rect 4618 17992 4674 18048
rect 3790 17720 3846 17776
rect 4199 17434 4255 17436
rect 4279 17434 4335 17436
rect 4359 17434 4415 17436
rect 4439 17434 4495 17436
rect 4199 17382 4245 17434
rect 4245 17382 4255 17434
rect 4279 17382 4309 17434
rect 4309 17382 4321 17434
rect 4321 17382 4335 17434
rect 4359 17382 4373 17434
rect 4373 17382 4385 17434
rect 4385 17382 4415 17434
rect 4439 17382 4449 17434
rect 4449 17382 4495 17434
rect 4199 17380 4255 17382
rect 4279 17380 4335 17382
rect 4359 17380 4415 17382
rect 4439 17380 4495 17382
rect 4066 16496 4122 16552
rect 4199 16346 4255 16348
rect 4279 16346 4335 16348
rect 4359 16346 4415 16348
rect 4439 16346 4495 16348
rect 4199 16294 4245 16346
rect 4245 16294 4255 16346
rect 4279 16294 4309 16346
rect 4309 16294 4321 16346
rect 4321 16294 4335 16346
rect 4359 16294 4373 16346
rect 4373 16294 4385 16346
rect 4385 16294 4415 16346
rect 4439 16294 4449 16346
rect 4449 16294 4495 16346
rect 4199 16292 4255 16294
rect 4279 16292 4335 16294
rect 4359 16292 4415 16294
rect 4439 16292 4495 16294
rect 4199 15258 4255 15260
rect 4279 15258 4335 15260
rect 4359 15258 4415 15260
rect 4439 15258 4495 15260
rect 4199 15206 4245 15258
rect 4245 15206 4255 15258
rect 4279 15206 4309 15258
rect 4309 15206 4321 15258
rect 4321 15206 4335 15258
rect 4359 15206 4373 15258
rect 4373 15206 4385 15258
rect 4385 15206 4415 15258
rect 4439 15206 4449 15258
rect 4449 15206 4495 15258
rect 4199 15204 4255 15206
rect 4279 15204 4335 15206
rect 4359 15204 4415 15206
rect 4439 15204 4495 15206
rect 4199 14170 4255 14172
rect 4279 14170 4335 14172
rect 4359 14170 4415 14172
rect 4439 14170 4495 14172
rect 4199 14118 4245 14170
rect 4245 14118 4255 14170
rect 4279 14118 4309 14170
rect 4309 14118 4321 14170
rect 4321 14118 4335 14170
rect 4359 14118 4373 14170
rect 4373 14118 4385 14170
rect 4385 14118 4415 14170
rect 4439 14118 4449 14170
rect 4449 14118 4495 14170
rect 4199 14116 4255 14118
rect 4279 14116 4335 14118
rect 4359 14116 4415 14118
rect 4439 14116 4495 14118
rect 4199 13082 4255 13084
rect 4279 13082 4335 13084
rect 4359 13082 4415 13084
rect 4439 13082 4495 13084
rect 4199 13030 4245 13082
rect 4245 13030 4255 13082
rect 4279 13030 4309 13082
rect 4309 13030 4321 13082
rect 4321 13030 4335 13082
rect 4359 13030 4373 13082
rect 4373 13030 4385 13082
rect 4385 13030 4415 13082
rect 4439 13030 4449 13082
rect 4449 13030 4495 13082
rect 4199 13028 4255 13030
rect 4279 13028 4335 13030
rect 4359 13028 4415 13030
rect 4439 13028 4495 13030
rect 4802 14320 4858 14376
rect 3238 11464 3294 11520
rect 3422 11328 3478 11384
rect 2134 5072 2190 5128
rect 2318 6860 2374 6896
rect 2318 6840 2320 6860
rect 2320 6840 2372 6860
rect 2372 6840 2374 6860
rect 2502 8372 2504 8392
rect 2504 8372 2556 8392
rect 2556 8372 2558 8392
rect 2502 8336 2558 8372
rect 2502 5616 2558 5672
rect 2686 7384 2742 7440
rect 2686 6024 2742 6080
rect 2318 4800 2374 4856
rect 3054 8064 3110 8120
rect 2870 4936 2926 4992
rect 2778 3984 2834 4040
rect 3146 6704 3202 6760
rect 3606 10648 3662 10704
rect 3698 10240 3754 10296
rect 3882 11464 3938 11520
rect 4199 11994 4255 11996
rect 4279 11994 4335 11996
rect 4359 11994 4415 11996
rect 4439 11994 4495 11996
rect 4199 11942 4245 11994
rect 4245 11942 4255 11994
rect 4279 11942 4309 11994
rect 4309 11942 4321 11994
rect 4321 11942 4335 11994
rect 4359 11942 4373 11994
rect 4373 11942 4385 11994
rect 4385 11942 4415 11994
rect 4439 11942 4449 11994
rect 4449 11942 4495 11994
rect 4199 11940 4255 11942
rect 4279 11940 4335 11942
rect 4359 11940 4415 11942
rect 4439 11940 4495 11942
rect 3974 10512 4030 10568
rect 3974 10240 4030 10296
rect 4802 11328 4858 11384
rect 4710 11056 4766 11112
rect 4199 10906 4255 10908
rect 4279 10906 4335 10908
rect 4359 10906 4415 10908
rect 4439 10906 4495 10908
rect 4199 10854 4245 10906
rect 4245 10854 4255 10906
rect 4279 10854 4309 10906
rect 4309 10854 4321 10906
rect 4321 10854 4335 10906
rect 4359 10854 4373 10906
rect 4373 10854 4385 10906
rect 4385 10854 4415 10906
rect 4439 10854 4449 10906
rect 4449 10854 4495 10906
rect 4199 10852 4255 10854
rect 4279 10852 4335 10854
rect 4359 10852 4415 10854
rect 4439 10852 4495 10854
rect 3422 9288 3478 9344
rect 4199 9818 4255 9820
rect 4279 9818 4335 9820
rect 4359 9818 4415 9820
rect 4439 9818 4495 9820
rect 4199 9766 4245 9818
rect 4245 9766 4255 9818
rect 4279 9766 4309 9818
rect 4309 9766 4321 9818
rect 4321 9766 4335 9818
rect 4359 9766 4373 9818
rect 4373 9766 4385 9818
rect 4385 9766 4415 9818
rect 4439 9766 4449 9818
rect 4449 9766 4495 9818
rect 4199 9764 4255 9766
rect 4279 9764 4335 9766
rect 4359 9764 4415 9766
rect 4439 9764 4495 9766
rect 4434 9288 4490 9344
rect 4526 9152 4582 9208
rect 4199 8730 4255 8732
rect 4279 8730 4335 8732
rect 4359 8730 4415 8732
rect 4439 8730 4495 8732
rect 4199 8678 4245 8730
rect 4245 8678 4255 8730
rect 4279 8678 4309 8730
rect 4309 8678 4321 8730
rect 4321 8678 4335 8730
rect 4359 8678 4373 8730
rect 4373 8678 4385 8730
rect 4385 8678 4415 8730
rect 4439 8678 4449 8730
rect 4449 8678 4495 8730
rect 4199 8676 4255 8678
rect 4279 8676 4335 8678
rect 4359 8676 4415 8678
rect 4439 8676 4495 8678
rect 3514 7828 3516 7848
rect 3516 7828 3568 7848
rect 3568 7828 3570 7848
rect 3514 7792 3570 7828
rect 3146 5480 3202 5536
rect 3422 5208 3478 5264
rect 4158 7828 4160 7848
rect 4160 7828 4212 7848
rect 4212 7828 4214 7848
rect 4158 7792 4214 7828
rect 4199 7642 4255 7644
rect 4279 7642 4335 7644
rect 4359 7642 4415 7644
rect 4439 7642 4495 7644
rect 4199 7590 4245 7642
rect 4245 7590 4255 7642
rect 4279 7590 4309 7642
rect 4309 7590 4321 7642
rect 4321 7590 4335 7642
rect 4359 7590 4373 7642
rect 4373 7590 4385 7642
rect 4385 7590 4415 7642
rect 4439 7590 4449 7642
rect 4449 7590 4495 7642
rect 4199 7588 4255 7590
rect 4279 7588 4335 7590
rect 4359 7588 4415 7590
rect 4439 7588 4495 7590
rect 4158 6840 4214 6896
rect 3974 6296 4030 6352
rect 4199 6554 4255 6556
rect 4279 6554 4335 6556
rect 4359 6554 4415 6556
rect 4439 6554 4495 6556
rect 4199 6502 4245 6554
rect 4245 6502 4255 6554
rect 4279 6502 4309 6554
rect 4309 6502 4321 6554
rect 4321 6502 4335 6554
rect 4359 6502 4373 6554
rect 4373 6502 4385 6554
rect 4385 6502 4415 6554
rect 4439 6502 4449 6554
rect 4449 6502 4495 6554
rect 4199 6500 4255 6502
rect 4279 6500 4335 6502
rect 4359 6500 4415 6502
rect 4439 6500 4495 6502
rect 3330 3848 3386 3904
rect 1858 2488 1914 2544
rect 2134 1400 2190 1456
rect 2042 1300 2044 1320
rect 2044 1300 2096 1320
rect 2096 1300 2098 1320
rect 2042 1264 2098 1300
rect 1674 876 1730 912
rect 1674 856 1676 876
rect 1676 856 1728 876
rect 1728 856 1730 876
rect 1490 720 1546 776
rect 4199 5466 4255 5468
rect 4279 5466 4335 5468
rect 4359 5466 4415 5468
rect 4439 5466 4495 5468
rect 4199 5414 4245 5466
rect 4245 5414 4255 5466
rect 4279 5414 4309 5466
rect 4309 5414 4321 5466
rect 4321 5414 4335 5466
rect 4359 5414 4373 5466
rect 4373 5414 4385 5466
rect 4385 5414 4415 5466
rect 4439 5414 4449 5466
rect 4449 5414 4495 5466
rect 4199 5412 4255 5414
rect 4279 5412 4335 5414
rect 4359 5412 4415 5414
rect 4439 5412 4495 5414
rect 3974 5344 4030 5400
rect 4434 4936 4490 4992
rect 4199 4378 4255 4380
rect 4279 4378 4335 4380
rect 4359 4378 4415 4380
rect 4439 4378 4495 4380
rect 4199 4326 4245 4378
rect 4245 4326 4255 4378
rect 4279 4326 4309 4378
rect 4309 4326 4321 4378
rect 4321 4326 4335 4378
rect 4359 4326 4373 4378
rect 4373 4326 4385 4378
rect 4385 4326 4415 4378
rect 4439 4326 4449 4378
rect 4449 4326 4495 4378
rect 4199 4324 4255 4326
rect 4279 4324 4335 4326
rect 4359 4324 4415 4326
rect 4439 4324 4495 4326
rect 3882 2896 3938 2952
rect 4250 3596 4306 3632
rect 4250 3576 4252 3596
rect 4252 3576 4304 3596
rect 4304 3576 4306 3596
rect 4199 3290 4255 3292
rect 4279 3290 4335 3292
rect 4359 3290 4415 3292
rect 4439 3290 4495 3292
rect 4199 3238 4245 3290
rect 4245 3238 4255 3290
rect 4279 3238 4309 3290
rect 4309 3238 4321 3290
rect 4321 3238 4335 3290
rect 4359 3238 4373 3290
rect 4373 3238 4385 3290
rect 4385 3238 4415 3290
rect 4439 3238 4449 3290
rect 4449 3238 4495 3290
rect 4199 3236 4255 3238
rect 4279 3236 4335 3238
rect 4359 3236 4415 3238
rect 4439 3236 4495 3238
rect 3974 2352 4030 2408
rect 5078 18844 5080 18864
rect 5080 18844 5132 18864
rect 5132 18844 5134 18864
rect 5078 18808 5134 18844
rect 4986 12144 5042 12200
rect 5446 20304 5502 20360
rect 5446 18672 5502 18728
rect 5354 18148 5410 18184
rect 5354 18128 5356 18148
rect 5356 18128 5408 18148
rect 5408 18128 5410 18148
rect 5906 21392 5962 21448
rect 5630 19352 5686 19408
rect 6182 19896 6238 19952
rect 5446 16904 5502 16960
rect 5630 16244 5686 16280
rect 5630 16224 5632 16244
rect 5632 16224 5684 16244
rect 5684 16224 5686 16244
rect 6274 19488 6330 19544
rect 6182 16632 6238 16688
rect 6458 18944 6514 19000
rect 6734 20712 6790 20768
rect 6918 19896 6974 19952
rect 6918 19388 6920 19408
rect 6920 19388 6972 19408
rect 6972 19388 6974 19408
rect 6918 19352 6974 19388
rect 6734 17992 6790 18048
rect 7010 16904 7066 16960
rect 6274 15544 6330 15600
rect 6182 15136 6238 15192
rect 6090 14864 6146 14920
rect 5538 14048 5594 14104
rect 5630 11328 5686 11384
rect 5354 10920 5410 10976
rect 5354 10668 5410 10704
rect 5354 10648 5356 10668
rect 5356 10648 5408 10668
rect 5408 10648 5410 10668
rect 5170 9832 5226 9888
rect 5354 9696 5410 9752
rect 5538 7384 5594 7440
rect 5262 6432 5318 6488
rect 6366 14184 6422 14240
rect 6090 12688 6146 12744
rect 6458 13504 6514 13560
rect 6458 13096 6514 13152
rect 5814 10648 5870 10704
rect 5814 9288 5870 9344
rect 5814 8200 5870 8256
rect 5814 7384 5870 7440
rect 6734 16496 6790 16552
rect 7562 20340 7564 20360
rect 7564 20340 7616 20360
rect 7616 20340 7618 20360
rect 7562 20304 7618 20340
rect 7562 18944 7618 19000
rect 7470 15408 7526 15464
rect 7286 14864 7342 14920
rect 7010 12416 7066 12472
rect 7102 12008 7158 12064
rect 6826 11328 6882 11384
rect 6090 7520 6146 7576
rect 5998 7420 6000 7440
rect 6000 7420 6052 7440
rect 6052 7420 6054 7440
rect 5998 7384 6054 7420
rect 6182 7112 6238 7168
rect 5630 6180 5686 6216
rect 5630 6160 5632 6180
rect 5632 6160 5684 6180
rect 5684 6160 5686 6180
rect 5538 5616 5594 5672
rect 5078 5480 5134 5536
rect 4710 4528 4766 4584
rect 4199 2202 4255 2204
rect 4279 2202 4335 2204
rect 4359 2202 4415 2204
rect 4439 2202 4495 2204
rect 4199 2150 4245 2202
rect 4245 2150 4255 2202
rect 4279 2150 4309 2202
rect 4309 2150 4321 2202
rect 4321 2150 4335 2202
rect 4359 2150 4373 2202
rect 4373 2150 4385 2202
rect 4385 2150 4415 2202
rect 4439 2150 4449 2202
rect 4449 2150 4495 2202
rect 4199 2148 4255 2150
rect 4279 2148 4335 2150
rect 4359 2148 4415 2150
rect 4439 2148 4495 2150
rect 5170 4936 5226 4992
rect 5078 4664 5134 4720
rect 4802 3984 4858 4040
rect 4199 1114 4255 1116
rect 4279 1114 4335 1116
rect 4359 1114 4415 1116
rect 4439 1114 4495 1116
rect 4199 1062 4245 1114
rect 4245 1062 4255 1114
rect 4279 1062 4309 1114
rect 4309 1062 4321 1114
rect 4321 1062 4335 1114
rect 4359 1062 4373 1114
rect 4373 1062 4385 1114
rect 4385 1062 4415 1114
rect 4439 1062 4449 1114
rect 4449 1062 4495 1114
rect 4199 1060 4255 1062
rect 4279 1060 4335 1062
rect 4359 1060 4415 1062
rect 4439 1060 4495 1062
rect 4894 620 4896 640
rect 4896 620 4948 640
rect 4948 620 4950 640
rect 4894 584 4950 620
rect 4802 176 4858 232
rect 5630 3476 5632 3496
rect 5632 3476 5684 3496
rect 5684 3476 5686 3496
rect 5630 3440 5686 3476
rect 6550 11056 6606 11112
rect 6642 9560 6698 9616
rect 6550 9288 6606 9344
rect 7010 9832 7066 9888
rect 6550 7656 6606 7712
rect 7470 12688 7526 12744
rect 7378 12552 7434 12608
rect 7654 12144 7710 12200
rect 6918 7928 6974 7984
rect 7010 7792 7066 7848
rect 6826 7540 6882 7576
rect 6826 7520 6828 7540
rect 6828 7520 6880 7540
rect 6880 7520 6882 7540
rect 7010 7384 7066 7440
rect 6918 6840 6974 6896
rect 7102 6976 7158 7032
rect 6734 6060 6736 6080
rect 6736 6060 6788 6080
rect 6788 6060 6790 6080
rect 6734 6024 6790 6060
rect 6182 5616 6238 5672
rect 6458 4800 6514 4856
rect 5998 2372 6054 2408
rect 5998 2352 6000 2372
rect 6000 2352 6052 2372
rect 6052 2352 6054 2372
rect 6918 5516 6920 5536
rect 6920 5516 6972 5536
rect 6972 5516 6974 5536
rect 6918 5480 6974 5516
rect 6734 5228 6790 5264
rect 6734 5208 6736 5228
rect 6736 5208 6788 5228
rect 6788 5208 6790 5228
rect 7286 8608 7342 8664
rect 7562 9152 7618 9208
rect 7994 21242 8050 21244
rect 8074 21242 8130 21244
rect 8154 21242 8210 21244
rect 8234 21242 8290 21244
rect 7994 21190 8040 21242
rect 8040 21190 8050 21242
rect 8074 21190 8104 21242
rect 8104 21190 8116 21242
rect 8116 21190 8130 21242
rect 8154 21190 8168 21242
rect 8168 21190 8180 21242
rect 8180 21190 8210 21242
rect 8234 21190 8244 21242
rect 8244 21190 8290 21242
rect 7994 21188 8050 21190
rect 8074 21188 8130 21190
rect 8154 21188 8210 21190
rect 8234 21188 8290 21190
rect 7838 20304 7894 20360
rect 7994 20154 8050 20156
rect 8074 20154 8130 20156
rect 8154 20154 8210 20156
rect 8234 20154 8290 20156
rect 7994 20102 8040 20154
rect 8040 20102 8050 20154
rect 8074 20102 8104 20154
rect 8104 20102 8116 20154
rect 8116 20102 8130 20154
rect 8154 20102 8168 20154
rect 8168 20102 8180 20154
rect 8180 20102 8210 20154
rect 8234 20102 8244 20154
rect 8244 20102 8290 20154
rect 7994 20100 8050 20102
rect 8074 20100 8130 20102
rect 8154 20100 8210 20102
rect 8234 20100 8290 20102
rect 7838 19080 7894 19136
rect 7994 19066 8050 19068
rect 8074 19066 8130 19068
rect 8154 19066 8210 19068
rect 8234 19066 8290 19068
rect 7994 19014 8040 19066
rect 8040 19014 8050 19066
rect 8074 19014 8104 19066
rect 8104 19014 8116 19066
rect 8116 19014 8130 19066
rect 8154 19014 8168 19066
rect 8168 19014 8180 19066
rect 8180 19014 8210 19066
rect 8234 19014 8244 19066
rect 8244 19014 8290 19066
rect 7994 19012 8050 19014
rect 8074 19012 8130 19014
rect 8154 19012 8210 19014
rect 8234 19012 8290 19014
rect 7838 18672 7894 18728
rect 9402 21392 9458 21448
rect 8942 20984 8998 21040
rect 8942 20576 8998 20632
rect 8850 20304 8906 20360
rect 8482 19080 8538 19136
rect 8574 18536 8630 18592
rect 8206 18300 8208 18320
rect 8208 18300 8260 18320
rect 8260 18300 8262 18320
rect 8206 18264 8262 18300
rect 8482 18264 8538 18320
rect 7994 17978 8050 17980
rect 8074 17978 8130 17980
rect 8154 17978 8210 17980
rect 8234 17978 8290 17980
rect 7994 17926 8040 17978
rect 8040 17926 8050 17978
rect 8074 17926 8104 17978
rect 8104 17926 8116 17978
rect 8116 17926 8130 17978
rect 8154 17926 8168 17978
rect 8168 17926 8180 17978
rect 8180 17926 8210 17978
rect 8234 17926 8244 17978
rect 8244 17926 8290 17978
rect 7994 17924 8050 17926
rect 8074 17924 8130 17926
rect 8154 17924 8210 17926
rect 8234 17924 8290 17926
rect 8390 17448 8446 17504
rect 8390 17196 8446 17232
rect 8758 17584 8814 17640
rect 8390 17176 8392 17196
rect 8392 17176 8444 17196
rect 8444 17176 8446 17196
rect 8482 17040 8538 17096
rect 7994 16890 8050 16892
rect 8074 16890 8130 16892
rect 8154 16890 8210 16892
rect 8234 16890 8290 16892
rect 7994 16838 8040 16890
rect 8040 16838 8050 16890
rect 8074 16838 8104 16890
rect 8104 16838 8116 16890
rect 8116 16838 8130 16890
rect 8154 16838 8168 16890
rect 8168 16838 8180 16890
rect 8180 16838 8210 16890
rect 8234 16838 8244 16890
rect 8244 16838 8290 16890
rect 7994 16836 8050 16838
rect 8074 16836 8130 16838
rect 8154 16836 8210 16838
rect 8234 16836 8290 16838
rect 9218 19352 9274 19408
rect 8942 18536 8998 18592
rect 8942 18264 8998 18320
rect 8942 18128 8998 18184
rect 9678 19216 9734 19272
rect 9678 19080 9734 19136
rect 9862 19080 9918 19136
rect 9126 17448 9182 17504
rect 7994 15802 8050 15804
rect 8074 15802 8130 15804
rect 8154 15802 8210 15804
rect 8234 15802 8290 15804
rect 7994 15750 8040 15802
rect 8040 15750 8050 15802
rect 8074 15750 8104 15802
rect 8104 15750 8116 15802
rect 8116 15750 8130 15802
rect 8154 15750 8168 15802
rect 8168 15750 8180 15802
rect 8180 15750 8210 15802
rect 8234 15750 8244 15802
rect 8244 15750 8290 15802
rect 7994 15748 8050 15750
rect 8074 15748 8130 15750
rect 8154 15748 8210 15750
rect 8234 15748 8290 15750
rect 8298 15564 8354 15600
rect 8298 15544 8300 15564
rect 8300 15544 8352 15564
rect 8352 15544 8354 15564
rect 8206 15136 8262 15192
rect 8482 14864 8538 14920
rect 7994 14714 8050 14716
rect 8074 14714 8130 14716
rect 8154 14714 8210 14716
rect 8234 14714 8290 14716
rect 7994 14662 8040 14714
rect 8040 14662 8050 14714
rect 8074 14662 8104 14714
rect 8104 14662 8116 14714
rect 8116 14662 8130 14714
rect 8154 14662 8168 14714
rect 8168 14662 8180 14714
rect 8180 14662 8210 14714
rect 8234 14662 8244 14714
rect 8244 14662 8290 14714
rect 7994 14660 8050 14662
rect 8074 14660 8130 14662
rect 8154 14660 8210 14662
rect 8234 14660 8290 14662
rect 7994 13626 8050 13628
rect 8074 13626 8130 13628
rect 8154 13626 8210 13628
rect 8234 13626 8290 13628
rect 7994 13574 8040 13626
rect 8040 13574 8050 13626
rect 8074 13574 8104 13626
rect 8104 13574 8116 13626
rect 8116 13574 8130 13626
rect 8154 13574 8168 13626
rect 8168 13574 8180 13626
rect 8180 13574 8210 13626
rect 8234 13574 8244 13626
rect 8244 13574 8290 13626
rect 7994 13572 8050 13574
rect 8074 13572 8130 13574
rect 8154 13572 8210 13574
rect 8234 13572 8290 13574
rect 9034 16496 9090 16552
rect 9218 16652 9274 16688
rect 9218 16632 9220 16652
rect 9220 16632 9272 16652
rect 9272 16632 9274 16652
rect 8574 14184 8630 14240
rect 7930 13132 7932 13152
rect 7932 13132 7984 13152
rect 7984 13132 7986 13152
rect 7930 13096 7986 13132
rect 7838 12960 7894 13016
rect 7994 12538 8050 12540
rect 8074 12538 8130 12540
rect 8154 12538 8210 12540
rect 8234 12538 8290 12540
rect 7994 12486 8040 12538
rect 8040 12486 8050 12538
rect 8074 12486 8104 12538
rect 8104 12486 8116 12538
rect 8116 12486 8130 12538
rect 8154 12486 8168 12538
rect 8168 12486 8180 12538
rect 8180 12486 8210 12538
rect 8234 12486 8244 12538
rect 8244 12486 8290 12538
rect 7994 12484 8050 12486
rect 8074 12484 8130 12486
rect 8154 12484 8210 12486
rect 8234 12484 8290 12486
rect 8482 11872 8538 11928
rect 7994 11450 8050 11452
rect 8074 11450 8130 11452
rect 8154 11450 8210 11452
rect 8234 11450 8290 11452
rect 7994 11398 8040 11450
rect 8040 11398 8050 11450
rect 8074 11398 8104 11450
rect 8104 11398 8116 11450
rect 8116 11398 8130 11450
rect 8154 11398 8168 11450
rect 8168 11398 8180 11450
rect 8180 11398 8210 11450
rect 8234 11398 8244 11450
rect 8244 11398 8290 11450
rect 7994 11396 8050 11398
rect 8074 11396 8130 11398
rect 8154 11396 8210 11398
rect 8234 11396 8290 11398
rect 8666 11328 8722 11384
rect 7746 9696 7802 9752
rect 7994 10362 8050 10364
rect 8074 10362 8130 10364
rect 8154 10362 8210 10364
rect 8234 10362 8290 10364
rect 7994 10310 8040 10362
rect 8040 10310 8050 10362
rect 8074 10310 8104 10362
rect 8104 10310 8116 10362
rect 8116 10310 8130 10362
rect 8154 10310 8168 10362
rect 8168 10310 8180 10362
rect 8180 10310 8210 10362
rect 8234 10310 8244 10362
rect 8244 10310 8290 10362
rect 7994 10308 8050 10310
rect 8074 10308 8130 10310
rect 8154 10308 8210 10310
rect 8234 10308 8290 10310
rect 8482 10920 8538 10976
rect 8942 13640 8998 13696
rect 8850 12588 8852 12608
rect 8852 12588 8904 12608
rect 8904 12588 8906 12608
rect 8850 12552 8906 12588
rect 9126 14320 9182 14376
rect 9586 17448 9642 17504
rect 9494 16088 9550 16144
rect 10874 20848 10930 20904
rect 10414 18672 10470 18728
rect 9678 14048 9734 14104
rect 10138 15136 10194 15192
rect 10414 16224 10470 16280
rect 10414 15000 10470 15056
rect 9678 13132 9680 13152
rect 9680 13132 9732 13152
rect 9732 13132 9734 13152
rect 9678 13096 9734 13132
rect 9494 12688 9550 12744
rect 8758 11056 8814 11112
rect 8574 10376 8630 10432
rect 7994 9274 8050 9276
rect 8074 9274 8130 9276
rect 8154 9274 8210 9276
rect 8234 9274 8290 9276
rect 7994 9222 8040 9274
rect 8040 9222 8050 9274
rect 8074 9222 8104 9274
rect 8104 9222 8116 9274
rect 8116 9222 8130 9274
rect 8154 9222 8168 9274
rect 8168 9222 8180 9274
rect 8180 9222 8210 9274
rect 8234 9222 8244 9274
rect 8244 9222 8290 9274
rect 7994 9220 8050 9222
rect 8074 9220 8130 9222
rect 8154 9220 8210 9222
rect 8234 9220 8290 9222
rect 7562 8336 7618 8392
rect 9862 12552 9918 12608
rect 9770 12280 9826 12336
rect 9034 11092 9036 11112
rect 9036 11092 9088 11112
rect 9088 11092 9090 11112
rect 9034 11056 9090 11092
rect 9862 11464 9918 11520
rect 9218 10412 9220 10432
rect 9220 10412 9272 10432
rect 9272 10412 9274 10432
rect 9218 10376 9274 10412
rect 9954 11056 10010 11112
rect 9586 10784 9642 10840
rect 10322 13640 10378 13696
rect 12530 21800 12586 21856
rect 11789 21786 11845 21788
rect 11869 21786 11925 21788
rect 11949 21786 12005 21788
rect 12029 21786 12085 21788
rect 11789 21734 11835 21786
rect 11835 21734 11845 21786
rect 11869 21734 11899 21786
rect 11899 21734 11911 21786
rect 11911 21734 11925 21786
rect 11949 21734 11963 21786
rect 11963 21734 11975 21786
rect 11975 21734 12005 21786
rect 12029 21734 12039 21786
rect 12039 21734 12085 21786
rect 11789 21732 11845 21734
rect 11869 21732 11925 21734
rect 11949 21732 12005 21734
rect 12029 21732 12085 21734
rect 11426 20440 11482 20496
rect 11242 19760 11298 19816
rect 10966 18164 10968 18184
rect 10968 18164 11020 18184
rect 11020 18164 11022 18184
rect 10966 18128 11022 18164
rect 10966 17992 11022 18048
rect 11058 16632 11114 16688
rect 10782 15816 10838 15872
rect 10230 13504 10286 13560
rect 10322 12960 10378 13016
rect 10782 13096 10838 13152
rect 9218 10104 9274 10160
rect 8666 8608 8722 8664
rect 7470 6432 7526 6488
rect 7654 6196 7656 6216
rect 7656 6196 7708 6216
rect 7708 6196 7710 6216
rect 7654 6160 7710 6196
rect 7562 5616 7618 5672
rect 7286 3188 7342 3224
rect 7286 3168 7288 3188
rect 7288 3168 7340 3188
rect 7340 3168 7342 3188
rect 7994 8186 8050 8188
rect 8074 8186 8130 8188
rect 8154 8186 8210 8188
rect 8234 8186 8290 8188
rect 7994 8134 8040 8186
rect 8040 8134 8050 8186
rect 8074 8134 8104 8186
rect 8104 8134 8116 8186
rect 8116 8134 8130 8186
rect 8154 8134 8168 8186
rect 8168 8134 8180 8186
rect 8180 8134 8210 8186
rect 8234 8134 8244 8186
rect 8244 8134 8290 8186
rect 7994 8132 8050 8134
rect 8074 8132 8130 8134
rect 8154 8132 8210 8134
rect 8234 8132 8290 8134
rect 7994 7098 8050 7100
rect 8074 7098 8130 7100
rect 8154 7098 8210 7100
rect 8234 7098 8290 7100
rect 7994 7046 8040 7098
rect 8040 7046 8050 7098
rect 8074 7046 8104 7098
rect 8104 7046 8116 7098
rect 8116 7046 8130 7098
rect 8154 7046 8168 7098
rect 8168 7046 8180 7098
rect 8180 7046 8210 7098
rect 8234 7046 8244 7098
rect 8244 7046 8290 7098
rect 7994 7044 8050 7046
rect 8074 7044 8130 7046
rect 8154 7044 8210 7046
rect 8234 7044 8290 7046
rect 7994 6010 8050 6012
rect 8074 6010 8130 6012
rect 8154 6010 8210 6012
rect 8234 6010 8290 6012
rect 7994 5958 8040 6010
rect 8040 5958 8050 6010
rect 8074 5958 8104 6010
rect 8104 5958 8116 6010
rect 8116 5958 8130 6010
rect 8154 5958 8168 6010
rect 8168 5958 8180 6010
rect 8180 5958 8210 6010
rect 8234 5958 8244 6010
rect 8244 5958 8290 6010
rect 7994 5956 8050 5958
rect 8074 5956 8130 5958
rect 8154 5956 8210 5958
rect 8234 5956 8290 5958
rect 7994 4922 8050 4924
rect 8074 4922 8130 4924
rect 8154 4922 8210 4924
rect 8234 4922 8290 4924
rect 7994 4870 8040 4922
rect 8040 4870 8050 4922
rect 8074 4870 8104 4922
rect 8104 4870 8116 4922
rect 8116 4870 8130 4922
rect 8154 4870 8168 4922
rect 8168 4870 8180 4922
rect 8180 4870 8210 4922
rect 8234 4870 8244 4922
rect 8244 4870 8290 4922
rect 7994 4868 8050 4870
rect 8074 4868 8130 4870
rect 8154 4868 8210 4870
rect 8234 4868 8290 4870
rect 7994 3834 8050 3836
rect 8074 3834 8130 3836
rect 8154 3834 8210 3836
rect 8234 3834 8290 3836
rect 7994 3782 8040 3834
rect 8040 3782 8050 3834
rect 8074 3782 8104 3834
rect 8104 3782 8116 3834
rect 8116 3782 8130 3834
rect 8154 3782 8168 3834
rect 8168 3782 8180 3834
rect 8180 3782 8210 3834
rect 8234 3782 8244 3834
rect 8244 3782 8290 3834
rect 7994 3780 8050 3782
rect 8074 3780 8130 3782
rect 8154 3780 8210 3782
rect 8234 3780 8290 3782
rect 7994 2746 8050 2748
rect 8074 2746 8130 2748
rect 8154 2746 8210 2748
rect 8234 2746 8290 2748
rect 7994 2694 8040 2746
rect 8040 2694 8050 2746
rect 8074 2694 8104 2746
rect 8104 2694 8116 2746
rect 8116 2694 8130 2746
rect 8154 2694 8168 2746
rect 8168 2694 8180 2746
rect 8180 2694 8210 2746
rect 8234 2694 8244 2746
rect 8244 2694 8290 2746
rect 7994 2692 8050 2694
rect 8074 2692 8130 2694
rect 8154 2692 8210 2694
rect 8234 2692 8290 2694
rect 7838 2352 7894 2408
rect 8390 1672 8446 1728
rect 7994 1658 8050 1660
rect 8074 1658 8130 1660
rect 8154 1658 8210 1660
rect 8234 1658 8290 1660
rect 7994 1606 8040 1658
rect 8040 1606 8050 1658
rect 8074 1606 8104 1658
rect 8104 1606 8116 1658
rect 8116 1606 8130 1658
rect 8154 1606 8168 1658
rect 8168 1606 8180 1658
rect 8180 1606 8210 1658
rect 8234 1606 8244 1658
rect 8244 1606 8290 1658
rect 7994 1604 8050 1606
rect 8074 1604 8130 1606
rect 8154 1604 8210 1606
rect 8234 1604 8290 1606
rect 6090 1128 6146 1184
rect 6182 584 6238 640
rect 9126 7828 9128 7848
rect 9128 7828 9180 7848
rect 9180 7828 9182 7848
rect 9126 7792 9182 7828
rect 9126 7112 9182 7168
rect 9126 6704 9182 6760
rect 10414 9016 10470 9072
rect 10598 9036 10654 9072
rect 10598 9016 10600 9036
rect 10600 9016 10652 9036
rect 10652 9016 10654 9036
rect 10506 7520 10562 7576
rect 9954 7112 10010 7168
rect 9218 3032 9274 3088
rect 8666 1536 8722 1592
rect 11334 14048 11390 14104
rect 11242 12960 11298 13016
rect 11058 12144 11114 12200
rect 14002 21528 14058 21584
rect 11789 20698 11845 20700
rect 11869 20698 11925 20700
rect 11949 20698 12005 20700
rect 12029 20698 12085 20700
rect 11789 20646 11835 20698
rect 11835 20646 11845 20698
rect 11869 20646 11899 20698
rect 11899 20646 11911 20698
rect 11911 20646 11925 20698
rect 11949 20646 11963 20698
rect 11963 20646 11975 20698
rect 11975 20646 12005 20698
rect 12029 20646 12039 20698
rect 12039 20646 12085 20698
rect 11789 20644 11845 20646
rect 11869 20644 11925 20646
rect 11949 20644 12005 20646
rect 12029 20644 12085 20646
rect 11789 19610 11845 19612
rect 11869 19610 11925 19612
rect 11949 19610 12005 19612
rect 12029 19610 12085 19612
rect 11789 19558 11835 19610
rect 11835 19558 11845 19610
rect 11869 19558 11899 19610
rect 11899 19558 11911 19610
rect 11911 19558 11925 19610
rect 11949 19558 11963 19610
rect 11963 19558 11975 19610
rect 11975 19558 12005 19610
rect 12029 19558 12039 19610
rect 12039 19558 12085 19610
rect 11789 19556 11845 19558
rect 11869 19556 11925 19558
rect 11949 19556 12005 19558
rect 12029 19556 12085 19558
rect 11794 18692 11850 18728
rect 11794 18672 11796 18692
rect 11796 18672 11848 18692
rect 11848 18672 11850 18692
rect 11789 18522 11845 18524
rect 11869 18522 11925 18524
rect 11949 18522 12005 18524
rect 12029 18522 12085 18524
rect 11789 18470 11835 18522
rect 11835 18470 11845 18522
rect 11869 18470 11899 18522
rect 11899 18470 11911 18522
rect 11911 18470 11925 18522
rect 11949 18470 11963 18522
rect 11963 18470 11975 18522
rect 11975 18470 12005 18522
rect 12029 18470 12039 18522
rect 12039 18470 12085 18522
rect 11789 18468 11845 18470
rect 11869 18468 11925 18470
rect 11949 18468 12005 18470
rect 12029 18468 12085 18470
rect 12346 18672 12402 18728
rect 12254 17876 12310 17912
rect 12254 17856 12256 17876
rect 12256 17856 12308 17876
rect 12308 17856 12310 17876
rect 11789 17434 11845 17436
rect 11869 17434 11925 17436
rect 11949 17434 12005 17436
rect 12029 17434 12085 17436
rect 11789 17382 11835 17434
rect 11835 17382 11845 17434
rect 11869 17382 11899 17434
rect 11899 17382 11911 17434
rect 11911 17382 11925 17434
rect 11949 17382 11963 17434
rect 11963 17382 11975 17434
rect 11975 17382 12005 17434
rect 12029 17382 12039 17434
rect 12039 17382 12085 17434
rect 11789 17380 11845 17382
rect 11869 17380 11925 17382
rect 11949 17380 12005 17382
rect 12029 17380 12085 17382
rect 11702 16768 11758 16824
rect 11886 16788 11942 16824
rect 11886 16768 11888 16788
rect 11888 16768 11940 16788
rect 11940 16768 11942 16788
rect 11794 16632 11850 16688
rect 11789 16346 11845 16348
rect 11869 16346 11925 16348
rect 11949 16346 12005 16348
rect 12029 16346 12085 16348
rect 11789 16294 11835 16346
rect 11835 16294 11845 16346
rect 11869 16294 11899 16346
rect 11899 16294 11911 16346
rect 11911 16294 11925 16346
rect 11949 16294 11963 16346
rect 11963 16294 11975 16346
rect 11975 16294 12005 16346
rect 12029 16294 12039 16346
rect 12039 16294 12085 16346
rect 11789 16292 11845 16294
rect 11869 16292 11925 16294
rect 11949 16292 12005 16294
rect 12029 16292 12085 16294
rect 11702 16088 11758 16144
rect 11789 15258 11845 15260
rect 11869 15258 11925 15260
rect 11949 15258 12005 15260
rect 12029 15258 12085 15260
rect 11789 15206 11835 15258
rect 11835 15206 11845 15258
rect 11869 15206 11899 15258
rect 11899 15206 11911 15258
rect 11911 15206 11925 15258
rect 11949 15206 11963 15258
rect 11963 15206 11975 15258
rect 11975 15206 12005 15258
rect 12029 15206 12039 15258
rect 12039 15206 12085 15258
rect 11789 15204 11845 15206
rect 11869 15204 11925 15206
rect 11949 15204 12005 15206
rect 12029 15204 12085 15206
rect 11794 14356 11796 14376
rect 11796 14356 11848 14376
rect 11848 14356 11850 14376
rect 11794 14320 11850 14356
rect 11789 14170 11845 14172
rect 11869 14170 11925 14172
rect 11949 14170 12005 14172
rect 12029 14170 12085 14172
rect 11789 14118 11835 14170
rect 11835 14118 11845 14170
rect 11869 14118 11899 14170
rect 11899 14118 11911 14170
rect 11911 14118 11925 14170
rect 11949 14118 11963 14170
rect 11963 14118 11975 14170
rect 11975 14118 12005 14170
rect 12029 14118 12039 14170
rect 12039 14118 12085 14170
rect 11789 14116 11845 14118
rect 11869 14116 11925 14118
rect 11949 14116 12005 14118
rect 12029 14116 12085 14118
rect 11058 11328 11114 11384
rect 11518 12300 11574 12336
rect 11518 12280 11520 12300
rect 11520 12280 11572 12300
rect 11572 12280 11574 12300
rect 13726 20576 13782 20632
rect 12530 14048 12586 14104
rect 11789 13082 11845 13084
rect 11869 13082 11925 13084
rect 11949 13082 12005 13084
rect 12029 13082 12085 13084
rect 11789 13030 11835 13082
rect 11835 13030 11845 13082
rect 11869 13030 11899 13082
rect 11899 13030 11911 13082
rect 11911 13030 11925 13082
rect 11949 13030 11963 13082
rect 11963 13030 11975 13082
rect 11975 13030 12005 13082
rect 12029 13030 12039 13082
rect 12039 13030 12085 13082
rect 11789 13028 11845 13030
rect 11869 13028 11925 13030
rect 11949 13028 12005 13030
rect 12029 13028 12085 13030
rect 12346 12960 12402 13016
rect 11610 12008 11666 12064
rect 11518 11736 11574 11792
rect 11789 11994 11845 11996
rect 11869 11994 11925 11996
rect 11949 11994 12005 11996
rect 12029 11994 12085 11996
rect 11789 11942 11835 11994
rect 11835 11942 11845 11994
rect 11869 11942 11899 11994
rect 11899 11942 11911 11994
rect 11911 11942 11925 11994
rect 11949 11942 11963 11994
rect 11963 11942 11975 11994
rect 11975 11942 12005 11994
rect 12029 11942 12039 11994
rect 12039 11942 12085 11994
rect 11789 11940 11845 11942
rect 11869 11940 11925 11942
rect 11949 11940 12005 11942
rect 12029 11940 12085 11942
rect 12162 11872 12218 11928
rect 12530 12280 12586 12336
rect 12070 11464 12126 11520
rect 12346 11600 12402 11656
rect 11150 8900 11206 8936
rect 11150 8880 11152 8900
rect 11152 8880 11204 8900
rect 11204 8880 11206 8900
rect 11058 7248 11114 7304
rect 11789 10906 11845 10908
rect 11869 10906 11925 10908
rect 11949 10906 12005 10908
rect 12029 10906 12085 10908
rect 11789 10854 11835 10906
rect 11835 10854 11845 10906
rect 11869 10854 11899 10906
rect 11899 10854 11911 10906
rect 11911 10854 11925 10906
rect 11949 10854 11963 10906
rect 11963 10854 11975 10906
rect 11975 10854 12005 10906
rect 12029 10854 12039 10906
rect 12039 10854 12085 10906
rect 11789 10852 11845 10854
rect 11869 10852 11925 10854
rect 11949 10852 12005 10854
rect 12029 10852 12085 10854
rect 11789 9818 11845 9820
rect 11869 9818 11925 9820
rect 11949 9818 12005 9820
rect 12029 9818 12085 9820
rect 11789 9766 11835 9818
rect 11835 9766 11845 9818
rect 11869 9766 11899 9818
rect 11899 9766 11911 9818
rect 11911 9766 11925 9818
rect 11949 9766 11963 9818
rect 11963 9766 11975 9818
rect 11975 9766 12005 9818
rect 12029 9766 12039 9818
rect 12039 9766 12085 9818
rect 11789 9764 11845 9766
rect 11869 9764 11925 9766
rect 11949 9764 12005 9766
rect 12029 9764 12085 9766
rect 10690 5480 10746 5536
rect 11789 8730 11845 8732
rect 11869 8730 11925 8732
rect 11949 8730 12005 8732
rect 12029 8730 12085 8732
rect 11789 8678 11835 8730
rect 11835 8678 11845 8730
rect 11869 8678 11899 8730
rect 11899 8678 11911 8730
rect 11911 8678 11925 8730
rect 11949 8678 11963 8730
rect 11963 8678 11975 8730
rect 11975 8678 12005 8730
rect 12029 8678 12039 8730
rect 12039 8678 12085 8730
rect 11789 8676 11845 8678
rect 11869 8676 11925 8678
rect 11949 8676 12005 8678
rect 12029 8676 12085 8678
rect 11518 8200 11574 8256
rect 11426 6296 11482 6352
rect 11334 5616 11390 5672
rect 9586 1128 9642 1184
rect 7994 570 8050 572
rect 8074 570 8130 572
rect 8154 570 8210 572
rect 8234 570 8290 572
rect 7994 518 8040 570
rect 8040 518 8050 570
rect 8074 518 8104 570
rect 8104 518 8116 570
rect 8116 518 8130 570
rect 8154 518 8168 570
rect 8168 518 8180 570
rect 8180 518 8210 570
rect 8234 518 8244 570
rect 8244 518 8290 570
rect 7994 516 8050 518
rect 8074 516 8130 518
rect 8154 516 8210 518
rect 8234 516 8290 518
rect 11150 3848 11206 3904
rect 10598 2488 10654 2544
rect 11150 3168 11206 3224
rect 11789 7642 11845 7644
rect 11869 7642 11925 7644
rect 11949 7642 12005 7644
rect 12029 7642 12085 7644
rect 11789 7590 11835 7642
rect 11835 7590 11845 7642
rect 11869 7590 11899 7642
rect 11899 7590 11911 7642
rect 11911 7590 11925 7642
rect 11949 7590 11963 7642
rect 11963 7590 11975 7642
rect 11975 7590 12005 7642
rect 12029 7590 12039 7642
rect 12039 7590 12085 7642
rect 11789 7588 11845 7590
rect 11869 7588 11925 7590
rect 11949 7588 12005 7590
rect 12029 7588 12085 7590
rect 12990 16904 13046 16960
rect 13358 19216 13414 19272
rect 13266 17212 13268 17232
rect 13268 17212 13320 17232
rect 13320 17212 13322 17232
rect 13266 17176 13322 17212
rect 12990 13504 13046 13560
rect 13358 16396 13360 16416
rect 13360 16396 13412 16416
rect 13412 16396 13414 16416
rect 13358 16360 13414 16396
rect 14186 21392 14242 21448
rect 15584 21242 15640 21244
rect 15664 21242 15720 21244
rect 15744 21242 15800 21244
rect 15824 21242 15880 21244
rect 15584 21190 15630 21242
rect 15630 21190 15640 21242
rect 15664 21190 15694 21242
rect 15694 21190 15706 21242
rect 15706 21190 15720 21242
rect 15744 21190 15758 21242
rect 15758 21190 15770 21242
rect 15770 21190 15800 21242
rect 15824 21190 15834 21242
rect 15834 21190 15880 21242
rect 15584 21188 15640 21190
rect 15664 21188 15720 21190
rect 15744 21188 15800 21190
rect 15824 21188 15880 21190
rect 15106 20984 15162 21040
rect 14462 19352 14518 19408
rect 15584 20154 15640 20156
rect 15664 20154 15720 20156
rect 15744 20154 15800 20156
rect 15824 20154 15880 20156
rect 15584 20102 15630 20154
rect 15630 20102 15640 20154
rect 15664 20102 15694 20154
rect 15694 20102 15706 20154
rect 15706 20102 15720 20154
rect 15744 20102 15758 20154
rect 15758 20102 15770 20154
rect 15770 20102 15800 20154
rect 15824 20102 15834 20154
rect 15834 20102 15880 20154
rect 15584 20100 15640 20102
rect 15664 20100 15720 20102
rect 15744 20100 15800 20102
rect 15824 20100 15880 20102
rect 13634 17040 13690 17096
rect 14094 17076 14096 17096
rect 14096 17076 14148 17096
rect 14148 17076 14150 17096
rect 13634 16224 13690 16280
rect 13542 15680 13598 15736
rect 13450 15544 13506 15600
rect 14094 17040 14150 17076
rect 14554 18828 14610 18864
rect 14554 18808 14556 18828
rect 14556 18808 14608 18828
rect 14608 18808 14610 18828
rect 15106 19216 15162 19272
rect 15584 19066 15640 19068
rect 15664 19066 15720 19068
rect 15744 19066 15800 19068
rect 15824 19066 15880 19068
rect 15584 19014 15630 19066
rect 15630 19014 15640 19066
rect 15664 19014 15694 19066
rect 15694 19014 15706 19066
rect 15706 19014 15720 19066
rect 15744 19014 15758 19066
rect 15758 19014 15770 19066
rect 15770 19014 15800 19066
rect 15824 19014 15834 19066
rect 15834 19014 15880 19066
rect 15584 19012 15640 19014
rect 15664 19012 15720 19014
rect 15744 19012 15800 19014
rect 15824 19012 15880 19014
rect 14554 16904 14610 16960
rect 15106 16768 15162 16824
rect 13910 15816 13966 15872
rect 14922 16496 14978 16552
rect 15584 17978 15640 17980
rect 15664 17978 15720 17980
rect 15744 17978 15800 17980
rect 15824 17978 15880 17980
rect 15584 17926 15630 17978
rect 15630 17926 15640 17978
rect 15664 17926 15694 17978
rect 15694 17926 15706 17978
rect 15706 17926 15720 17978
rect 15744 17926 15758 17978
rect 15758 17926 15770 17978
rect 15770 17926 15800 17978
rect 15824 17926 15834 17978
rect 15834 17926 15880 17978
rect 15584 17924 15640 17926
rect 15664 17924 15720 17926
rect 15744 17924 15800 17926
rect 15824 17924 15880 17926
rect 13450 14864 13506 14920
rect 14278 14320 14334 14376
rect 14094 14184 14150 14240
rect 14278 13912 14334 13968
rect 13358 13640 13414 13696
rect 13726 13640 13782 13696
rect 13174 11872 13230 11928
rect 13174 11500 13176 11520
rect 13176 11500 13228 11520
rect 13228 11500 13230 11520
rect 13174 11464 13230 11500
rect 12990 10240 13046 10296
rect 14462 14356 14464 14376
rect 14464 14356 14516 14376
rect 14516 14356 14518 14376
rect 14462 14320 14518 14356
rect 14554 12688 14610 12744
rect 14278 12280 14334 12336
rect 13910 11328 13966 11384
rect 12438 9016 12494 9072
rect 11789 6554 11845 6556
rect 11869 6554 11925 6556
rect 11949 6554 12005 6556
rect 12029 6554 12085 6556
rect 11789 6502 11835 6554
rect 11835 6502 11845 6554
rect 11869 6502 11899 6554
rect 11899 6502 11911 6554
rect 11911 6502 11925 6554
rect 11949 6502 11963 6554
rect 11963 6502 11975 6554
rect 11975 6502 12005 6554
rect 12029 6502 12039 6554
rect 12039 6502 12085 6554
rect 11789 6500 11845 6502
rect 11869 6500 11925 6502
rect 11949 6500 12005 6502
rect 12029 6500 12085 6502
rect 12806 8880 12862 8936
rect 11789 5466 11845 5468
rect 11869 5466 11925 5468
rect 11949 5466 12005 5468
rect 12029 5466 12085 5468
rect 11789 5414 11835 5466
rect 11835 5414 11845 5466
rect 11869 5414 11899 5466
rect 11899 5414 11911 5466
rect 11911 5414 11925 5466
rect 11949 5414 11963 5466
rect 11963 5414 11975 5466
rect 11975 5414 12005 5466
rect 12029 5414 12039 5466
rect 12039 5414 12085 5466
rect 11789 5412 11845 5414
rect 11869 5412 11925 5414
rect 11949 5412 12005 5414
rect 12029 5412 12085 5414
rect 12254 5752 12310 5808
rect 11789 4378 11845 4380
rect 11869 4378 11925 4380
rect 11949 4378 12005 4380
rect 12029 4378 12085 4380
rect 11789 4326 11835 4378
rect 11835 4326 11845 4378
rect 11869 4326 11899 4378
rect 11899 4326 11911 4378
rect 11911 4326 11925 4378
rect 11949 4326 11963 4378
rect 11963 4326 11975 4378
rect 11975 4326 12005 4378
rect 12029 4326 12039 4378
rect 12039 4326 12085 4378
rect 11789 4324 11845 4326
rect 11869 4324 11925 4326
rect 11949 4324 12005 4326
rect 12029 4324 12085 4326
rect 14094 11464 14150 11520
rect 14002 9968 14058 10024
rect 15106 14864 15162 14920
rect 15198 13776 15254 13832
rect 12438 5752 12494 5808
rect 13450 5344 13506 5400
rect 13266 5208 13322 5264
rect 12254 3848 12310 3904
rect 11789 3290 11845 3292
rect 11869 3290 11925 3292
rect 11949 3290 12005 3292
rect 12029 3290 12085 3292
rect 11789 3238 11835 3290
rect 11835 3238 11845 3290
rect 11869 3238 11899 3290
rect 11899 3238 11911 3290
rect 11911 3238 11925 3290
rect 11949 3238 11963 3290
rect 11963 3238 11975 3290
rect 11975 3238 12005 3290
rect 12029 3238 12039 3290
rect 12039 3238 12085 3290
rect 11789 3236 11845 3238
rect 11869 3236 11925 3238
rect 11949 3236 12005 3238
rect 12029 3236 12085 3238
rect 12254 3032 12310 3088
rect 11058 1400 11114 1456
rect 11789 2202 11845 2204
rect 11869 2202 11925 2204
rect 11949 2202 12005 2204
rect 12029 2202 12085 2204
rect 11789 2150 11835 2202
rect 11835 2150 11845 2202
rect 11869 2150 11899 2202
rect 11899 2150 11911 2202
rect 11911 2150 11925 2202
rect 11949 2150 11963 2202
rect 11963 2150 11975 2202
rect 11975 2150 12005 2202
rect 12029 2150 12039 2202
rect 12039 2150 12085 2202
rect 11789 2148 11845 2150
rect 11869 2148 11925 2150
rect 11949 2148 12005 2150
rect 12029 2148 12085 2150
rect 11426 1672 11482 1728
rect 11426 1400 11482 1456
rect 11610 620 11612 640
rect 11612 620 11664 640
rect 11664 620 11666 640
rect 11610 584 11666 620
rect 11789 1114 11845 1116
rect 11869 1114 11925 1116
rect 11949 1114 12005 1116
rect 12029 1114 12085 1116
rect 11789 1062 11835 1114
rect 11835 1062 11845 1114
rect 11869 1062 11899 1114
rect 11899 1062 11911 1114
rect 11911 1062 11925 1114
rect 11949 1062 11963 1114
rect 11963 1062 11975 1114
rect 11975 1062 12005 1114
rect 12029 1062 12039 1114
rect 12039 1062 12085 1114
rect 11789 1060 11845 1062
rect 11869 1060 11925 1062
rect 11949 1060 12005 1062
rect 12029 1060 12085 1062
rect 13634 4020 13636 4040
rect 13636 4020 13688 4040
rect 13688 4020 13690 4040
rect 13634 3984 13690 4020
rect 12162 312 12218 368
rect 13818 1400 13874 1456
rect 14830 7520 14886 7576
rect 14462 3984 14518 4040
rect 14462 2488 14518 2544
rect 14462 1536 14518 1592
rect 16026 17720 16082 17776
rect 15584 16890 15640 16892
rect 15664 16890 15720 16892
rect 15744 16890 15800 16892
rect 15824 16890 15880 16892
rect 15584 16838 15630 16890
rect 15630 16838 15640 16890
rect 15664 16838 15694 16890
rect 15694 16838 15706 16890
rect 15706 16838 15720 16890
rect 15744 16838 15758 16890
rect 15758 16838 15770 16890
rect 15770 16838 15800 16890
rect 15824 16838 15834 16890
rect 15834 16838 15880 16890
rect 15584 16836 15640 16838
rect 15664 16836 15720 16838
rect 15744 16836 15800 16838
rect 15824 16836 15880 16838
rect 15934 16632 15990 16688
rect 15474 16244 15530 16280
rect 15474 16224 15476 16244
rect 15476 16224 15528 16244
rect 15528 16224 15530 16244
rect 15584 15802 15640 15804
rect 15664 15802 15720 15804
rect 15744 15802 15800 15804
rect 15824 15802 15880 15804
rect 15584 15750 15630 15802
rect 15630 15750 15640 15802
rect 15664 15750 15694 15802
rect 15694 15750 15706 15802
rect 15706 15750 15720 15802
rect 15744 15750 15758 15802
rect 15758 15750 15770 15802
rect 15770 15750 15800 15802
rect 15824 15750 15834 15802
rect 15834 15750 15880 15802
rect 15584 15748 15640 15750
rect 15664 15748 15720 15750
rect 15744 15748 15800 15750
rect 15824 15748 15880 15750
rect 15382 13640 15438 13696
rect 15584 14714 15640 14716
rect 15664 14714 15720 14716
rect 15744 14714 15800 14716
rect 15824 14714 15880 14716
rect 15584 14662 15630 14714
rect 15630 14662 15640 14714
rect 15664 14662 15694 14714
rect 15694 14662 15706 14714
rect 15706 14662 15720 14714
rect 15744 14662 15758 14714
rect 15758 14662 15770 14714
rect 15770 14662 15800 14714
rect 15824 14662 15834 14714
rect 15834 14662 15880 14714
rect 15584 14660 15640 14662
rect 15664 14660 15720 14662
rect 15744 14660 15800 14662
rect 15824 14660 15880 14662
rect 15584 13626 15640 13628
rect 15664 13626 15720 13628
rect 15744 13626 15800 13628
rect 15824 13626 15880 13628
rect 15584 13574 15630 13626
rect 15630 13574 15640 13626
rect 15664 13574 15694 13626
rect 15694 13574 15706 13626
rect 15706 13574 15720 13626
rect 15744 13574 15758 13626
rect 15758 13574 15770 13626
rect 15770 13574 15800 13626
rect 15824 13574 15834 13626
rect 15834 13574 15880 13626
rect 15584 13572 15640 13574
rect 15664 13572 15720 13574
rect 15744 13572 15800 13574
rect 15824 13572 15880 13574
rect 16670 21392 16726 21448
rect 16578 20984 16634 21040
rect 16670 19352 16726 19408
rect 16302 19216 16358 19272
rect 16486 19216 16542 19272
rect 16302 18128 16358 18184
rect 16486 17176 16542 17232
rect 16302 16768 16358 16824
rect 16302 16124 16304 16144
rect 16304 16124 16356 16144
rect 16356 16124 16358 16144
rect 16302 16088 16358 16124
rect 17130 21528 17186 21584
rect 18510 21412 18566 21448
rect 18510 21392 18512 21412
rect 18512 21392 18564 21412
rect 18564 21392 18566 21412
rect 17866 20984 17922 21040
rect 19379 21786 19435 21788
rect 19459 21786 19515 21788
rect 19539 21786 19595 21788
rect 19619 21786 19675 21788
rect 19379 21734 19425 21786
rect 19425 21734 19435 21786
rect 19459 21734 19489 21786
rect 19489 21734 19501 21786
rect 19501 21734 19515 21786
rect 19539 21734 19553 21786
rect 19553 21734 19565 21786
rect 19565 21734 19595 21786
rect 19619 21734 19629 21786
rect 19629 21734 19675 21786
rect 19379 21732 19435 21734
rect 19459 21732 19515 21734
rect 19539 21732 19595 21734
rect 19619 21732 19675 21734
rect 19379 20698 19435 20700
rect 19459 20698 19515 20700
rect 19539 20698 19595 20700
rect 19619 20698 19675 20700
rect 19379 20646 19425 20698
rect 19425 20646 19435 20698
rect 19459 20646 19489 20698
rect 19489 20646 19501 20698
rect 19501 20646 19515 20698
rect 19539 20646 19553 20698
rect 19553 20646 19565 20698
rect 19565 20646 19595 20698
rect 19619 20646 19629 20698
rect 19629 20646 19675 20698
rect 19379 20644 19435 20646
rect 19459 20644 19515 20646
rect 19539 20644 19595 20646
rect 19619 20644 19675 20646
rect 18694 20460 18750 20496
rect 18694 20440 18696 20460
rect 18696 20440 18748 20460
rect 18748 20440 18750 20460
rect 17682 19304 17738 19348
rect 17682 19292 17684 19304
rect 17684 19292 17736 19304
rect 17736 19292 17738 19304
rect 17038 17992 17094 18048
rect 16854 17040 16910 17096
rect 16394 15000 16450 15056
rect 17130 15952 17186 16008
rect 18970 17584 19026 17640
rect 16854 15428 16910 15464
rect 16854 15408 16856 15428
rect 16856 15408 16908 15428
rect 16908 15408 16910 15428
rect 16670 13912 16726 13968
rect 15584 12538 15640 12540
rect 15664 12538 15720 12540
rect 15744 12538 15800 12540
rect 15824 12538 15880 12540
rect 15584 12486 15630 12538
rect 15630 12486 15640 12538
rect 15664 12486 15694 12538
rect 15694 12486 15706 12538
rect 15706 12486 15720 12538
rect 15744 12486 15758 12538
rect 15758 12486 15770 12538
rect 15770 12486 15800 12538
rect 15824 12486 15834 12538
rect 15834 12486 15880 12538
rect 15584 12484 15640 12486
rect 15664 12484 15720 12486
rect 15744 12484 15800 12486
rect 15824 12484 15880 12486
rect 15566 11736 15622 11792
rect 15584 11450 15640 11452
rect 15664 11450 15720 11452
rect 15744 11450 15800 11452
rect 15824 11450 15880 11452
rect 15584 11398 15630 11450
rect 15630 11398 15640 11450
rect 15664 11398 15694 11450
rect 15694 11398 15706 11450
rect 15706 11398 15720 11450
rect 15744 11398 15758 11450
rect 15758 11398 15770 11450
rect 15770 11398 15800 11450
rect 15824 11398 15834 11450
rect 15834 11398 15880 11450
rect 15584 11396 15640 11398
rect 15664 11396 15720 11398
rect 15744 11396 15800 11398
rect 15824 11396 15880 11398
rect 15290 10512 15346 10568
rect 15584 10362 15640 10364
rect 15664 10362 15720 10364
rect 15744 10362 15800 10364
rect 15824 10362 15880 10364
rect 15584 10310 15630 10362
rect 15630 10310 15640 10362
rect 15664 10310 15694 10362
rect 15694 10310 15706 10362
rect 15706 10310 15720 10362
rect 15744 10310 15758 10362
rect 15758 10310 15770 10362
rect 15770 10310 15800 10362
rect 15824 10310 15834 10362
rect 15834 10310 15880 10362
rect 15584 10308 15640 10310
rect 15664 10308 15720 10310
rect 15744 10308 15800 10310
rect 15824 10308 15880 10310
rect 15584 9274 15640 9276
rect 15664 9274 15720 9276
rect 15744 9274 15800 9276
rect 15824 9274 15880 9276
rect 15584 9222 15630 9274
rect 15630 9222 15640 9274
rect 15664 9222 15694 9274
rect 15694 9222 15706 9274
rect 15706 9222 15720 9274
rect 15744 9222 15758 9274
rect 15758 9222 15770 9274
rect 15770 9222 15800 9274
rect 15824 9222 15834 9274
rect 15834 9222 15880 9274
rect 15584 9220 15640 9222
rect 15664 9220 15720 9222
rect 15744 9220 15800 9222
rect 15824 9220 15880 9222
rect 15584 8186 15640 8188
rect 15664 8186 15720 8188
rect 15744 8186 15800 8188
rect 15824 8186 15880 8188
rect 15584 8134 15630 8186
rect 15630 8134 15640 8186
rect 15664 8134 15694 8186
rect 15694 8134 15706 8186
rect 15706 8134 15720 8186
rect 15744 8134 15758 8186
rect 15758 8134 15770 8186
rect 15770 8134 15800 8186
rect 15824 8134 15834 8186
rect 15834 8134 15880 8186
rect 15584 8132 15640 8134
rect 15664 8132 15720 8134
rect 15744 8132 15800 8134
rect 15824 8132 15880 8134
rect 15658 7812 15714 7848
rect 15658 7792 15660 7812
rect 15660 7792 15712 7812
rect 15712 7792 15714 7812
rect 15584 7098 15640 7100
rect 15664 7098 15720 7100
rect 15744 7098 15800 7100
rect 15824 7098 15880 7100
rect 15584 7046 15630 7098
rect 15630 7046 15640 7098
rect 15664 7046 15694 7098
rect 15694 7046 15706 7098
rect 15706 7046 15720 7098
rect 15744 7046 15758 7098
rect 15758 7046 15770 7098
rect 15770 7046 15800 7098
rect 15824 7046 15834 7098
rect 15834 7046 15880 7098
rect 15584 7044 15640 7046
rect 15664 7044 15720 7046
rect 15744 7044 15800 7046
rect 15824 7044 15880 7046
rect 15290 5072 15346 5128
rect 15106 3052 15162 3088
rect 15106 3032 15108 3052
rect 15108 3032 15160 3052
rect 15160 3032 15162 3052
rect 11978 176 12034 232
rect 15584 6010 15640 6012
rect 15664 6010 15720 6012
rect 15744 6010 15800 6012
rect 15824 6010 15880 6012
rect 15584 5958 15630 6010
rect 15630 5958 15640 6010
rect 15664 5958 15694 6010
rect 15694 5958 15706 6010
rect 15706 5958 15720 6010
rect 15744 5958 15758 6010
rect 15758 5958 15770 6010
rect 15770 5958 15800 6010
rect 15824 5958 15834 6010
rect 15834 5958 15880 6010
rect 15584 5956 15640 5958
rect 15664 5956 15720 5958
rect 15744 5956 15800 5958
rect 15824 5956 15880 5958
rect 16578 13268 16580 13288
rect 16580 13268 16632 13288
rect 16632 13268 16634 13288
rect 16578 13232 16634 13268
rect 16302 12688 16358 12744
rect 16762 12960 16818 13016
rect 18326 15000 18382 15056
rect 19379 19610 19435 19612
rect 19459 19610 19515 19612
rect 19539 19610 19595 19612
rect 19619 19610 19675 19612
rect 19379 19558 19425 19610
rect 19425 19558 19435 19610
rect 19459 19558 19489 19610
rect 19489 19558 19501 19610
rect 19501 19558 19515 19610
rect 19539 19558 19553 19610
rect 19553 19558 19565 19610
rect 19565 19558 19595 19610
rect 19619 19558 19629 19610
rect 19629 19558 19675 19610
rect 19379 19556 19435 19558
rect 19459 19556 19515 19558
rect 19539 19556 19595 19558
rect 19619 19556 19675 19558
rect 20994 19932 20996 19952
rect 20996 19932 21048 19952
rect 21048 19932 21050 19952
rect 20994 19896 21050 19932
rect 19379 18522 19435 18524
rect 19459 18522 19515 18524
rect 19539 18522 19595 18524
rect 19619 18522 19675 18524
rect 19379 18470 19425 18522
rect 19425 18470 19435 18522
rect 19459 18470 19489 18522
rect 19489 18470 19501 18522
rect 19501 18470 19515 18522
rect 19539 18470 19553 18522
rect 19553 18470 19565 18522
rect 19565 18470 19595 18522
rect 19619 18470 19629 18522
rect 19629 18470 19675 18522
rect 19379 18468 19435 18470
rect 19459 18468 19515 18470
rect 19539 18468 19595 18470
rect 19619 18468 19675 18470
rect 19246 17992 19302 18048
rect 19982 17448 20038 17504
rect 19379 17434 19435 17436
rect 19459 17434 19515 17436
rect 19539 17434 19595 17436
rect 19619 17434 19675 17436
rect 19379 17382 19425 17434
rect 19425 17382 19435 17434
rect 19459 17382 19489 17434
rect 19489 17382 19501 17434
rect 19501 17382 19515 17434
rect 19539 17382 19553 17434
rect 19553 17382 19565 17434
rect 19565 17382 19595 17434
rect 19619 17382 19629 17434
rect 19629 17382 19675 17434
rect 19379 17380 19435 17382
rect 19459 17380 19515 17382
rect 19539 17380 19595 17382
rect 19619 17380 19675 17382
rect 19338 16496 19394 16552
rect 19379 16346 19435 16348
rect 19459 16346 19515 16348
rect 19539 16346 19595 16348
rect 19619 16346 19675 16348
rect 19379 16294 19425 16346
rect 19425 16294 19435 16346
rect 19459 16294 19489 16346
rect 19489 16294 19501 16346
rect 19501 16294 19515 16346
rect 19539 16294 19553 16346
rect 19553 16294 19565 16346
rect 19565 16294 19595 16346
rect 19619 16294 19629 16346
rect 19629 16294 19675 16346
rect 19379 16292 19435 16294
rect 19459 16292 19515 16294
rect 19539 16292 19595 16294
rect 19619 16292 19675 16294
rect 19062 14864 19118 14920
rect 19062 14728 19118 14784
rect 18970 14340 19026 14376
rect 18970 14320 18972 14340
rect 18972 14320 19024 14340
rect 19024 14320 19026 14340
rect 18970 14048 19026 14104
rect 19614 15680 19670 15736
rect 19706 15564 19762 15600
rect 19706 15544 19708 15564
rect 19708 15544 19760 15564
rect 19760 15544 19762 15564
rect 19379 15258 19435 15260
rect 19459 15258 19515 15260
rect 19539 15258 19595 15260
rect 19619 15258 19675 15260
rect 19379 15206 19425 15258
rect 19425 15206 19435 15258
rect 19459 15206 19489 15258
rect 19489 15206 19501 15258
rect 19501 15206 19515 15258
rect 19539 15206 19553 15258
rect 19553 15206 19565 15258
rect 19565 15206 19595 15258
rect 19619 15206 19629 15258
rect 19629 15206 19675 15258
rect 19379 15204 19435 15206
rect 19459 15204 19515 15206
rect 19539 15204 19595 15206
rect 19619 15204 19675 15206
rect 19379 14170 19435 14172
rect 19459 14170 19515 14172
rect 19539 14170 19595 14172
rect 19619 14170 19675 14172
rect 19379 14118 19425 14170
rect 19425 14118 19435 14170
rect 19459 14118 19489 14170
rect 19489 14118 19501 14170
rect 19501 14118 19515 14170
rect 19539 14118 19553 14170
rect 19553 14118 19565 14170
rect 19565 14118 19595 14170
rect 19619 14118 19629 14170
rect 19629 14118 19675 14170
rect 19379 14116 19435 14118
rect 19459 14116 19515 14118
rect 19539 14116 19595 14118
rect 19619 14116 19675 14118
rect 16578 10668 16634 10704
rect 16578 10648 16580 10668
rect 16580 10648 16632 10668
rect 16632 10648 16634 10668
rect 16486 10104 16542 10160
rect 16578 9580 16634 9616
rect 16578 9560 16580 9580
rect 16580 9560 16632 9580
rect 16632 9560 16634 9580
rect 16394 7928 16450 7984
rect 16302 7384 16358 7440
rect 16210 6704 16266 6760
rect 15584 4922 15640 4924
rect 15664 4922 15720 4924
rect 15744 4922 15800 4924
rect 15824 4922 15880 4924
rect 15584 4870 15630 4922
rect 15630 4870 15640 4922
rect 15664 4870 15694 4922
rect 15694 4870 15706 4922
rect 15706 4870 15720 4922
rect 15744 4870 15758 4922
rect 15758 4870 15770 4922
rect 15770 4870 15800 4922
rect 15824 4870 15834 4922
rect 15834 4870 15880 4922
rect 15584 4868 15640 4870
rect 15664 4868 15720 4870
rect 15744 4868 15800 4870
rect 15824 4868 15880 4870
rect 15584 3834 15640 3836
rect 15664 3834 15720 3836
rect 15744 3834 15800 3836
rect 15824 3834 15880 3836
rect 15584 3782 15630 3834
rect 15630 3782 15640 3834
rect 15664 3782 15694 3834
rect 15694 3782 15706 3834
rect 15706 3782 15720 3834
rect 15744 3782 15758 3834
rect 15758 3782 15770 3834
rect 15770 3782 15800 3834
rect 15824 3782 15834 3834
rect 15834 3782 15880 3834
rect 15584 3780 15640 3782
rect 15664 3780 15720 3782
rect 15744 3780 15800 3782
rect 15824 3780 15880 3782
rect 15584 2746 15640 2748
rect 15664 2746 15720 2748
rect 15744 2746 15800 2748
rect 15824 2746 15880 2748
rect 15584 2694 15630 2746
rect 15630 2694 15640 2746
rect 15664 2694 15694 2746
rect 15694 2694 15706 2746
rect 15706 2694 15720 2746
rect 15744 2694 15758 2746
rect 15758 2694 15770 2746
rect 15770 2694 15800 2746
rect 15824 2694 15834 2746
rect 15834 2694 15880 2746
rect 15584 2692 15640 2694
rect 15664 2692 15720 2694
rect 15744 2692 15800 2694
rect 15824 2692 15880 2694
rect 15584 1658 15640 1660
rect 15664 1658 15720 1660
rect 15744 1658 15800 1660
rect 15824 1658 15880 1660
rect 15584 1606 15630 1658
rect 15630 1606 15640 1658
rect 15664 1606 15694 1658
rect 15694 1606 15706 1658
rect 15706 1606 15720 1658
rect 15744 1606 15758 1658
rect 15758 1606 15770 1658
rect 15770 1606 15800 1658
rect 15824 1606 15834 1658
rect 15834 1606 15880 1658
rect 15584 1604 15640 1606
rect 15664 1604 15720 1606
rect 15744 1604 15800 1606
rect 15824 1604 15880 1606
rect 17130 10240 17186 10296
rect 16670 7928 16726 7984
rect 16670 7792 16726 7848
rect 16670 6452 16726 6488
rect 16670 6432 16672 6452
rect 16672 6432 16724 6452
rect 16724 6432 16726 6452
rect 16394 4120 16450 4176
rect 17590 9424 17646 9480
rect 17314 7520 17370 7576
rect 17222 7148 17224 7168
rect 17224 7148 17276 7168
rect 17276 7148 17278 7168
rect 17222 7112 17278 7148
rect 16946 5364 17002 5400
rect 16946 5344 16948 5364
rect 16948 5344 17000 5364
rect 17000 5344 17002 5364
rect 16854 3304 16910 3360
rect 17498 6976 17554 7032
rect 17406 6296 17462 6352
rect 20718 16088 20774 16144
rect 21270 19760 21326 19816
rect 20534 15136 20590 15192
rect 19890 14592 19946 14648
rect 20166 14320 20222 14376
rect 19379 13082 19435 13084
rect 19459 13082 19515 13084
rect 19539 13082 19595 13084
rect 19619 13082 19675 13084
rect 19379 13030 19425 13082
rect 19425 13030 19435 13082
rect 19459 13030 19489 13082
rect 19489 13030 19501 13082
rect 19501 13030 19515 13082
rect 19539 13030 19553 13082
rect 19553 13030 19565 13082
rect 19565 13030 19595 13082
rect 19619 13030 19629 13082
rect 19629 13030 19675 13082
rect 19379 13028 19435 13030
rect 19459 13028 19515 13030
rect 19539 13028 19595 13030
rect 19619 13028 19675 13030
rect 20626 14320 20682 14376
rect 20534 14184 20590 14240
rect 20626 13232 20682 13288
rect 21086 17720 21142 17776
rect 21270 17584 21326 17640
rect 21822 19896 21878 19952
rect 22006 18400 22062 18456
rect 23174 21242 23230 21244
rect 23254 21242 23310 21244
rect 23334 21242 23390 21244
rect 23414 21242 23470 21244
rect 23174 21190 23220 21242
rect 23220 21190 23230 21242
rect 23254 21190 23284 21242
rect 23284 21190 23296 21242
rect 23296 21190 23310 21242
rect 23334 21190 23348 21242
rect 23348 21190 23360 21242
rect 23360 21190 23390 21242
rect 23414 21190 23424 21242
rect 23424 21190 23470 21242
rect 23174 21188 23230 21190
rect 23254 21188 23310 21190
rect 23334 21188 23390 21190
rect 23414 21188 23470 21190
rect 23174 20154 23230 20156
rect 23254 20154 23310 20156
rect 23334 20154 23390 20156
rect 23414 20154 23470 20156
rect 23174 20102 23220 20154
rect 23220 20102 23230 20154
rect 23254 20102 23284 20154
rect 23284 20102 23296 20154
rect 23296 20102 23310 20154
rect 23334 20102 23348 20154
rect 23348 20102 23360 20154
rect 23360 20102 23390 20154
rect 23414 20102 23424 20154
rect 23424 20102 23470 20154
rect 23174 20100 23230 20102
rect 23254 20100 23310 20102
rect 23334 20100 23390 20102
rect 23414 20100 23470 20102
rect 23570 19236 23626 19272
rect 23570 19216 23572 19236
rect 23572 19216 23624 19236
rect 23624 19216 23626 19236
rect 23174 19066 23230 19068
rect 23254 19066 23310 19068
rect 23334 19066 23390 19068
rect 23414 19066 23470 19068
rect 23174 19014 23220 19066
rect 23220 19014 23230 19066
rect 23254 19014 23284 19066
rect 23284 19014 23296 19066
rect 23296 19014 23310 19066
rect 23334 19014 23348 19066
rect 23348 19014 23360 19066
rect 23360 19014 23390 19066
rect 23414 19014 23424 19066
rect 23424 19014 23470 19066
rect 23174 19012 23230 19014
rect 23254 19012 23310 19014
rect 23334 19012 23390 19014
rect 23414 19012 23470 19014
rect 23846 19760 23902 19816
rect 24398 20440 24454 20496
rect 24214 20168 24270 20224
rect 25134 21120 25190 21176
rect 24674 20032 24730 20088
rect 24122 18808 24178 18864
rect 24582 18944 24638 19000
rect 23846 18264 23902 18320
rect 22926 18164 22928 18184
rect 22928 18164 22980 18184
rect 22980 18164 22982 18184
rect 21638 16632 21694 16688
rect 21270 14592 21326 14648
rect 22926 18128 22982 18164
rect 22558 17992 22614 18048
rect 21914 17312 21970 17368
rect 22282 17448 22338 17504
rect 22466 17448 22522 17504
rect 22466 17040 22522 17096
rect 21822 16360 21878 16416
rect 21730 15680 21786 15736
rect 22006 14864 22062 14920
rect 19379 11994 19435 11996
rect 19459 11994 19515 11996
rect 19539 11994 19595 11996
rect 19619 11994 19675 11996
rect 19379 11942 19425 11994
rect 19425 11942 19435 11994
rect 19459 11942 19489 11994
rect 19489 11942 19501 11994
rect 19501 11942 19515 11994
rect 19539 11942 19553 11994
rect 19553 11942 19565 11994
rect 19565 11942 19595 11994
rect 19619 11942 19629 11994
rect 19629 11942 19675 11994
rect 19379 11940 19435 11942
rect 19459 11940 19515 11942
rect 19539 11940 19595 11942
rect 19619 11940 19675 11942
rect 19379 10906 19435 10908
rect 19459 10906 19515 10908
rect 19539 10906 19595 10908
rect 19619 10906 19675 10908
rect 19379 10854 19425 10906
rect 19425 10854 19435 10906
rect 19459 10854 19489 10906
rect 19489 10854 19501 10906
rect 19501 10854 19515 10906
rect 19539 10854 19553 10906
rect 19553 10854 19565 10906
rect 19565 10854 19595 10906
rect 19619 10854 19629 10906
rect 19629 10854 19675 10906
rect 19379 10852 19435 10854
rect 19459 10852 19515 10854
rect 19539 10852 19595 10854
rect 19619 10852 19675 10854
rect 18510 8880 18566 8936
rect 19379 9818 19435 9820
rect 19459 9818 19515 9820
rect 19539 9818 19595 9820
rect 19619 9818 19675 9820
rect 19379 9766 19425 9818
rect 19425 9766 19435 9818
rect 19459 9766 19489 9818
rect 19489 9766 19501 9818
rect 19501 9766 19515 9818
rect 19539 9766 19553 9818
rect 19553 9766 19565 9818
rect 19565 9766 19595 9818
rect 19619 9766 19629 9818
rect 19629 9766 19675 9818
rect 19379 9764 19435 9766
rect 19459 9764 19515 9766
rect 19539 9764 19595 9766
rect 19619 9764 19675 9766
rect 22466 15408 22522 15464
rect 22650 16788 22706 16824
rect 22650 16768 22652 16788
rect 22652 16768 22704 16788
rect 22704 16768 22706 16788
rect 23018 17992 23074 18048
rect 23174 17978 23230 17980
rect 23254 17978 23310 17980
rect 23334 17978 23390 17980
rect 23414 17978 23470 17980
rect 23174 17926 23220 17978
rect 23220 17926 23230 17978
rect 23254 17926 23284 17978
rect 23284 17926 23296 17978
rect 23296 17926 23310 17978
rect 23334 17926 23348 17978
rect 23348 17926 23360 17978
rect 23360 17926 23390 17978
rect 23414 17926 23424 17978
rect 23424 17926 23470 17978
rect 23174 17924 23230 17926
rect 23254 17924 23310 17926
rect 23334 17924 23390 17926
rect 23414 17924 23470 17926
rect 23938 18128 23994 18184
rect 23174 16890 23230 16892
rect 23254 16890 23310 16892
rect 23334 16890 23390 16892
rect 23414 16890 23470 16892
rect 23174 16838 23220 16890
rect 23220 16838 23230 16890
rect 23254 16838 23284 16890
rect 23284 16838 23296 16890
rect 23296 16838 23310 16890
rect 23334 16838 23348 16890
rect 23348 16838 23360 16890
rect 23360 16838 23390 16890
rect 23414 16838 23424 16890
rect 23424 16838 23470 16890
rect 23174 16836 23230 16838
rect 23254 16836 23310 16838
rect 23334 16836 23390 16838
rect 23414 16836 23470 16838
rect 23846 17040 23902 17096
rect 23662 16632 23718 16688
rect 22650 16088 22706 16144
rect 22834 15952 22890 16008
rect 23174 15802 23230 15804
rect 23254 15802 23310 15804
rect 23334 15802 23390 15804
rect 23414 15802 23470 15804
rect 23174 15750 23220 15802
rect 23220 15750 23230 15802
rect 23254 15750 23284 15802
rect 23284 15750 23296 15802
rect 23296 15750 23310 15802
rect 23334 15750 23348 15802
rect 23348 15750 23360 15802
rect 23360 15750 23390 15802
rect 23414 15750 23424 15802
rect 23424 15750 23470 15802
rect 23174 15748 23230 15750
rect 23254 15748 23310 15750
rect 23334 15748 23390 15750
rect 23414 15748 23470 15750
rect 23754 15272 23810 15328
rect 23662 15136 23718 15192
rect 22558 12144 22614 12200
rect 23174 14714 23230 14716
rect 23254 14714 23310 14716
rect 23334 14714 23390 14716
rect 23414 14714 23470 14716
rect 23174 14662 23220 14714
rect 23220 14662 23230 14714
rect 23254 14662 23284 14714
rect 23284 14662 23296 14714
rect 23296 14662 23310 14714
rect 23334 14662 23348 14714
rect 23348 14662 23360 14714
rect 23360 14662 23390 14714
rect 23414 14662 23424 14714
rect 23424 14662 23470 14714
rect 23174 14660 23230 14662
rect 23254 14660 23310 14662
rect 23334 14660 23390 14662
rect 23414 14660 23470 14662
rect 23570 14592 23626 14648
rect 23846 14728 23902 14784
rect 23570 14184 23626 14240
rect 23174 13626 23230 13628
rect 23254 13626 23310 13628
rect 23334 13626 23390 13628
rect 23414 13626 23470 13628
rect 23174 13574 23220 13626
rect 23220 13574 23230 13626
rect 23254 13574 23284 13626
rect 23284 13574 23296 13626
rect 23296 13574 23310 13626
rect 23334 13574 23348 13626
rect 23348 13574 23360 13626
rect 23360 13574 23390 13626
rect 23414 13574 23424 13626
rect 23424 13574 23470 13626
rect 23174 13572 23230 13574
rect 23254 13572 23310 13574
rect 23334 13572 23390 13574
rect 23414 13572 23470 13574
rect 23174 12538 23230 12540
rect 23254 12538 23310 12540
rect 23334 12538 23390 12540
rect 23414 12538 23470 12540
rect 23174 12486 23220 12538
rect 23220 12486 23230 12538
rect 23254 12486 23284 12538
rect 23284 12486 23296 12538
rect 23296 12486 23310 12538
rect 23334 12486 23348 12538
rect 23348 12486 23360 12538
rect 23360 12486 23390 12538
rect 23414 12486 23424 12538
rect 23424 12486 23470 12538
rect 23174 12484 23230 12486
rect 23254 12484 23310 12486
rect 23334 12484 23390 12486
rect 23414 12484 23470 12486
rect 22282 11600 22338 11656
rect 20442 10140 20444 10160
rect 20444 10140 20496 10160
rect 20496 10140 20498 10160
rect 20442 10104 20498 10140
rect 19379 8730 19435 8732
rect 19459 8730 19515 8732
rect 19539 8730 19595 8732
rect 19619 8730 19675 8732
rect 19379 8678 19425 8730
rect 19425 8678 19435 8730
rect 19459 8678 19489 8730
rect 19489 8678 19501 8730
rect 19501 8678 19515 8730
rect 19539 8678 19553 8730
rect 19553 8678 19565 8730
rect 19565 8678 19595 8730
rect 19619 8678 19629 8730
rect 19629 8678 19675 8730
rect 19379 8676 19435 8678
rect 19459 8676 19515 8678
rect 19539 8676 19595 8678
rect 19619 8676 19675 8678
rect 17958 7248 18014 7304
rect 19706 7928 19762 7984
rect 19379 7642 19435 7644
rect 19459 7642 19515 7644
rect 19539 7642 19595 7644
rect 19619 7642 19675 7644
rect 19379 7590 19425 7642
rect 19425 7590 19435 7642
rect 19459 7590 19489 7642
rect 19489 7590 19501 7642
rect 19501 7590 19515 7642
rect 19539 7590 19553 7642
rect 19553 7590 19565 7642
rect 19565 7590 19595 7642
rect 19619 7590 19629 7642
rect 19629 7590 19675 7642
rect 19379 7588 19435 7590
rect 19459 7588 19515 7590
rect 19539 7588 19595 7590
rect 19619 7588 19675 7590
rect 17774 5072 17830 5128
rect 16762 2760 16818 2816
rect 15382 584 15438 640
rect 15584 570 15640 572
rect 15664 570 15720 572
rect 15744 570 15800 572
rect 15824 570 15880 572
rect 15584 518 15630 570
rect 15630 518 15640 570
rect 15664 518 15694 570
rect 15694 518 15706 570
rect 15706 518 15720 570
rect 15744 518 15758 570
rect 15758 518 15770 570
rect 15770 518 15800 570
rect 15824 518 15834 570
rect 15834 518 15880 570
rect 15584 516 15640 518
rect 15664 516 15720 518
rect 15744 516 15800 518
rect 15824 516 15880 518
rect 17866 3576 17922 3632
rect 17958 2352 18014 2408
rect 18970 7248 19026 7304
rect 19154 6840 19210 6896
rect 18786 6296 18842 6352
rect 19379 6554 19435 6556
rect 19459 6554 19515 6556
rect 19539 6554 19595 6556
rect 19619 6554 19675 6556
rect 19379 6502 19425 6554
rect 19425 6502 19435 6554
rect 19459 6502 19489 6554
rect 19489 6502 19501 6554
rect 19501 6502 19515 6554
rect 19539 6502 19553 6554
rect 19553 6502 19565 6554
rect 19565 6502 19595 6554
rect 19619 6502 19629 6554
rect 19629 6502 19675 6554
rect 19379 6500 19435 6502
rect 19459 6500 19515 6502
rect 19539 6500 19595 6502
rect 19619 6500 19675 6502
rect 19062 3712 19118 3768
rect 18694 2896 18750 2952
rect 17866 1808 17922 1864
rect 18786 2388 18788 2408
rect 18788 2388 18840 2408
rect 18840 2388 18842 2408
rect 18786 2352 18842 2388
rect 19379 5466 19435 5468
rect 19459 5466 19515 5468
rect 19539 5466 19595 5468
rect 19619 5466 19675 5468
rect 19379 5414 19425 5466
rect 19425 5414 19435 5466
rect 19459 5414 19489 5466
rect 19489 5414 19501 5466
rect 19501 5414 19515 5466
rect 19539 5414 19553 5466
rect 19553 5414 19565 5466
rect 19565 5414 19595 5466
rect 19619 5414 19629 5466
rect 19629 5414 19675 5466
rect 19379 5412 19435 5414
rect 19459 5412 19515 5414
rect 19539 5412 19595 5414
rect 19619 5412 19675 5414
rect 19379 4378 19435 4380
rect 19459 4378 19515 4380
rect 19539 4378 19595 4380
rect 19619 4378 19675 4380
rect 19379 4326 19425 4378
rect 19425 4326 19435 4378
rect 19459 4326 19489 4378
rect 19489 4326 19501 4378
rect 19501 4326 19515 4378
rect 19539 4326 19553 4378
rect 19553 4326 19565 4378
rect 19565 4326 19595 4378
rect 19619 4326 19629 4378
rect 19629 4326 19675 4378
rect 19379 4324 19435 4326
rect 19459 4324 19515 4326
rect 19539 4324 19595 4326
rect 19619 4324 19675 4326
rect 20074 4528 20130 4584
rect 19379 3290 19435 3292
rect 19459 3290 19515 3292
rect 19539 3290 19595 3292
rect 19619 3290 19675 3292
rect 19379 3238 19425 3290
rect 19425 3238 19435 3290
rect 19459 3238 19489 3290
rect 19489 3238 19501 3290
rect 19501 3238 19515 3290
rect 19539 3238 19553 3290
rect 19553 3238 19565 3290
rect 19565 3238 19595 3290
rect 19619 3238 19629 3290
rect 19629 3238 19675 3290
rect 19379 3236 19435 3238
rect 19459 3236 19515 3238
rect 19539 3236 19595 3238
rect 19619 3236 19675 3238
rect 20902 8472 20958 8528
rect 20626 6160 20682 6216
rect 21270 10124 21326 10160
rect 21270 10104 21272 10124
rect 21272 10104 21324 10124
rect 21324 10104 21326 10124
rect 21086 9424 21142 9480
rect 20902 4684 20958 4720
rect 20902 4664 20904 4684
rect 20904 4664 20956 4684
rect 20956 4664 20958 4684
rect 20626 3984 20682 4040
rect 19379 2202 19435 2204
rect 19459 2202 19515 2204
rect 19539 2202 19595 2204
rect 19619 2202 19675 2204
rect 19379 2150 19425 2202
rect 19425 2150 19435 2202
rect 19459 2150 19489 2202
rect 19489 2150 19501 2202
rect 19501 2150 19515 2202
rect 19539 2150 19553 2202
rect 19553 2150 19565 2202
rect 19565 2150 19595 2202
rect 19619 2150 19629 2202
rect 19629 2150 19675 2202
rect 19379 2148 19435 2150
rect 19459 2148 19515 2150
rect 19539 2148 19595 2150
rect 19619 2148 19675 2150
rect 20534 2080 20590 2136
rect 20074 1128 20130 1184
rect 19379 1114 19435 1116
rect 19459 1114 19515 1116
rect 19539 1114 19595 1116
rect 19619 1114 19675 1116
rect 19379 1062 19425 1114
rect 19425 1062 19435 1114
rect 19459 1062 19489 1114
rect 19489 1062 19501 1114
rect 19501 1062 19515 1114
rect 19539 1062 19553 1114
rect 19553 1062 19565 1114
rect 19565 1062 19595 1114
rect 19619 1062 19629 1114
rect 19629 1062 19675 1114
rect 19379 1060 19435 1062
rect 19459 1060 19515 1062
rect 19539 1060 19595 1062
rect 19619 1060 19675 1062
rect 18234 720 18290 776
rect 21362 8336 21418 8392
rect 23174 11450 23230 11452
rect 23254 11450 23310 11452
rect 23334 11450 23390 11452
rect 23414 11450 23470 11452
rect 23174 11398 23220 11450
rect 23220 11398 23230 11450
rect 23254 11398 23284 11450
rect 23284 11398 23296 11450
rect 23296 11398 23310 11450
rect 23334 11398 23348 11450
rect 23348 11398 23360 11450
rect 23360 11398 23390 11450
rect 23414 11398 23424 11450
rect 23424 11398 23470 11450
rect 23174 11396 23230 11398
rect 23254 11396 23310 11398
rect 23334 11396 23390 11398
rect 23414 11396 23470 11398
rect 23174 10362 23230 10364
rect 23254 10362 23310 10364
rect 23334 10362 23390 10364
rect 23414 10362 23470 10364
rect 23174 10310 23220 10362
rect 23220 10310 23230 10362
rect 23254 10310 23284 10362
rect 23284 10310 23296 10362
rect 23296 10310 23310 10362
rect 23334 10310 23348 10362
rect 23348 10310 23360 10362
rect 23360 10310 23390 10362
rect 23414 10310 23424 10362
rect 23424 10310 23470 10362
rect 23174 10308 23230 10310
rect 23254 10308 23310 10310
rect 23334 10308 23390 10310
rect 23414 10308 23470 10310
rect 24122 16224 24178 16280
rect 24398 18536 24454 18592
rect 24398 16496 24454 16552
rect 24306 16088 24362 16144
rect 24398 15408 24454 15464
rect 25594 20168 25650 20224
rect 24858 17992 24914 18048
rect 24674 16360 24730 16416
rect 24858 15952 24914 16008
rect 25686 18808 25742 18864
rect 25594 17312 25650 17368
rect 26969 21786 27025 21788
rect 27049 21786 27105 21788
rect 27129 21786 27185 21788
rect 27209 21786 27265 21788
rect 26969 21734 27015 21786
rect 27015 21734 27025 21786
rect 27049 21734 27079 21786
rect 27079 21734 27091 21786
rect 27091 21734 27105 21786
rect 27129 21734 27143 21786
rect 27143 21734 27155 21786
rect 27155 21734 27185 21786
rect 27209 21734 27219 21786
rect 27219 21734 27265 21786
rect 26969 21732 27025 21734
rect 27049 21732 27105 21734
rect 27129 21732 27185 21734
rect 27209 21732 27265 21734
rect 26054 20576 26110 20632
rect 24674 15816 24730 15872
rect 25502 15544 25558 15600
rect 24674 15000 24730 15056
rect 24214 14048 24270 14104
rect 23938 13776 23994 13832
rect 23846 13640 23902 13696
rect 23938 12688 23994 12744
rect 24306 11192 24362 11248
rect 23846 11092 23848 11112
rect 23848 11092 23900 11112
rect 23900 11092 23902 11112
rect 23846 11056 23902 11092
rect 23754 10104 23810 10160
rect 22006 9016 22062 9072
rect 22466 8744 22522 8800
rect 22282 8372 22284 8392
rect 22284 8372 22336 8392
rect 22336 8372 22338 8392
rect 22282 8336 22338 8372
rect 21822 6432 21878 6488
rect 21546 5752 21602 5808
rect 22006 4392 22062 4448
rect 22282 4120 22338 4176
rect 23174 9274 23230 9276
rect 23254 9274 23310 9276
rect 23334 9274 23390 9276
rect 23414 9274 23470 9276
rect 23174 9222 23220 9274
rect 23220 9222 23230 9274
rect 23254 9222 23284 9274
rect 23284 9222 23296 9274
rect 23296 9222 23310 9274
rect 23334 9222 23348 9274
rect 23348 9222 23360 9274
rect 23360 9222 23390 9274
rect 23414 9222 23424 9274
rect 23424 9222 23470 9274
rect 23174 9220 23230 9222
rect 23254 9220 23310 9222
rect 23334 9220 23390 9222
rect 23414 9220 23470 9222
rect 23174 8186 23230 8188
rect 23254 8186 23310 8188
rect 23334 8186 23390 8188
rect 23414 8186 23470 8188
rect 23174 8134 23220 8186
rect 23220 8134 23230 8186
rect 23254 8134 23284 8186
rect 23284 8134 23296 8186
rect 23296 8134 23310 8186
rect 23334 8134 23348 8186
rect 23348 8134 23360 8186
rect 23360 8134 23390 8186
rect 23414 8134 23424 8186
rect 23424 8134 23470 8186
rect 23174 8132 23230 8134
rect 23254 8132 23310 8134
rect 23334 8132 23390 8134
rect 23414 8132 23470 8134
rect 23174 7098 23230 7100
rect 23254 7098 23310 7100
rect 23334 7098 23390 7100
rect 23414 7098 23470 7100
rect 23174 7046 23220 7098
rect 23220 7046 23230 7098
rect 23254 7046 23284 7098
rect 23284 7046 23296 7098
rect 23296 7046 23310 7098
rect 23334 7046 23348 7098
rect 23348 7046 23360 7098
rect 23360 7046 23390 7098
rect 23414 7046 23424 7098
rect 23424 7046 23470 7098
rect 23174 7044 23230 7046
rect 23254 7044 23310 7046
rect 23334 7044 23390 7046
rect 23414 7044 23470 7046
rect 23754 9016 23810 9072
rect 25042 14048 25098 14104
rect 24858 13640 24914 13696
rect 25686 14320 25742 14376
rect 24766 11736 24822 11792
rect 24122 9460 24124 9480
rect 24124 9460 24176 9480
rect 24176 9460 24178 9480
rect 24122 9424 24178 9460
rect 24214 8472 24270 8528
rect 23174 6010 23230 6012
rect 23254 6010 23310 6012
rect 23334 6010 23390 6012
rect 23414 6010 23470 6012
rect 23174 5958 23220 6010
rect 23220 5958 23230 6010
rect 23254 5958 23284 6010
rect 23284 5958 23296 6010
rect 23296 5958 23310 6010
rect 23334 5958 23348 6010
rect 23348 5958 23360 6010
rect 23360 5958 23390 6010
rect 23414 5958 23424 6010
rect 23424 5958 23470 6010
rect 23174 5956 23230 5958
rect 23254 5956 23310 5958
rect 23334 5956 23390 5958
rect 23414 5956 23470 5958
rect 22650 5480 22706 5536
rect 23570 5652 23572 5672
rect 23572 5652 23624 5672
rect 23624 5652 23626 5672
rect 23570 5616 23626 5652
rect 23386 5208 23442 5264
rect 23662 5208 23718 5264
rect 22834 4392 22890 4448
rect 23174 4922 23230 4924
rect 23254 4922 23310 4924
rect 23334 4922 23390 4924
rect 23414 4922 23470 4924
rect 23174 4870 23220 4922
rect 23220 4870 23230 4922
rect 23254 4870 23284 4922
rect 23284 4870 23296 4922
rect 23296 4870 23310 4922
rect 23334 4870 23348 4922
rect 23348 4870 23360 4922
rect 23360 4870 23390 4922
rect 23414 4870 23424 4922
rect 23424 4870 23470 4922
rect 23174 4868 23230 4870
rect 23254 4868 23310 4870
rect 23334 4868 23390 4870
rect 23414 4868 23470 4870
rect 23174 3834 23230 3836
rect 23254 3834 23310 3836
rect 23334 3834 23390 3836
rect 23414 3834 23470 3836
rect 23174 3782 23220 3834
rect 23220 3782 23230 3834
rect 23254 3782 23284 3834
rect 23284 3782 23296 3834
rect 23296 3782 23310 3834
rect 23334 3782 23348 3834
rect 23348 3782 23360 3834
rect 23360 3782 23390 3834
rect 23414 3782 23424 3834
rect 23424 3782 23470 3834
rect 23174 3780 23230 3782
rect 23254 3780 23310 3782
rect 23334 3780 23390 3782
rect 23414 3780 23470 3782
rect 22742 3032 22798 3088
rect 22650 1400 22706 1456
rect 23174 2746 23230 2748
rect 23254 2746 23310 2748
rect 23334 2746 23390 2748
rect 23414 2746 23470 2748
rect 23174 2694 23220 2746
rect 23220 2694 23230 2746
rect 23254 2694 23284 2746
rect 23284 2694 23296 2746
rect 23296 2694 23310 2746
rect 23334 2694 23348 2746
rect 23348 2694 23360 2746
rect 23360 2694 23390 2746
rect 23414 2694 23424 2746
rect 23424 2694 23470 2746
rect 23174 2692 23230 2694
rect 23254 2692 23310 2694
rect 23334 2692 23390 2694
rect 23414 2692 23470 2694
rect 25042 6976 25098 7032
rect 24398 6432 24454 6488
rect 23662 2216 23718 2272
rect 24674 5652 24676 5672
rect 24676 5652 24728 5672
rect 24728 5652 24730 5672
rect 24674 5616 24730 5652
rect 23174 1658 23230 1660
rect 23254 1658 23310 1660
rect 23334 1658 23390 1660
rect 23414 1658 23470 1660
rect 23174 1606 23220 1658
rect 23220 1606 23230 1658
rect 23254 1606 23284 1658
rect 23284 1606 23296 1658
rect 23296 1606 23310 1658
rect 23334 1606 23348 1658
rect 23348 1606 23360 1658
rect 23360 1606 23390 1658
rect 23414 1606 23424 1658
rect 23424 1606 23470 1658
rect 23174 1604 23230 1606
rect 23254 1604 23310 1606
rect 23334 1604 23390 1606
rect 23414 1604 23470 1606
rect 21454 756 21456 776
rect 21456 756 21508 776
rect 21508 756 21510 776
rect 21454 720 21510 756
rect 24582 4392 24638 4448
rect 24858 4684 24914 4720
rect 24858 4664 24860 4684
rect 24860 4664 24912 4684
rect 24912 4664 24914 4684
rect 23938 756 23940 776
rect 23940 756 23992 776
rect 23992 756 23994 776
rect 23938 720 23994 756
rect 24306 2080 24362 2136
rect 24306 1420 24362 1456
rect 24306 1400 24308 1420
rect 24308 1400 24360 1420
rect 24360 1400 24362 1420
rect 23174 570 23230 572
rect 23254 570 23310 572
rect 23334 570 23390 572
rect 23414 570 23470 572
rect 23174 518 23220 570
rect 23220 518 23230 570
rect 23254 518 23284 570
rect 23284 518 23296 570
rect 23296 518 23310 570
rect 23334 518 23348 570
rect 23348 518 23360 570
rect 23360 518 23390 570
rect 23414 518 23424 570
rect 23424 518 23470 570
rect 23174 516 23230 518
rect 23254 516 23310 518
rect 23334 516 23390 518
rect 23414 516 23470 518
rect 25870 16108 25926 16144
rect 25870 16088 25872 16108
rect 25872 16088 25924 16108
rect 25924 16088 25926 16108
rect 26054 15408 26110 15464
rect 26514 18944 26570 19000
rect 26698 18808 26754 18864
rect 26698 17584 26754 17640
rect 26606 17312 26662 17368
rect 26238 15952 26294 16008
rect 26238 15272 26294 15328
rect 26514 15136 26570 15192
rect 26969 20698 27025 20700
rect 27049 20698 27105 20700
rect 27129 20698 27185 20700
rect 27209 20698 27265 20700
rect 26969 20646 27015 20698
rect 27015 20646 27025 20698
rect 27049 20646 27079 20698
rect 27079 20646 27091 20698
rect 27091 20646 27105 20698
rect 27129 20646 27143 20698
rect 27143 20646 27155 20698
rect 27155 20646 27185 20698
rect 27209 20646 27219 20698
rect 27219 20646 27265 20698
rect 26969 20644 27025 20646
rect 27049 20644 27105 20646
rect 27129 20644 27185 20646
rect 27209 20644 27265 20646
rect 26969 19610 27025 19612
rect 27049 19610 27105 19612
rect 27129 19610 27185 19612
rect 27209 19610 27265 19612
rect 26969 19558 27015 19610
rect 27015 19558 27025 19610
rect 27049 19558 27079 19610
rect 27079 19558 27091 19610
rect 27091 19558 27105 19610
rect 27129 19558 27143 19610
rect 27143 19558 27155 19610
rect 27155 19558 27185 19610
rect 27209 19558 27219 19610
rect 27219 19558 27265 19610
rect 26969 19556 27025 19558
rect 27049 19556 27105 19558
rect 27129 19556 27185 19558
rect 27209 19556 27265 19558
rect 27158 18808 27214 18864
rect 26969 18522 27025 18524
rect 27049 18522 27105 18524
rect 27129 18522 27185 18524
rect 27209 18522 27265 18524
rect 26969 18470 27015 18522
rect 27015 18470 27025 18522
rect 27049 18470 27079 18522
rect 27079 18470 27091 18522
rect 27091 18470 27105 18522
rect 27129 18470 27143 18522
rect 27143 18470 27155 18522
rect 27155 18470 27185 18522
rect 27209 18470 27219 18522
rect 27219 18470 27265 18522
rect 26969 18468 27025 18470
rect 27049 18468 27105 18470
rect 27129 18468 27185 18470
rect 27209 18468 27265 18470
rect 27158 17720 27214 17776
rect 26969 17434 27025 17436
rect 27049 17434 27105 17436
rect 27129 17434 27185 17436
rect 27209 17434 27265 17436
rect 26969 17382 27015 17434
rect 27015 17382 27025 17434
rect 27049 17382 27079 17434
rect 27079 17382 27091 17434
rect 27091 17382 27105 17434
rect 27129 17382 27143 17434
rect 27143 17382 27155 17434
rect 27155 17382 27185 17434
rect 27209 17382 27219 17434
rect 27219 17382 27265 17434
rect 26969 17380 27025 17382
rect 27049 17380 27105 17382
rect 27129 17380 27185 17382
rect 27209 17380 27265 17382
rect 26969 16346 27025 16348
rect 27049 16346 27105 16348
rect 27129 16346 27185 16348
rect 27209 16346 27265 16348
rect 26969 16294 27015 16346
rect 27015 16294 27025 16346
rect 27049 16294 27079 16346
rect 27079 16294 27091 16346
rect 27091 16294 27105 16346
rect 27129 16294 27143 16346
rect 27143 16294 27155 16346
rect 27155 16294 27185 16346
rect 27209 16294 27219 16346
rect 27219 16294 27265 16346
rect 26969 16292 27025 16294
rect 27049 16292 27105 16294
rect 27129 16292 27185 16294
rect 27209 16292 27265 16294
rect 26606 13368 26662 13424
rect 26969 15258 27025 15260
rect 27049 15258 27105 15260
rect 27129 15258 27185 15260
rect 27209 15258 27265 15260
rect 26969 15206 27015 15258
rect 27015 15206 27025 15258
rect 27049 15206 27079 15258
rect 27079 15206 27091 15258
rect 27091 15206 27105 15258
rect 27129 15206 27143 15258
rect 27143 15206 27155 15258
rect 27155 15206 27185 15258
rect 27209 15206 27219 15258
rect 27219 15206 27265 15258
rect 26969 15204 27025 15206
rect 27049 15204 27105 15206
rect 27129 15204 27185 15206
rect 27209 15204 27265 15206
rect 27066 14592 27122 14648
rect 26969 14170 27025 14172
rect 27049 14170 27105 14172
rect 27129 14170 27185 14172
rect 27209 14170 27265 14172
rect 26969 14118 27015 14170
rect 27015 14118 27025 14170
rect 27049 14118 27079 14170
rect 27079 14118 27091 14170
rect 27091 14118 27105 14170
rect 27129 14118 27143 14170
rect 27143 14118 27155 14170
rect 27155 14118 27185 14170
rect 27209 14118 27219 14170
rect 27219 14118 27265 14170
rect 26969 14116 27025 14118
rect 27049 14116 27105 14118
rect 27129 14116 27185 14118
rect 27209 14116 27265 14118
rect 27618 14864 27674 14920
rect 28078 18808 28134 18864
rect 27894 15408 27950 15464
rect 28078 15816 28134 15872
rect 27802 14592 27858 14648
rect 25134 3576 25190 3632
rect 26422 11056 26478 11112
rect 26514 8336 26570 8392
rect 26969 13082 27025 13084
rect 27049 13082 27105 13084
rect 27129 13082 27185 13084
rect 27209 13082 27265 13084
rect 26969 13030 27015 13082
rect 27015 13030 27025 13082
rect 27049 13030 27079 13082
rect 27079 13030 27091 13082
rect 27091 13030 27105 13082
rect 27129 13030 27143 13082
rect 27143 13030 27155 13082
rect 27155 13030 27185 13082
rect 27209 13030 27219 13082
rect 27219 13030 27265 13082
rect 26969 13028 27025 13030
rect 27049 13028 27105 13030
rect 27129 13028 27185 13030
rect 27209 13028 27265 13030
rect 26969 11994 27025 11996
rect 27049 11994 27105 11996
rect 27129 11994 27185 11996
rect 27209 11994 27265 11996
rect 26969 11942 27015 11994
rect 27015 11942 27025 11994
rect 27049 11942 27079 11994
rect 27079 11942 27091 11994
rect 27091 11942 27105 11994
rect 27129 11942 27143 11994
rect 27143 11942 27155 11994
rect 27155 11942 27185 11994
rect 27209 11942 27219 11994
rect 27219 11942 27265 11994
rect 26969 11940 27025 11942
rect 27049 11940 27105 11942
rect 27129 11940 27185 11942
rect 27209 11940 27265 11942
rect 28538 20032 28594 20088
rect 28354 19916 28410 19952
rect 28354 19896 28356 19916
rect 28356 19896 28408 19916
rect 28408 19896 28410 19916
rect 28354 17212 28356 17232
rect 28356 17212 28408 17232
rect 28408 17212 28410 17232
rect 28354 17176 28410 17212
rect 27986 13232 28042 13288
rect 26969 10906 27025 10908
rect 27049 10906 27105 10908
rect 27129 10906 27185 10908
rect 27209 10906 27265 10908
rect 26969 10854 27015 10906
rect 27015 10854 27025 10906
rect 27049 10854 27079 10906
rect 27079 10854 27091 10906
rect 27091 10854 27105 10906
rect 27129 10854 27143 10906
rect 27143 10854 27155 10906
rect 27155 10854 27185 10906
rect 27209 10854 27219 10906
rect 27219 10854 27265 10906
rect 26969 10852 27025 10854
rect 27049 10852 27105 10854
rect 27129 10852 27185 10854
rect 27209 10852 27265 10854
rect 28630 16088 28686 16144
rect 28538 13796 28594 13832
rect 28538 13776 28540 13796
rect 28540 13776 28592 13796
rect 28592 13776 28594 13796
rect 28722 14728 28778 14784
rect 28722 14612 28778 14648
rect 28722 14592 28724 14612
rect 28724 14592 28776 14612
rect 28776 14592 28778 14612
rect 26969 9818 27025 9820
rect 27049 9818 27105 9820
rect 27129 9818 27185 9820
rect 27209 9818 27265 9820
rect 26969 9766 27015 9818
rect 27015 9766 27025 9818
rect 27049 9766 27079 9818
rect 27079 9766 27091 9818
rect 27091 9766 27105 9818
rect 27129 9766 27143 9818
rect 27143 9766 27155 9818
rect 27155 9766 27185 9818
rect 27209 9766 27219 9818
rect 27219 9766 27265 9818
rect 26969 9764 27025 9766
rect 27049 9764 27105 9766
rect 27129 9764 27185 9766
rect 27209 9764 27265 9766
rect 26790 8880 26846 8936
rect 25778 7248 25834 7304
rect 26238 6316 26294 6352
rect 26238 6296 26240 6316
rect 26240 6296 26292 6316
rect 26292 6296 26294 6316
rect 25870 5480 25926 5536
rect 26330 5480 26386 5536
rect 26969 8730 27025 8732
rect 27049 8730 27105 8732
rect 27129 8730 27185 8732
rect 27209 8730 27265 8732
rect 26969 8678 27015 8730
rect 27015 8678 27025 8730
rect 27049 8678 27079 8730
rect 27079 8678 27091 8730
rect 27091 8678 27105 8730
rect 27129 8678 27143 8730
rect 27143 8678 27155 8730
rect 27155 8678 27185 8730
rect 27209 8678 27219 8730
rect 27219 8678 27265 8730
rect 26969 8676 27025 8678
rect 27049 8676 27105 8678
rect 27129 8676 27185 8678
rect 27209 8676 27265 8678
rect 26969 7642 27025 7644
rect 27049 7642 27105 7644
rect 27129 7642 27185 7644
rect 27209 7642 27265 7644
rect 26969 7590 27015 7642
rect 27015 7590 27025 7642
rect 27049 7590 27079 7642
rect 27079 7590 27091 7642
rect 27091 7590 27105 7642
rect 27129 7590 27143 7642
rect 27143 7590 27155 7642
rect 27155 7590 27185 7642
rect 27209 7590 27219 7642
rect 27219 7590 27265 7642
rect 26969 7588 27025 7590
rect 27049 7588 27105 7590
rect 27129 7588 27185 7590
rect 27209 7588 27265 7590
rect 26969 6554 27025 6556
rect 27049 6554 27105 6556
rect 27129 6554 27185 6556
rect 27209 6554 27265 6556
rect 26969 6502 27015 6554
rect 27015 6502 27025 6554
rect 27049 6502 27079 6554
rect 27079 6502 27091 6554
rect 27091 6502 27105 6554
rect 27129 6502 27143 6554
rect 27143 6502 27155 6554
rect 27155 6502 27185 6554
rect 27209 6502 27219 6554
rect 27219 6502 27265 6554
rect 26969 6500 27025 6502
rect 27049 6500 27105 6502
rect 27129 6500 27185 6502
rect 27209 6500 27265 6502
rect 26422 2216 26478 2272
rect 25962 1420 26018 1456
rect 25962 1400 25964 1420
rect 25964 1400 26016 1420
rect 26016 1400 26018 1420
rect 25778 720 25834 776
rect 26969 5466 27025 5468
rect 27049 5466 27105 5468
rect 27129 5466 27185 5468
rect 27209 5466 27265 5468
rect 26969 5414 27015 5466
rect 27015 5414 27025 5466
rect 27049 5414 27079 5466
rect 27079 5414 27091 5466
rect 27091 5414 27105 5466
rect 27129 5414 27143 5466
rect 27143 5414 27155 5466
rect 27155 5414 27185 5466
rect 27209 5414 27219 5466
rect 27219 5414 27265 5466
rect 26969 5412 27025 5414
rect 27049 5412 27105 5414
rect 27129 5412 27185 5414
rect 27209 5412 27265 5414
rect 27618 5752 27674 5808
rect 27342 5208 27398 5264
rect 26969 4378 27025 4380
rect 27049 4378 27105 4380
rect 27129 4378 27185 4380
rect 27209 4378 27265 4380
rect 26969 4326 27015 4378
rect 27015 4326 27025 4378
rect 27049 4326 27079 4378
rect 27079 4326 27091 4378
rect 27091 4326 27105 4378
rect 27129 4326 27143 4378
rect 27143 4326 27155 4378
rect 27155 4326 27185 4378
rect 27209 4326 27219 4378
rect 27219 4326 27265 4378
rect 26969 4324 27025 4326
rect 27049 4324 27105 4326
rect 27129 4324 27185 4326
rect 27209 4324 27265 4326
rect 26969 3290 27025 3292
rect 27049 3290 27105 3292
rect 27129 3290 27185 3292
rect 27209 3290 27265 3292
rect 26969 3238 27015 3290
rect 27015 3238 27025 3290
rect 27049 3238 27079 3290
rect 27079 3238 27091 3290
rect 27091 3238 27105 3290
rect 27129 3238 27143 3290
rect 27143 3238 27155 3290
rect 27155 3238 27185 3290
rect 27209 3238 27219 3290
rect 27219 3238 27265 3290
rect 26969 3236 27025 3238
rect 27049 3236 27105 3238
rect 27129 3236 27185 3238
rect 27209 3236 27265 3238
rect 27066 2896 27122 2952
rect 27618 4528 27674 4584
rect 27710 4120 27766 4176
rect 26969 2202 27025 2204
rect 27049 2202 27105 2204
rect 27129 2202 27185 2204
rect 27209 2202 27265 2204
rect 26969 2150 27015 2202
rect 27015 2150 27025 2202
rect 27049 2150 27079 2202
rect 27079 2150 27091 2202
rect 27091 2150 27105 2202
rect 27129 2150 27143 2202
rect 27143 2150 27155 2202
rect 27155 2150 27185 2202
rect 27209 2150 27219 2202
rect 27219 2150 27265 2202
rect 26969 2148 27025 2150
rect 27049 2148 27105 2150
rect 27129 2148 27185 2150
rect 27209 2148 27265 2150
rect 26974 1420 27030 1456
rect 27434 1944 27490 2000
rect 26974 1400 26976 1420
rect 26976 1400 27028 1420
rect 27028 1400 27030 1420
rect 26882 1264 26938 1320
rect 26330 1128 26386 1184
rect 26969 1114 27025 1116
rect 27049 1114 27105 1116
rect 27129 1114 27185 1116
rect 27209 1114 27265 1116
rect 26969 1062 27015 1114
rect 27015 1062 27025 1114
rect 27049 1062 27079 1114
rect 27079 1062 27091 1114
rect 27091 1062 27105 1114
rect 27129 1062 27143 1114
rect 27143 1062 27155 1114
rect 27155 1062 27185 1114
rect 27209 1062 27219 1114
rect 27219 1062 27265 1114
rect 26969 1060 27025 1062
rect 27049 1060 27105 1062
rect 27129 1060 27185 1062
rect 27209 1060 27265 1062
rect 26238 856 26294 912
rect 27894 3440 27950 3496
rect 29274 16768 29330 16824
rect 29182 16496 29238 16552
rect 29090 16360 29146 16416
rect 28998 16244 29054 16280
rect 28998 16224 29000 16244
rect 29000 16224 29052 16244
rect 29052 16224 29054 16244
rect 29366 16088 29422 16144
rect 29090 15680 29146 15736
rect 29090 14048 29146 14104
rect 28998 13948 29000 13968
rect 29000 13948 29052 13968
rect 29052 13948 29054 13968
rect 28998 13912 29054 13948
rect 29274 13812 29276 13832
rect 29276 13812 29328 13832
rect 29328 13812 29330 13832
rect 29274 13776 29330 13812
rect 29366 13640 29422 13696
rect 29274 13524 29330 13560
rect 29274 13504 29276 13524
rect 29276 13504 29328 13524
rect 29328 13504 29330 13524
rect 29274 13368 29330 13424
rect 29090 12980 29146 13016
rect 29090 12960 29092 12980
rect 29092 12960 29144 12980
rect 29144 12960 29146 12980
rect 28998 12824 29054 12880
rect 28906 12300 28962 12336
rect 28906 12280 28908 12300
rect 28908 12280 28960 12300
rect 28960 12280 28962 12300
rect 29274 12708 29330 12744
rect 29274 12688 29276 12708
rect 29276 12688 29328 12708
rect 29328 12688 29330 12708
rect 29274 12416 29330 12472
rect 28630 6160 28686 6216
rect 28722 5072 28778 5128
rect 28538 3984 28594 4040
rect 29550 19352 29606 19408
rect 29550 17040 29606 17096
rect 29734 18672 29790 18728
rect 30102 18264 30158 18320
rect 30102 16652 30158 16688
rect 30102 16632 30104 16652
rect 30104 16632 30156 16652
rect 30156 16632 30158 16652
rect 30378 18028 30380 18048
rect 30380 18028 30432 18048
rect 30432 18028 30434 18048
rect 30378 17992 30434 18028
rect 30194 16224 30250 16280
rect 30010 15816 30066 15872
rect 29918 14476 29974 14512
rect 29918 14456 29920 14476
rect 29920 14456 29972 14476
rect 29972 14456 29974 14476
rect 30010 12724 30012 12744
rect 30012 12724 30064 12744
rect 30064 12724 30066 12744
rect 30010 12688 30066 12724
rect 29918 12144 29974 12200
rect 30764 21242 30820 21244
rect 30844 21242 30900 21244
rect 30924 21242 30980 21244
rect 31004 21242 31060 21244
rect 30764 21190 30810 21242
rect 30810 21190 30820 21242
rect 30844 21190 30874 21242
rect 30874 21190 30886 21242
rect 30886 21190 30900 21242
rect 30924 21190 30938 21242
rect 30938 21190 30950 21242
rect 30950 21190 30980 21242
rect 31004 21190 31014 21242
rect 31014 21190 31060 21242
rect 30764 21188 30820 21190
rect 30844 21188 30900 21190
rect 30924 21188 30980 21190
rect 31004 21188 31060 21190
rect 30764 20154 30820 20156
rect 30844 20154 30900 20156
rect 30924 20154 30980 20156
rect 31004 20154 31060 20156
rect 30764 20102 30810 20154
rect 30810 20102 30820 20154
rect 30844 20102 30874 20154
rect 30874 20102 30886 20154
rect 30886 20102 30900 20154
rect 30924 20102 30938 20154
rect 30938 20102 30950 20154
rect 30950 20102 30980 20154
rect 31004 20102 31014 20154
rect 31014 20102 31060 20154
rect 30764 20100 30820 20102
rect 30844 20100 30900 20102
rect 30924 20100 30980 20102
rect 31004 20100 31060 20102
rect 30764 19066 30820 19068
rect 30844 19066 30900 19068
rect 30924 19066 30980 19068
rect 31004 19066 31060 19068
rect 30764 19014 30810 19066
rect 30810 19014 30820 19066
rect 30844 19014 30874 19066
rect 30874 19014 30886 19066
rect 30886 19014 30900 19066
rect 30924 19014 30938 19066
rect 30938 19014 30950 19066
rect 30950 19014 30980 19066
rect 31004 19014 31014 19066
rect 31014 19014 31060 19066
rect 30764 19012 30820 19014
rect 30844 19012 30900 19014
rect 30924 19012 30980 19014
rect 31004 19012 31060 19014
rect 30654 18128 30710 18184
rect 30764 17978 30820 17980
rect 30844 17978 30900 17980
rect 30924 17978 30980 17980
rect 31004 17978 31060 17980
rect 30764 17926 30810 17978
rect 30810 17926 30820 17978
rect 30844 17926 30874 17978
rect 30874 17926 30886 17978
rect 30886 17926 30900 17978
rect 30924 17926 30938 17978
rect 30938 17926 30950 17978
rect 30950 17926 30980 17978
rect 31004 17926 31014 17978
rect 31014 17926 31060 17978
rect 30764 17924 30820 17926
rect 30844 17924 30900 17926
rect 30924 17924 30980 17926
rect 31004 17924 31060 17926
rect 30764 16890 30820 16892
rect 30844 16890 30900 16892
rect 30924 16890 30980 16892
rect 31004 16890 31060 16892
rect 30764 16838 30810 16890
rect 30810 16838 30820 16890
rect 30844 16838 30874 16890
rect 30874 16838 30886 16890
rect 30886 16838 30900 16890
rect 30924 16838 30938 16890
rect 30938 16838 30950 16890
rect 30950 16838 30980 16890
rect 31004 16838 31014 16890
rect 31014 16838 31060 16890
rect 30764 16836 30820 16838
rect 30844 16836 30900 16838
rect 30924 16836 30980 16838
rect 31004 16836 31060 16838
rect 31114 15952 31170 16008
rect 30764 15802 30820 15804
rect 30844 15802 30900 15804
rect 30924 15802 30980 15804
rect 31004 15802 31060 15804
rect 30764 15750 30810 15802
rect 30810 15750 30820 15802
rect 30844 15750 30874 15802
rect 30874 15750 30886 15802
rect 30886 15750 30900 15802
rect 30924 15750 30938 15802
rect 30938 15750 30950 15802
rect 30950 15750 30980 15802
rect 31004 15750 31014 15802
rect 31014 15750 31060 15802
rect 30764 15748 30820 15750
rect 30844 15748 30900 15750
rect 30924 15748 30980 15750
rect 31004 15748 31060 15750
rect 30286 13776 30342 13832
rect 30286 13640 30342 13696
rect 30764 14714 30820 14716
rect 30844 14714 30900 14716
rect 30924 14714 30980 14716
rect 31004 14714 31060 14716
rect 30764 14662 30810 14714
rect 30810 14662 30820 14714
rect 30844 14662 30874 14714
rect 30874 14662 30886 14714
rect 30886 14662 30900 14714
rect 30924 14662 30938 14714
rect 30938 14662 30950 14714
rect 30950 14662 30980 14714
rect 31004 14662 31014 14714
rect 31014 14662 31060 14714
rect 30764 14660 30820 14662
rect 30844 14660 30900 14662
rect 30924 14660 30980 14662
rect 31004 14660 31060 14662
rect 30764 13626 30820 13628
rect 30844 13626 30900 13628
rect 30924 13626 30980 13628
rect 31004 13626 31060 13628
rect 30764 13574 30810 13626
rect 30810 13574 30820 13626
rect 30844 13574 30874 13626
rect 30874 13574 30886 13626
rect 30886 13574 30900 13626
rect 30924 13574 30938 13626
rect 30938 13574 30950 13626
rect 30950 13574 30980 13626
rect 31004 13574 31014 13626
rect 31014 13574 31060 13626
rect 30764 13572 30820 13574
rect 30844 13572 30900 13574
rect 30924 13572 30980 13574
rect 31004 13572 31060 13574
rect 30764 12538 30820 12540
rect 30844 12538 30900 12540
rect 30924 12538 30980 12540
rect 31004 12538 31060 12540
rect 30764 12486 30810 12538
rect 30810 12486 30820 12538
rect 30844 12486 30874 12538
rect 30874 12486 30886 12538
rect 30886 12486 30900 12538
rect 30924 12486 30938 12538
rect 30938 12486 30950 12538
rect 30950 12486 30980 12538
rect 31004 12486 31014 12538
rect 31014 12486 31060 12538
rect 30764 12484 30820 12486
rect 30844 12484 30900 12486
rect 30924 12484 30980 12486
rect 31004 12484 31060 12486
rect 30286 11736 30342 11792
rect 30378 11600 30434 11656
rect 29182 1808 29238 1864
rect 31298 18672 31354 18728
rect 31390 15952 31446 16008
rect 31298 13368 31354 13424
rect 30764 11450 30820 11452
rect 30844 11450 30900 11452
rect 30924 11450 30980 11452
rect 31004 11450 31060 11452
rect 30764 11398 30810 11450
rect 30810 11398 30820 11450
rect 30844 11398 30874 11450
rect 30874 11398 30886 11450
rect 30886 11398 30900 11450
rect 30924 11398 30938 11450
rect 30938 11398 30950 11450
rect 30950 11398 30980 11450
rect 31004 11398 31014 11450
rect 31014 11398 31060 11450
rect 30764 11396 30820 11398
rect 30844 11396 30900 11398
rect 30924 11396 30980 11398
rect 31004 11396 31060 11398
rect 30764 10362 30820 10364
rect 30844 10362 30900 10364
rect 30924 10362 30980 10364
rect 31004 10362 31060 10364
rect 30764 10310 30810 10362
rect 30810 10310 30820 10362
rect 30844 10310 30874 10362
rect 30874 10310 30886 10362
rect 30886 10310 30900 10362
rect 30924 10310 30938 10362
rect 30938 10310 30950 10362
rect 30950 10310 30980 10362
rect 31004 10310 31014 10362
rect 31014 10310 31060 10362
rect 30764 10308 30820 10310
rect 30844 10308 30900 10310
rect 30924 10308 30980 10310
rect 31004 10308 31060 10310
rect 30764 9274 30820 9276
rect 30844 9274 30900 9276
rect 30924 9274 30980 9276
rect 31004 9274 31060 9276
rect 30764 9222 30810 9274
rect 30810 9222 30820 9274
rect 30844 9222 30874 9274
rect 30874 9222 30886 9274
rect 30886 9222 30900 9274
rect 30924 9222 30938 9274
rect 30938 9222 30950 9274
rect 30950 9222 30980 9274
rect 31004 9222 31014 9274
rect 31014 9222 31060 9274
rect 30764 9220 30820 9222
rect 30844 9220 30900 9222
rect 30924 9220 30980 9222
rect 31004 9220 31060 9222
rect 30764 8186 30820 8188
rect 30844 8186 30900 8188
rect 30924 8186 30980 8188
rect 31004 8186 31060 8188
rect 30764 8134 30810 8186
rect 30810 8134 30820 8186
rect 30844 8134 30874 8186
rect 30874 8134 30886 8186
rect 30886 8134 30900 8186
rect 30924 8134 30938 8186
rect 30938 8134 30950 8186
rect 30950 8134 30980 8186
rect 31004 8134 31014 8186
rect 31014 8134 31060 8186
rect 30764 8132 30820 8134
rect 30844 8132 30900 8134
rect 30924 8132 30980 8134
rect 31004 8132 31060 8134
rect 30764 7098 30820 7100
rect 30844 7098 30900 7100
rect 30924 7098 30980 7100
rect 31004 7098 31060 7100
rect 30764 7046 30810 7098
rect 30810 7046 30820 7098
rect 30844 7046 30874 7098
rect 30874 7046 30886 7098
rect 30886 7046 30900 7098
rect 30924 7046 30938 7098
rect 30938 7046 30950 7098
rect 30950 7046 30980 7098
rect 31004 7046 31014 7098
rect 31014 7046 31060 7098
rect 30764 7044 30820 7046
rect 30844 7044 30900 7046
rect 30924 7044 30980 7046
rect 31004 7044 31060 7046
rect 30764 6010 30820 6012
rect 30844 6010 30900 6012
rect 30924 6010 30980 6012
rect 31004 6010 31060 6012
rect 30764 5958 30810 6010
rect 30810 5958 30820 6010
rect 30844 5958 30874 6010
rect 30874 5958 30886 6010
rect 30886 5958 30900 6010
rect 30924 5958 30938 6010
rect 30938 5958 30950 6010
rect 30950 5958 30980 6010
rect 31004 5958 31014 6010
rect 31014 5958 31060 6010
rect 30764 5956 30820 5958
rect 30844 5956 30900 5958
rect 30924 5956 30980 5958
rect 31004 5956 31060 5958
rect 30764 4922 30820 4924
rect 30844 4922 30900 4924
rect 30924 4922 30980 4924
rect 31004 4922 31060 4924
rect 30764 4870 30810 4922
rect 30810 4870 30820 4922
rect 30844 4870 30874 4922
rect 30874 4870 30886 4922
rect 30886 4870 30900 4922
rect 30924 4870 30938 4922
rect 30938 4870 30950 4922
rect 30950 4870 30980 4922
rect 31004 4870 31014 4922
rect 31014 4870 31060 4922
rect 30764 4868 30820 4870
rect 30844 4868 30900 4870
rect 30924 4868 30980 4870
rect 31004 4868 31060 4870
rect 30764 3834 30820 3836
rect 30844 3834 30900 3836
rect 30924 3834 30980 3836
rect 31004 3834 31060 3836
rect 30764 3782 30810 3834
rect 30810 3782 30820 3834
rect 30844 3782 30874 3834
rect 30874 3782 30886 3834
rect 30886 3782 30900 3834
rect 30924 3782 30938 3834
rect 30938 3782 30950 3834
rect 30950 3782 30980 3834
rect 31004 3782 31014 3834
rect 31014 3782 31060 3834
rect 30764 3780 30820 3782
rect 30844 3780 30900 3782
rect 30924 3780 30980 3782
rect 31004 3780 31060 3782
rect 30764 2746 30820 2748
rect 30844 2746 30900 2748
rect 30924 2746 30980 2748
rect 31004 2746 31060 2748
rect 30764 2694 30810 2746
rect 30810 2694 30820 2746
rect 30844 2694 30874 2746
rect 30874 2694 30886 2746
rect 30886 2694 30900 2746
rect 30924 2694 30938 2746
rect 30938 2694 30950 2746
rect 30950 2694 30980 2746
rect 31004 2694 31014 2746
rect 31014 2694 31060 2746
rect 30764 2692 30820 2694
rect 30844 2692 30900 2694
rect 30924 2692 30980 2694
rect 31004 2692 31060 2694
rect 30764 1658 30820 1660
rect 30844 1658 30900 1660
rect 30924 1658 30980 1660
rect 31004 1658 31060 1660
rect 30764 1606 30810 1658
rect 30810 1606 30820 1658
rect 30844 1606 30874 1658
rect 30874 1606 30886 1658
rect 30886 1606 30900 1658
rect 30924 1606 30938 1658
rect 30938 1606 30950 1658
rect 30950 1606 30980 1658
rect 31004 1606 31014 1658
rect 31014 1606 31060 1658
rect 30764 1604 30820 1606
rect 30844 1604 30900 1606
rect 30924 1604 30980 1606
rect 31004 1604 31060 1606
rect 30764 570 30820 572
rect 30844 570 30900 572
rect 30924 570 30980 572
rect 31004 570 31060 572
rect 30764 518 30810 570
rect 30810 518 30820 570
rect 30844 518 30874 570
rect 30874 518 30886 570
rect 30886 518 30900 570
rect 30924 518 30938 570
rect 30938 518 30950 570
rect 30950 518 30980 570
rect 31004 518 31014 570
rect 31014 518 31060 570
rect 30764 516 30820 518
rect 30844 516 30900 518
rect 30924 516 30980 518
rect 31004 516 31060 518
rect 25318 312 25374 368
<< metal3 >>
rect 10726 22204 10732 22268
rect 10796 22266 10802 22268
rect 10961 22266 11027 22269
rect 10796 22264 11027 22266
rect 10796 22208 10966 22264
rect 11022 22208 11027 22264
rect 10796 22206 11027 22208
rect 10796 22204 10802 22206
rect 10961 22203 11027 22206
rect 12198 21796 12204 21860
rect 12268 21858 12274 21860
rect 12525 21858 12591 21861
rect 12268 21856 12591 21858
rect 12268 21800 12530 21856
rect 12586 21800 12591 21856
rect 12268 21798 12591 21800
rect 12268 21796 12274 21798
rect 12525 21795 12591 21798
rect 4189 21792 4505 21793
rect 4189 21728 4195 21792
rect 4259 21728 4275 21792
rect 4339 21728 4355 21792
rect 4419 21728 4435 21792
rect 4499 21728 4505 21792
rect 4189 21727 4505 21728
rect 11779 21792 12095 21793
rect 11779 21728 11785 21792
rect 11849 21728 11865 21792
rect 11929 21728 11945 21792
rect 12009 21728 12025 21792
rect 12089 21728 12095 21792
rect 11779 21727 12095 21728
rect 19369 21792 19685 21793
rect 19369 21728 19375 21792
rect 19439 21728 19455 21792
rect 19519 21728 19535 21792
rect 19599 21728 19615 21792
rect 19679 21728 19685 21792
rect 19369 21727 19685 21728
rect 26959 21792 27275 21793
rect 26959 21728 26965 21792
rect 27029 21728 27045 21792
rect 27109 21728 27125 21792
rect 27189 21728 27205 21792
rect 27269 21728 27275 21792
rect 26959 21727 27275 21728
rect 13670 21524 13676 21588
rect 13740 21586 13746 21588
rect 13997 21586 14063 21589
rect 13740 21584 14063 21586
rect 13740 21528 14002 21584
rect 14058 21528 14063 21584
rect 13740 21526 14063 21528
rect 13740 21524 13746 21526
rect 13997 21523 14063 21526
rect 16982 21524 16988 21588
rect 17052 21586 17058 21588
rect 17125 21586 17191 21589
rect 25446 21586 25452 21588
rect 17052 21584 17191 21586
rect 17052 21528 17130 21584
rect 17186 21528 17191 21584
rect 17052 21526 17191 21528
rect 17052 21524 17058 21526
rect 17125 21523 17191 21526
rect 17358 21526 25452 21586
rect 5901 21450 5967 21453
rect 9397 21450 9463 21453
rect 5901 21448 9463 21450
rect 5901 21392 5906 21448
rect 5962 21392 9402 21448
rect 9458 21392 9463 21448
rect 5901 21390 9463 21392
rect 5901 21387 5967 21390
rect 9397 21387 9463 21390
rect 13670 21388 13676 21452
rect 13740 21450 13746 21452
rect 14181 21450 14247 21453
rect 13740 21448 14247 21450
rect 13740 21392 14186 21448
rect 14242 21392 14247 21448
rect 13740 21390 14247 21392
rect 13740 21388 13746 21390
rect 14181 21387 14247 21390
rect 16665 21450 16731 21453
rect 17358 21450 17418 21526
rect 25446 21524 25452 21526
rect 25516 21524 25522 21588
rect 16665 21448 17418 21450
rect 16665 21392 16670 21448
rect 16726 21392 17418 21448
rect 16665 21390 17418 21392
rect 18505 21450 18571 21453
rect 28758 21450 28764 21452
rect 18505 21448 28764 21450
rect 18505 21392 18510 21448
rect 18566 21392 28764 21448
rect 18505 21390 28764 21392
rect 16665 21387 16731 21390
rect 18505 21387 18571 21390
rect 28758 21388 28764 21390
rect 28828 21388 28834 21452
rect 7984 21248 8300 21249
rect 7984 21184 7990 21248
rect 8054 21184 8070 21248
rect 8134 21184 8150 21248
rect 8214 21184 8230 21248
rect 8294 21184 8300 21248
rect 7984 21183 8300 21184
rect 15574 21248 15890 21249
rect 15574 21184 15580 21248
rect 15644 21184 15660 21248
rect 15724 21184 15740 21248
rect 15804 21184 15820 21248
rect 15884 21184 15890 21248
rect 15574 21183 15890 21184
rect 23164 21248 23480 21249
rect 23164 21184 23170 21248
rect 23234 21184 23250 21248
rect 23314 21184 23330 21248
rect 23394 21184 23410 21248
rect 23474 21184 23480 21248
rect 23164 21183 23480 21184
rect 30754 21248 31070 21249
rect 30754 21184 30760 21248
rect 30824 21184 30840 21248
rect 30904 21184 30920 21248
rect 30984 21184 31000 21248
rect 31064 21184 31070 21248
rect 30754 21183 31070 21184
rect 25129 21178 25195 21181
rect 26366 21178 26372 21180
rect 25129 21176 26372 21178
rect 25129 21120 25134 21176
rect 25190 21120 26372 21176
rect 25129 21118 26372 21120
rect 25129 21115 25195 21118
rect 26366 21116 26372 21118
rect 26436 21116 26442 21180
rect 1669 21042 1735 21045
rect 8937 21042 9003 21045
rect 11278 21042 11284 21044
rect 1669 21040 2790 21042
rect 1669 20984 1674 21040
rect 1730 20984 2790 21040
rect 1669 20982 2790 20984
rect 1669 20979 1735 20982
rect 2730 20906 2790 20982
rect 8937 21040 11284 21042
rect 8937 20984 8942 21040
rect 8998 20984 11284 21040
rect 8937 20982 11284 20984
rect 8937 20979 9003 20982
rect 11278 20980 11284 20982
rect 11348 20980 11354 21044
rect 15101 21042 15167 21045
rect 16573 21042 16639 21045
rect 15101 21040 16639 21042
rect 15101 20984 15106 21040
rect 15162 20984 16578 21040
rect 16634 20984 16639 21040
rect 15101 20982 16639 20984
rect 15101 20979 15167 20982
rect 16573 20979 16639 20982
rect 17861 21042 17927 21045
rect 24894 21042 24900 21044
rect 17861 21040 24900 21042
rect 17861 20984 17866 21040
rect 17922 20984 24900 21040
rect 17861 20982 24900 20984
rect 17861 20979 17927 20982
rect 24894 20980 24900 20982
rect 24964 20980 24970 21044
rect 10869 20906 10935 20909
rect 11462 20906 11468 20908
rect 2730 20846 10242 20906
rect 2957 20770 3023 20773
rect 3918 20770 3924 20772
rect 2957 20768 3924 20770
rect 2957 20712 2962 20768
rect 3018 20712 3924 20768
rect 2957 20710 3924 20712
rect 2957 20707 3023 20710
rect 3918 20708 3924 20710
rect 3988 20708 3994 20772
rect 6729 20770 6795 20773
rect 10182 20772 10242 20846
rect 10869 20904 11468 20906
rect 10869 20848 10874 20904
rect 10930 20848 11468 20904
rect 10869 20846 11468 20848
rect 10869 20843 10935 20846
rect 11462 20844 11468 20846
rect 11532 20844 11538 20908
rect 8886 20770 8892 20772
rect 6729 20768 8892 20770
rect 6729 20712 6734 20768
rect 6790 20712 8892 20768
rect 6729 20710 8892 20712
rect 6729 20707 6795 20710
rect 8886 20708 8892 20710
rect 8956 20708 8962 20772
rect 10174 20708 10180 20772
rect 10244 20708 10250 20772
rect 4189 20704 4505 20705
rect 4189 20640 4195 20704
rect 4259 20640 4275 20704
rect 4339 20640 4355 20704
rect 4419 20640 4435 20704
rect 4499 20640 4505 20704
rect 4189 20639 4505 20640
rect 11779 20704 12095 20705
rect 11779 20640 11785 20704
rect 11849 20640 11865 20704
rect 11929 20640 11945 20704
rect 12009 20640 12025 20704
rect 12089 20640 12095 20704
rect 11779 20639 12095 20640
rect 19369 20704 19685 20705
rect 19369 20640 19375 20704
rect 19439 20640 19455 20704
rect 19519 20640 19535 20704
rect 19599 20640 19615 20704
rect 19679 20640 19685 20704
rect 19369 20639 19685 20640
rect 26959 20704 27275 20705
rect 26959 20640 26965 20704
rect 27029 20640 27045 20704
rect 27109 20640 27125 20704
rect 27189 20640 27205 20704
rect 27269 20640 27275 20704
rect 26959 20639 27275 20640
rect 7598 20572 7604 20636
rect 7668 20634 7674 20636
rect 8937 20634 9003 20637
rect 7668 20632 9003 20634
rect 7668 20576 8942 20632
rect 8998 20576 9003 20632
rect 7668 20574 9003 20576
rect 7668 20572 7674 20574
rect 8937 20571 9003 20574
rect 13721 20634 13787 20637
rect 15142 20634 15148 20636
rect 13721 20632 15148 20634
rect 13721 20576 13726 20632
rect 13782 20576 15148 20632
rect 13721 20574 15148 20576
rect 13721 20571 13787 20574
rect 15142 20572 15148 20574
rect 15212 20572 15218 20636
rect 23606 20634 23612 20636
rect 22050 20574 23612 20634
rect 1669 20498 1735 20501
rect 11421 20498 11487 20501
rect 1669 20496 11487 20498
rect 1669 20440 1674 20496
rect 1730 20440 11426 20496
rect 11482 20440 11487 20496
rect 1669 20438 11487 20440
rect 1669 20435 1735 20438
rect 11421 20435 11487 20438
rect 18689 20498 18755 20501
rect 22050 20498 22110 20574
rect 23606 20572 23612 20574
rect 23676 20634 23682 20636
rect 26049 20634 26115 20637
rect 23676 20632 26115 20634
rect 23676 20576 26054 20632
rect 26110 20576 26115 20632
rect 23676 20574 26115 20576
rect 23676 20572 23682 20574
rect 26049 20571 26115 20574
rect 18689 20496 22110 20498
rect 18689 20440 18694 20496
rect 18750 20440 22110 20496
rect 18689 20438 22110 20440
rect 24393 20498 24459 20501
rect 27654 20498 27660 20500
rect 24393 20496 27660 20498
rect 24393 20440 24398 20496
rect 24454 20440 27660 20496
rect 24393 20438 27660 20440
rect 18689 20435 18755 20438
rect 24393 20435 24459 20438
rect 27654 20436 27660 20438
rect 27724 20436 27730 20500
rect 5441 20362 5507 20365
rect 7557 20362 7623 20365
rect 5441 20360 7623 20362
rect 5441 20304 5446 20360
rect 5502 20304 7562 20360
rect 7618 20304 7623 20360
rect 5441 20302 7623 20304
rect 5441 20299 5507 20302
rect 7557 20299 7623 20302
rect 7833 20362 7899 20365
rect 8845 20362 8911 20365
rect 7833 20360 8911 20362
rect 7833 20304 7838 20360
rect 7894 20304 8850 20360
rect 8906 20304 8911 20360
rect 7833 20302 8911 20304
rect 7833 20299 7899 20302
rect 8845 20299 8911 20302
rect 24209 20226 24275 20229
rect 25589 20226 25655 20229
rect 24209 20224 25655 20226
rect 24209 20168 24214 20224
rect 24270 20168 25594 20224
rect 25650 20168 25655 20224
rect 24209 20166 25655 20168
rect 24209 20163 24275 20166
rect 25589 20163 25655 20166
rect 7984 20160 8300 20161
rect 7984 20096 7990 20160
rect 8054 20096 8070 20160
rect 8134 20096 8150 20160
rect 8214 20096 8230 20160
rect 8294 20096 8300 20160
rect 7984 20095 8300 20096
rect 15574 20160 15890 20161
rect 15574 20096 15580 20160
rect 15644 20096 15660 20160
rect 15724 20096 15740 20160
rect 15804 20096 15820 20160
rect 15884 20096 15890 20160
rect 15574 20095 15890 20096
rect 23164 20160 23480 20161
rect 23164 20096 23170 20160
rect 23234 20096 23250 20160
rect 23314 20096 23330 20160
rect 23394 20096 23410 20160
rect 23474 20096 23480 20160
rect 23164 20095 23480 20096
rect 30754 20160 31070 20161
rect 30754 20096 30760 20160
rect 30824 20096 30840 20160
rect 30904 20096 30920 20160
rect 30984 20096 31000 20160
rect 31064 20096 31070 20160
rect 30754 20095 31070 20096
rect 24669 20090 24735 20093
rect 28533 20090 28599 20093
rect 24669 20088 28599 20090
rect 24669 20032 24674 20088
rect 24730 20032 28538 20088
rect 28594 20032 28599 20088
rect 24669 20030 28599 20032
rect 24669 20027 24735 20030
rect 28533 20027 28599 20030
rect 6177 19954 6243 19957
rect 6913 19954 6979 19957
rect 6177 19952 6979 19954
rect 6177 19896 6182 19952
rect 6238 19896 6918 19952
rect 6974 19896 6979 19952
rect 6177 19894 6979 19896
rect 6177 19891 6243 19894
rect 6913 19891 6979 19894
rect 20989 19954 21055 19957
rect 21817 19954 21883 19957
rect 20989 19952 21883 19954
rect 20989 19896 20994 19952
rect 21050 19896 21822 19952
rect 21878 19896 21883 19952
rect 20989 19894 21883 19896
rect 20989 19891 21055 19894
rect 21817 19891 21883 19894
rect 21950 19892 21956 19956
rect 22020 19954 22026 19956
rect 28349 19954 28415 19957
rect 22020 19952 28415 19954
rect 22020 19896 28354 19952
rect 28410 19896 28415 19952
rect 22020 19894 28415 19896
rect 22020 19892 22026 19894
rect 28349 19891 28415 19894
rect 3601 19818 3667 19821
rect 11237 19818 11303 19821
rect 3601 19816 11303 19818
rect 3601 19760 3606 19816
rect 3662 19760 11242 19816
rect 11298 19760 11303 19816
rect 3601 19758 11303 19760
rect 3601 19755 3667 19758
rect 11237 19755 11303 19758
rect 21265 19818 21331 19821
rect 23841 19818 23907 19821
rect 21265 19816 23907 19818
rect 21265 19760 21270 19816
rect 21326 19760 23846 19816
rect 23902 19760 23907 19816
rect 21265 19758 23907 19760
rect 21265 19755 21331 19758
rect 23841 19755 23907 19758
rect 4189 19616 4505 19617
rect 4189 19552 4195 19616
rect 4259 19552 4275 19616
rect 4339 19552 4355 19616
rect 4419 19552 4435 19616
rect 4499 19552 4505 19616
rect 4189 19551 4505 19552
rect 11779 19616 12095 19617
rect 11779 19552 11785 19616
rect 11849 19552 11865 19616
rect 11929 19552 11945 19616
rect 12009 19552 12025 19616
rect 12089 19552 12095 19616
rect 11779 19551 12095 19552
rect 19369 19616 19685 19617
rect 19369 19552 19375 19616
rect 19439 19552 19455 19616
rect 19519 19552 19535 19616
rect 19599 19552 19615 19616
rect 19679 19552 19685 19616
rect 19369 19551 19685 19552
rect 26959 19616 27275 19617
rect 26959 19552 26965 19616
rect 27029 19552 27045 19616
rect 27109 19552 27125 19616
rect 27189 19552 27205 19616
rect 27269 19552 27275 19616
rect 26959 19551 27275 19552
rect 6269 19546 6335 19549
rect 5398 19544 6335 19546
rect 5398 19488 6274 19544
rect 6330 19488 6335 19544
rect 5398 19486 6335 19488
rect 1669 19410 1735 19413
rect 5398 19410 5458 19486
rect 6269 19483 6335 19486
rect 1669 19408 5458 19410
rect 1669 19352 1674 19408
rect 1730 19352 5458 19408
rect 1669 19350 5458 19352
rect 5625 19410 5691 19413
rect 6913 19410 6979 19413
rect 5625 19408 6979 19410
rect 5625 19352 5630 19408
rect 5686 19352 6918 19408
rect 6974 19352 6979 19408
rect 5625 19350 6979 19352
rect 1669 19347 1735 19350
rect 5625 19347 5691 19350
rect 6913 19347 6979 19350
rect 9213 19410 9279 19413
rect 11462 19410 11468 19412
rect 9213 19408 11468 19410
rect 9213 19352 9218 19408
rect 9274 19352 11468 19408
rect 9213 19350 11468 19352
rect 9213 19347 9279 19350
rect 11462 19348 11468 19350
rect 11532 19348 11538 19412
rect 14457 19410 14523 19413
rect 16665 19410 16731 19413
rect 14457 19408 17786 19410
rect 14457 19352 14462 19408
rect 14518 19352 16670 19408
rect 16726 19352 17786 19408
rect 14457 19350 17786 19352
rect 14457 19347 14523 19350
rect 16665 19347 16731 19350
rect 17677 19348 17786 19350
rect 26550 19348 26556 19412
rect 26620 19410 26626 19412
rect 29545 19410 29611 19413
rect 26620 19408 29611 19410
rect 26620 19352 29550 19408
rect 29606 19352 29611 19408
rect 26620 19350 29611 19352
rect 26620 19348 26626 19350
rect 17677 19292 17682 19348
rect 17738 19292 17786 19348
rect 29545 19347 29611 19350
rect 17677 19290 17786 19292
rect 17677 19287 17743 19290
rect 9673 19274 9739 19277
rect 10910 19274 10916 19276
rect 2730 19214 9506 19274
rect 1393 18730 1459 18733
rect 2730 18730 2790 19214
rect 3877 19138 3943 19141
rect 7833 19138 7899 19141
rect 3877 19136 7899 19138
rect 3877 19080 3882 19136
rect 3938 19080 7838 19136
rect 7894 19080 7899 19136
rect 3877 19078 7899 19080
rect 3877 19075 3943 19078
rect 7833 19075 7899 19078
rect 8477 19138 8543 19141
rect 8702 19138 8708 19140
rect 8477 19136 8708 19138
rect 8477 19080 8482 19136
rect 8538 19080 8708 19136
rect 8477 19078 8708 19080
rect 8477 19075 8543 19078
rect 8702 19076 8708 19078
rect 8772 19076 8778 19140
rect 9446 19138 9506 19214
rect 9673 19272 10916 19274
rect 9673 19216 9678 19272
rect 9734 19216 10916 19272
rect 9673 19214 10916 19216
rect 9673 19211 9739 19214
rect 10910 19212 10916 19214
rect 10980 19212 10986 19276
rect 12566 19212 12572 19276
rect 12636 19274 12642 19276
rect 13353 19274 13419 19277
rect 12636 19272 13419 19274
rect 12636 19216 13358 19272
rect 13414 19216 13419 19272
rect 12636 19214 13419 19216
rect 12636 19212 12642 19214
rect 13353 19211 13419 19214
rect 14774 19212 14780 19276
rect 14844 19274 14850 19276
rect 15101 19274 15167 19277
rect 14844 19272 15167 19274
rect 14844 19216 15106 19272
rect 15162 19216 15167 19272
rect 14844 19214 15167 19216
rect 14844 19212 14850 19214
rect 15101 19211 15167 19214
rect 16062 19212 16068 19276
rect 16132 19274 16138 19276
rect 16297 19274 16363 19277
rect 16481 19276 16547 19277
rect 16132 19272 16363 19274
rect 16132 19216 16302 19272
rect 16358 19216 16363 19272
rect 16132 19214 16363 19216
rect 16132 19212 16138 19214
rect 16297 19211 16363 19214
rect 16430 19212 16436 19276
rect 16500 19274 16547 19276
rect 23565 19274 23631 19277
rect 24710 19274 24716 19276
rect 16500 19272 16592 19274
rect 16542 19216 16592 19272
rect 16500 19214 16592 19216
rect 23565 19272 24716 19274
rect 23565 19216 23570 19272
rect 23626 19216 24716 19272
rect 23565 19214 24716 19216
rect 16500 19212 16547 19214
rect 16481 19211 16547 19212
rect 23565 19211 23631 19214
rect 24710 19212 24716 19214
rect 24780 19212 24786 19276
rect 9673 19138 9739 19141
rect 9857 19140 9923 19141
rect 9446 19136 9739 19138
rect 9446 19080 9678 19136
rect 9734 19080 9739 19136
rect 9446 19078 9739 19080
rect 9673 19075 9739 19078
rect 9806 19076 9812 19140
rect 9876 19138 9923 19140
rect 9876 19136 9968 19138
rect 9918 19080 9968 19136
rect 9876 19078 9968 19080
rect 9876 19076 9923 19078
rect 9857 19075 9923 19076
rect 7984 19072 8300 19073
rect 7984 19008 7990 19072
rect 8054 19008 8070 19072
rect 8134 19008 8150 19072
rect 8214 19008 8230 19072
rect 8294 19008 8300 19072
rect 7984 19007 8300 19008
rect 15574 19072 15890 19073
rect 15574 19008 15580 19072
rect 15644 19008 15660 19072
rect 15724 19008 15740 19072
rect 15804 19008 15820 19072
rect 15884 19008 15890 19072
rect 15574 19007 15890 19008
rect 23164 19072 23480 19073
rect 23164 19008 23170 19072
rect 23234 19008 23250 19072
rect 23314 19008 23330 19072
rect 23394 19008 23410 19072
rect 23474 19008 23480 19072
rect 23164 19007 23480 19008
rect 30754 19072 31070 19073
rect 30754 19008 30760 19072
rect 30824 19008 30840 19072
rect 30904 19008 30920 19072
rect 30984 19008 31000 19072
rect 31064 19008 31070 19072
rect 30754 19007 31070 19008
rect 6453 19002 6519 19005
rect 7557 19002 7623 19005
rect 6453 19000 7623 19002
rect 6453 18944 6458 19000
rect 6514 18944 7562 19000
rect 7618 18944 7623 19000
rect 6453 18942 7623 18944
rect 6453 18939 6519 18942
rect 7557 18939 7623 18942
rect 24577 19002 24643 19005
rect 26509 19002 26575 19005
rect 24577 19000 26575 19002
rect 24577 18944 24582 19000
rect 24638 18944 26514 19000
rect 26570 18944 26575 19000
rect 24577 18942 26575 18944
rect 24577 18939 24643 18942
rect 26509 18939 26575 18942
rect 5073 18866 5139 18869
rect 9254 18866 9260 18868
rect 5073 18864 9260 18866
rect 5073 18808 5078 18864
rect 5134 18808 9260 18864
rect 5073 18806 9260 18808
rect 5073 18803 5139 18806
rect 9254 18804 9260 18806
rect 9324 18804 9330 18868
rect 14549 18866 14615 18869
rect 23974 18866 23980 18868
rect 14549 18864 23980 18866
rect 14549 18808 14554 18864
rect 14610 18808 23980 18864
rect 14549 18806 23980 18808
rect 14549 18803 14615 18806
rect 23974 18804 23980 18806
rect 24044 18804 24050 18868
rect 24117 18866 24183 18869
rect 25681 18866 25747 18869
rect 26693 18866 26759 18869
rect 24117 18864 26759 18866
rect 24117 18808 24122 18864
rect 24178 18808 25686 18864
rect 25742 18808 26698 18864
rect 26754 18808 26759 18864
rect 24117 18806 26759 18808
rect 24117 18803 24183 18806
rect 25681 18803 25747 18806
rect 26693 18803 26759 18806
rect 27153 18866 27219 18869
rect 28073 18866 28139 18869
rect 27153 18864 28139 18866
rect 27153 18808 27158 18864
rect 27214 18808 28078 18864
rect 28134 18808 28139 18864
rect 27153 18806 28139 18808
rect 27153 18803 27219 18806
rect 28073 18803 28139 18806
rect 5441 18732 5507 18733
rect 5390 18730 5396 18732
rect 1393 18728 2790 18730
rect 1393 18672 1398 18728
rect 1454 18672 2790 18728
rect 1393 18670 2790 18672
rect 5350 18670 5396 18730
rect 5460 18728 5507 18732
rect 5502 18672 5507 18728
rect 1393 18667 1459 18670
rect 5390 18668 5396 18670
rect 5460 18668 5507 18672
rect 5441 18667 5507 18668
rect 7833 18730 7899 18733
rect 8702 18730 8708 18732
rect 7833 18728 8708 18730
rect 7833 18672 7838 18728
rect 7894 18672 8708 18728
rect 7833 18670 8708 18672
rect 7833 18667 7899 18670
rect 8702 18668 8708 18670
rect 8772 18730 8778 18732
rect 10409 18730 10475 18733
rect 8772 18728 10475 18730
rect 8772 18672 10414 18728
rect 10470 18672 10475 18728
rect 8772 18670 10475 18672
rect 8772 18668 8778 18670
rect 10409 18667 10475 18670
rect 11789 18730 11855 18733
rect 12341 18730 12407 18733
rect 29729 18730 29795 18733
rect 31293 18730 31359 18733
rect 11789 18728 12407 18730
rect 11789 18672 11794 18728
rect 11850 18672 12346 18728
rect 12402 18672 12407 18728
rect 11789 18670 12407 18672
rect 11789 18667 11855 18670
rect 12341 18667 12407 18670
rect 24534 18728 31359 18730
rect 24534 18672 29734 18728
rect 29790 18672 31298 18728
rect 31354 18672 31359 18728
rect 24534 18670 31359 18672
rect 8569 18594 8635 18597
rect 8937 18594 9003 18597
rect 24393 18594 24459 18597
rect 24534 18594 24594 18670
rect 29729 18667 29795 18670
rect 31293 18667 31359 18670
rect 8569 18592 9003 18594
rect 8569 18536 8574 18592
rect 8630 18536 8942 18592
rect 8998 18536 9003 18592
rect 8569 18534 9003 18536
rect 8569 18531 8635 18534
rect 8937 18531 9003 18534
rect 22050 18592 24594 18594
rect 22050 18536 24398 18592
rect 24454 18536 24594 18592
rect 22050 18534 24594 18536
rect 4189 18528 4505 18529
rect 4189 18464 4195 18528
rect 4259 18464 4275 18528
rect 4339 18464 4355 18528
rect 4419 18464 4435 18528
rect 4499 18464 4505 18528
rect 4189 18463 4505 18464
rect 11779 18528 12095 18529
rect 11779 18464 11785 18528
rect 11849 18464 11865 18528
rect 11929 18464 11945 18528
rect 12009 18464 12025 18528
rect 12089 18464 12095 18528
rect 11779 18463 12095 18464
rect 19369 18528 19685 18529
rect 19369 18464 19375 18528
rect 19439 18464 19455 18528
rect 19519 18464 19535 18528
rect 19599 18464 19615 18528
rect 19679 18464 19685 18528
rect 19369 18463 19685 18464
rect 22050 18461 22110 18534
rect 24393 18531 24459 18534
rect 26959 18528 27275 18529
rect 26959 18464 26965 18528
rect 27029 18464 27045 18528
rect 27109 18464 27125 18528
rect 27189 18464 27205 18528
rect 27269 18464 27275 18528
rect 26959 18463 27275 18464
rect 4613 18460 4679 18461
rect 4613 18456 4660 18460
rect 4724 18458 4730 18460
rect 4613 18400 4618 18456
rect 4613 18396 4660 18400
rect 4724 18398 4770 18458
rect 4724 18396 4730 18398
rect 5206 18396 5212 18460
rect 5276 18458 5282 18460
rect 10542 18458 10548 18460
rect 5276 18398 10548 18458
rect 5276 18396 5282 18398
rect 10542 18396 10548 18398
rect 10612 18396 10618 18460
rect 22001 18456 22110 18461
rect 22001 18400 22006 18456
rect 22062 18400 22110 18456
rect 22001 18398 22110 18400
rect 4613 18395 4679 18396
rect 22001 18395 22067 18398
rect 7046 18260 7052 18324
rect 7116 18322 7122 18324
rect 8201 18322 8267 18325
rect 7116 18320 8267 18322
rect 7116 18264 8206 18320
rect 8262 18264 8267 18320
rect 7116 18262 8267 18264
rect 7116 18260 7122 18262
rect 8201 18259 8267 18262
rect 8477 18322 8543 18325
rect 8937 18322 9003 18325
rect 8477 18320 9003 18322
rect 8477 18264 8482 18320
rect 8538 18264 8942 18320
rect 8998 18264 9003 18320
rect 8477 18262 9003 18264
rect 8477 18259 8543 18262
rect 8937 18259 9003 18262
rect 23841 18322 23907 18325
rect 30097 18322 30163 18325
rect 23841 18320 30163 18322
rect 23841 18264 23846 18320
rect 23902 18264 30102 18320
rect 30158 18264 30163 18320
rect 23841 18262 30163 18264
rect 23841 18259 23907 18262
rect 30097 18259 30163 18262
rect 1301 18186 1367 18189
rect 5349 18186 5415 18189
rect 1301 18184 5415 18186
rect 1301 18128 1306 18184
rect 1362 18128 5354 18184
rect 5410 18128 5415 18184
rect 1301 18126 5415 18128
rect 1301 18123 1367 18126
rect 5349 18123 5415 18126
rect 6494 18124 6500 18188
rect 6564 18186 6570 18188
rect 8937 18186 9003 18189
rect 6564 18184 9003 18186
rect 6564 18128 8942 18184
rect 8998 18128 9003 18184
rect 6564 18126 9003 18128
rect 6564 18124 6570 18126
rect 8937 18123 9003 18126
rect 10961 18186 11027 18189
rect 16297 18186 16363 18189
rect 10961 18184 16363 18186
rect 10961 18128 10966 18184
rect 11022 18128 16302 18184
rect 16358 18128 16363 18184
rect 10961 18126 16363 18128
rect 10961 18123 11027 18126
rect 16297 18123 16363 18126
rect 22921 18186 22987 18189
rect 23933 18186 23999 18189
rect 24158 18186 24164 18188
rect 22921 18184 23858 18186
rect 22921 18128 22926 18184
rect 22982 18128 23858 18184
rect 22921 18126 23858 18128
rect 22921 18123 22987 18126
rect 4613 18050 4679 18053
rect 6729 18052 6795 18053
rect 5390 18050 5396 18052
rect 4613 18048 5396 18050
rect 4613 17992 4618 18048
rect 4674 17992 5396 18048
rect 4613 17990 5396 17992
rect 4613 17987 4679 17990
rect 5390 17988 5396 17990
rect 5460 17988 5466 18052
rect 6678 18050 6684 18052
rect 6638 17990 6684 18050
rect 6748 18048 6795 18052
rect 6790 17992 6795 18048
rect 6678 17988 6684 17990
rect 6748 17988 6795 17992
rect 6729 17987 6795 17988
rect 10961 18050 11027 18053
rect 17033 18050 17099 18053
rect 19241 18050 19307 18053
rect 22553 18052 22619 18053
rect 22502 18050 22508 18052
rect 10961 18048 12266 18050
rect 10961 17992 10966 18048
rect 11022 17992 12266 18048
rect 10961 17990 12266 17992
rect 10961 17987 11027 17990
rect 7984 17984 8300 17985
rect 7984 17920 7990 17984
rect 8054 17920 8070 17984
rect 8134 17920 8150 17984
rect 8214 17920 8230 17984
rect 8294 17920 8300 17984
rect 7984 17919 8300 17920
rect 12206 17917 12266 17990
rect 17033 18048 19307 18050
rect 17033 17992 17038 18048
rect 17094 17992 19246 18048
rect 19302 17992 19307 18048
rect 17033 17990 19307 17992
rect 22462 17990 22508 18050
rect 22572 18048 22619 18052
rect 22614 17992 22619 18048
rect 17033 17987 17099 17990
rect 19241 17987 19307 17990
rect 22502 17988 22508 17990
rect 22572 17988 22619 17992
rect 22870 17988 22876 18052
rect 22940 18050 22946 18052
rect 23013 18050 23079 18053
rect 22940 18048 23079 18050
rect 22940 17992 23018 18048
rect 23074 17992 23079 18048
rect 22940 17990 23079 17992
rect 23798 18050 23858 18126
rect 23933 18184 24164 18186
rect 23933 18128 23938 18184
rect 23994 18128 24164 18184
rect 23933 18126 24164 18128
rect 23933 18123 23999 18126
rect 24158 18124 24164 18126
rect 24228 18124 24234 18188
rect 30649 18186 30715 18189
rect 24718 18184 30715 18186
rect 24718 18128 30654 18184
rect 30710 18128 30715 18184
rect 24718 18126 30715 18128
rect 24718 18050 24778 18126
rect 30649 18123 30715 18126
rect 23798 17990 24778 18050
rect 24853 18050 24919 18053
rect 30373 18050 30439 18053
rect 24853 18048 30439 18050
rect 24853 17992 24858 18048
rect 24914 17992 30378 18048
rect 30434 17992 30439 18048
rect 24853 17990 30439 17992
rect 22940 17988 22946 17990
rect 22553 17987 22619 17988
rect 23013 17987 23079 17990
rect 24853 17987 24919 17990
rect 30373 17987 30439 17990
rect 15574 17984 15890 17985
rect 15574 17920 15580 17984
rect 15644 17920 15660 17984
rect 15724 17920 15740 17984
rect 15804 17920 15820 17984
rect 15884 17920 15890 17984
rect 15574 17919 15890 17920
rect 23164 17984 23480 17985
rect 23164 17920 23170 17984
rect 23234 17920 23250 17984
rect 23314 17920 23330 17984
rect 23394 17920 23410 17984
rect 23474 17920 23480 17984
rect 23164 17919 23480 17920
rect 30754 17984 31070 17985
rect 30754 17920 30760 17984
rect 30824 17920 30840 17984
rect 30904 17920 30920 17984
rect 30984 17920 31000 17984
rect 31064 17920 31070 17984
rect 30754 17919 31070 17920
rect 12206 17912 12315 17917
rect 12206 17856 12254 17912
rect 12310 17856 12315 17912
rect 12206 17854 12315 17856
rect 12249 17851 12315 17854
rect 3785 17778 3851 17781
rect 16021 17778 16087 17781
rect 3785 17776 16087 17778
rect 3785 17720 3790 17776
rect 3846 17720 16026 17776
rect 16082 17720 16087 17776
rect 3785 17718 16087 17720
rect 3785 17715 3851 17718
rect 16021 17715 16087 17718
rect 21081 17778 21147 17781
rect 27153 17778 27219 17781
rect 21081 17776 27219 17778
rect 21081 17720 21086 17776
rect 21142 17720 27158 17776
rect 27214 17720 27219 17776
rect 21081 17718 27219 17720
rect 21081 17715 21147 17718
rect 27153 17715 27219 17718
rect 8753 17642 8819 17645
rect 18965 17642 19031 17645
rect 8753 17640 19031 17642
rect 8753 17584 8758 17640
rect 8814 17584 18970 17640
rect 19026 17584 19031 17640
rect 8753 17582 19031 17584
rect 8753 17579 8819 17582
rect 18965 17579 19031 17582
rect 21265 17642 21331 17645
rect 26693 17642 26759 17645
rect 21265 17640 26759 17642
rect 21265 17584 21270 17640
rect 21326 17584 26698 17640
rect 26754 17584 26759 17640
rect 21265 17582 26759 17584
rect 21265 17579 21331 17582
rect 26693 17579 26759 17582
rect 8385 17506 8451 17509
rect 9121 17506 9187 17509
rect 9581 17506 9647 17509
rect 8385 17504 9187 17506
rect 8385 17448 8390 17504
rect 8446 17448 9126 17504
rect 9182 17448 9187 17504
rect 8385 17446 9187 17448
rect 8385 17443 8451 17446
rect 9121 17443 9187 17446
rect 9262 17504 9647 17506
rect 9262 17448 9586 17504
rect 9642 17448 9647 17504
rect 9262 17446 9647 17448
rect 4189 17440 4505 17441
rect 4189 17376 4195 17440
rect 4259 17376 4275 17440
rect 4339 17376 4355 17440
rect 4419 17376 4435 17440
rect 4499 17376 4505 17440
rect 4189 17375 4505 17376
rect 5942 17308 5948 17372
rect 6012 17370 6018 17372
rect 9262 17370 9322 17446
rect 9581 17443 9647 17446
rect 19977 17506 20043 17509
rect 22277 17506 22343 17509
rect 19977 17504 22343 17506
rect 19977 17448 19982 17504
rect 20038 17448 22282 17504
rect 22338 17448 22343 17504
rect 19977 17446 22343 17448
rect 19977 17443 20043 17446
rect 22277 17443 22343 17446
rect 22461 17506 22527 17509
rect 22461 17504 25882 17506
rect 22461 17448 22466 17504
rect 22522 17448 25882 17504
rect 22461 17446 25882 17448
rect 22461 17443 22527 17446
rect 11779 17440 12095 17441
rect 11779 17376 11785 17440
rect 11849 17376 11865 17440
rect 11929 17376 11945 17440
rect 12009 17376 12025 17440
rect 12089 17376 12095 17440
rect 11779 17375 12095 17376
rect 19369 17440 19685 17441
rect 19369 17376 19375 17440
rect 19439 17376 19455 17440
rect 19519 17376 19535 17440
rect 19599 17376 19615 17440
rect 19679 17376 19685 17440
rect 19369 17375 19685 17376
rect 6012 17310 9322 17370
rect 21909 17370 21975 17373
rect 25589 17370 25655 17373
rect 21909 17368 25655 17370
rect 21909 17312 21914 17368
rect 21970 17312 25594 17368
rect 25650 17312 25655 17368
rect 21909 17310 25655 17312
rect 25822 17370 25882 17446
rect 26959 17440 27275 17441
rect 26959 17376 26965 17440
rect 27029 17376 27045 17440
rect 27109 17376 27125 17440
rect 27189 17376 27205 17440
rect 27269 17376 27275 17440
rect 26959 17375 27275 17376
rect 26601 17370 26667 17373
rect 25822 17368 26667 17370
rect 25822 17312 26606 17368
rect 26662 17312 26667 17368
rect 25822 17310 26667 17312
rect 6012 17308 6018 17310
rect 21909 17307 21975 17310
rect 25589 17307 25655 17310
rect 26601 17307 26667 17310
rect 8385 17234 8451 17237
rect 13261 17234 13327 17237
rect 16481 17234 16547 17237
rect 28349 17234 28415 17237
rect 8385 17232 13327 17234
rect 8385 17176 8390 17232
rect 8446 17176 13266 17232
rect 13322 17176 13327 17232
rect 8385 17174 13327 17176
rect 8385 17171 8451 17174
rect 13261 17171 13327 17174
rect 15334 17232 28415 17234
rect 15334 17176 16486 17232
rect 16542 17176 28354 17232
rect 28410 17176 28415 17232
rect 15334 17174 28415 17176
rect 8477 17098 8543 17101
rect 13629 17098 13695 17101
rect 14089 17098 14155 17101
rect 8477 17096 14155 17098
rect 8477 17040 8482 17096
rect 8538 17040 13634 17096
rect 13690 17040 14094 17096
rect 14150 17040 14155 17096
rect 8477 17038 14155 17040
rect 8477 17035 8543 17038
rect 13629 17035 13695 17038
rect 14089 17035 14155 17038
rect 5441 16962 5507 16965
rect 7005 16962 7071 16965
rect 5441 16960 7071 16962
rect 5441 16904 5446 16960
rect 5502 16904 7010 16960
rect 7066 16904 7071 16960
rect 5441 16902 7071 16904
rect 5441 16899 5507 16902
rect 7005 16899 7071 16902
rect 12985 16962 13051 16965
rect 14549 16962 14615 16965
rect 12985 16960 14615 16962
rect 12985 16904 12990 16960
rect 13046 16904 14554 16960
rect 14610 16904 14615 16960
rect 12985 16902 14615 16904
rect 12985 16899 13051 16902
rect 14549 16899 14615 16902
rect 7984 16896 8300 16897
rect 7984 16832 7990 16896
rect 8054 16832 8070 16896
rect 8134 16832 8150 16896
rect 8214 16832 8230 16896
rect 8294 16832 8300 16896
rect 7984 16831 8300 16832
rect 1761 16826 1827 16829
rect 1761 16824 6562 16826
rect 1761 16768 1766 16824
rect 1822 16768 6562 16824
rect 1761 16766 6562 16768
rect 1761 16763 1827 16766
rect 5942 16628 5948 16692
rect 6012 16690 6018 16692
rect 6177 16690 6243 16693
rect 6012 16688 6243 16690
rect 6012 16632 6182 16688
rect 6238 16632 6243 16688
rect 6012 16630 6243 16632
rect 6502 16690 6562 16766
rect 8518 16764 8524 16828
rect 8588 16764 8594 16828
rect 11697 16826 11763 16829
rect 11056 16824 11763 16826
rect 11056 16768 11702 16824
rect 11758 16768 11763 16824
rect 11056 16766 11763 16768
rect 8526 16690 8586 16764
rect 11056 16693 11116 16766
rect 11697 16763 11763 16766
rect 11881 16826 11947 16829
rect 15101 16826 15167 16829
rect 15334 16826 15394 17174
rect 16481 17171 16547 17174
rect 28349 17171 28415 17174
rect 16849 17098 16915 17101
rect 22461 17098 22527 17101
rect 23841 17098 23907 17101
rect 29545 17100 29611 17101
rect 29494 17098 29500 17100
rect 16849 17096 22527 17098
rect 16849 17040 16854 17096
rect 16910 17040 22466 17096
rect 22522 17040 22527 17096
rect 16849 17038 22527 17040
rect 16849 17035 16915 17038
rect 22461 17035 22527 17038
rect 22878 17096 23907 17098
rect 22878 17040 23846 17096
rect 23902 17040 23907 17096
rect 22878 17038 23907 17040
rect 29454 17038 29500 17098
rect 29564 17096 29611 17100
rect 29606 17040 29611 17096
rect 22878 16962 22938 17038
rect 23841 17035 23907 17038
rect 29494 17036 29500 17038
rect 29564 17036 29611 17040
rect 29545 17035 29611 17036
rect 22050 16902 22938 16962
rect 15574 16896 15890 16897
rect 15574 16832 15580 16896
rect 15644 16832 15660 16896
rect 15724 16832 15740 16896
rect 15804 16832 15820 16896
rect 15884 16832 15890 16896
rect 15574 16831 15890 16832
rect 11881 16824 15394 16826
rect 11881 16768 11886 16824
rect 11942 16768 15106 16824
rect 15162 16768 15394 16824
rect 11881 16766 15394 16768
rect 16297 16826 16363 16829
rect 22050 16826 22110 16902
rect 23164 16896 23480 16897
rect 23164 16832 23170 16896
rect 23234 16832 23250 16896
rect 23314 16832 23330 16896
rect 23394 16832 23410 16896
rect 23474 16832 23480 16896
rect 23164 16831 23480 16832
rect 30754 16896 31070 16897
rect 30754 16832 30760 16896
rect 30824 16832 30840 16896
rect 30904 16832 30920 16896
rect 30984 16832 31000 16896
rect 31064 16832 31070 16896
rect 30754 16831 31070 16832
rect 22645 16826 22711 16829
rect 29269 16828 29335 16829
rect 29269 16826 29316 16828
rect 16297 16824 22110 16826
rect 16297 16768 16302 16824
rect 16358 16768 22110 16824
rect 16297 16766 22110 16768
rect 22510 16824 22711 16826
rect 22510 16768 22650 16824
rect 22706 16768 22711 16824
rect 22510 16766 22711 16768
rect 29224 16824 29316 16826
rect 29224 16768 29274 16824
rect 29224 16766 29316 16768
rect 11881 16763 11947 16766
rect 15101 16763 15167 16766
rect 16297 16763 16363 16766
rect 6502 16630 8586 16690
rect 9213 16690 9279 16693
rect 11053 16690 11119 16693
rect 9213 16688 11119 16690
rect 9213 16632 9218 16688
rect 9274 16632 11058 16688
rect 11114 16632 11119 16688
rect 9213 16630 11119 16632
rect 6012 16628 6018 16630
rect 6177 16627 6243 16630
rect 9213 16627 9279 16630
rect 11053 16627 11119 16630
rect 11789 16690 11855 16693
rect 15929 16690 15995 16693
rect 11789 16688 15995 16690
rect 11789 16632 11794 16688
rect 11850 16632 15934 16688
rect 15990 16632 15995 16688
rect 11789 16630 15995 16632
rect 11789 16627 11855 16630
rect 15929 16627 15995 16630
rect 21633 16690 21699 16693
rect 22510 16690 22570 16766
rect 22645 16763 22711 16766
rect 29269 16764 29316 16766
rect 29380 16764 29386 16828
rect 29269 16763 29335 16764
rect 21633 16688 22570 16690
rect 21633 16632 21638 16688
rect 21694 16632 22570 16688
rect 21633 16630 22570 16632
rect 23657 16690 23723 16693
rect 30097 16690 30163 16693
rect 23657 16688 30163 16690
rect 23657 16632 23662 16688
rect 23718 16632 30102 16688
rect 30158 16632 30163 16688
rect 23657 16630 30163 16632
rect 21633 16627 21699 16630
rect 23657 16627 23723 16630
rect 30097 16627 30163 16630
rect 4061 16554 4127 16557
rect 6729 16554 6795 16557
rect 4061 16552 6795 16554
rect 4061 16496 4066 16552
rect 4122 16496 6734 16552
rect 6790 16496 6795 16552
rect 4061 16494 6795 16496
rect 4061 16491 4127 16494
rect 6729 16491 6795 16494
rect 9029 16554 9095 16557
rect 14917 16554 14983 16557
rect 9029 16552 14983 16554
rect 9029 16496 9034 16552
rect 9090 16496 14922 16552
rect 14978 16496 14983 16552
rect 9029 16494 14983 16496
rect 9029 16491 9095 16494
rect 14917 16491 14983 16494
rect 19333 16554 19399 16557
rect 24393 16554 24459 16557
rect 29177 16556 29243 16557
rect 29126 16554 29132 16556
rect 19333 16552 24459 16554
rect 19333 16496 19338 16552
rect 19394 16496 24398 16552
rect 24454 16496 24459 16552
rect 19333 16494 24459 16496
rect 29086 16494 29132 16554
rect 29196 16552 29243 16556
rect 29238 16496 29243 16552
rect 19333 16491 19399 16494
rect 24393 16491 24459 16494
rect 29126 16492 29132 16494
rect 29196 16492 29243 16496
rect 29177 16491 29243 16492
rect 13353 16418 13419 16421
rect 14222 16418 14228 16420
rect 13353 16416 14228 16418
rect 13353 16360 13358 16416
rect 13414 16360 14228 16416
rect 13353 16358 14228 16360
rect 13353 16355 13419 16358
rect 14222 16356 14228 16358
rect 14292 16356 14298 16420
rect 21817 16418 21883 16421
rect 24669 16418 24735 16421
rect 21817 16416 24735 16418
rect 21817 16360 21822 16416
rect 21878 16360 24674 16416
rect 24730 16360 24735 16416
rect 21817 16358 24735 16360
rect 21817 16355 21883 16358
rect 24669 16355 24735 16358
rect 29085 16418 29151 16421
rect 29678 16418 29684 16420
rect 29085 16416 29684 16418
rect 29085 16360 29090 16416
rect 29146 16360 29684 16416
rect 29085 16358 29684 16360
rect 29085 16355 29151 16358
rect 29678 16356 29684 16358
rect 29748 16356 29754 16420
rect 4189 16352 4505 16353
rect 4189 16288 4195 16352
rect 4259 16288 4275 16352
rect 4339 16288 4355 16352
rect 4419 16288 4435 16352
rect 4499 16288 4505 16352
rect 4189 16287 4505 16288
rect 11779 16352 12095 16353
rect 11779 16288 11785 16352
rect 11849 16288 11865 16352
rect 11929 16288 11945 16352
rect 12009 16288 12025 16352
rect 12089 16288 12095 16352
rect 11779 16287 12095 16288
rect 19369 16352 19685 16353
rect 19369 16288 19375 16352
rect 19439 16288 19455 16352
rect 19519 16288 19535 16352
rect 19599 16288 19615 16352
rect 19679 16288 19685 16352
rect 19369 16287 19685 16288
rect 26959 16352 27275 16353
rect 26959 16288 26965 16352
rect 27029 16288 27045 16352
rect 27109 16288 27125 16352
rect 27189 16288 27205 16352
rect 27269 16288 27275 16352
rect 26959 16287 27275 16288
rect 5625 16282 5691 16285
rect 10409 16282 10475 16285
rect 5625 16280 10475 16282
rect 5625 16224 5630 16280
rect 5686 16224 10414 16280
rect 10470 16224 10475 16280
rect 5625 16222 10475 16224
rect 5625 16219 5691 16222
rect 10409 16219 10475 16222
rect 13629 16282 13695 16285
rect 15469 16282 15535 16285
rect 24117 16282 24183 16285
rect 28993 16282 29059 16285
rect 30189 16282 30255 16285
rect 13629 16280 15535 16282
rect 13629 16224 13634 16280
rect 13690 16224 15474 16280
rect 15530 16224 15535 16280
rect 13629 16222 15535 16224
rect 13629 16219 13695 16222
rect 15469 16219 15535 16222
rect 22050 16280 26802 16282
rect 22050 16224 24122 16280
rect 24178 16224 26802 16280
rect 22050 16222 26802 16224
rect 2681 16146 2747 16149
rect 9489 16146 9555 16149
rect 2681 16144 9555 16146
rect 2681 16088 2686 16144
rect 2742 16088 9494 16144
rect 9550 16088 9555 16144
rect 2681 16086 9555 16088
rect 2681 16083 2747 16086
rect 9489 16083 9555 16086
rect 11697 16146 11763 16149
rect 16297 16146 16363 16149
rect 11697 16144 16363 16146
rect 11697 16088 11702 16144
rect 11758 16088 16302 16144
rect 16358 16088 16363 16144
rect 11697 16086 16363 16088
rect 11697 16083 11763 16086
rect 16297 16083 16363 16086
rect 20713 16146 20779 16149
rect 22050 16146 22110 16222
rect 24117 16219 24183 16222
rect 20713 16144 22110 16146
rect 20713 16088 20718 16144
rect 20774 16088 22110 16144
rect 20713 16086 22110 16088
rect 22645 16146 22711 16149
rect 24301 16146 24367 16149
rect 25865 16146 25931 16149
rect 22645 16144 25931 16146
rect 22645 16088 22650 16144
rect 22706 16088 24306 16144
rect 24362 16088 25870 16144
rect 25926 16088 25931 16144
rect 22645 16086 25931 16088
rect 26742 16146 26802 16222
rect 28993 16280 30255 16282
rect 28993 16224 28998 16280
rect 29054 16224 30194 16280
rect 30250 16224 30255 16280
rect 28993 16222 30255 16224
rect 28993 16219 29059 16222
rect 30189 16219 30255 16222
rect 28625 16146 28691 16149
rect 26742 16144 28691 16146
rect 26742 16088 28630 16144
rect 28686 16088 28691 16144
rect 26742 16086 28691 16088
rect 20713 16083 20779 16086
rect 22645 16083 22711 16086
rect 24301 16083 24367 16086
rect 25865 16083 25931 16086
rect 28625 16083 28691 16086
rect 29361 16146 29427 16149
rect 29494 16146 29500 16148
rect 29361 16144 29500 16146
rect 29361 16088 29366 16144
rect 29422 16088 29500 16144
rect 29361 16086 29500 16088
rect 29361 16083 29427 16086
rect 29494 16084 29500 16086
rect 29564 16084 29570 16148
rect 2129 16010 2195 16013
rect 17125 16010 17191 16013
rect 2129 16008 17191 16010
rect 2129 15952 2134 16008
rect 2190 15952 17130 16008
rect 17186 15952 17191 16008
rect 2129 15950 17191 15952
rect 2129 15947 2195 15950
rect 17125 15947 17191 15950
rect 22829 16010 22895 16013
rect 24853 16010 24919 16013
rect 22829 16008 24919 16010
rect 22829 15952 22834 16008
rect 22890 15952 24858 16008
rect 24914 15952 24919 16008
rect 22829 15950 24919 15952
rect 22829 15947 22895 15950
rect 24853 15947 24919 15950
rect 26233 16010 26299 16013
rect 31109 16010 31175 16013
rect 31385 16010 31451 16013
rect 26233 16008 31451 16010
rect 26233 15952 26238 16008
rect 26294 15952 31114 16008
rect 31170 15952 31390 16008
rect 31446 15952 31451 16008
rect 26233 15950 31451 15952
rect 26233 15947 26299 15950
rect 31109 15947 31175 15950
rect 31385 15947 31451 15950
rect 10777 15874 10843 15877
rect 13905 15874 13971 15877
rect 10777 15872 13971 15874
rect 10777 15816 10782 15872
rect 10838 15816 13910 15872
rect 13966 15816 13971 15872
rect 10777 15814 13971 15816
rect 10777 15811 10843 15814
rect 13905 15811 13971 15814
rect 24669 15874 24735 15877
rect 28073 15874 28139 15877
rect 30005 15874 30071 15877
rect 24669 15872 30071 15874
rect 24669 15816 24674 15872
rect 24730 15816 28078 15872
rect 28134 15816 30010 15872
rect 30066 15816 30071 15872
rect 24669 15814 30071 15816
rect 24669 15811 24735 15814
rect 28073 15811 28139 15814
rect 30005 15811 30071 15814
rect 7984 15808 8300 15809
rect 7984 15744 7990 15808
rect 8054 15744 8070 15808
rect 8134 15744 8150 15808
rect 8214 15744 8230 15808
rect 8294 15744 8300 15808
rect 7984 15743 8300 15744
rect 15574 15808 15890 15809
rect 15574 15744 15580 15808
rect 15644 15744 15660 15808
rect 15724 15744 15740 15808
rect 15804 15744 15820 15808
rect 15884 15744 15890 15808
rect 15574 15743 15890 15744
rect 23164 15808 23480 15809
rect 23164 15744 23170 15808
rect 23234 15744 23250 15808
rect 23314 15744 23330 15808
rect 23394 15744 23410 15808
rect 23474 15744 23480 15808
rect 23164 15743 23480 15744
rect 30754 15808 31070 15809
rect 30754 15744 30760 15808
rect 30824 15744 30840 15808
rect 30904 15744 30920 15808
rect 30984 15744 31000 15808
rect 31064 15744 31070 15808
rect 30754 15743 31070 15744
rect 12566 15676 12572 15740
rect 12636 15738 12642 15740
rect 13537 15738 13603 15741
rect 12636 15736 13603 15738
rect 12636 15680 13542 15736
rect 13598 15680 13603 15736
rect 12636 15678 13603 15680
rect 12636 15676 12642 15678
rect 13537 15675 13603 15678
rect 19609 15738 19675 15741
rect 21725 15738 21791 15741
rect 19609 15736 21791 15738
rect 19609 15680 19614 15736
rect 19670 15680 21730 15736
rect 21786 15680 21791 15736
rect 19609 15678 21791 15680
rect 19609 15675 19675 15678
rect 21725 15675 21791 15678
rect 29085 15738 29151 15741
rect 29310 15738 29316 15740
rect 29085 15736 29316 15738
rect 29085 15680 29090 15736
rect 29146 15680 29316 15736
rect 29085 15678 29316 15680
rect 29085 15675 29151 15678
rect 29310 15676 29316 15678
rect 29380 15676 29386 15740
rect 6269 15602 6335 15605
rect 8293 15602 8359 15605
rect 13445 15602 13511 15605
rect 6269 15600 7666 15602
rect 6269 15544 6274 15600
rect 6330 15544 7666 15600
rect 6269 15542 7666 15544
rect 6269 15539 6335 15542
rect 2037 15466 2103 15469
rect 7465 15466 7531 15469
rect 2037 15464 7531 15466
rect 2037 15408 2042 15464
rect 2098 15408 7470 15464
rect 7526 15408 7531 15464
rect 2037 15406 7531 15408
rect 7606 15466 7666 15542
rect 8293 15600 13511 15602
rect 8293 15544 8298 15600
rect 8354 15544 13450 15600
rect 13506 15544 13511 15600
rect 8293 15542 13511 15544
rect 8293 15539 8359 15542
rect 13445 15539 13511 15542
rect 19701 15602 19767 15605
rect 25497 15602 25563 15605
rect 19701 15600 25563 15602
rect 19701 15544 19706 15600
rect 19762 15544 25502 15600
rect 25558 15544 25563 15600
rect 19701 15542 25563 15544
rect 19701 15539 19767 15542
rect 25497 15539 25563 15542
rect 16849 15466 16915 15469
rect 7606 15464 16915 15466
rect 7606 15408 16854 15464
rect 16910 15408 16915 15464
rect 7606 15406 16915 15408
rect 2037 15403 2103 15406
rect 7465 15403 7531 15406
rect 16849 15403 16915 15406
rect 22461 15466 22527 15469
rect 24393 15466 24459 15469
rect 22461 15464 24459 15466
rect 22461 15408 22466 15464
rect 22522 15408 24398 15464
rect 24454 15408 24459 15464
rect 22461 15406 24459 15408
rect 22461 15403 22527 15406
rect 24393 15403 24459 15406
rect 26049 15466 26115 15469
rect 27889 15466 27955 15469
rect 26049 15464 27955 15466
rect 26049 15408 26054 15464
rect 26110 15408 27894 15464
rect 27950 15408 27955 15464
rect 26049 15406 27955 15408
rect 26049 15403 26115 15406
rect 27889 15403 27955 15406
rect 23749 15330 23815 15333
rect 26233 15330 26299 15333
rect 23749 15328 26299 15330
rect 23749 15272 23754 15328
rect 23810 15272 26238 15328
rect 26294 15272 26299 15328
rect 23749 15270 26299 15272
rect 23749 15267 23815 15270
rect 26233 15267 26299 15270
rect 4189 15264 4505 15265
rect 4189 15200 4195 15264
rect 4259 15200 4275 15264
rect 4339 15200 4355 15264
rect 4419 15200 4435 15264
rect 4499 15200 4505 15264
rect 4189 15199 4505 15200
rect 11779 15264 12095 15265
rect 11779 15200 11785 15264
rect 11849 15200 11865 15264
rect 11929 15200 11945 15264
rect 12009 15200 12025 15264
rect 12089 15200 12095 15264
rect 11779 15199 12095 15200
rect 19369 15264 19685 15265
rect 19369 15200 19375 15264
rect 19439 15200 19455 15264
rect 19519 15200 19535 15264
rect 19599 15200 19615 15264
rect 19679 15200 19685 15264
rect 19369 15199 19685 15200
rect 26959 15264 27275 15265
rect 26959 15200 26965 15264
rect 27029 15200 27045 15264
rect 27109 15200 27125 15264
rect 27189 15200 27205 15264
rect 27269 15200 27275 15264
rect 26959 15199 27275 15200
rect 6177 15194 6243 15197
rect 8201 15194 8267 15197
rect 6177 15192 8267 15194
rect 6177 15136 6182 15192
rect 6238 15136 8206 15192
rect 8262 15136 8267 15192
rect 6177 15134 8267 15136
rect 6177 15131 6243 15134
rect 8201 15131 8267 15134
rect 8518 15132 8524 15196
rect 8588 15194 8594 15196
rect 10133 15194 10199 15197
rect 8588 15192 10199 15194
rect 8588 15136 10138 15192
rect 10194 15136 10199 15192
rect 8588 15134 10199 15136
rect 8588 15132 8594 15134
rect 10133 15131 10199 15134
rect 20529 15194 20595 15197
rect 23657 15194 23723 15197
rect 26509 15196 26575 15197
rect 26509 15194 26556 15196
rect 20529 15192 23723 15194
rect 20529 15136 20534 15192
rect 20590 15136 23662 15192
rect 23718 15136 23723 15192
rect 20529 15134 23723 15136
rect 26464 15192 26556 15194
rect 26464 15136 26514 15192
rect 26464 15134 26556 15136
rect 20529 15131 20595 15134
rect 23657 15131 23723 15134
rect 26509 15132 26556 15134
rect 26620 15132 26626 15196
rect 26509 15131 26575 15132
rect 2129 15058 2195 15061
rect 10409 15058 10475 15061
rect 2129 15056 10475 15058
rect 2129 15000 2134 15056
rect 2190 15000 10414 15056
rect 10470 15000 10475 15056
rect 2129 14998 10475 15000
rect 2129 14995 2195 14998
rect 10409 14995 10475 14998
rect 16389 15058 16455 15061
rect 18321 15058 18387 15061
rect 24669 15058 24735 15061
rect 16389 15056 18387 15058
rect 16389 15000 16394 15056
rect 16450 15000 18326 15056
rect 18382 15000 18387 15056
rect 16389 14998 18387 15000
rect 16389 14995 16455 14998
rect 18321 14995 18387 14998
rect 19198 15056 24735 15058
rect 19198 15000 24674 15056
rect 24730 15000 24735 15056
rect 19198 14998 24735 15000
rect 6085 14922 6151 14925
rect 7281 14922 7347 14925
rect 6085 14920 7347 14922
rect 6085 14864 6090 14920
rect 6146 14864 7286 14920
rect 7342 14864 7347 14920
rect 6085 14862 7347 14864
rect 6085 14859 6151 14862
rect 7281 14859 7347 14862
rect 8477 14922 8543 14925
rect 13445 14922 13511 14925
rect 8477 14920 13511 14922
rect 8477 14864 8482 14920
rect 8538 14864 13450 14920
rect 13506 14864 13511 14920
rect 8477 14862 13511 14864
rect 8477 14859 8543 14862
rect 13445 14859 13511 14862
rect 15101 14922 15167 14925
rect 19057 14922 19123 14925
rect 15101 14920 19123 14922
rect 15101 14864 15106 14920
rect 15162 14864 19062 14920
rect 19118 14864 19123 14920
rect 15101 14862 19123 14864
rect 15101 14859 15167 14862
rect 19057 14859 19123 14862
rect 19057 14786 19123 14789
rect 19198 14786 19258 14998
rect 24669 14995 24735 14998
rect 22001 14922 22067 14925
rect 27613 14922 27679 14925
rect 22001 14920 27679 14922
rect 22001 14864 22006 14920
rect 22062 14864 27618 14920
rect 27674 14864 27679 14920
rect 22001 14862 27679 14864
rect 22001 14859 22067 14862
rect 27613 14859 27679 14862
rect 19057 14784 19258 14786
rect 19057 14728 19062 14784
rect 19118 14728 19258 14784
rect 19057 14726 19258 14728
rect 23841 14786 23907 14789
rect 28717 14786 28783 14789
rect 23841 14784 28783 14786
rect 23841 14728 23846 14784
rect 23902 14728 28722 14784
rect 28778 14728 28783 14784
rect 23841 14726 28783 14728
rect 19057 14723 19123 14726
rect 23841 14723 23907 14726
rect 28717 14723 28783 14726
rect 7984 14720 8300 14721
rect 7984 14656 7990 14720
rect 8054 14656 8070 14720
rect 8134 14656 8150 14720
rect 8214 14656 8230 14720
rect 8294 14656 8300 14720
rect 7984 14655 8300 14656
rect 15574 14720 15890 14721
rect 15574 14656 15580 14720
rect 15644 14656 15660 14720
rect 15724 14656 15740 14720
rect 15804 14656 15820 14720
rect 15884 14656 15890 14720
rect 15574 14655 15890 14656
rect 23164 14720 23480 14721
rect 23164 14656 23170 14720
rect 23234 14656 23250 14720
rect 23314 14656 23330 14720
rect 23394 14656 23410 14720
rect 23474 14656 23480 14720
rect 23164 14655 23480 14656
rect 30754 14720 31070 14721
rect 30754 14656 30760 14720
rect 30824 14656 30840 14720
rect 30904 14656 30920 14720
rect 30984 14656 31000 14720
rect 31064 14656 31070 14720
rect 30754 14655 31070 14656
rect 19885 14650 19951 14653
rect 21265 14650 21331 14653
rect 19885 14648 21331 14650
rect 19885 14592 19890 14648
rect 19946 14592 21270 14648
rect 21326 14592 21331 14648
rect 19885 14590 21331 14592
rect 19885 14587 19951 14590
rect 21265 14587 21331 14590
rect 23565 14650 23631 14653
rect 27061 14650 27127 14653
rect 23565 14648 27127 14650
rect 23565 14592 23570 14648
rect 23626 14592 27066 14648
rect 27122 14592 27127 14648
rect 23565 14590 27127 14592
rect 23565 14587 23631 14590
rect 27061 14587 27127 14590
rect 27797 14650 27863 14653
rect 28717 14650 28783 14653
rect 27797 14648 28783 14650
rect 27797 14592 27802 14648
rect 27858 14592 28722 14648
rect 28778 14592 28783 14648
rect 27797 14590 28783 14592
rect 27797 14587 27863 14590
rect 28717 14587 28783 14590
rect 2037 14514 2103 14517
rect 29913 14514 29979 14517
rect 2037 14512 29979 14514
rect 2037 14456 2042 14512
rect 2098 14456 29918 14512
rect 29974 14456 29979 14512
rect 2037 14454 29979 14456
rect 2037 14451 2103 14454
rect 29913 14451 29979 14454
rect 4797 14378 4863 14381
rect 9121 14378 9187 14381
rect 4797 14376 9187 14378
rect 4797 14320 4802 14376
rect 4858 14320 9126 14376
rect 9182 14320 9187 14376
rect 4797 14318 9187 14320
rect 4797 14315 4863 14318
rect 9121 14315 9187 14318
rect 11789 14378 11855 14381
rect 14273 14378 14339 14381
rect 11789 14376 14339 14378
rect 11789 14320 11794 14376
rect 11850 14320 14278 14376
rect 14334 14320 14339 14376
rect 11789 14318 14339 14320
rect 11789 14315 11855 14318
rect 14273 14315 14339 14318
rect 14457 14378 14523 14381
rect 18965 14378 19031 14381
rect 20161 14378 20227 14381
rect 14457 14376 19031 14378
rect 14457 14320 14462 14376
rect 14518 14320 18970 14376
rect 19026 14320 19031 14376
rect 14457 14318 19031 14320
rect 14457 14315 14523 14318
rect 18965 14315 19031 14318
rect 19198 14376 20227 14378
rect 19198 14320 20166 14376
rect 20222 14320 20227 14376
rect 19198 14318 20227 14320
rect 6361 14242 6427 14245
rect 8569 14242 8635 14245
rect 6361 14240 8635 14242
rect 6361 14184 6366 14240
rect 6422 14184 8574 14240
rect 8630 14184 8635 14240
rect 6361 14182 8635 14184
rect 6361 14179 6427 14182
rect 8569 14179 8635 14182
rect 14089 14242 14155 14245
rect 19198 14242 19258 14318
rect 20161 14315 20227 14318
rect 20621 14378 20687 14381
rect 25681 14378 25747 14381
rect 20621 14376 25747 14378
rect 20621 14320 20626 14376
rect 20682 14320 25686 14376
rect 25742 14320 25747 14376
rect 20621 14318 25747 14320
rect 20621 14315 20687 14318
rect 25681 14315 25747 14318
rect 14089 14240 19258 14242
rect 14089 14184 14094 14240
rect 14150 14184 19258 14240
rect 14089 14182 19258 14184
rect 20529 14242 20595 14245
rect 23565 14242 23631 14245
rect 20529 14240 23631 14242
rect 20529 14184 20534 14240
rect 20590 14184 23570 14240
rect 23626 14184 23631 14240
rect 20529 14182 23631 14184
rect 14089 14179 14155 14182
rect 20529 14179 20595 14182
rect 23565 14179 23631 14182
rect 4189 14176 4505 14177
rect 4189 14112 4195 14176
rect 4259 14112 4275 14176
rect 4339 14112 4355 14176
rect 4419 14112 4435 14176
rect 4499 14112 4505 14176
rect 4189 14111 4505 14112
rect 11779 14176 12095 14177
rect 11779 14112 11785 14176
rect 11849 14112 11865 14176
rect 11929 14112 11945 14176
rect 12009 14112 12025 14176
rect 12089 14112 12095 14176
rect 11779 14111 12095 14112
rect 19369 14176 19685 14177
rect 19369 14112 19375 14176
rect 19439 14112 19455 14176
rect 19519 14112 19535 14176
rect 19599 14112 19615 14176
rect 19679 14112 19685 14176
rect 19369 14111 19685 14112
rect 26959 14176 27275 14177
rect 26959 14112 26965 14176
rect 27029 14112 27045 14176
rect 27109 14112 27125 14176
rect 27189 14112 27205 14176
rect 27269 14112 27275 14176
rect 26959 14111 27275 14112
rect 5533 14106 5599 14109
rect 9673 14106 9739 14109
rect 11329 14106 11395 14109
rect 5533 14104 11395 14106
rect 5533 14048 5538 14104
rect 5594 14048 9678 14104
rect 9734 14048 11334 14104
rect 11390 14048 11395 14104
rect 5533 14046 11395 14048
rect 5533 14043 5599 14046
rect 9673 14043 9739 14046
rect 11329 14043 11395 14046
rect 12525 14106 12591 14109
rect 18965 14106 19031 14109
rect 12525 14104 19031 14106
rect 12525 14048 12530 14104
rect 12586 14048 18970 14104
rect 19026 14048 19031 14104
rect 12525 14046 19031 14048
rect 12525 14043 12591 14046
rect 18965 14043 19031 14046
rect 24209 14106 24275 14109
rect 25037 14106 25103 14109
rect 24209 14104 25103 14106
rect 24209 14048 24214 14104
rect 24270 14048 25042 14104
rect 25098 14048 25103 14104
rect 24209 14046 25103 14048
rect 24209 14043 24275 14046
rect 25037 14043 25103 14046
rect 29085 14106 29151 14109
rect 29085 14104 29194 14106
rect 29085 14048 29090 14104
rect 29146 14048 29194 14104
rect 29085 14043 29194 14048
rect 5390 13908 5396 13972
rect 5460 13970 5466 13972
rect 14273 13970 14339 13973
rect 5460 13968 14339 13970
rect 5460 13912 14278 13968
rect 14334 13912 14339 13968
rect 5460 13910 14339 13912
rect 5460 13908 5466 13910
rect 14273 13907 14339 13910
rect 16665 13970 16731 13973
rect 28993 13970 29059 13973
rect 16665 13968 29059 13970
rect 16665 13912 16670 13968
rect 16726 13912 28998 13968
rect 29054 13912 29059 13968
rect 16665 13910 29059 13912
rect 16665 13907 16731 13910
rect 28993 13907 29059 13910
rect 3049 13834 3115 13837
rect 15193 13834 15259 13837
rect 3049 13832 15259 13834
rect 3049 13776 3054 13832
rect 3110 13776 15198 13832
rect 15254 13776 15259 13832
rect 3049 13774 15259 13776
rect 3049 13771 3115 13774
rect 15193 13771 15259 13774
rect 23933 13834 23999 13837
rect 28533 13834 28599 13837
rect 23933 13832 28599 13834
rect 23933 13776 23938 13832
rect 23994 13776 28538 13832
rect 28594 13776 28599 13832
rect 23933 13774 28599 13776
rect 23933 13771 23999 13774
rect 28533 13771 28599 13774
rect 8937 13700 9003 13701
rect 8886 13636 8892 13700
rect 8956 13698 9003 13700
rect 10317 13698 10383 13701
rect 13353 13698 13419 13701
rect 8956 13696 9048 13698
rect 8998 13640 9048 13696
rect 8956 13638 9048 13640
rect 10317 13696 13419 13698
rect 10317 13640 10322 13696
rect 10378 13640 13358 13696
rect 13414 13640 13419 13696
rect 10317 13638 13419 13640
rect 8956 13636 9003 13638
rect 8937 13635 9003 13636
rect 10317 13635 10383 13638
rect 13353 13635 13419 13638
rect 13721 13698 13787 13701
rect 15377 13698 15443 13701
rect 13721 13696 15443 13698
rect 13721 13640 13726 13696
rect 13782 13640 15382 13696
rect 15438 13640 15443 13696
rect 13721 13638 15443 13640
rect 13721 13635 13787 13638
rect 15377 13635 15443 13638
rect 23841 13698 23907 13701
rect 24853 13698 24919 13701
rect 23841 13696 24919 13698
rect 23841 13640 23846 13696
rect 23902 13640 24858 13696
rect 24914 13640 24919 13696
rect 23841 13638 24919 13640
rect 29134 13698 29194 14043
rect 29269 13834 29335 13837
rect 30281 13834 30347 13837
rect 29269 13832 30347 13834
rect 29269 13776 29274 13832
rect 29330 13776 30286 13832
rect 30342 13776 30347 13832
rect 29269 13774 30347 13776
rect 29269 13771 29335 13774
rect 30281 13771 30347 13774
rect 29361 13698 29427 13701
rect 29134 13696 29427 13698
rect 29134 13640 29366 13696
rect 29422 13640 29427 13696
rect 29134 13638 29427 13640
rect 23841 13635 23907 13638
rect 24853 13635 24919 13638
rect 29361 13635 29427 13638
rect 29678 13636 29684 13700
rect 29748 13698 29754 13700
rect 30281 13698 30347 13701
rect 29748 13696 30347 13698
rect 29748 13640 30286 13696
rect 30342 13640 30347 13696
rect 29748 13638 30347 13640
rect 29748 13636 29754 13638
rect 30281 13635 30347 13638
rect 7984 13632 8300 13633
rect 7984 13568 7990 13632
rect 8054 13568 8070 13632
rect 8134 13568 8150 13632
rect 8214 13568 8230 13632
rect 8294 13568 8300 13632
rect 7984 13567 8300 13568
rect 15574 13632 15890 13633
rect 15574 13568 15580 13632
rect 15644 13568 15660 13632
rect 15724 13568 15740 13632
rect 15804 13568 15820 13632
rect 15884 13568 15890 13632
rect 15574 13567 15890 13568
rect 23164 13632 23480 13633
rect 23164 13568 23170 13632
rect 23234 13568 23250 13632
rect 23314 13568 23330 13632
rect 23394 13568 23410 13632
rect 23474 13568 23480 13632
rect 23164 13567 23480 13568
rect 30754 13632 31070 13633
rect 30754 13568 30760 13632
rect 30824 13568 30840 13632
rect 30904 13568 30920 13632
rect 30984 13568 31000 13632
rect 31064 13568 31070 13632
rect 30754 13567 31070 13568
rect 2405 13562 2471 13565
rect 6453 13562 6519 13565
rect 2405 13560 6519 13562
rect 2405 13504 2410 13560
rect 2466 13504 6458 13560
rect 6514 13504 6519 13560
rect 2405 13502 6519 13504
rect 2405 13499 2471 13502
rect 6453 13499 6519 13502
rect 10225 13562 10291 13565
rect 12985 13562 13051 13565
rect 10225 13560 13051 13562
rect 10225 13504 10230 13560
rect 10286 13504 12990 13560
rect 13046 13504 13051 13560
rect 10225 13502 13051 13504
rect 10225 13499 10291 13502
rect 12985 13499 13051 13502
rect 23974 13500 23980 13564
rect 24044 13562 24050 13564
rect 29269 13562 29335 13565
rect 24044 13560 29335 13562
rect 24044 13504 29274 13560
rect 29330 13504 29335 13560
rect 24044 13502 29335 13504
rect 24044 13500 24050 13502
rect 29269 13499 29335 13502
rect 1945 13426 2011 13429
rect 26601 13426 26667 13429
rect 1945 13424 26667 13426
rect 1945 13368 1950 13424
rect 2006 13368 26606 13424
rect 26662 13368 26667 13424
rect 1945 13366 26667 13368
rect 1945 13363 2011 13366
rect 26601 13363 26667 13366
rect 29269 13426 29335 13429
rect 31293 13426 31359 13429
rect 29269 13424 31359 13426
rect 29269 13368 29274 13424
rect 29330 13368 31298 13424
rect 31354 13368 31359 13424
rect 29269 13366 31359 13368
rect 29269 13363 29335 13366
rect 31293 13363 31359 13366
rect 2773 13290 2839 13293
rect 16573 13290 16639 13293
rect 2773 13288 16639 13290
rect 2773 13232 2778 13288
rect 2834 13232 16578 13288
rect 16634 13232 16639 13288
rect 2773 13230 16639 13232
rect 2773 13227 2839 13230
rect 16573 13227 16639 13230
rect 20621 13290 20687 13293
rect 27981 13290 28047 13293
rect 20621 13288 28047 13290
rect 20621 13232 20626 13288
rect 20682 13232 27986 13288
rect 28042 13232 28047 13288
rect 20621 13230 28047 13232
rect 20621 13227 20687 13230
rect 27981 13227 28047 13230
rect 6453 13154 6519 13157
rect 7925 13154 7991 13157
rect 6453 13152 7991 13154
rect 6453 13096 6458 13152
rect 6514 13096 7930 13152
rect 7986 13096 7991 13152
rect 6453 13094 7991 13096
rect 6453 13091 6519 13094
rect 7925 13091 7991 13094
rect 9673 13154 9739 13157
rect 10777 13154 10843 13157
rect 9673 13152 10843 13154
rect 9673 13096 9678 13152
rect 9734 13096 10782 13152
rect 10838 13096 10843 13152
rect 9673 13094 10843 13096
rect 9673 13091 9739 13094
rect 10777 13091 10843 13094
rect 4189 13088 4505 13089
rect 4189 13024 4195 13088
rect 4259 13024 4275 13088
rect 4339 13024 4355 13088
rect 4419 13024 4435 13088
rect 4499 13024 4505 13088
rect 4189 13023 4505 13024
rect 11779 13088 12095 13089
rect 11779 13024 11785 13088
rect 11849 13024 11865 13088
rect 11929 13024 11945 13088
rect 12009 13024 12025 13088
rect 12089 13024 12095 13088
rect 11779 13023 12095 13024
rect 19369 13088 19685 13089
rect 19369 13024 19375 13088
rect 19439 13024 19455 13088
rect 19519 13024 19535 13088
rect 19599 13024 19615 13088
rect 19679 13024 19685 13088
rect 19369 13023 19685 13024
rect 26959 13088 27275 13089
rect 26959 13024 26965 13088
rect 27029 13024 27045 13088
rect 27109 13024 27125 13088
rect 27189 13024 27205 13088
rect 27269 13024 27275 13088
rect 26959 13023 27275 13024
rect 7833 13018 7899 13021
rect 10317 13018 10383 13021
rect 7833 13016 10383 13018
rect 7833 12960 7838 13016
rect 7894 12960 10322 13016
rect 10378 12960 10383 13016
rect 7833 12958 10383 12960
rect 7833 12955 7899 12958
rect 10317 12955 10383 12958
rect 10542 12956 10548 13020
rect 10612 13018 10618 13020
rect 11237 13018 11303 13021
rect 10612 13016 11303 13018
rect 10612 12960 11242 13016
rect 11298 12960 11303 13016
rect 10612 12958 11303 12960
rect 10612 12956 10618 12958
rect 11237 12955 11303 12958
rect 12341 13018 12407 13021
rect 16757 13018 16823 13021
rect 29085 13020 29151 13021
rect 29085 13018 29132 13020
rect 12341 13016 16823 13018
rect 12341 12960 12346 13016
rect 12402 12960 16762 13016
rect 16818 12960 16823 13016
rect 12341 12958 16823 12960
rect 29040 13016 29132 13018
rect 29040 12960 29090 13016
rect 29040 12958 29132 12960
rect 12341 12955 12407 12958
rect 16757 12955 16823 12958
rect 29085 12956 29132 12958
rect 29196 12956 29202 13020
rect 29085 12955 29151 12956
rect 2129 12882 2195 12885
rect 28993 12882 29059 12885
rect 2129 12880 29059 12882
rect 2129 12824 2134 12880
rect 2190 12824 28998 12880
rect 29054 12824 29059 12880
rect 2129 12822 29059 12824
rect 2129 12819 2195 12822
rect 28993 12819 29059 12822
rect 6085 12746 6151 12749
rect 6310 12746 6316 12748
rect 6085 12744 6316 12746
rect 6085 12688 6090 12744
rect 6146 12688 6316 12744
rect 6085 12686 6316 12688
rect 6085 12683 6151 12686
rect 6310 12684 6316 12686
rect 6380 12746 6386 12748
rect 7465 12746 7531 12749
rect 6380 12744 7531 12746
rect 6380 12688 7470 12744
rect 7526 12688 7531 12744
rect 6380 12686 7531 12688
rect 6380 12684 6386 12686
rect 7465 12683 7531 12686
rect 7782 12684 7788 12748
rect 7852 12746 7858 12748
rect 9489 12746 9555 12749
rect 14549 12746 14615 12749
rect 7852 12744 9555 12746
rect 7852 12688 9494 12744
rect 9550 12688 9555 12744
rect 7852 12686 9555 12688
rect 7852 12684 7858 12686
rect 9489 12683 9555 12686
rect 11470 12744 14615 12746
rect 11470 12688 14554 12744
rect 14610 12688 14615 12744
rect 11470 12686 14615 12688
rect 7373 12608 7439 12613
rect 7373 12552 7378 12608
rect 7434 12552 7439 12608
rect 7373 12547 7439 12552
rect 8845 12610 8911 12613
rect 9857 12610 9923 12613
rect 8845 12608 9923 12610
rect 8845 12552 8850 12608
rect 8906 12552 9862 12608
rect 9918 12552 9923 12608
rect 8845 12550 9923 12552
rect 8845 12547 8911 12550
rect 9857 12547 9923 12550
rect 2313 12474 2379 12477
rect 2814 12474 2820 12476
rect 2313 12472 2820 12474
rect 2313 12416 2318 12472
rect 2374 12416 2820 12472
rect 2313 12414 2820 12416
rect 2313 12411 2379 12414
rect 2814 12412 2820 12414
rect 2884 12412 2890 12476
rect 7005 12474 7071 12477
rect 7376 12474 7436 12547
rect 7984 12544 8300 12545
rect 7984 12480 7990 12544
rect 8054 12480 8070 12544
rect 8134 12480 8150 12544
rect 8214 12480 8230 12544
rect 8294 12480 8300 12544
rect 7984 12479 8300 12480
rect 11470 12474 11530 12686
rect 14549 12683 14615 12686
rect 16297 12746 16363 12749
rect 23933 12746 23999 12749
rect 16297 12744 23999 12746
rect 16297 12688 16302 12744
rect 16358 12688 23938 12744
rect 23994 12688 23999 12744
rect 16297 12686 23999 12688
rect 16297 12683 16363 12686
rect 23933 12683 23999 12686
rect 29269 12746 29335 12749
rect 30005 12746 30071 12749
rect 29269 12744 30071 12746
rect 29269 12688 29274 12744
rect 29330 12688 30010 12744
rect 30066 12688 30071 12744
rect 29269 12686 30071 12688
rect 29269 12683 29335 12686
rect 30005 12683 30071 12686
rect 15574 12544 15890 12545
rect 15574 12480 15580 12544
rect 15644 12480 15660 12544
rect 15724 12480 15740 12544
rect 15804 12480 15820 12544
rect 15884 12480 15890 12544
rect 15574 12479 15890 12480
rect 23164 12544 23480 12545
rect 23164 12480 23170 12544
rect 23234 12480 23250 12544
rect 23314 12480 23330 12544
rect 23394 12480 23410 12544
rect 23474 12480 23480 12544
rect 23164 12479 23480 12480
rect 30754 12544 31070 12545
rect 30754 12480 30760 12544
rect 30824 12480 30840 12544
rect 30904 12480 30920 12544
rect 30984 12480 31000 12544
rect 31064 12480 31070 12544
rect 30754 12479 31070 12480
rect 7005 12472 7436 12474
rect 7005 12416 7010 12472
rect 7066 12416 7436 12472
rect 7005 12414 7436 12416
rect 9630 12414 11530 12474
rect 7005 12411 7071 12414
rect 1761 12338 1827 12341
rect 2221 12338 2287 12341
rect 9630 12338 9690 12414
rect 27654 12412 27660 12476
rect 27724 12474 27730 12476
rect 29269 12474 29335 12477
rect 27724 12472 29335 12474
rect 27724 12416 29274 12472
rect 29330 12416 29335 12472
rect 27724 12414 29335 12416
rect 27724 12412 27730 12414
rect 29269 12411 29335 12414
rect 1761 12336 9690 12338
rect 1761 12280 1766 12336
rect 1822 12280 2226 12336
rect 2282 12280 9690 12336
rect 1761 12278 9690 12280
rect 9765 12338 9831 12341
rect 11513 12338 11579 12341
rect 9765 12336 11579 12338
rect 9765 12280 9770 12336
rect 9826 12280 11518 12336
rect 11574 12280 11579 12336
rect 9765 12278 11579 12280
rect 1761 12275 1827 12278
rect 2221 12275 2287 12278
rect 9765 12275 9831 12278
rect 11513 12275 11579 12278
rect 12525 12338 12591 12341
rect 14273 12338 14339 12341
rect 12525 12336 14339 12338
rect 12525 12280 12530 12336
rect 12586 12280 14278 12336
rect 14334 12280 14339 12336
rect 12525 12278 14339 12280
rect 12525 12275 12591 12278
rect 14273 12275 14339 12278
rect 28758 12276 28764 12340
rect 28828 12338 28834 12340
rect 28901 12338 28967 12341
rect 28828 12336 28967 12338
rect 28828 12280 28906 12336
rect 28962 12280 28967 12336
rect 28828 12278 28967 12280
rect 28828 12276 28834 12278
rect 28901 12275 28967 12278
rect 1209 12202 1275 12205
rect 4981 12202 5047 12205
rect 1209 12200 5047 12202
rect 1209 12144 1214 12200
rect 1270 12144 4986 12200
rect 5042 12144 5047 12200
rect 1209 12142 5047 12144
rect 1209 12139 1275 12142
rect 4981 12139 5047 12142
rect 7649 12202 7715 12205
rect 11053 12202 11119 12205
rect 12566 12202 12572 12204
rect 7649 12200 11119 12202
rect 7649 12144 7654 12200
rect 7710 12144 11058 12200
rect 11114 12144 11119 12200
rect 7649 12142 11119 12144
rect 7649 12139 7715 12142
rect 11053 12139 11119 12142
rect 11286 12142 12572 12202
rect 7097 12066 7163 12069
rect 11286 12066 11346 12142
rect 12566 12140 12572 12142
rect 12636 12140 12642 12204
rect 22553 12202 22619 12205
rect 29913 12202 29979 12205
rect 22553 12200 29979 12202
rect 22553 12144 22558 12200
rect 22614 12144 29918 12200
rect 29974 12144 29979 12200
rect 22553 12142 29979 12144
rect 22553 12139 22619 12142
rect 29913 12139 29979 12142
rect 7097 12064 11346 12066
rect 7097 12008 7102 12064
rect 7158 12008 11346 12064
rect 7097 12006 11346 12008
rect 7097 12003 7163 12006
rect 11462 12004 11468 12068
rect 11532 12066 11538 12068
rect 11605 12066 11671 12069
rect 11532 12064 11671 12066
rect 11532 12008 11610 12064
rect 11666 12008 11671 12064
rect 11532 12006 11671 12008
rect 11532 12004 11538 12006
rect 11605 12003 11671 12006
rect 4189 12000 4505 12001
rect 4189 11936 4195 12000
rect 4259 11936 4275 12000
rect 4339 11936 4355 12000
rect 4419 11936 4435 12000
rect 4499 11936 4505 12000
rect 4189 11935 4505 11936
rect 11779 12000 12095 12001
rect 11779 11936 11785 12000
rect 11849 11936 11865 12000
rect 11929 11936 11945 12000
rect 12009 11936 12025 12000
rect 12089 11936 12095 12000
rect 11779 11935 12095 11936
rect 19369 12000 19685 12001
rect 19369 11936 19375 12000
rect 19439 11936 19455 12000
rect 19519 11936 19535 12000
rect 19599 11936 19615 12000
rect 19679 11936 19685 12000
rect 19369 11935 19685 11936
rect 26959 12000 27275 12001
rect 26959 11936 26965 12000
rect 27029 11936 27045 12000
rect 27109 11936 27125 12000
rect 27189 11936 27205 12000
rect 27269 11936 27275 12000
rect 26959 11935 27275 11936
rect 8477 11930 8543 11933
rect 12157 11930 12223 11933
rect 13169 11930 13235 11933
rect 8477 11928 11714 11930
rect 8477 11872 8482 11928
rect 8538 11872 11714 11928
rect 8477 11870 11714 11872
rect 8477 11867 8543 11870
rect 11278 11732 11284 11796
rect 11348 11794 11354 11796
rect 11513 11794 11579 11797
rect 11348 11792 11579 11794
rect 11348 11736 11518 11792
rect 11574 11736 11579 11792
rect 11348 11734 11579 11736
rect 11654 11794 11714 11870
rect 12157 11928 13235 11930
rect 12157 11872 12162 11928
rect 12218 11872 13174 11928
rect 13230 11872 13235 11928
rect 12157 11870 13235 11872
rect 12157 11867 12223 11870
rect 13169 11867 13235 11870
rect 15561 11794 15627 11797
rect 11654 11792 15627 11794
rect 11654 11736 15566 11792
rect 15622 11736 15627 11792
rect 11654 11734 15627 11736
rect 11348 11732 11354 11734
rect 11513 11731 11579 11734
rect 15561 11731 15627 11734
rect 24761 11794 24827 11797
rect 30281 11794 30347 11797
rect 24761 11792 30347 11794
rect 24761 11736 24766 11792
rect 24822 11736 30286 11792
rect 30342 11736 30347 11792
rect 24761 11734 30347 11736
rect 24761 11731 24827 11734
rect 30281 11731 30347 11734
rect 6678 11596 6684 11660
rect 6748 11658 6754 11660
rect 12341 11658 12407 11661
rect 6748 11656 12407 11658
rect 6748 11600 12346 11656
rect 12402 11600 12407 11656
rect 6748 11598 12407 11600
rect 6748 11596 6754 11598
rect 12341 11595 12407 11598
rect 22277 11658 22343 11661
rect 30373 11658 30439 11661
rect 22277 11656 30439 11658
rect 22277 11600 22282 11656
rect 22338 11600 30378 11656
rect 30434 11600 30439 11656
rect 22277 11598 30439 11600
rect 22277 11595 22343 11598
rect 30373 11595 30439 11598
rect 3233 11522 3299 11525
rect 3877 11522 3943 11525
rect 3233 11520 3943 11522
rect 3233 11464 3238 11520
rect 3294 11464 3882 11520
rect 3938 11464 3943 11520
rect 3233 11462 3943 11464
rect 3233 11459 3299 11462
rect 3877 11459 3943 11462
rect 9857 11522 9923 11525
rect 12065 11522 12131 11525
rect 9857 11520 12131 11522
rect 9857 11464 9862 11520
rect 9918 11464 12070 11520
rect 12126 11464 12131 11520
rect 9857 11462 12131 11464
rect 9857 11459 9923 11462
rect 12065 11459 12131 11462
rect 13169 11522 13235 11525
rect 14089 11522 14155 11525
rect 13169 11520 14155 11522
rect 13169 11464 13174 11520
rect 13230 11464 14094 11520
rect 14150 11464 14155 11520
rect 13169 11462 14155 11464
rect 13169 11459 13235 11462
rect 14089 11459 14155 11462
rect 7984 11456 8300 11457
rect 7984 11392 7990 11456
rect 8054 11392 8070 11456
rect 8134 11392 8150 11456
rect 8214 11392 8230 11456
rect 8294 11392 8300 11456
rect 7984 11391 8300 11392
rect 15574 11456 15890 11457
rect 15574 11392 15580 11456
rect 15644 11392 15660 11456
rect 15724 11392 15740 11456
rect 15804 11392 15820 11456
rect 15884 11392 15890 11456
rect 15574 11391 15890 11392
rect 23164 11456 23480 11457
rect 23164 11392 23170 11456
rect 23234 11392 23250 11456
rect 23314 11392 23330 11456
rect 23394 11392 23410 11456
rect 23474 11392 23480 11456
rect 23164 11391 23480 11392
rect 30754 11456 31070 11457
rect 30754 11392 30760 11456
rect 30824 11392 30840 11456
rect 30904 11392 30920 11456
rect 30984 11392 31000 11456
rect 31064 11392 31070 11456
rect 30754 11391 31070 11392
rect 3417 11386 3483 11389
rect 4797 11386 4863 11389
rect 5625 11386 5691 11389
rect 6821 11386 6887 11389
rect 8661 11388 8727 11389
rect 8661 11386 8708 11388
rect 3417 11384 6887 11386
rect 3417 11328 3422 11384
rect 3478 11328 4802 11384
rect 4858 11328 5630 11384
rect 5686 11328 6826 11384
rect 6882 11328 6887 11384
rect 3417 11326 6887 11328
rect 8616 11384 8708 11386
rect 8616 11328 8666 11384
rect 8616 11326 8708 11328
rect 3417 11323 3483 11326
rect 4797 11323 4863 11326
rect 5625 11323 5691 11326
rect 6821 11323 6887 11326
rect 8661 11324 8708 11326
rect 8772 11324 8778 11388
rect 11053 11386 11119 11389
rect 13905 11386 13971 11389
rect 11053 11384 13971 11386
rect 11053 11328 11058 11384
rect 11114 11328 13910 11384
rect 13966 11328 13971 11384
rect 11053 11326 13971 11328
rect 8661 11323 8727 11324
rect 11053 11323 11119 11326
rect 13905 11323 13971 11326
rect 1945 11250 2011 11253
rect 24301 11250 24367 11253
rect 1945 11248 24367 11250
rect 1945 11192 1950 11248
rect 2006 11192 24306 11248
rect 24362 11192 24367 11248
rect 1945 11190 24367 11192
rect 1945 11187 2011 11190
rect 24301 11187 24367 11190
rect 4705 11114 4771 11117
rect 6545 11114 6611 11117
rect 4705 11112 6611 11114
rect 4705 11056 4710 11112
rect 4766 11056 6550 11112
rect 6606 11056 6611 11112
rect 4705 11054 6611 11056
rect 4705 11051 4771 11054
rect 6545 11051 6611 11054
rect 7046 11052 7052 11116
rect 7116 11114 7122 11116
rect 8753 11114 8819 11117
rect 7116 11112 8819 11114
rect 7116 11056 8758 11112
rect 8814 11056 8819 11112
rect 7116 11054 8819 11056
rect 7116 11052 7122 11054
rect 8753 11051 8819 11054
rect 9029 11114 9095 11117
rect 9949 11114 10015 11117
rect 9029 11112 10015 11114
rect 9029 11056 9034 11112
rect 9090 11056 9954 11112
rect 10010 11056 10015 11112
rect 9029 11054 10015 11056
rect 9029 11051 9095 11054
rect 9949 11051 10015 11054
rect 23841 11114 23907 11117
rect 26417 11114 26483 11117
rect 23841 11112 26483 11114
rect 23841 11056 23846 11112
rect 23902 11056 26422 11112
rect 26478 11056 26483 11112
rect 23841 11054 26483 11056
rect 23841 11051 23907 11054
rect 26417 11051 26483 11054
rect 1853 10978 1919 10981
rect 2998 10978 3004 10980
rect 1853 10976 3004 10978
rect 1853 10920 1858 10976
rect 1914 10920 3004 10976
rect 1853 10918 3004 10920
rect 1853 10915 1919 10918
rect 2998 10916 3004 10918
rect 3068 10916 3074 10980
rect 5349 10978 5415 10981
rect 8477 10978 8543 10981
rect 5349 10976 8543 10978
rect 5349 10920 5354 10976
rect 5410 10920 8482 10976
rect 8538 10920 8543 10976
rect 5349 10918 8543 10920
rect 5349 10915 5415 10918
rect 8477 10915 8543 10918
rect 4189 10912 4505 10913
rect 4189 10848 4195 10912
rect 4259 10848 4275 10912
rect 4339 10848 4355 10912
rect 4419 10848 4435 10912
rect 4499 10848 4505 10912
rect 4189 10847 4505 10848
rect 11779 10912 12095 10913
rect 11779 10848 11785 10912
rect 11849 10848 11865 10912
rect 11929 10848 11945 10912
rect 12009 10848 12025 10912
rect 12089 10848 12095 10912
rect 11779 10847 12095 10848
rect 19369 10912 19685 10913
rect 19369 10848 19375 10912
rect 19439 10848 19455 10912
rect 19519 10848 19535 10912
rect 19599 10848 19615 10912
rect 19679 10848 19685 10912
rect 19369 10847 19685 10848
rect 26959 10912 27275 10913
rect 26959 10848 26965 10912
rect 27029 10848 27045 10912
rect 27109 10848 27125 10912
rect 27189 10848 27205 10912
rect 27269 10848 27275 10912
rect 26959 10847 27275 10848
rect 9581 10842 9647 10845
rect 4616 10840 9647 10842
rect 4616 10784 9586 10840
rect 9642 10784 9647 10840
rect 4616 10782 9647 10784
rect 3601 10706 3667 10709
rect 4616 10706 4676 10782
rect 9581 10779 9647 10782
rect 3601 10704 4676 10706
rect 3601 10648 3606 10704
rect 3662 10648 4676 10704
rect 3601 10646 4676 10648
rect 5349 10706 5415 10709
rect 5809 10706 5875 10709
rect 5349 10704 5875 10706
rect 5349 10648 5354 10704
rect 5410 10648 5814 10704
rect 5870 10648 5875 10704
rect 5349 10646 5875 10648
rect 3601 10643 3667 10646
rect 5349 10643 5415 10646
rect 5809 10643 5875 10646
rect 6678 10644 6684 10708
rect 6748 10706 6754 10708
rect 16573 10706 16639 10709
rect 6748 10704 16639 10706
rect 6748 10648 16578 10704
rect 16634 10648 16639 10704
rect 6748 10646 16639 10648
rect 6748 10644 6754 10646
rect 16573 10643 16639 10646
rect 3969 10570 4035 10573
rect 15285 10570 15351 10573
rect 3969 10568 15351 10570
rect 3969 10512 3974 10568
rect 4030 10512 15290 10568
rect 15346 10512 15351 10568
rect 3969 10510 15351 10512
rect 3969 10507 4035 10510
rect 15285 10507 15351 10510
rect 8569 10434 8635 10437
rect 9213 10434 9279 10437
rect 8569 10432 9279 10434
rect 8569 10376 8574 10432
rect 8630 10376 9218 10432
rect 9274 10376 9279 10432
rect 8569 10374 9279 10376
rect 8569 10371 8635 10374
rect 9213 10371 9279 10374
rect 7984 10368 8300 10369
rect 7984 10304 7990 10368
rect 8054 10304 8070 10368
rect 8134 10304 8150 10368
rect 8214 10304 8230 10368
rect 8294 10304 8300 10368
rect 7984 10303 8300 10304
rect 15574 10368 15890 10369
rect 15574 10304 15580 10368
rect 15644 10304 15660 10368
rect 15724 10304 15740 10368
rect 15804 10304 15820 10368
rect 15884 10304 15890 10368
rect 15574 10303 15890 10304
rect 23164 10368 23480 10369
rect 23164 10304 23170 10368
rect 23234 10304 23250 10368
rect 23314 10304 23330 10368
rect 23394 10304 23410 10368
rect 23474 10304 23480 10368
rect 23164 10303 23480 10304
rect 30754 10368 31070 10369
rect 30754 10304 30760 10368
rect 30824 10304 30840 10368
rect 30904 10304 30920 10368
rect 30984 10304 31000 10368
rect 31064 10304 31070 10368
rect 30754 10303 31070 10304
rect 3693 10298 3759 10301
rect 3969 10298 4035 10301
rect 12985 10298 13051 10301
rect 3693 10296 4035 10298
rect 3693 10240 3698 10296
rect 3754 10240 3974 10296
rect 4030 10240 4035 10296
rect 3693 10238 4035 10240
rect 3693 10235 3759 10238
rect 3969 10235 4035 10238
rect 8526 10296 13051 10298
rect 8526 10240 12990 10296
rect 13046 10240 13051 10296
rect 8526 10238 13051 10240
rect 1485 10162 1551 10165
rect 8526 10162 8586 10238
rect 12985 10235 13051 10238
rect 17125 10298 17191 10301
rect 17902 10298 17908 10300
rect 17125 10296 17908 10298
rect 17125 10240 17130 10296
rect 17186 10240 17908 10296
rect 17125 10238 17908 10240
rect 17125 10235 17191 10238
rect 17902 10236 17908 10238
rect 17972 10236 17978 10300
rect 1485 10160 8586 10162
rect 1485 10104 1490 10160
rect 1546 10104 8586 10160
rect 1485 10102 8586 10104
rect 9213 10162 9279 10165
rect 16481 10162 16547 10165
rect 9213 10160 16547 10162
rect 9213 10104 9218 10160
rect 9274 10104 16486 10160
rect 16542 10104 16547 10160
rect 9213 10102 16547 10104
rect 1485 10099 1551 10102
rect 9213 10099 9279 10102
rect 16481 10099 16547 10102
rect 20437 10162 20503 10165
rect 21265 10162 21331 10165
rect 23749 10162 23815 10165
rect 20437 10160 23815 10162
rect 20437 10104 20442 10160
rect 20498 10104 21270 10160
rect 21326 10104 23754 10160
rect 23810 10104 23815 10160
rect 20437 10102 23815 10104
rect 20437 10099 20503 10102
rect 21265 10099 21331 10102
rect 23749 10099 23815 10102
rect 1669 10026 1735 10029
rect 13997 10026 14063 10029
rect 1669 10024 14063 10026
rect 1669 9968 1674 10024
rect 1730 9968 14002 10024
rect 14058 9968 14063 10024
rect 1669 9966 14063 9968
rect 1669 9963 1735 9966
rect 13997 9963 14063 9966
rect 5165 9890 5231 9893
rect 7005 9890 7071 9893
rect 5165 9888 7071 9890
rect 5165 9832 5170 9888
rect 5226 9832 7010 9888
rect 7066 9832 7071 9888
rect 5165 9830 7071 9832
rect 5165 9827 5231 9830
rect 7005 9827 7071 9830
rect 4189 9824 4505 9825
rect 4189 9760 4195 9824
rect 4259 9760 4275 9824
rect 4339 9760 4355 9824
rect 4419 9760 4435 9824
rect 4499 9760 4505 9824
rect 4189 9759 4505 9760
rect 11779 9824 12095 9825
rect 11779 9760 11785 9824
rect 11849 9760 11865 9824
rect 11929 9760 11945 9824
rect 12009 9760 12025 9824
rect 12089 9760 12095 9824
rect 11779 9759 12095 9760
rect 19369 9824 19685 9825
rect 19369 9760 19375 9824
rect 19439 9760 19455 9824
rect 19519 9760 19535 9824
rect 19599 9760 19615 9824
rect 19679 9760 19685 9824
rect 19369 9759 19685 9760
rect 26959 9824 27275 9825
rect 26959 9760 26965 9824
rect 27029 9760 27045 9824
rect 27109 9760 27125 9824
rect 27189 9760 27205 9824
rect 27269 9760 27275 9824
rect 26959 9759 27275 9760
rect 5349 9754 5415 9757
rect 6126 9754 6132 9756
rect 5349 9752 6132 9754
rect 5349 9696 5354 9752
rect 5410 9696 6132 9752
rect 5349 9694 6132 9696
rect 5349 9691 5415 9694
rect 6126 9692 6132 9694
rect 6196 9692 6202 9756
rect 6862 9692 6868 9756
rect 6932 9754 6938 9756
rect 7741 9754 7807 9757
rect 6932 9752 7807 9754
rect 6932 9696 7746 9752
rect 7802 9696 7807 9752
rect 6932 9694 7807 9696
rect 6932 9692 6938 9694
rect 7741 9691 7807 9694
rect 6310 9556 6316 9620
rect 6380 9618 6386 9620
rect 6637 9618 6703 9621
rect 6380 9616 6703 9618
rect 6380 9560 6642 9616
rect 6698 9560 6703 9616
rect 6380 9558 6703 9560
rect 6380 9556 6386 9558
rect 6637 9555 6703 9558
rect 7230 9556 7236 9620
rect 7300 9618 7306 9620
rect 16573 9618 16639 9621
rect 7300 9616 16639 9618
rect 7300 9560 16578 9616
rect 16634 9560 16639 9616
rect 7300 9558 16639 9560
rect 7300 9556 7306 9558
rect 16573 9555 16639 9558
rect 5022 9420 5028 9484
rect 5092 9482 5098 9484
rect 17585 9482 17651 9485
rect 5092 9480 17651 9482
rect 5092 9424 17590 9480
rect 17646 9424 17651 9480
rect 5092 9422 17651 9424
rect 5092 9420 5098 9422
rect 17585 9419 17651 9422
rect 21081 9482 21147 9485
rect 24117 9482 24183 9485
rect 21081 9480 24183 9482
rect 21081 9424 21086 9480
rect 21142 9424 24122 9480
rect 24178 9424 24183 9480
rect 21081 9422 24183 9424
rect 21081 9419 21147 9422
rect 24117 9419 24183 9422
rect 3417 9346 3483 9349
rect 4429 9346 4495 9349
rect 3417 9344 4495 9346
rect 3417 9288 3422 9344
rect 3478 9288 4434 9344
rect 4490 9288 4495 9344
rect 3417 9286 4495 9288
rect 3417 9283 3483 9286
rect 4429 9283 4495 9286
rect 5809 9346 5875 9349
rect 6545 9346 6611 9349
rect 5809 9344 6611 9346
rect 5809 9288 5814 9344
rect 5870 9288 6550 9344
rect 6606 9288 6611 9344
rect 5809 9286 6611 9288
rect 5809 9283 5875 9286
rect 6545 9283 6611 9286
rect 7984 9280 8300 9281
rect 7984 9216 7990 9280
rect 8054 9216 8070 9280
rect 8134 9216 8150 9280
rect 8214 9216 8230 9280
rect 8294 9216 8300 9280
rect 7984 9215 8300 9216
rect 15574 9280 15890 9281
rect 15574 9216 15580 9280
rect 15644 9216 15660 9280
rect 15724 9216 15740 9280
rect 15804 9216 15820 9280
rect 15884 9216 15890 9280
rect 15574 9215 15890 9216
rect 23164 9280 23480 9281
rect 23164 9216 23170 9280
rect 23234 9216 23250 9280
rect 23314 9216 23330 9280
rect 23394 9216 23410 9280
rect 23474 9216 23480 9280
rect 23164 9215 23480 9216
rect 30754 9280 31070 9281
rect 30754 9216 30760 9280
rect 30824 9216 30840 9280
rect 30904 9216 30920 9280
rect 30984 9216 31000 9280
rect 31064 9216 31070 9280
rect 30754 9215 31070 9216
rect 4521 9210 4587 9213
rect 7557 9210 7623 9213
rect 4521 9208 7623 9210
rect 4521 9152 4526 9208
rect 4582 9152 7562 9208
rect 7618 9152 7623 9208
rect 4521 9150 7623 9152
rect 4521 9147 4587 9150
rect 7557 9147 7623 9150
rect 1761 9074 1827 9077
rect 10409 9074 10475 9077
rect 1761 9072 10475 9074
rect 1761 9016 1766 9072
rect 1822 9016 10414 9072
rect 10470 9016 10475 9072
rect 1761 9014 10475 9016
rect 1761 9011 1827 9014
rect 10409 9011 10475 9014
rect 10593 9074 10659 9077
rect 12433 9074 12499 9077
rect 10593 9072 12499 9074
rect 10593 9016 10598 9072
rect 10654 9016 12438 9072
rect 12494 9016 12499 9072
rect 10593 9014 12499 9016
rect 10593 9011 10659 9014
rect 12433 9011 12499 9014
rect 22001 9074 22067 9077
rect 23749 9074 23815 9077
rect 22001 9072 23815 9074
rect 22001 9016 22006 9072
rect 22062 9016 23754 9072
rect 23810 9016 23815 9072
rect 22001 9014 23815 9016
rect 22001 9011 22067 9014
rect 23749 9011 23815 9014
rect 11145 8938 11211 8941
rect 12801 8938 12867 8941
rect 11145 8936 12867 8938
rect 11145 8880 11150 8936
rect 11206 8880 12806 8936
rect 12862 8880 12867 8936
rect 11145 8878 12867 8880
rect 11145 8875 11211 8878
rect 12801 8875 12867 8878
rect 18505 8938 18571 8941
rect 24710 8938 24716 8940
rect 18505 8936 24716 8938
rect 18505 8880 18510 8936
rect 18566 8880 24716 8936
rect 18505 8878 24716 8880
rect 18505 8875 18571 8878
rect 24710 8876 24716 8878
rect 24780 8876 24786 8940
rect 26785 8938 26851 8941
rect 26742 8936 26851 8938
rect 26742 8880 26790 8936
rect 26846 8880 26851 8936
rect 26742 8875 26851 8880
rect 22461 8802 22527 8805
rect 26742 8802 26802 8875
rect 22461 8800 26802 8802
rect 22461 8744 22466 8800
rect 22522 8744 26802 8800
rect 22461 8742 26802 8744
rect 22461 8739 22527 8742
rect 4189 8736 4505 8737
rect 4189 8672 4195 8736
rect 4259 8672 4275 8736
rect 4339 8672 4355 8736
rect 4419 8672 4435 8736
rect 4499 8672 4505 8736
rect 4189 8671 4505 8672
rect 11779 8736 12095 8737
rect 11779 8672 11785 8736
rect 11849 8672 11865 8736
rect 11929 8672 11945 8736
rect 12009 8672 12025 8736
rect 12089 8672 12095 8736
rect 11779 8671 12095 8672
rect 19369 8736 19685 8737
rect 19369 8672 19375 8736
rect 19439 8672 19455 8736
rect 19519 8672 19535 8736
rect 19599 8672 19615 8736
rect 19679 8672 19685 8736
rect 19369 8671 19685 8672
rect 7281 8666 7347 8669
rect 8661 8666 8727 8669
rect 7281 8664 8727 8666
rect 7281 8608 7286 8664
rect 7342 8608 8666 8664
rect 8722 8608 8727 8664
rect 7281 8606 8727 8608
rect 7281 8603 7347 8606
rect 8661 8603 8727 8606
rect 20897 8530 20963 8533
rect 24209 8530 24275 8533
rect 20897 8528 24275 8530
rect 20897 8472 20902 8528
rect 20958 8472 24214 8528
rect 24270 8472 24275 8528
rect 20897 8470 24275 8472
rect 20897 8467 20963 8470
rect 24209 8467 24275 8470
rect 26558 8397 26618 8742
rect 26959 8736 27275 8737
rect 26959 8672 26965 8736
rect 27029 8672 27045 8736
rect 27109 8672 27125 8736
rect 27189 8672 27205 8736
rect 27269 8672 27275 8736
rect 26959 8671 27275 8672
rect 2497 8394 2563 8397
rect 7557 8394 7623 8397
rect 2497 8392 7623 8394
rect 2497 8336 2502 8392
rect 2558 8336 7562 8392
rect 7618 8336 7623 8392
rect 2497 8334 7623 8336
rect 2497 8331 2563 8334
rect 7557 8331 7623 8334
rect 21357 8394 21423 8397
rect 22277 8394 22343 8397
rect 21357 8392 22343 8394
rect 21357 8336 21362 8392
rect 21418 8336 22282 8392
rect 22338 8336 22343 8392
rect 21357 8334 22343 8336
rect 21357 8331 21423 8334
rect 22277 8331 22343 8334
rect 26509 8392 26618 8397
rect 26509 8336 26514 8392
rect 26570 8336 26618 8392
rect 26509 8334 26618 8336
rect 26509 8331 26575 8334
rect 5809 8258 5875 8261
rect 5942 8258 5948 8260
rect 5809 8256 5948 8258
rect 5809 8200 5814 8256
rect 5870 8200 5948 8256
rect 5809 8198 5948 8200
rect 5809 8195 5875 8198
rect 5942 8196 5948 8198
rect 6012 8196 6018 8260
rect 7046 8196 7052 8260
rect 7116 8196 7122 8260
rect 10174 8196 10180 8260
rect 10244 8258 10250 8260
rect 11513 8258 11579 8261
rect 10244 8256 11579 8258
rect 10244 8200 11518 8256
rect 11574 8200 11579 8256
rect 10244 8198 11579 8200
rect 10244 8196 10250 8198
rect 3049 8122 3115 8125
rect 7054 8122 7114 8196
rect 11513 8195 11579 8198
rect 7984 8192 8300 8193
rect 7984 8128 7990 8192
rect 8054 8128 8070 8192
rect 8134 8128 8150 8192
rect 8214 8128 8230 8192
rect 8294 8128 8300 8192
rect 7984 8127 8300 8128
rect 15574 8192 15890 8193
rect 15574 8128 15580 8192
rect 15644 8128 15660 8192
rect 15724 8128 15740 8192
rect 15804 8128 15820 8192
rect 15884 8128 15890 8192
rect 15574 8127 15890 8128
rect 23164 8192 23480 8193
rect 23164 8128 23170 8192
rect 23234 8128 23250 8192
rect 23314 8128 23330 8192
rect 23394 8128 23410 8192
rect 23474 8128 23480 8192
rect 23164 8127 23480 8128
rect 30754 8192 31070 8193
rect 30754 8128 30760 8192
rect 30824 8128 30840 8192
rect 30904 8128 30920 8192
rect 30984 8128 31000 8192
rect 31064 8128 31070 8192
rect 30754 8127 31070 8128
rect 3049 8120 7114 8122
rect 3049 8064 3054 8120
rect 3110 8064 7114 8120
rect 3049 8062 7114 8064
rect 3049 8059 3115 8062
rect 6913 7986 6979 7989
rect 16389 7986 16455 7989
rect 16665 7986 16731 7989
rect 6913 7984 15946 7986
rect 6913 7928 6918 7984
rect 6974 7928 15946 7984
rect 6913 7926 15946 7928
rect 6913 7923 6979 7926
rect 1485 7850 1551 7853
rect 3509 7850 3575 7853
rect 1485 7848 3575 7850
rect 1485 7792 1490 7848
rect 1546 7792 3514 7848
rect 3570 7792 3575 7848
rect 1485 7790 3575 7792
rect 1485 7787 1551 7790
rect 3509 7787 3575 7790
rect 4153 7850 4219 7853
rect 7005 7850 7071 7853
rect 4153 7848 7071 7850
rect 4153 7792 4158 7848
rect 4214 7792 7010 7848
rect 7066 7792 7071 7848
rect 4153 7790 7071 7792
rect 4153 7787 4219 7790
rect 7005 7787 7071 7790
rect 9121 7850 9187 7853
rect 15653 7850 15719 7853
rect 9121 7848 15719 7850
rect 9121 7792 9126 7848
rect 9182 7792 15658 7848
rect 15714 7792 15719 7848
rect 9121 7790 15719 7792
rect 15886 7850 15946 7926
rect 16389 7984 16731 7986
rect 16389 7928 16394 7984
rect 16450 7928 16670 7984
rect 16726 7928 16731 7984
rect 16389 7926 16731 7928
rect 16389 7923 16455 7926
rect 16665 7923 16731 7926
rect 19701 7986 19767 7989
rect 26182 7986 26188 7988
rect 19701 7984 26188 7986
rect 19701 7928 19706 7984
rect 19762 7928 26188 7984
rect 19701 7926 26188 7928
rect 19701 7923 19767 7926
rect 26182 7924 26188 7926
rect 26252 7924 26258 7988
rect 16665 7850 16731 7853
rect 15886 7848 16731 7850
rect 15886 7792 16670 7848
rect 16726 7792 16731 7848
rect 15886 7790 16731 7792
rect 9121 7787 9187 7790
rect 15653 7787 15719 7790
rect 16665 7787 16731 7790
rect 6545 7714 6611 7717
rect 6545 7712 11530 7714
rect 6545 7656 6550 7712
rect 6606 7656 11530 7712
rect 6545 7654 11530 7656
rect 6545 7651 6611 7654
rect 4189 7648 4505 7649
rect 4189 7584 4195 7648
rect 4259 7584 4275 7648
rect 4339 7584 4355 7648
rect 4419 7584 4435 7648
rect 4499 7584 4505 7648
rect 4189 7583 4505 7584
rect 6085 7578 6151 7581
rect 5812 7576 6151 7578
rect 5812 7520 6090 7576
rect 6146 7520 6151 7576
rect 5812 7518 6151 7520
rect 5812 7445 5872 7518
rect 6085 7515 6151 7518
rect 6821 7578 6887 7581
rect 10501 7578 10567 7581
rect 6821 7576 10567 7578
rect 6821 7520 6826 7576
rect 6882 7520 10506 7576
rect 10562 7520 10567 7576
rect 6821 7518 10567 7520
rect 6821 7515 6887 7518
rect 10501 7515 10567 7518
rect 2681 7442 2747 7445
rect 5533 7442 5599 7445
rect 2681 7440 5599 7442
rect 2681 7384 2686 7440
rect 2742 7384 5538 7440
rect 5594 7384 5599 7440
rect 2681 7382 5599 7384
rect 2681 7379 2747 7382
rect 5533 7379 5599 7382
rect 5809 7440 5875 7445
rect 5809 7384 5814 7440
rect 5870 7384 5875 7440
rect 5809 7379 5875 7384
rect 5993 7442 6059 7445
rect 6862 7442 6868 7444
rect 5993 7440 6868 7442
rect 5993 7384 5998 7440
rect 6054 7384 6868 7440
rect 5993 7382 6868 7384
rect 5993 7379 6059 7382
rect 6862 7380 6868 7382
rect 6932 7380 6938 7444
rect 7005 7442 7071 7445
rect 11470 7442 11530 7654
rect 11779 7648 12095 7649
rect 11779 7584 11785 7648
rect 11849 7584 11865 7648
rect 11929 7584 11945 7648
rect 12009 7584 12025 7648
rect 12089 7584 12095 7648
rect 11779 7583 12095 7584
rect 19369 7648 19685 7649
rect 19369 7584 19375 7648
rect 19439 7584 19455 7648
rect 19519 7584 19535 7648
rect 19599 7584 19615 7648
rect 19679 7584 19685 7648
rect 19369 7583 19685 7584
rect 26959 7648 27275 7649
rect 26959 7584 26965 7648
rect 27029 7584 27045 7648
rect 27109 7584 27125 7648
rect 27189 7584 27205 7648
rect 27269 7584 27275 7648
rect 26959 7583 27275 7584
rect 14825 7578 14891 7581
rect 17309 7578 17375 7581
rect 14825 7576 17375 7578
rect 14825 7520 14830 7576
rect 14886 7520 17314 7576
rect 17370 7520 17375 7576
rect 14825 7518 17375 7520
rect 14825 7515 14891 7518
rect 17309 7515 17375 7518
rect 16297 7442 16363 7445
rect 7005 7440 11346 7442
rect 7005 7384 7010 7440
rect 7066 7384 11346 7440
rect 7005 7382 11346 7384
rect 11470 7440 16363 7442
rect 11470 7384 16302 7440
rect 16358 7384 16363 7440
rect 11470 7382 16363 7384
rect 7005 7379 7071 7382
rect 1761 7306 1827 7309
rect 11053 7306 11119 7309
rect 1761 7304 11119 7306
rect 1761 7248 1766 7304
rect 1822 7248 11058 7304
rect 11114 7248 11119 7304
rect 1761 7246 11119 7248
rect 11286 7306 11346 7382
rect 16297 7379 16363 7382
rect 17953 7306 18019 7309
rect 11286 7304 18019 7306
rect 11286 7248 17958 7304
rect 18014 7248 18019 7304
rect 11286 7246 18019 7248
rect 1761 7243 1827 7246
rect 11053 7243 11119 7246
rect 17953 7243 18019 7246
rect 18965 7306 19031 7309
rect 25773 7306 25839 7309
rect 18965 7304 25839 7306
rect 18965 7248 18970 7304
rect 19026 7248 25778 7304
rect 25834 7248 25839 7304
rect 18965 7246 25839 7248
rect 18965 7243 19031 7246
rect 25773 7243 25839 7246
rect 1117 7170 1183 7173
rect 6177 7170 6243 7173
rect 1117 7168 6243 7170
rect 1117 7112 1122 7168
rect 1178 7112 6182 7168
rect 6238 7112 6243 7168
rect 1117 7110 6243 7112
rect 1117 7107 1183 7110
rect 6177 7107 6243 7110
rect 9121 7170 9187 7173
rect 9949 7170 10015 7173
rect 9121 7168 10015 7170
rect 9121 7112 9126 7168
rect 9182 7112 9954 7168
rect 10010 7112 10015 7168
rect 9121 7110 10015 7112
rect 9121 7107 9187 7110
rect 9949 7107 10015 7110
rect 16798 7108 16804 7172
rect 16868 7170 16874 7172
rect 17217 7170 17283 7173
rect 16868 7168 17283 7170
rect 16868 7112 17222 7168
rect 17278 7112 17283 7168
rect 16868 7110 17283 7112
rect 16868 7108 16874 7110
rect 17217 7107 17283 7110
rect 7984 7104 8300 7105
rect 7984 7040 7990 7104
rect 8054 7040 8070 7104
rect 8134 7040 8150 7104
rect 8214 7040 8230 7104
rect 8294 7040 8300 7104
rect 7984 7039 8300 7040
rect 15574 7104 15890 7105
rect 15574 7040 15580 7104
rect 15644 7040 15660 7104
rect 15724 7040 15740 7104
rect 15804 7040 15820 7104
rect 15884 7040 15890 7104
rect 15574 7039 15890 7040
rect 23164 7104 23480 7105
rect 23164 7040 23170 7104
rect 23234 7040 23250 7104
rect 23314 7040 23330 7104
rect 23394 7040 23410 7104
rect 23474 7040 23480 7104
rect 23164 7039 23480 7040
rect 30754 7104 31070 7105
rect 30754 7040 30760 7104
rect 30824 7040 30840 7104
rect 30904 7040 30920 7104
rect 30984 7040 31000 7104
rect 31064 7040 31070 7104
rect 30754 7039 31070 7040
rect 6126 6972 6132 7036
rect 6196 7034 6202 7036
rect 7097 7034 7163 7037
rect 6196 7032 7163 7034
rect 6196 6976 7102 7032
rect 7158 6976 7163 7032
rect 6196 6974 7163 6976
rect 6196 6972 6202 6974
rect 7097 6971 7163 6974
rect 16614 6972 16620 7036
rect 16684 7034 16690 7036
rect 17493 7034 17559 7037
rect 25037 7034 25103 7037
rect 16684 7032 17559 7034
rect 16684 6976 17498 7032
rect 17554 6976 17559 7032
rect 16684 6974 17559 6976
rect 16684 6972 16690 6974
rect 17493 6971 17559 6974
rect 24902 7032 25103 7034
rect 24902 6976 25042 7032
rect 25098 6976 25103 7032
rect 24902 6974 25103 6976
rect 2313 6898 2379 6901
rect 4153 6898 4219 6901
rect 2313 6896 4219 6898
rect 2313 6840 2318 6896
rect 2374 6840 4158 6896
rect 4214 6840 4219 6896
rect 2313 6838 4219 6840
rect 2313 6835 2379 6838
rect 4153 6835 4219 6838
rect 6913 6898 6979 6901
rect 19149 6898 19215 6901
rect 24902 6898 24962 6974
rect 25037 6971 25103 6974
rect 6913 6896 16498 6898
rect 6913 6840 6918 6896
rect 6974 6840 16498 6896
rect 6913 6838 16498 6840
rect 6913 6835 6979 6838
rect 3141 6762 3207 6765
rect 6678 6762 6684 6764
rect 3141 6760 6684 6762
rect 3141 6704 3146 6760
rect 3202 6704 6684 6760
rect 3141 6702 6684 6704
rect 3141 6699 3207 6702
rect 6678 6700 6684 6702
rect 6748 6700 6754 6764
rect 9121 6762 9187 6765
rect 16205 6762 16271 6765
rect 9121 6760 16271 6762
rect 9121 6704 9126 6760
rect 9182 6704 16210 6760
rect 16266 6704 16271 6760
rect 9121 6702 16271 6704
rect 9121 6699 9187 6702
rect 16205 6699 16271 6702
rect 4189 6560 4505 6561
rect 4189 6496 4195 6560
rect 4259 6496 4275 6560
rect 4339 6496 4355 6560
rect 4419 6496 4435 6560
rect 4499 6496 4505 6560
rect 4189 6495 4505 6496
rect 11779 6560 12095 6561
rect 11779 6496 11785 6560
rect 11849 6496 11865 6560
rect 11929 6496 11945 6560
rect 12009 6496 12025 6560
rect 12089 6496 12095 6560
rect 11779 6495 12095 6496
rect 5257 6490 5323 6493
rect 7465 6490 7531 6493
rect 5257 6488 7531 6490
rect 5257 6432 5262 6488
rect 5318 6432 7470 6488
rect 7526 6432 7531 6488
rect 5257 6430 7531 6432
rect 16438 6490 16498 6838
rect 19149 6896 24962 6898
rect 19149 6840 19154 6896
rect 19210 6840 24962 6896
rect 19149 6838 24962 6840
rect 19149 6835 19215 6838
rect 19369 6560 19685 6561
rect 19369 6496 19375 6560
rect 19439 6496 19455 6560
rect 19519 6496 19535 6560
rect 19599 6496 19615 6560
rect 19679 6496 19685 6560
rect 19369 6495 19685 6496
rect 26959 6560 27275 6561
rect 26959 6496 26965 6560
rect 27029 6496 27045 6560
rect 27109 6496 27125 6560
rect 27189 6496 27205 6560
rect 27269 6496 27275 6560
rect 26959 6495 27275 6496
rect 16665 6490 16731 6493
rect 16438 6488 16731 6490
rect 16438 6432 16670 6488
rect 16726 6432 16731 6488
rect 16438 6430 16731 6432
rect 5257 6427 5323 6430
rect 7465 6427 7531 6430
rect 16665 6427 16731 6430
rect 21817 6490 21883 6493
rect 24393 6490 24459 6493
rect 21817 6488 24459 6490
rect 21817 6432 21822 6488
rect 21878 6432 24398 6488
rect 24454 6432 24459 6488
rect 21817 6430 24459 6432
rect 21817 6427 21883 6430
rect 24393 6427 24459 6430
rect 1577 6354 1643 6357
rect 3969 6354 4035 6357
rect 1577 6352 4035 6354
rect 1577 6296 1582 6352
rect 1638 6296 3974 6352
rect 4030 6296 4035 6352
rect 1577 6294 4035 6296
rect 1577 6291 1643 6294
rect 3969 6291 4035 6294
rect 11421 6354 11487 6357
rect 17401 6354 17467 6357
rect 11421 6352 17467 6354
rect 11421 6296 11426 6352
rect 11482 6296 17406 6352
rect 17462 6296 17467 6352
rect 11421 6294 17467 6296
rect 11421 6291 11487 6294
rect 17401 6291 17467 6294
rect 18781 6354 18847 6357
rect 26233 6354 26299 6357
rect 18781 6352 26299 6354
rect 18781 6296 18786 6352
rect 18842 6296 26238 6352
rect 26294 6296 26299 6352
rect 18781 6294 26299 6296
rect 18781 6291 18847 6294
rect 26233 6291 26299 6294
rect 5625 6218 5691 6221
rect 7649 6218 7715 6221
rect 5625 6216 7715 6218
rect 5625 6160 5630 6216
rect 5686 6160 7654 6216
rect 7710 6160 7715 6216
rect 5625 6158 7715 6160
rect 5625 6155 5691 6158
rect 7649 6155 7715 6158
rect 20621 6218 20687 6221
rect 28625 6218 28691 6221
rect 20621 6216 28691 6218
rect 20621 6160 20626 6216
rect 20682 6160 28630 6216
rect 28686 6160 28691 6216
rect 20621 6158 28691 6160
rect 20621 6155 20687 6158
rect 28625 6155 28691 6158
rect 2681 6082 2747 6085
rect 6729 6082 6795 6085
rect 2681 6080 6795 6082
rect 2681 6024 2686 6080
rect 2742 6024 6734 6080
rect 6790 6024 6795 6080
rect 2681 6022 6795 6024
rect 2681 6019 2747 6022
rect 6729 6019 6795 6022
rect 7984 6016 8300 6017
rect 7984 5952 7990 6016
rect 8054 5952 8070 6016
rect 8134 5952 8150 6016
rect 8214 5952 8230 6016
rect 8294 5952 8300 6016
rect 7984 5951 8300 5952
rect 15574 6016 15890 6017
rect 15574 5952 15580 6016
rect 15644 5952 15660 6016
rect 15724 5952 15740 6016
rect 15804 5952 15820 6016
rect 15884 5952 15890 6016
rect 15574 5951 15890 5952
rect 23164 6016 23480 6017
rect 23164 5952 23170 6016
rect 23234 5952 23250 6016
rect 23314 5952 23330 6016
rect 23394 5952 23410 6016
rect 23474 5952 23480 6016
rect 23164 5951 23480 5952
rect 30754 6016 31070 6017
rect 30754 5952 30760 6016
rect 30824 5952 30840 6016
rect 30904 5952 30920 6016
rect 30984 5952 31000 6016
rect 31064 5952 31070 6016
rect 30754 5951 31070 5952
rect 12249 5810 12315 5813
rect 12433 5810 12499 5813
rect 12249 5808 12499 5810
rect 12249 5752 12254 5808
rect 12310 5752 12438 5808
rect 12494 5752 12499 5808
rect 12249 5750 12499 5752
rect 12249 5747 12315 5750
rect 12433 5747 12499 5750
rect 21541 5810 21607 5813
rect 27613 5810 27679 5813
rect 21541 5808 27679 5810
rect 21541 5752 21546 5808
rect 21602 5752 27618 5808
rect 27674 5752 27679 5808
rect 21541 5750 27679 5752
rect 21541 5747 21607 5750
rect 27613 5747 27679 5750
rect 2497 5674 2563 5677
rect 5533 5674 5599 5677
rect 2497 5672 5599 5674
rect 2497 5616 2502 5672
rect 2558 5616 5538 5672
rect 5594 5616 5599 5672
rect 2497 5614 5599 5616
rect 2497 5611 2563 5614
rect 5533 5611 5599 5614
rect 6177 5674 6243 5677
rect 7557 5674 7623 5677
rect 11329 5674 11395 5677
rect 6177 5672 11395 5674
rect 6177 5616 6182 5672
rect 6238 5616 7562 5672
rect 7618 5616 11334 5672
rect 11390 5616 11395 5672
rect 6177 5614 11395 5616
rect 6177 5611 6243 5614
rect 7557 5611 7623 5614
rect 11329 5611 11395 5614
rect 23565 5674 23631 5677
rect 24669 5674 24735 5677
rect 23565 5672 24735 5674
rect 23565 5616 23570 5672
rect 23626 5616 24674 5672
rect 24730 5616 24735 5672
rect 23565 5614 24735 5616
rect 23565 5611 23631 5614
rect 24669 5611 24735 5614
rect 2998 5476 3004 5540
rect 3068 5538 3074 5540
rect 3141 5538 3207 5541
rect 3068 5536 3207 5538
rect 3068 5480 3146 5536
rect 3202 5480 3207 5536
rect 3068 5478 3207 5480
rect 3068 5476 3074 5478
rect 3141 5475 3207 5478
rect 5073 5538 5139 5541
rect 6913 5538 6979 5541
rect 5073 5536 6979 5538
rect 5073 5480 5078 5536
rect 5134 5480 6918 5536
rect 6974 5480 6979 5536
rect 5073 5478 6979 5480
rect 5073 5475 5139 5478
rect 6913 5475 6979 5478
rect 8518 5476 8524 5540
rect 8588 5538 8594 5540
rect 10685 5538 10751 5541
rect 8588 5536 10751 5538
rect 8588 5480 10690 5536
rect 10746 5480 10751 5536
rect 8588 5478 10751 5480
rect 8588 5476 8594 5478
rect 10685 5475 10751 5478
rect 22645 5538 22711 5541
rect 25865 5538 25931 5541
rect 22645 5536 25931 5538
rect 22645 5480 22650 5536
rect 22706 5480 25870 5536
rect 25926 5480 25931 5536
rect 22645 5478 25931 5480
rect 22645 5475 22711 5478
rect 25865 5475 25931 5478
rect 26182 5476 26188 5540
rect 26252 5538 26258 5540
rect 26325 5538 26391 5541
rect 26252 5536 26391 5538
rect 26252 5480 26330 5536
rect 26386 5480 26391 5536
rect 26252 5478 26391 5480
rect 26252 5476 26258 5478
rect 26325 5475 26391 5478
rect 4189 5472 4505 5473
rect 4189 5408 4195 5472
rect 4259 5408 4275 5472
rect 4339 5408 4355 5472
rect 4419 5408 4435 5472
rect 4499 5408 4505 5472
rect 4189 5407 4505 5408
rect 11779 5472 12095 5473
rect 11779 5408 11785 5472
rect 11849 5408 11865 5472
rect 11929 5408 11945 5472
rect 12009 5408 12025 5472
rect 12089 5408 12095 5472
rect 11779 5407 12095 5408
rect 19369 5472 19685 5473
rect 19369 5408 19375 5472
rect 19439 5408 19455 5472
rect 19519 5408 19535 5472
rect 19599 5408 19615 5472
rect 19679 5408 19685 5472
rect 19369 5407 19685 5408
rect 26959 5472 27275 5473
rect 26959 5408 26965 5472
rect 27029 5408 27045 5472
rect 27109 5408 27125 5472
rect 27189 5408 27205 5472
rect 27269 5408 27275 5472
rect 26959 5407 27275 5408
rect 1393 5402 1459 5405
rect 3969 5402 4035 5405
rect 1393 5400 4035 5402
rect 1393 5344 1398 5400
rect 1454 5344 3974 5400
rect 4030 5344 4035 5400
rect 1393 5342 4035 5344
rect 1393 5339 1459 5342
rect 3969 5339 4035 5342
rect 13445 5402 13511 5405
rect 16941 5402 17007 5405
rect 13445 5400 17007 5402
rect 13445 5344 13450 5400
rect 13506 5344 16946 5400
rect 17002 5344 17007 5400
rect 13445 5342 17007 5344
rect 13445 5339 13511 5342
rect 16941 5339 17007 5342
rect 3417 5266 3483 5269
rect 6729 5266 6795 5269
rect 3417 5264 6795 5266
rect 3417 5208 3422 5264
rect 3478 5208 6734 5264
rect 6790 5208 6795 5264
rect 3417 5206 6795 5208
rect 3417 5203 3483 5206
rect 6729 5203 6795 5206
rect 13261 5266 13327 5269
rect 23381 5266 23447 5269
rect 13261 5264 23447 5266
rect 13261 5208 13266 5264
rect 13322 5208 23386 5264
rect 23442 5208 23447 5264
rect 13261 5206 23447 5208
rect 13261 5203 13327 5206
rect 23381 5203 23447 5206
rect 23657 5266 23723 5269
rect 27337 5266 27403 5269
rect 23657 5264 27403 5266
rect 23657 5208 23662 5264
rect 23718 5208 27342 5264
rect 27398 5208 27403 5264
rect 23657 5206 27403 5208
rect 23657 5203 23723 5206
rect 27337 5203 27403 5206
rect 2129 5130 2195 5133
rect 15285 5130 15351 5133
rect 2129 5128 15351 5130
rect 2129 5072 2134 5128
rect 2190 5072 15290 5128
rect 15346 5072 15351 5128
rect 2129 5070 15351 5072
rect 2129 5067 2195 5070
rect 15285 5067 15351 5070
rect 17769 5130 17835 5133
rect 28717 5130 28783 5133
rect 17769 5128 28783 5130
rect 17769 5072 17774 5128
rect 17830 5072 28722 5128
rect 28778 5072 28783 5128
rect 17769 5070 28783 5072
rect 17769 5067 17835 5070
rect 28717 5067 28783 5070
rect 2865 4994 2931 4997
rect 4429 4994 4495 4997
rect 5165 4994 5231 4997
rect 2865 4992 5231 4994
rect 2865 4936 2870 4992
rect 2926 4936 4434 4992
rect 4490 4936 5170 4992
rect 5226 4936 5231 4992
rect 2865 4934 5231 4936
rect 2865 4931 2931 4934
rect 4429 4931 4495 4934
rect 5165 4931 5231 4934
rect 7984 4928 8300 4929
rect 7984 4864 7990 4928
rect 8054 4864 8070 4928
rect 8134 4864 8150 4928
rect 8214 4864 8230 4928
rect 8294 4864 8300 4928
rect 7984 4863 8300 4864
rect 15574 4928 15890 4929
rect 15574 4864 15580 4928
rect 15644 4864 15660 4928
rect 15724 4864 15740 4928
rect 15804 4864 15820 4928
rect 15884 4864 15890 4928
rect 15574 4863 15890 4864
rect 23164 4928 23480 4929
rect 23164 4864 23170 4928
rect 23234 4864 23250 4928
rect 23314 4864 23330 4928
rect 23394 4864 23410 4928
rect 23474 4864 23480 4928
rect 23164 4863 23480 4864
rect 30754 4928 31070 4929
rect 30754 4864 30760 4928
rect 30824 4864 30840 4928
rect 30904 4864 30920 4928
rect 30984 4864 31000 4928
rect 31064 4864 31070 4928
rect 30754 4863 31070 4864
rect 2313 4858 2379 4861
rect 6453 4858 6519 4861
rect 2313 4856 6519 4858
rect 2313 4800 2318 4856
rect 2374 4800 6458 4856
rect 6514 4800 6519 4856
rect 2313 4798 6519 4800
rect 2313 4795 2379 4798
rect 6453 4795 6519 4798
rect 5073 4722 5139 4725
rect 16614 4722 16620 4724
rect 5073 4720 16620 4722
rect 5073 4664 5078 4720
rect 5134 4664 16620 4720
rect 5073 4662 16620 4664
rect 5073 4659 5139 4662
rect 16614 4660 16620 4662
rect 16684 4660 16690 4724
rect 20897 4722 20963 4725
rect 24853 4722 24919 4725
rect 20897 4720 24919 4722
rect 20897 4664 20902 4720
rect 20958 4664 24858 4720
rect 24914 4664 24919 4720
rect 20897 4662 24919 4664
rect 20897 4659 20963 4662
rect 24853 4659 24919 4662
rect 4705 4586 4771 4589
rect 16798 4586 16804 4588
rect 4705 4584 16804 4586
rect 4705 4528 4710 4584
rect 4766 4528 16804 4584
rect 4705 4526 16804 4528
rect 4705 4523 4771 4526
rect 16798 4524 16804 4526
rect 16868 4524 16874 4588
rect 20069 4586 20135 4589
rect 27613 4586 27679 4589
rect 20069 4584 27679 4586
rect 20069 4528 20074 4584
rect 20130 4528 27618 4584
rect 27674 4528 27679 4584
rect 20069 4526 27679 4528
rect 20069 4523 20135 4526
rect 27613 4523 27679 4526
rect 22001 4450 22067 4453
rect 22829 4450 22895 4453
rect 24577 4450 24643 4453
rect 22001 4448 24643 4450
rect 22001 4392 22006 4448
rect 22062 4392 22834 4448
rect 22890 4392 24582 4448
rect 24638 4392 24643 4448
rect 22001 4390 24643 4392
rect 22001 4387 22067 4390
rect 22829 4387 22895 4390
rect 24577 4387 24643 4390
rect 4189 4384 4505 4385
rect 4189 4320 4195 4384
rect 4259 4320 4275 4384
rect 4339 4320 4355 4384
rect 4419 4320 4435 4384
rect 4499 4320 4505 4384
rect 4189 4319 4505 4320
rect 11779 4384 12095 4385
rect 11779 4320 11785 4384
rect 11849 4320 11865 4384
rect 11929 4320 11945 4384
rect 12009 4320 12025 4384
rect 12089 4320 12095 4384
rect 11779 4319 12095 4320
rect 19369 4384 19685 4385
rect 19369 4320 19375 4384
rect 19439 4320 19455 4384
rect 19519 4320 19535 4384
rect 19599 4320 19615 4384
rect 19679 4320 19685 4384
rect 19369 4319 19685 4320
rect 26959 4384 27275 4385
rect 26959 4320 26965 4384
rect 27029 4320 27045 4384
rect 27109 4320 27125 4384
rect 27189 4320 27205 4384
rect 27269 4320 27275 4384
rect 26959 4319 27275 4320
rect 22050 4254 22570 4314
rect 16389 4178 16455 4181
rect 9630 4176 16455 4178
rect 9630 4120 16394 4176
rect 16450 4120 16455 4176
rect 9630 4118 16455 4120
rect 2773 4044 2839 4045
rect 2773 4040 2820 4044
rect 2884 4042 2890 4044
rect 4797 4042 4863 4045
rect 9630 4042 9690 4118
rect 16389 4115 16455 4118
rect 17902 4116 17908 4180
rect 17972 4178 17978 4180
rect 22050 4178 22110 4254
rect 17972 4118 22110 4178
rect 22277 4178 22343 4181
rect 22510 4178 22570 4254
rect 27705 4178 27771 4181
rect 22277 4176 22386 4178
rect 22277 4120 22282 4176
rect 22338 4120 22386 4176
rect 17972 4116 17978 4118
rect 22277 4115 22386 4120
rect 22510 4176 27771 4178
rect 22510 4120 27710 4176
rect 27766 4120 27771 4176
rect 22510 4118 27771 4120
rect 27705 4115 27771 4118
rect 2773 3984 2778 4040
rect 2773 3980 2820 3984
rect 2884 3982 2930 4042
rect 4797 4040 9690 4042
rect 4797 3984 4802 4040
rect 4858 3984 9690 4040
rect 4797 3982 9690 3984
rect 13629 4042 13695 4045
rect 14457 4042 14523 4045
rect 13629 4040 14523 4042
rect 13629 3984 13634 4040
rect 13690 3984 14462 4040
rect 14518 3984 14523 4040
rect 13629 3982 14523 3984
rect 2884 3980 2890 3982
rect 2773 3979 2839 3980
rect 4797 3979 4863 3982
rect 13629 3979 13695 3982
rect 14457 3979 14523 3982
rect 3325 3906 3391 3909
rect 7230 3906 7236 3908
rect 3325 3904 7236 3906
rect 3325 3848 3330 3904
rect 3386 3848 7236 3904
rect 3325 3846 7236 3848
rect 3325 3843 3391 3846
rect 7230 3844 7236 3846
rect 7300 3844 7306 3908
rect 11145 3906 11211 3909
rect 12249 3906 12315 3909
rect 11145 3904 12315 3906
rect 11145 3848 11150 3904
rect 11206 3848 12254 3904
rect 12310 3848 12315 3904
rect 11145 3846 12315 3848
rect 11145 3843 11211 3846
rect 12249 3843 12315 3846
rect 7984 3840 8300 3841
rect 7984 3776 7990 3840
rect 8054 3776 8070 3840
rect 8134 3776 8150 3840
rect 8214 3776 8230 3840
rect 8294 3776 8300 3840
rect 7984 3775 8300 3776
rect 15574 3840 15890 3841
rect 15574 3776 15580 3840
rect 15644 3776 15660 3840
rect 15724 3776 15740 3840
rect 15804 3776 15820 3840
rect 15884 3776 15890 3840
rect 15574 3775 15890 3776
rect 16392 3770 16452 4115
rect 20621 4042 20687 4045
rect 22326 4042 22386 4115
rect 20621 4040 22386 4042
rect 20621 3984 20626 4040
rect 20682 3984 22386 4040
rect 20621 3982 22386 3984
rect 20621 3979 20687 3982
rect 24710 3980 24716 4044
rect 24780 4042 24786 4044
rect 28533 4042 28599 4045
rect 24780 4040 28599 4042
rect 24780 3984 28538 4040
rect 28594 3984 28599 4040
rect 24780 3982 28599 3984
rect 24780 3980 24786 3982
rect 28533 3979 28599 3982
rect 23164 3840 23480 3841
rect 23164 3776 23170 3840
rect 23234 3776 23250 3840
rect 23314 3776 23330 3840
rect 23394 3776 23410 3840
rect 23474 3776 23480 3840
rect 23164 3775 23480 3776
rect 30754 3840 31070 3841
rect 30754 3776 30760 3840
rect 30824 3776 30840 3840
rect 30904 3776 30920 3840
rect 30984 3776 31000 3840
rect 31064 3776 31070 3840
rect 30754 3775 31070 3776
rect 19057 3770 19123 3773
rect 16392 3768 19350 3770
rect 16392 3712 19062 3768
rect 19118 3712 19350 3768
rect 16392 3710 19350 3712
rect 19057 3707 19123 3710
rect 4245 3634 4311 3637
rect 17861 3634 17927 3637
rect 4245 3632 17927 3634
rect 4245 3576 4250 3632
rect 4306 3576 17866 3632
rect 17922 3576 17927 3632
rect 4245 3574 17927 3576
rect 19290 3634 19350 3710
rect 25129 3634 25195 3637
rect 19290 3632 25195 3634
rect 19290 3576 25134 3632
rect 25190 3576 25195 3632
rect 19290 3574 25195 3576
rect 4245 3571 4311 3574
rect 17861 3571 17927 3574
rect 25129 3571 25195 3574
rect 5625 3498 5691 3501
rect 27889 3498 27955 3501
rect 5625 3496 27955 3498
rect 5625 3440 5630 3496
rect 5686 3440 27894 3496
rect 27950 3440 27955 3496
rect 5625 3438 27955 3440
rect 5625 3435 5691 3438
rect 27889 3435 27955 3438
rect 16849 3362 16915 3365
rect 12390 3360 16915 3362
rect 12390 3304 16854 3360
rect 16910 3304 16915 3360
rect 12390 3302 16915 3304
rect 4189 3296 4505 3297
rect 4189 3232 4195 3296
rect 4259 3232 4275 3296
rect 4339 3232 4355 3296
rect 4419 3232 4435 3296
rect 4499 3232 4505 3296
rect 4189 3231 4505 3232
rect 11779 3296 12095 3297
rect 11779 3232 11785 3296
rect 11849 3232 11865 3296
rect 11929 3232 11945 3296
rect 12009 3232 12025 3296
rect 12089 3232 12095 3296
rect 11779 3231 12095 3232
rect 7281 3226 7347 3229
rect 11145 3226 11211 3229
rect 7281 3224 11211 3226
rect 7281 3168 7286 3224
rect 7342 3168 11150 3224
rect 11206 3168 11211 3224
rect 7281 3166 11211 3168
rect 7281 3163 7347 3166
rect 11145 3163 11211 3166
rect 1669 3090 1735 3093
rect 8518 3090 8524 3092
rect 1669 3088 8524 3090
rect 1669 3032 1674 3088
rect 1730 3032 8524 3088
rect 1669 3030 8524 3032
rect 1669 3027 1735 3030
rect 8518 3028 8524 3030
rect 8588 3028 8594 3092
rect 9213 3090 9279 3093
rect 12249 3090 12315 3093
rect 12390 3090 12450 3302
rect 16849 3299 16915 3302
rect 19369 3296 19685 3297
rect 19369 3232 19375 3296
rect 19439 3232 19455 3296
rect 19519 3232 19535 3296
rect 19599 3232 19615 3296
rect 19679 3232 19685 3296
rect 19369 3231 19685 3232
rect 26959 3296 27275 3297
rect 26959 3232 26965 3296
rect 27029 3232 27045 3296
rect 27109 3232 27125 3296
rect 27189 3232 27205 3296
rect 27269 3232 27275 3296
rect 26959 3231 27275 3232
rect 9213 3088 12450 3090
rect 9213 3032 9218 3088
rect 9274 3032 12254 3088
rect 12310 3032 12450 3088
rect 9213 3030 12450 3032
rect 15101 3090 15167 3093
rect 22737 3090 22803 3093
rect 15101 3088 22803 3090
rect 15101 3032 15106 3088
rect 15162 3032 22742 3088
rect 22798 3032 22803 3088
rect 15101 3030 22803 3032
rect 9213 3027 9279 3030
rect 12249 3027 12315 3030
rect 15101 3027 15167 3030
rect 22737 3027 22803 3030
rect 3877 2954 3943 2957
rect 18689 2954 18755 2957
rect 27061 2954 27127 2957
rect 3877 2952 18755 2954
rect 3877 2896 3882 2952
rect 3938 2896 18694 2952
rect 18750 2896 18755 2952
rect 3877 2894 18755 2896
rect 3877 2891 3943 2894
rect 18689 2891 18755 2894
rect 22050 2952 27127 2954
rect 22050 2896 27066 2952
rect 27122 2896 27127 2952
rect 22050 2894 27127 2896
rect 16757 2818 16823 2821
rect 22050 2818 22110 2894
rect 27061 2891 27127 2894
rect 16757 2816 22110 2818
rect 16757 2760 16762 2816
rect 16818 2760 22110 2816
rect 16757 2758 22110 2760
rect 16757 2755 16823 2758
rect 7984 2752 8300 2753
rect 7984 2688 7990 2752
rect 8054 2688 8070 2752
rect 8134 2688 8150 2752
rect 8214 2688 8230 2752
rect 8294 2688 8300 2752
rect 7984 2687 8300 2688
rect 15574 2752 15890 2753
rect 15574 2688 15580 2752
rect 15644 2688 15660 2752
rect 15724 2688 15740 2752
rect 15804 2688 15820 2752
rect 15884 2688 15890 2752
rect 15574 2687 15890 2688
rect 23164 2752 23480 2753
rect 23164 2688 23170 2752
rect 23234 2688 23250 2752
rect 23314 2688 23330 2752
rect 23394 2688 23410 2752
rect 23474 2688 23480 2752
rect 23164 2687 23480 2688
rect 30754 2752 31070 2753
rect 30754 2688 30760 2752
rect 30824 2688 30840 2752
rect 30904 2688 30920 2752
rect 30984 2688 31000 2752
rect 31064 2688 31070 2752
rect 30754 2687 31070 2688
rect 1853 2546 1919 2549
rect 5022 2546 5028 2548
rect 1853 2544 5028 2546
rect 1853 2488 1858 2544
rect 1914 2488 5028 2544
rect 1853 2486 5028 2488
rect 1853 2483 1919 2486
rect 5022 2484 5028 2486
rect 5092 2484 5098 2548
rect 10593 2546 10659 2549
rect 14457 2546 14523 2549
rect 10593 2544 14523 2546
rect 10593 2488 10598 2544
rect 10654 2488 14462 2544
rect 14518 2488 14523 2544
rect 10593 2486 14523 2488
rect 10593 2483 10659 2486
rect 14457 2483 14523 2486
rect 3969 2412 4035 2413
rect 3918 2410 3924 2412
rect 3878 2350 3924 2410
rect 3988 2408 4035 2412
rect 4030 2352 4035 2408
rect 3918 2348 3924 2350
rect 3988 2348 4035 2352
rect 3969 2347 4035 2348
rect 5993 2410 6059 2413
rect 7833 2410 7899 2413
rect 5993 2408 7899 2410
rect 5993 2352 5998 2408
rect 6054 2352 7838 2408
rect 7894 2352 7899 2408
rect 5993 2350 7899 2352
rect 5993 2347 6059 2350
rect 7833 2347 7899 2350
rect 17953 2410 18019 2413
rect 18781 2410 18847 2413
rect 17953 2408 18847 2410
rect 17953 2352 17958 2408
rect 18014 2352 18786 2408
rect 18842 2352 18847 2408
rect 17953 2350 18847 2352
rect 17953 2347 18019 2350
rect 18781 2347 18847 2350
rect 23657 2274 23723 2277
rect 26417 2274 26483 2277
rect 23657 2272 26483 2274
rect 23657 2216 23662 2272
rect 23718 2216 26422 2272
rect 26478 2216 26483 2272
rect 23657 2214 26483 2216
rect 23657 2211 23723 2214
rect 26417 2211 26483 2214
rect 4189 2208 4505 2209
rect 4189 2144 4195 2208
rect 4259 2144 4275 2208
rect 4339 2144 4355 2208
rect 4419 2144 4435 2208
rect 4499 2144 4505 2208
rect 4189 2143 4505 2144
rect 11779 2208 12095 2209
rect 11779 2144 11785 2208
rect 11849 2144 11865 2208
rect 11929 2144 11945 2208
rect 12009 2144 12025 2208
rect 12089 2144 12095 2208
rect 11779 2143 12095 2144
rect 19369 2208 19685 2209
rect 19369 2144 19375 2208
rect 19439 2144 19455 2208
rect 19519 2144 19535 2208
rect 19599 2144 19615 2208
rect 19679 2144 19685 2208
rect 19369 2143 19685 2144
rect 26959 2208 27275 2209
rect 26959 2144 26965 2208
rect 27029 2144 27045 2208
rect 27109 2144 27125 2208
rect 27189 2144 27205 2208
rect 27269 2144 27275 2208
rect 26959 2143 27275 2144
rect 20529 2138 20595 2141
rect 24301 2138 24367 2141
rect 20529 2136 24367 2138
rect 20529 2080 20534 2136
rect 20590 2080 24306 2136
rect 24362 2080 24367 2136
rect 20529 2078 24367 2080
rect 20529 2075 20595 2078
rect 24301 2075 24367 2078
rect 1669 2002 1735 2005
rect 27429 2002 27495 2005
rect 1669 2000 27495 2002
rect 1669 1944 1674 2000
rect 1730 1944 27434 2000
rect 27490 1944 27495 2000
rect 1669 1942 27495 1944
rect 1669 1939 1735 1942
rect 27429 1939 27495 1942
rect 17861 1866 17927 1869
rect 29177 1866 29243 1869
rect 17861 1864 29243 1866
rect 17861 1808 17866 1864
rect 17922 1808 29182 1864
rect 29238 1808 29243 1864
rect 17861 1806 29243 1808
rect 17861 1803 17927 1806
rect 29177 1803 29243 1806
rect 8385 1730 8451 1733
rect 11421 1730 11487 1733
rect 8385 1728 11487 1730
rect 8385 1672 8390 1728
rect 8446 1672 11426 1728
rect 11482 1672 11487 1728
rect 8385 1670 11487 1672
rect 8385 1667 8451 1670
rect 11421 1667 11487 1670
rect 7984 1664 8300 1665
rect 7984 1600 7990 1664
rect 8054 1600 8070 1664
rect 8134 1600 8150 1664
rect 8214 1600 8230 1664
rect 8294 1600 8300 1664
rect 7984 1599 8300 1600
rect 15574 1664 15890 1665
rect 15574 1600 15580 1664
rect 15644 1600 15660 1664
rect 15724 1600 15740 1664
rect 15804 1600 15820 1664
rect 15884 1600 15890 1664
rect 15574 1599 15890 1600
rect 23164 1664 23480 1665
rect 23164 1600 23170 1664
rect 23234 1600 23250 1664
rect 23314 1600 23330 1664
rect 23394 1600 23410 1664
rect 23474 1600 23480 1664
rect 23164 1599 23480 1600
rect 30754 1664 31070 1665
rect 30754 1600 30760 1664
rect 30824 1600 30840 1664
rect 30904 1600 30920 1664
rect 30984 1600 31000 1664
rect 31064 1600 31070 1664
rect 30754 1599 31070 1600
rect 8661 1594 8727 1597
rect 14457 1594 14523 1597
rect 8661 1592 14523 1594
rect 8661 1536 8666 1592
rect 8722 1536 14462 1592
rect 14518 1536 14523 1592
rect 8661 1534 14523 1536
rect 8661 1531 8727 1534
rect 14457 1531 14523 1534
rect 2129 1458 2195 1461
rect 11053 1458 11119 1461
rect 2129 1456 11119 1458
rect 2129 1400 2134 1456
rect 2190 1400 11058 1456
rect 11114 1400 11119 1456
rect 2129 1398 11119 1400
rect 2129 1395 2195 1398
rect 11053 1395 11119 1398
rect 11421 1458 11487 1461
rect 13813 1458 13879 1461
rect 11421 1456 13879 1458
rect 11421 1400 11426 1456
rect 11482 1400 13818 1456
rect 13874 1400 13879 1456
rect 11421 1398 13879 1400
rect 11421 1395 11487 1398
rect 13813 1395 13879 1398
rect 22645 1458 22711 1461
rect 24301 1458 24367 1461
rect 22645 1456 24367 1458
rect 22645 1400 22650 1456
rect 22706 1400 24306 1456
rect 24362 1400 24367 1456
rect 22645 1398 24367 1400
rect 22645 1395 22711 1398
rect 24301 1395 24367 1398
rect 25957 1458 26023 1461
rect 26969 1458 27035 1461
rect 25957 1456 27035 1458
rect 25957 1400 25962 1456
rect 26018 1400 26974 1456
rect 27030 1400 27035 1456
rect 25957 1398 27035 1400
rect 25957 1395 26023 1398
rect 26969 1395 27035 1398
rect 2037 1322 2103 1325
rect 26877 1322 26943 1325
rect 2037 1320 26943 1322
rect 2037 1264 2042 1320
rect 2098 1264 26882 1320
rect 26938 1264 26943 1320
rect 2037 1262 26943 1264
rect 2037 1259 2103 1262
rect 26877 1259 26943 1262
rect 6085 1186 6151 1189
rect 9581 1186 9647 1189
rect 6085 1184 9647 1186
rect 6085 1128 6090 1184
rect 6146 1128 9586 1184
rect 9642 1128 9647 1184
rect 6085 1126 9647 1128
rect 6085 1123 6151 1126
rect 9581 1123 9647 1126
rect 20069 1186 20135 1189
rect 26325 1186 26391 1189
rect 20069 1184 26391 1186
rect 20069 1128 20074 1184
rect 20130 1128 26330 1184
rect 26386 1128 26391 1184
rect 20069 1126 26391 1128
rect 20069 1123 20135 1126
rect 26325 1123 26391 1126
rect 4189 1120 4505 1121
rect 4189 1056 4195 1120
rect 4259 1056 4275 1120
rect 4339 1056 4355 1120
rect 4419 1056 4435 1120
rect 4499 1056 4505 1120
rect 4189 1055 4505 1056
rect 11779 1120 12095 1121
rect 11779 1056 11785 1120
rect 11849 1056 11865 1120
rect 11929 1056 11945 1120
rect 12009 1056 12025 1120
rect 12089 1056 12095 1120
rect 11779 1055 12095 1056
rect 19369 1120 19685 1121
rect 19369 1056 19375 1120
rect 19439 1056 19455 1120
rect 19519 1056 19535 1120
rect 19599 1056 19615 1120
rect 19679 1056 19685 1120
rect 19369 1055 19685 1056
rect 26959 1120 27275 1121
rect 26959 1056 26965 1120
rect 27029 1056 27045 1120
rect 27109 1056 27125 1120
rect 27189 1056 27205 1120
rect 27269 1056 27275 1120
rect 26959 1055 27275 1056
rect 1669 914 1735 917
rect 26233 914 26299 917
rect 1669 912 26299 914
rect 1669 856 1674 912
rect 1730 856 26238 912
rect 26294 856 26299 912
rect 1669 854 26299 856
rect 1669 851 1735 854
rect 26233 851 26299 854
rect 1485 778 1551 781
rect 18229 778 18295 781
rect 1485 776 18295 778
rect 1485 720 1490 776
rect 1546 720 18234 776
rect 18290 720 18295 776
rect 1485 718 18295 720
rect 1485 715 1551 718
rect 18229 715 18295 718
rect 21449 778 21515 781
rect 23933 778 23999 781
rect 25773 778 25839 781
rect 21449 776 25839 778
rect 21449 720 21454 776
rect 21510 720 23938 776
rect 23994 720 25778 776
rect 25834 720 25839 776
rect 21449 718 25839 720
rect 21449 715 21515 718
rect 23933 715 23999 718
rect 25773 715 25839 718
rect 4889 642 4955 645
rect 6177 642 6243 645
rect 4889 640 6243 642
rect 4889 584 4894 640
rect 4950 584 6182 640
rect 6238 584 6243 640
rect 4889 582 6243 584
rect 4889 579 4955 582
rect 6177 579 6243 582
rect 11605 642 11671 645
rect 15377 642 15443 645
rect 11605 640 15443 642
rect 11605 584 11610 640
rect 11666 584 15382 640
rect 15438 584 15443 640
rect 11605 582 15443 584
rect 11605 579 11671 582
rect 15377 579 15443 582
rect 7984 576 8300 577
rect 7984 512 7990 576
rect 8054 512 8070 576
rect 8134 512 8150 576
rect 8214 512 8230 576
rect 8294 512 8300 576
rect 7984 511 8300 512
rect 15574 576 15890 577
rect 15574 512 15580 576
rect 15644 512 15660 576
rect 15724 512 15740 576
rect 15804 512 15820 576
rect 15884 512 15890 576
rect 15574 511 15890 512
rect 23164 576 23480 577
rect 23164 512 23170 576
rect 23234 512 23250 576
rect 23314 512 23330 576
rect 23394 512 23410 576
rect 23474 512 23480 576
rect 23164 511 23480 512
rect 30754 576 31070 577
rect 30754 512 30760 576
rect 30824 512 30840 576
rect 30904 512 30920 576
rect 30984 512 31000 576
rect 31064 512 31070 576
rect 30754 511 31070 512
rect 12157 370 12223 373
rect 25313 370 25379 373
rect 12157 368 25379 370
rect 12157 312 12162 368
rect 12218 312 25318 368
rect 25374 312 25379 368
rect 12157 310 25379 312
rect 12157 307 12223 310
rect 25313 307 25379 310
rect 4797 234 4863 237
rect 11973 234 12039 237
rect 4797 232 12039 234
rect 4797 176 4802 232
rect 4858 176 11978 232
rect 12034 176 12039 232
rect 4797 174 12039 176
rect 4797 171 4863 174
rect 11973 171 12039 174
<< via3 >>
rect 10732 22204 10796 22268
rect 12204 21796 12268 21860
rect 4195 21788 4259 21792
rect 4195 21732 4199 21788
rect 4199 21732 4255 21788
rect 4255 21732 4259 21788
rect 4195 21728 4259 21732
rect 4275 21788 4339 21792
rect 4275 21732 4279 21788
rect 4279 21732 4335 21788
rect 4335 21732 4339 21788
rect 4275 21728 4339 21732
rect 4355 21788 4419 21792
rect 4355 21732 4359 21788
rect 4359 21732 4415 21788
rect 4415 21732 4419 21788
rect 4355 21728 4419 21732
rect 4435 21788 4499 21792
rect 4435 21732 4439 21788
rect 4439 21732 4495 21788
rect 4495 21732 4499 21788
rect 4435 21728 4499 21732
rect 11785 21788 11849 21792
rect 11785 21732 11789 21788
rect 11789 21732 11845 21788
rect 11845 21732 11849 21788
rect 11785 21728 11849 21732
rect 11865 21788 11929 21792
rect 11865 21732 11869 21788
rect 11869 21732 11925 21788
rect 11925 21732 11929 21788
rect 11865 21728 11929 21732
rect 11945 21788 12009 21792
rect 11945 21732 11949 21788
rect 11949 21732 12005 21788
rect 12005 21732 12009 21788
rect 11945 21728 12009 21732
rect 12025 21788 12089 21792
rect 12025 21732 12029 21788
rect 12029 21732 12085 21788
rect 12085 21732 12089 21788
rect 12025 21728 12089 21732
rect 19375 21788 19439 21792
rect 19375 21732 19379 21788
rect 19379 21732 19435 21788
rect 19435 21732 19439 21788
rect 19375 21728 19439 21732
rect 19455 21788 19519 21792
rect 19455 21732 19459 21788
rect 19459 21732 19515 21788
rect 19515 21732 19519 21788
rect 19455 21728 19519 21732
rect 19535 21788 19599 21792
rect 19535 21732 19539 21788
rect 19539 21732 19595 21788
rect 19595 21732 19599 21788
rect 19535 21728 19599 21732
rect 19615 21788 19679 21792
rect 19615 21732 19619 21788
rect 19619 21732 19675 21788
rect 19675 21732 19679 21788
rect 19615 21728 19679 21732
rect 26965 21788 27029 21792
rect 26965 21732 26969 21788
rect 26969 21732 27025 21788
rect 27025 21732 27029 21788
rect 26965 21728 27029 21732
rect 27045 21788 27109 21792
rect 27045 21732 27049 21788
rect 27049 21732 27105 21788
rect 27105 21732 27109 21788
rect 27045 21728 27109 21732
rect 27125 21788 27189 21792
rect 27125 21732 27129 21788
rect 27129 21732 27185 21788
rect 27185 21732 27189 21788
rect 27125 21728 27189 21732
rect 27205 21788 27269 21792
rect 27205 21732 27209 21788
rect 27209 21732 27265 21788
rect 27265 21732 27269 21788
rect 27205 21728 27269 21732
rect 13676 21524 13740 21588
rect 16988 21524 17052 21588
rect 13676 21388 13740 21452
rect 25452 21524 25516 21588
rect 28764 21388 28828 21452
rect 7990 21244 8054 21248
rect 7990 21188 7994 21244
rect 7994 21188 8050 21244
rect 8050 21188 8054 21244
rect 7990 21184 8054 21188
rect 8070 21244 8134 21248
rect 8070 21188 8074 21244
rect 8074 21188 8130 21244
rect 8130 21188 8134 21244
rect 8070 21184 8134 21188
rect 8150 21244 8214 21248
rect 8150 21188 8154 21244
rect 8154 21188 8210 21244
rect 8210 21188 8214 21244
rect 8150 21184 8214 21188
rect 8230 21244 8294 21248
rect 8230 21188 8234 21244
rect 8234 21188 8290 21244
rect 8290 21188 8294 21244
rect 8230 21184 8294 21188
rect 15580 21244 15644 21248
rect 15580 21188 15584 21244
rect 15584 21188 15640 21244
rect 15640 21188 15644 21244
rect 15580 21184 15644 21188
rect 15660 21244 15724 21248
rect 15660 21188 15664 21244
rect 15664 21188 15720 21244
rect 15720 21188 15724 21244
rect 15660 21184 15724 21188
rect 15740 21244 15804 21248
rect 15740 21188 15744 21244
rect 15744 21188 15800 21244
rect 15800 21188 15804 21244
rect 15740 21184 15804 21188
rect 15820 21244 15884 21248
rect 15820 21188 15824 21244
rect 15824 21188 15880 21244
rect 15880 21188 15884 21244
rect 15820 21184 15884 21188
rect 23170 21244 23234 21248
rect 23170 21188 23174 21244
rect 23174 21188 23230 21244
rect 23230 21188 23234 21244
rect 23170 21184 23234 21188
rect 23250 21244 23314 21248
rect 23250 21188 23254 21244
rect 23254 21188 23310 21244
rect 23310 21188 23314 21244
rect 23250 21184 23314 21188
rect 23330 21244 23394 21248
rect 23330 21188 23334 21244
rect 23334 21188 23390 21244
rect 23390 21188 23394 21244
rect 23330 21184 23394 21188
rect 23410 21244 23474 21248
rect 23410 21188 23414 21244
rect 23414 21188 23470 21244
rect 23470 21188 23474 21244
rect 23410 21184 23474 21188
rect 30760 21244 30824 21248
rect 30760 21188 30764 21244
rect 30764 21188 30820 21244
rect 30820 21188 30824 21244
rect 30760 21184 30824 21188
rect 30840 21244 30904 21248
rect 30840 21188 30844 21244
rect 30844 21188 30900 21244
rect 30900 21188 30904 21244
rect 30840 21184 30904 21188
rect 30920 21244 30984 21248
rect 30920 21188 30924 21244
rect 30924 21188 30980 21244
rect 30980 21188 30984 21244
rect 30920 21184 30984 21188
rect 31000 21244 31064 21248
rect 31000 21188 31004 21244
rect 31004 21188 31060 21244
rect 31060 21188 31064 21244
rect 31000 21184 31064 21188
rect 26372 21116 26436 21180
rect 11284 20980 11348 21044
rect 24900 20980 24964 21044
rect 3924 20708 3988 20772
rect 11468 20844 11532 20908
rect 8892 20708 8956 20772
rect 10180 20708 10244 20772
rect 4195 20700 4259 20704
rect 4195 20644 4199 20700
rect 4199 20644 4255 20700
rect 4255 20644 4259 20700
rect 4195 20640 4259 20644
rect 4275 20700 4339 20704
rect 4275 20644 4279 20700
rect 4279 20644 4335 20700
rect 4335 20644 4339 20700
rect 4275 20640 4339 20644
rect 4355 20700 4419 20704
rect 4355 20644 4359 20700
rect 4359 20644 4415 20700
rect 4415 20644 4419 20700
rect 4355 20640 4419 20644
rect 4435 20700 4499 20704
rect 4435 20644 4439 20700
rect 4439 20644 4495 20700
rect 4495 20644 4499 20700
rect 4435 20640 4499 20644
rect 11785 20700 11849 20704
rect 11785 20644 11789 20700
rect 11789 20644 11845 20700
rect 11845 20644 11849 20700
rect 11785 20640 11849 20644
rect 11865 20700 11929 20704
rect 11865 20644 11869 20700
rect 11869 20644 11925 20700
rect 11925 20644 11929 20700
rect 11865 20640 11929 20644
rect 11945 20700 12009 20704
rect 11945 20644 11949 20700
rect 11949 20644 12005 20700
rect 12005 20644 12009 20700
rect 11945 20640 12009 20644
rect 12025 20700 12089 20704
rect 12025 20644 12029 20700
rect 12029 20644 12085 20700
rect 12085 20644 12089 20700
rect 12025 20640 12089 20644
rect 19375 20700 19439 20704
rect 19375 20644 19379 20700
rect 19379 20644 19435 20700
rect 19435 20644 19439 20700
rect 19375 20640 19439 20644
rect 19455 20700 19519 20704
rect 19455 20644 19459 20700
rect 19459 20644 19515 20700
rect 19515 20644 19519 20700
rect 19455 20640 19519 20644
rect 19535 20700 19599 20704
rect 19535 20644 19539 20700
rect 19539 20644 19595 20700
rect 19595 20644 19599 20700
rect 19535 20640 19599 20644
rect 19615 20700 19679 20704
rect 19615 20644 19619 20700
rect 19619 20644 19675 20700
rect 19675 20644 19679 20700
rect 19615 20640 19679 20644
rect 26965 20700 27029 20704
rect 26965 20644 26969 20700
rect 26969 20644 27025 20700
rect 27025 20644 27029 20700
rect 26965 20640 27029 20644
rect 27045 20700 27109 20704
rect 27045 20644 27049 20700
rect 27049 20644 27105 20700
rect 27105 20644 27109 20700
rect 27045 20640 27109 20644
rect 27125 20700 27189 20704
rect 27125 20644 27129 20700
rect 27129 20644 27185 20700
rect 27185 20644 27189 20700
rect 27125 20640 27189 20644
rect 27205 20700 27269 20704
rect 27205 20644 27209 20700
rect 27209 20644 27265 20700
rect 27265 20644 27269 20700
rect 27205 20640 27269 20644
rect 7604 20572 7668 20636
rect 15148 20572 15212 20636
rect 23612 20572 23676 20636
rect 27660 20436 27724 20500
rect 7990 20156 8054 20160
rect 7990 20100 7994 20156
rect 7994 20100 8050 20156
rect 8050 20100 8054 20156
rect 7990 20096 8054 20100
rect 8070 20156 8134 20160
rect 8070 20100 8074 20156
rect 8074 20100 8130 20156
rect 8130 20100 8134 20156
rect 8070 20096 8134 20100
rect 8150 20156 8214 20160
rect 8150 20100 8154 20156
rect 8154 20100 8210 20156
rect 8210 20100 8214 20156
rect 8150 20096 8214 20100
rect 8230 20156 8294 20160
rect 8230 20100 8234 20156
rect 8234 20100 8290 20156
rect 8290 20100 8294 20156
rect 8230 20096 8294 20100
rect 15580 20156 15644 20160
rect 15580 20100 15584 20156
rect 15584 20100 15640 20156
rect 15640 20100 15644 20156
rect 15580 20096 15644 20100
rect 15660 20156 15724 20160
rect 15660 20100 15664 20156
rect 15664 20100 15720 20156
rect 15720 20100 15724 20156
rect 15660 20096 15724 20100
rect 15740 20156 15804 20160
rect 15740 20100 15744 20156
rect 15744 20100 15800 20156
rect 15800 20100 15804 20156
rect 15740 20096 15804 20100
rect 15820 20156 15884 20160
rect 15820 20100 15824 20156
rect 15824 20100 15880 20156
rect 15880 20100 15884 20156
rect 15820 20096 15884 20100
rect 23170 20156 23234 20160
rect 23170 20100 23174 20156
rect 23174 20100 23230 20156
rect 23230 20100 23234 20156
rect 23170 20096 23234 20100
rect 23250 20156 23314 20160
rect 23250 20100 23254 20156
rect 23254 20100 23310 20156
rect 23310 20100 23314 20156
rect 23250 20096 23314 20100
rect 23330 20156 23394 20160
rect 23330 20100 23334 20156
rect 23334 20100 23390 20156
rect 23390 20100 23394 20156
rect 23330 20096 23394 20100
rect 23410 20156 23474 20160
rect 23410 20100 23414 20156
rect 23414 20100 23470 20156
rect 23470 20100 23474 20156
rect 23410 20096 23474 20100
rect 30760 20156 30824 20160
rect 30760 20100 30764 20156
rect 30764 20100 30820 20156
rect 30820 20100 30824 20156
rect 30760 20096 30824 20100
rect 30840 20156 30904 20160
rect 30840 20100 30844 20156
rect 30844 20100 30900 20156
rect 30900 20100 30904 20156
rect 30840 20096 30904 20100
rect 30920 20156 30984 20160
rect 30920 20100 30924 20156
rect 30924 20100 30980 20156
rect 30980 20100 30984 20156
rect 30920 20096 30984 20100
rect 31000 20156 31064 20160
rect 31000 20100 31004 20156
rect 31004 20100 31060 20156
rect 31060 20100 31064 20156
rect 31000 20096 31064 20100
rect 21956 19892 22020 19956
rect 4195 19612 4259 19616
rect 4195 19556 4199 19612
rect 4199 19556 4255 19612
rect 4255 19556 4259 19612
rect 4195 19552 4259 19556
rect 4275 19612 4339 19616
rect 4275 19556 4279 19612
rect 4279 19556 4335 19612
rect 4335 19556 4339 19612
rect 4275 19552 4339 19556
rect 4355 19612 4419 19616
rect 4355 19556 4359 19612
rect 4359 19556 4415 19612
rect 4415 19556 4419 19612
rect 4355 19552 4419 19556
rect 4435 19612 4499 19616
rect 4435 19556 4439 19612
rect 4439 19556 4495 19612
rect 4495 19556 4499 19612
rect 4435 19552 4499 19556
rect 11785 19612 11849 19616
rect 11785 19556 11789 19612
rect 11789 19556 11845 19612
rect 11845 19556 11849 19612
rect 11785 19552 11849 19556
rect 11865 19612 11929 19616
rect 11865 19556 11869 19612
rect 11869 19556 11925 19612
rect 11925 19556 11929 19612
rect 11865 19552 11929 19556
rect 11945 19612 12009 19616
rect 11945 19556 11949 19612
rect 11949 19556 12005 19612
rect 12005 19556 12009 19612
rect 11945 19552 12009 19556
rect 12025 19612 12089 19616
rect 12025 19556 12029 19612
rect 12029 19556 12085 19612
rect 12085 19556 12089 19612
rect 12025 19552 12089 19556
rect 19375 19612 19439 19616
rect 19375 19556 19379 19612
rect 19379 19556 19435 19612
rect 19435 19556 19439 19612
rect 19375 19552 19439 19556
rect 19455 19612 19519 19616
rect 19455 19556 19459 19612
rect 19459 19556 19515 19612
rect 19515 19556 19519 19612
rect 19455 19552 19519 19556
rect 19535 19612 19599 19616
rect 19535 19556 19539 19612
rect 19539 19556 19595 19612
rect 19595 19556 19599 19612
rect 19535 19552 19599 19556
rect 19615 19612 19679 19616
rect 19615 19556 19619 19612
rect 19619 19556 19675 19612
rect 19675 19556 19679 19612
rect 19615 19552 19679 19556
rect 26965 19612 27029 19616
rect 26965 19556 26969 19612
rect 26969 19556 27025 19612
rect 27025 19556 27029 19612
rect 26965 19552 27029 19556
rect 27045 19612 27109 19616
rect 27045 19556 27049 19612
rect 27049 19556 27105 19612
rect 27105 19556 27109 19612
rect 27045 19552 27109 19556
rect 27125 19612 27189 19616
rect 27125 19556 27129 19612
rect 27129 19556 27185 19612
rect 27185 19556 27189 19612
rect 27125 19552 27189 19556
rect 27205 19612 27269 19616
rect 27205 19556 27209 19612
rect 27209 19556 27265 19612
rect 27265 19556 27269 19612
rect 27205 19552 27269 19556
rect 11468 19348 11532 19412
rect 26556 19348 26620 19412
rect 8708 19076 8772 19140
rect 10916 19212 10980 19276
rect 12572 19212 12636 19276
rect 14780 19212 14844 19276
rect 16068 19212 16132 19276
rect 16436 19272 16500 19276
rect 16436 19216 16486 19272
rect 16486 19216 16500 19272
rect 16436 19212 16500 19216
rect 24716 19212 24780 19276
rect 9812 19136 9876 19140
rect 9812 19080 9862 19136
rect 9862 19080 9876 19136
rect 9812 19076 9876 19080
rect 7990 19068 8054 19072
rect 7990 19012 7994 19068
rect 7994 19012 8050 19068
rect 8050 19012 8054 19068
rect 7990 19008 8054 19012
rect 8070 19068 8134 19072
rect 8070 19012 8074 19068
rect 8074 19012 8130 19068
rect 8130 19012 8134 19068
rect 8070 19008 8134 19012
rect 8150 19068 8214 19072
rect 8150 19012 8154 19068
rect 8154 19012 8210 19068
rect 8210 19012 8214 19068
rect 8150 19008 8214 19012
rect 8230 19068 8294 19072
rect 8230 19012 8234 19068
rect 8234 19012 8290 19068
rect 8290 19012 8294 19068
rect 8230 19008 8294 19012
rect 15580 19068 15644 19072
rect 15580 19012 15584 19068
rect 15584 19012 15640 19068
rect 15640 19012 15644 19068
rect 15580 19008 15644 19012
rect 15660 19068 15724 19072
rect 15660 19012 15664 19068
rect 15664 19012 15720 19068
rect 15720 19012 15724 19068
rect 15660 19008 15724 19012
rect 15740 19068 15804 19072
rect 15740 19012 15744 19068
rect 15744 19012 15800 19068
rect 15800 19012 15804 19068
rect 15740 19008 15804 19012
rect 15820 19068 15884 19072
rect 15820 19012 15824 19068
rect 15824 19012 15880 19068
rect 15880 19012 15884 19068
rect 15820 19008 15884 19012
rect 23170 19068 23234 19072
rect 23170 19012 23174 19068
rect 23174 19012 23230 19068
rect 23230 19012 23234 19068
rect 23170 19008 23234 19012
rect 23250 19068 23314 19072
rect 23250 19012 23254 19068
rect 23254 19012 23310 19068
rect 23310 19012 23314 19068
rect 23250 19008 23314 19012
rect 23330 19068 23394 19072
rect 23330 19012 23334 19068
rect 23334 19012 23390 19068
rect 23390 19012 23394 19068
rect 23330 19008 23394 19012
rect 23410 19068 23474 19072
rect 23410 19012 23414 19068
rect 23414 19012 23470 19068
rect 23470 19012 23474 19068
rect 23410 19008 23474 19012
rect 30760 19068 30824 19072
rect 30760 19012 30764 19068
rect 30764 19012 30820 19068
rect 30820 19012 30824 19068
rect 30760 19008 30824 19012
rect 30840 19068 30904 19072
rect 30840 19012 30844 19068
rect 30844 19012 30900 19068
rect 30900 19012 30904 19068
rect 30840 19008 30904 19012
rect 30920 19068 30984 19072
rect 30920 19012 30924 19068
rect 30924 19012 30980 19068
rect 30980 19012 30984 19068
rect 30920 19008 30984 19012
rect 31000 19068 31064 19072
rect 31000 19012 31004 19068
rect 31004 19012 31060 19068
rect 31060 19012 31064 19068
rect 31000 19008 31064 19012
rect 9260 18804 9324 18868
rect 23980 18804 24044 18868
rect 5396 18728 5460 18732
rect 5396 18672 5446 18728
rect 5446 18672 5460 18728
rect 5396 18668 5460 18672
rect 8708 18668 8772 18732
rect 4195 18524 4259 18528
rect 4195 18468 4199 18524
rect 4199 18468 4255 18524
rect 4255 18468 4259 18524
rect 4195 18464 4259 18468
rect 4275 18524 4339 18528
rect 4275 18468 4279 18524
rect 4279 18468 4335 18524
rect 4335 18468 4339 18524
rect 4275 18464 4339 18468
rect 4355 18524 4419 18528
rect 4355 18468 4359 18524
rect 4359 18468 4415 18524
rect 4415 18468 4419 18524
rect 4355 18464 4419 18468
rect 4435 18524 4499 18528
rect 4435 18468 4439 18524
rect 4439 18468 4495 18524
rect 4495 18468 4499 18524
rect 4435 18464 4499 18468
rect 11785 18524 11849 18528
rect 11785 18468 11789 18524
rect 11789 18468 11845 18524
rect 11845 18468 11849 18524
rect 11785 18464 11849 18468
rect 11865 18524 11929 18528
rect 11865 18468 11869 18524
rect 11869 18468 11925 18524
rect 11925 18468 11929 18524
rect 11865 18464 11929 18468
rect 11945 18524 12009 18528
rect 11945 18468 11949 18524
rect 11949 18468 12005 18524
rect 12005 18468 12009 18524
rect 11945 18464 12009 18468
rect 12025 18524 12089 18528
rect 12025 18468 12029 18524
rect 12029 18468 12085 18524
rect 12085 18468 12089 18524
rect 12025 18464 12089 18468
rect 19375 18524 19439 18528
rect 19375 18468 19379 18524
rect 19379 18468 19435 18524
rect 19435 18468 19439 18524
rect 19375 18464 19439 18468
rect 19455 18524 19519 18528
rect 19455 18468 19459 18524
rect 19459 18468 19515 18524
rect 19515 18468 19519 18524
rect 19455 18464 19519 18468
rect 19535 18524 19599 18528
rect 19535 18468 19539 18524
rect 19539 18468 19595 18524
rect 19595 18468 19599 18524
rect 19535 18464 19599 18468
rect 19615 18524 19679 18528
rect 19615 18468 19619 18524
rect 19619 18468 19675 18524
rect 19675 18468 19679 18524
rect 19615 18464 19679 18468
rect 26965 18524 27029 18528
rect 26965 18468 26969 18524
rect 26969 18468 27025 18524
rect 27025 18468 27029 18524
rect 26965 18464 27029 18468
rect 27045 18524 27109 18528
rect 27045 18468 27049 18524
rect 27049 18468 27105 18524
rect 27105 18468 27109 18524
rect 27045 18464 27109 18468
rect 27125 18524 27189 18528
rect 27125 18468 27129 18524
rect 27129 18468 27185 18524
rect 27185 18468 27189 18524
rect 27125 18464 27189 18468
rect 27205 18524 27269 18528
rect 27205 18468 27209 18524
rect 27209 18468 27265 18524
rect 27265 18468 27269 18524
rect 27205 18464 27269 18468
rect 4660 18456 4724 18460
rect 4660 18400 4674 18456
rect 4674 18400 4724 18456
rect 4660 18396 4724 18400
rect 5212 18396 5276 18460
rect 10548 18396 10612 18460
rect 7052 18260 7116 18324
rect 6500 18124 6564 18188
rect 5396 17988 5460 18052
rect 6684 18048 6748 18052
rect 6684 17992 6734 18048
rect 6734 17992 6748 18048
rect 6684 17988 6748 17992
rect 7990 17980 8054 17984
rect 7990 17924 7994 17980
rect 7994 17924 8050 17980
rect 8050 17924 8054 17980
rect 7990 17920 8054 17924
rect 8070 17980 8134 17984
rect 8070 17924 8074 17980
rect 8074 17924 8130 17980
rect 8130 17924 8134 17980
rect 8070 17920 8134 17924
rect 8150 17980 8214 17984
rect 8150 17924 8154 17980
rect 8154 17924 8210 17980
rect 8210 17924 8214 17980
rect 8150 17920 8214 17924
rect 8230 17980 8294 17984
rect 8230 17924 8234 17980
rect 8234 17924 8290 17980
rect 8290 17924 8294 17980
rect 8230 17920 8294 17924
rect 22508 18048 22572 18052
rect 22508 17992 22558 18048
rect 22558 17992 22572 18048
rect 22508 17988 22572 17992
rect 22876 17988 22940 18052
rect 24164 18124 24228 18188
rect 15580 17980 15644 17984
rect 15580 17924 15584 17980
rect 15584 17924 15640 17980
rect 15640 17924 15644 17980
rect 15580 17920 15644 17924
rect 15660 17980 15724 17984
rect 15660 17924 15664 17980
rect 15664 17924 15720 17980
rect 15720 17924 15724 17980
rect 15660 17920 15724 17924
rect 15740 17980 15804 17984
rect 15740 17924 15744 17980
rect 15744 17924 15800 17980
rect 15800 17924 15804 17980
rect 15740 17920 15804 17924
rect 15820 17980 15884 17984
rect 15820 17924 15824 17980
rect 15824 17924 15880 17980
rect 15880 17924 15884 17980
rect 15820 17920 15884 17924
rect 23170 17980 23234 17984
rect 23170 17924 23174 17980
rect 23174 17924 23230 17980
rect 23230 17924 23234 17980
rect 23170 17920 23234 17924
rect 23250 17980 23314 17984
rect 23250 17924 23254 17980
rect 23254 17924 23310 17980
rect 23310 17924 23314 17980
rect 23250 17920 23314 17924
rect 23330 17980 23394 17984
rect 23330 17924 23334 17980
rect 23334 17924 23390 17980
rect 23390 17924 23394 17980
rect 23330 17920 23394 17924
rect 23410 17980 23474 17984
rect 23410 17924 23414 17980
rect 23414 17924 23470 17980
rect 23470 17924 23474 17980
rect 23410 17920 23474 17924
rect 30760 17980 30824 17984
rect 30760 17924 30764 17980
rect 30764 17924 30820 17980
rect 30820 17924 30824 17980
rect 30760 17920 30824 17924
rect 30840 17980 30904 17984
rect 30840 17924 30844 17980
rect 30844 17924 30900 17980
rect 30900 17924 30904 17980
rect 30840 17920 30904 17924
rect 30920 17980 30984 17984
rect 30920 17924 30924 17980
rect 30924 17924 30980 17980
rect 30980 17924 30984 17980
rect 30920 17920 30984 17924
rect 31000 17980 31064 17984
rect 31000 17924 31004 17980
rect 31004 17924 31060 17980
rect 31060 17924 31064 17980
rect 31000 17920 31064 17924
rect 4195 17436 4259 17440
rect 4195 17380 4199 17436
rect 4199 17380 4255 17436
rect 4255 17380 4259 17436
rect 4195 17376 4259 17380
rect 4275 17436 4339 17440
rect 4275 17380 4279 17436
rect 4279 17380 4335 17436
rect 4335 17380 4339 17436
rect 4275 17376 4339 17380
rect 4355 17436 4419 17440
rect 4355 17380 4359 17436
rect 4359 17380 4415 17436
rect 4415 17380 4419 17436
rect 4355 17376 4419 17380
rect 4435 17436 4499 17440
rect 4435 17380 4439 17436
rect 4439 17380 4495 17436
rect 4495 17380 4499 17436
rect 4435 17376 4499 17380
rect 5948 17308 6012 17372
rect 11785 17436 11849 17440
rect 11785 17380 11789 17436
rect 11789 17380 11845 17436
rect 11845 17380 11849 17436
rect 11785 17376 11849 17380
rect 11865 17436 11929 17440
rect 11865 17380 11869 17436
rect 11869 17380 11925 17436
rect 11925 17380 11929 17436
rect 11865 17376 11929 17380
rect 11945 17436 12009 17440
rect 11945 17380 11949 17436
rect 11949 17380 12005 17436
rect 12005 17380 12009 17436
rect 11945 17376 12009 17380
rect 12025 17436 12089 17440
rect 12025 17380 12029 17436
rect 12029 17380 12085 17436
rect 12085 17380 12089 17436
rect 12025 17376 12089 17380
rect 19375 17436 19439 17440
rect 19375 17380 19379 17436
rect 19379 17380 19435 17436
rect 19435 17380 19439 17436
rect 19375 17376 19439 17380
rect 19455 17436 19519 17440
rect 19455 17380 19459 17436
rect 19459 17380 19515 17436
rect 19515 17380 19519 17436
rect 19455 17376 19519 17380
rect 19535 17436 19599 17440
rect 19535 17380 19539 17436
rect 19539 17380 19595 17436
rect 19595 17380 19599 17436
rect 19535 17376 19599 17380
rect 19615 17436 19679 17440
rect 19615 17380 19619 17436
rect 19619 17380 19675 17436
rect 19675 17380 19679 17436
rect 19615 17376 19679 17380
rect 26965 17436 27029 17440
rect 26965 17380 26969 17436
rect 26969 17380 27025 17436
rect 27025 17380 27029 17436
rect 26965 17376 27029 17380
rect 27045 17436 27109 17440
rect 27045 17380 27049 17436
rect 27049 17380 27105 17436
rect 27105 17380 27109 17436
rect 27045 17376 27109 17380
rect 27125 17436 27189 17440
rect 27125 17380 27129 17436
rect 27129 17380 27185 17436
rect 27185 17380 27189 17436
rect 27125 17376 27189 17380
rect 27205 17436 27269 17440
rect 27205 17380 27209 17436
rect 27209 17380 27265 17436
rect 27265 17380 27269 17436
rect 27205 17376 27269 17380
rect 7990 16892 8054 16896
rect 7990 16836 7994 16892
rect 7994 16836 8050 16892
rect 8050 16836 8054 16892
rect 7990 16832 8054 16836
rect 8070 16892 8134 16896
rect 8070 16836 8074 16892
rect 8074 16836 8130 16892
rect 8130 16836 8134 16892
rect 8070 16832 8134 16836
rect 8150 16892 8214 16896
rect 8150 16836 8154 16892
rect 8154 16836 8210 16892
rect 8210 16836 8214 16892
rect 8150 16832 8214 16836
rect 8230 16892 8294 16896
rect 8230 16836 8234 16892
rect 8234 16836 8290 16892
rect 8290 16836 8294 16892
rect 8230 16832 8294 16836
rect 5948 16628 6012 16692
rect 8524 16764 8588 16828
rect 29500 17096 29564 17100
rect 29500 17040 29550 17096
rect 29550 17040 29564 17096
rect 29500 17036 29564 17040
rect 15580 16892 15644 16896
rect 15580 16836 15584 16892
rect 15584 16836 15640 16892
rect 15640 16836 15644 16892
rect 15580 16832 15644 16836
rect 15660 16892 15724 16896
rect 15660 16836 15664 16892
rect 15664 16836 15720 16892
rect 15720 16836 15724 16892
rect 15660 16832 15724 16836
rect 15740 16892 15804 16896
rect 15740 16836 15744 16892
rect 15744 16836 15800 16892
rect 15800 16836 15804 16892
rect 15740 16832 15804 16836
rect 15820 16892 15884 16896
rect 15820 16836 15824 16892
rect 15824 16836 15880 16892
rect 15880 16836 15884 16892
rect 15820 16832 15884 16836
rect 23170 16892 23234 16896
rect 23170 16836 23174 16892
rect 23174 16836 23230 16892
rect 23230 16836 23234 16892
rect 23170 16832 23234 16836
rect 23250 16892 23314 16896
rect 23250 16836 23254 16892
rect 23254 16836 23310 16892
rect 23310 16836 23314 16892
rect 23250 16832 23314 16836
rect 23330 16892 23394 16896
rect 23330 16836 23334 16892
rect 23334 16836 23390 16892
rect 23390 16836 23394 16892
rect 23330 16832 23394 16836
rect 23410 16892 23474 16896
rect 23410 16836 23414 16892
rect 23414 16836 23470 16892
rect 23470 16836 23474 16892
rect 23410 16832 23474 16836
rect 30760 16892 30824 16896
rect 30760 16836 30764 16892
rect 30764 16836 30820 16892
rect 30820 16836 30824 16892
rect 30760 16832 30824 16836
rect 30840 16892 30904 16896
rect 30840 16836 30844 16892
rect 30844 16836 30900 16892
rect 30900 16836 30904 16892
rect 30840 16832 30904 16836
rect 30920 16892 30984 16896
rect 30920 16836 30924 16892
rect 30924 16836 30980 16892
rect 30980 16836 30984 16892
rect 30920 16832 30984 16836
rect 31000 16892 31064 16896
rect 31000 16836 31004 16892
rect 31004 16836 31060 16892
rect 31060 16836 31064 16892
rect 31000 16832 31064 16836
rect 29316 16824 29380 16828
rect 29316 16768 29330 16824
rect 29330 16768 29380 16824
rect 29316 16764 29380 16768
rect 29132 16552 29196 16556
rect 29132 16496 29182 16552
rect 29182 16496 29196 16552
rect 29132 16492 29196 16496
rect 14228 16356 14292 16420
rect 29684 16356 29748 16420
rect 4195 16348 4259 16352
rect 4195 16292 4199 16348
rect 4199 16292 4255 16348
rect 4255 16292 4259 16348
rect 4195 16288 4259 16292
rect 4275 16348 4339 16352
rect 4275 16292 4279 16348
rect 4279 16292 4335 16348
rect 4335 16292 4339 16348
rect 4275 16288 4339 16292
rect 4355 16348 4419 16352
rect 4355 16292 4359 16348
rect 4359 16292 4415 16348
rect 4415 16292 4419 16348
rect 4355 16288 4419 16292
rect 4435 16348 4499 16352
rect 4435 16292 4439 16348
rect 4439 16292 4495 16348
rect 4495 16292 4499 16348
rect 4435 16288 4499 16292
rect 11785 16348 11849 16352
rect 11785 16292 11789 16348
rect 11789 16292 11845 16348
rect 11845 16292 11849 16348
rect 11785 16288 11849 16292
rect 11865 16348 11929 16352
rect 11865 16292 11869 16348
rect 11869 16292 11925 16348
rect 11925 16292 11929 16348
rect 11865 16288 11929 16292
rect 11945 16348 12009 16352
rect 11945 16292 11949 16348
rect 11949 16292 12005 16348
rect 12005 16292 12009 16348
rect 11945 16288 12009 16292
rect 12025 16348 12089 16352
rect 12025 16292 12029 16348
rect 12029 16292 12085 16348
rect 12085 16292 12089 16348
rect 12025 16288 12089 16292
rect 19375 16348 19439 16352
rect 19375 16292 19379 16348
rect 19379 16292 19435 16348
rect 19435 16292 19439 16348
rect 19375 16288 19439 16292
rect 19455 16348 19519 16352
rect 19455 16292 19459 16348
rect 19459 16292 19515 16348
rect 19515 16292 19519 16348
rect 19455 16288 19519 16292
rect 19535 16348 19599 16352
rect 19535 16292 19539 16348
rect 19539 16292 19595 16348
rect 19595 16292 19599 16348
rect 19535 16288 19599 16292
rect 19615 16348 19679 16352
rect 19615 16292 19619 16348
rect 19619 16292 19675 16348
rect 19675 16292 19679 16348
rect 19615 16288 19679 16292
rect 26965 16348 27029 16352
rect 26965 16292 26969 16348
rect 26969 16292 27025 16348
rect 27025 16292 27029 16348
rect 26965 16288 27029 16292
rect 27045 16348 27109 16352
rect 27045 16292 27049 16348
rect 27049 16292 27105 16348
rect 27105 16292 27109 16348
rect 27045 16288 27109 16292
rect 27125 16348 27189 16352
rect 27125 16292 27129 16348
rect 27129 16292 27185 16348
rect 27185 16292 27189 16348
rect 27125 16288 27189 16292
rect 27205 16348 27269 16352
rect 27205 16292 27209 16348
rect 27209 16292 27265 16348
rect 27265 16292 27269 16348
rect 27205 16288 27269 16292
rect 29500 16084 29564 16148
rect 7990 15804 8054 15808
rect 7990 15748 7994 15804
rect 7994 15748 8050 15804
rect 8050 15748 8054 15804
rect 7990 15744 8054 15748
rect 8070 15804 8134 15808
rect 8070 15748 8074 15804
rect 8074 15748 8130 15804
rect 8130 15748 8134 15804
rect 8070 15744 8134 15748
rect 8150 15804 8214 15808
rect 8150 15748 8154 15804
rect 8154 15748 8210 15804
rect 8210 15748 8214 15804
rect 8150 15744 8214 15748
rect 8230 15804 8294 15808
rect 8230 15748 8234 15804
rect 8234 15748 8290 15804
rect 8290 15748 8294 15804
rect 8230 15744 8294 15748
rect 15580 15804 15644 15808
rect 15580 15748 15584 15804
rect 15584 15748 15640 15804
rect 15640 15748 15644 15804
rect 15580 15744 15644 15748
rect 15660 15804 15724 15808
rect 15660 15748 15664 15804
rect 15664 15748 15720 15804
rect 15720 15748 15724 15804
rect 15660 15744 15724 15748
rect 15740 15804 15804 15808
rect 15740 15748 15744 15804
rect 15744 15748 15800 15804
rect 15800 15748 15804 15804
rect 15740 15744 15804 15748
rect 15820 15804 15884 15808
rect 15820 15748 15824 15804
rect 15824 15748 15880 15804
rect 15880 15748 15884 15804
rect 15820 15744 15884 15748
rect 23170 15804 23234 15808
rect 23170 15748 23174 15804
rect 23174 15748 23230 15804
rect 23230 15748 23234 15804
rect 23170 15744 23234 15748
rect 23250 15804 23314 15808
rect 23250 15748 23254 15804
rect 23254 15748 23310 15804
rect 23310 15748 23314 15804
rect 23250 15744 23314 15748
rect 23330 15804 23394 15808
rect 23330 15748 23334 15804
rect 23334 15748 23390 15804
rect 23390 15748 23394 15804
rect 23330 15744 23394 15748
rect 23410 15804 23474 15808
rect 23410 15748 23414 15804
rect 23414 15748 23470 15804
rect 23470 15748 23474 15804
rect 23410 15744 23474 15748
rect 30760 15804 30824 15808
rect 30760 15748 30764 15804
rect 30764 15748 30820 15804
rect 30820 15748 30824 15804
rect 30760 15744 30824 15748
rect 30840 15804 30904 15808
rect 30840 15748 30844 15804
rect 30844 15748 30900 15804
rect 30900 15748 30904 15804
rect 30840 15744 30904 15748
rect 30920 15804 30984 15808
rect 30920 15748 30924 15804
rect 30924 15748 30980 15804
rect 30980 15748 30984 15804
rect 30920 15744 30984 15748
rect 31000 15804 31064 15808
rect 31000 15748 31004 15804
rect 31004 15748 31060 15804
rect 31060 15748 31064 15804
rect 31000 15744 31064 15748
rect 12572 15676 12636 15740
rect 29316 15676 29380 15740
rect 4195 15260 4259 15264
rect 4195 15204 4199 15260
rect 4199 15204 4255 15260
rect 4255 15204 4259 15260
rect 4195 15200 4259 15204
rect 4275 15260 4339 15264
rect 4275 15204 4279 15260
rect 4279 15204 4335 15260
rect 4335 15204 4339 15260
rect 4275 15200 4339 15204
rect 4355 15260 4419 15264
rect 4355 15204 4359 15260
rect 4359 15204 4415 15260
rect 4415 15204 4419 15260
rect 4355 15200 4419 15204
rect 4435 15260 4499 15264
rect 4435 15204 4439 15260
rect 4439 15204 4495 15260
rect 4495 15204 4499 15260
rect 4435 15200 4499 15204
rect 11785 15260 11849 15264
rect 11785 15204 11789 15260
rect 11789 15204 11845 15260
rect 11845 15204 11849 15260
rect 11785 15200 11849 15204
rect 11865 15260 11929 15264
rect 11865 15204 11869 15260
rect 11869 15204 11925 15260
rect 11925 15204 11929 15260
rect 11865 15200 11929 15204
rect 11945 15260 12009 15264
rect 11945 15204 11949 15260
rect 11949 15204 12005 15260
rect 12005 15204 12009 15260
rect 11945 15200 12009 15204
rect 12025 15260 12089 15264
rect 12025 15204 12029 15260
rect 12029 15204 12085 15260
rect 12085 15204 12089 15260
rect 12025 15200 12089 15204
rect 19375 15260 19439 15264
rect 19375 15204 19379 15260
rect 19379 15204 19435 15260
rect 19435 15204 19439 15260
rect 19375 15200 19439 15204
rect 19455 15260 19519 15264
rect 19455 15204 19459 15260
rect 19459 15204 19515 15260
rect 19515 15204 19519 15260
rect 19455 15200 19519 15204
rect 19535 15260 19599 15264
rect 19535 15204 19539 15260
rect 19539 15204 19595 15260
rect 19595 15204 19599 15260
rect 19535 15200 19599 15204
rect 19615 15260 19679 15264
rect 19615 15204 19619 15260
rect 19619 15204 19675 15260
rect 19675 15204 19679 15260
rect 19615 15200 19679 15204
rect 26965 15260 27029 15264
rect 26965 15204 26969 15260
rect 26969 15204 27025 15260
rect 27025 15204 27029 15260
rect 26965 15200 27029 15204
rect 27045 15260 27109 15264
rect 27045 15204 27049 15260
rect 27049 15204 27105 15260
rect 27105 15204 27109 15260
rect 27045 15200 27109 15204
rect 27125 15260 27189 15264
rect 27125 15204 27129 15260
rect 27129 15204 27185 15260
rect 27185 15204 27189 15260
rect 27125 15200 27189 15204
rect 27205 15260 27269 15264
rect 27205 15204 27209 15260
rect 27209 15204 27265 15260
rect 27265 15204 27269 15260
rect 27205 15200 27269 15204
rect 8524 15132 8588 15196
rect 26556 15192 26620 15196
rect 26556 15136 26570 15192
rect 26570 15136 26620 15192
rect 26556 15132 26620 15136
rect 7990 14716 8054 14720
rect 7990 14660 7994 14716
rect 7994 14660 8050 14716
rect 8050 14660 8054 14716
rect 7990 14656 8054 14660
rect 8070 14716 8134 14720
rect 8070 14660 8074 14716
rect 8074 14660 8130 14716
rect 8130 14660 8134 14716
rect 8070 14656 8134 14660
rect 8150 14716 8214 14720
rect 8150 14660 8154 14716
rect 8154 14660 8210 14716
rect 8210 14660 8214 14716
rect 8150 14656 8214 14660
rect 8230 14716 8294 14720
rect 8230 14660 8234 14716
rect 8234 14660 8290 14716
rect 8290 14660 8294 14716
rect 8230 14656 8294 14660
rect 15580 14716 15644 14720
rect 15580 14660 15584 14716
rect 15584 14660 15640 14716
rect 15640 14660 15644 14716
rect 15580 14656 15644 14660
rect 15660 14716 15724 14720
rect 15660 14660 15664 14716
rect 15664 14660 15720 14716
rect 15720 14660 15724 14716
rect 15660 14656 15724 14660
rect 15740 14716 15804 14720
rect 15740 14660 15744 14716
rect 15744 14660 15800 14716
rect 15800 14660 15804 14716
rect 15740 14656 15804 14660
rect 15820 14716 15884 14720
rect 15820 14660 15824 14716
rect 15824 14660 15880 14716
rect 15880 14660 15884 14716
rect 15820 14656 15884 14660
rect 23170 14716 23234 14720
rect 23170 14660 23174 14716
rect 23174 14660 23230 14716
rect 23230 14660 23234 14716
rect 23170 14656 23234 14660
rect 23250 14716 23314 14720
rect 23250 14660 23254 14716
rect 23254 14660 23310 14716
rect 23310 14660 23314 14716
rect 23250 14656 23314 14660
rect 23330 14716 23394 14720
rect 23330 14660 23334 14716
rect 23334 14660 23390 14716
rect 23390 14660 23394 14716
rect 23330 14656 23394 14660
rect 23410 14716 23474 14720
rect 23410 14660 23414 14716
rect 23414 14660 23470 14716
rect 23470 14660 23474 14716
rect 23410 14656 23474 14660
rect 30760 14716 30824 14720
rect 30760 14660 30764 14716
rect 30764 14660 30820 14716
rect 30820 14660 30824 14716
rect 30760 14656 30824 14660
rect 30840 14716 30904 14720
rect 30840 14660 30844 14716
rect 30844 14660 30900 14716
rect 30900 14660 30904 14716
rect 30840 14656 30904 14660
rect 30920 14716 30984 14720
rect 30920 14660 30924 14716
rect 30924 14660 30980 14716
rect 30980 14660 30984 14716
rect 30920 14656 30984 14660
rect 31000 14716 31064 14720
rect 31000 14660 31004 14716
rect 31004 14660 31060 14716
rect 31060 14660 31064 14716
rect 31000 14656 31064 14660
rect 4195 14172 4259 14176
rect 4195 14116 4199 14172
rect 4199 14116 4255 14172
rect 4255 14116 4259 14172
rect 4195 14112 4259 14116
rect 4275 14172 4339 14176
rect 4275 14116 4279 14172
rect 4279 14116 4335 14172
rect 4335 14116 4339 14172
rect 4275 14112 4339 14116
rect 4355 14172 4419 14176
rect 4355 14116 4359 14172
rect 4359 14116 4415 14172
rect 4415 14116 4419 14172
rect 4355 14112 4419 14116
rect 4435 14172 4499 14176
rect 4435 14116 4439 14172
rect 4439 14116 4495 14172
rect 4495 14116 4499 14172
rect 4435 14112 4499 14116
rect 11785 14172 11849 14176
rect 11785 14116 11789 14172
rect 11789 14116 11845 14172
rect 11845 14116 11849 14172
rect 11785 14112 11849 14116
rect 11865 14172 11929 14176
rect 11865 14116 11869 14172
rect 11869 14116 11925 14172
rect 11925 14116 11929 14172
rect 11865 14112 11929 14116
rect 11945 14172 12009 14176
rect 11945 14116 11949 14172
rect 11949 14116 12005 14172
rect 12005 14116 12009 14172
rect 11945 14112 12009 14116
rect 12025 14172 12089 14176
rect 12025 14116 12029 14172
rect 12029 14116 12085 14172
rect 12085 14116 12089 14172
rect 12025 14112 12089 14116
rect 19375 14172 19439 14176
rect 19375 14116 19379 14172
rect 19379 14116 19435 14172
rect 19435 14116 19439 14172
rect 19375 14112 19439 14116
rect 19455 14172 19519 14176
rect 19455 14116 19459 14172
rect 19459 14116 19515 14172
rect 19515 14116 19519 14172
rect 19455 14112 19519 14116
rect 19535 14172 19599 14176
rect 19535 14116 19539 14172
rect 19539 14116 19595 14172
rect 19595 14116 19599 14172
rect 19535 14112 19599 14116
rect 19615 14172 19679 14176
rect 19615 14116 19619 14172
rect 19619 14116 19675 14172
rect 19675 14116 19679 14172
rect 19615 14112 19679 14116
rect 26965 14172 27029 14176
rect 26965 14116 26969 14172
rect 26969 14116 27025 14172
rect 27025 14116 27029 14172
rect 26965 14112 27029 14116
rect 27045 14172 27109 14176
rect 27045 14116 27049 14172
rect 27049 14116 27105 14172
rect 27105 14116 27109 14172
rect 27045 14112 27109 14116
rect 27125 14172 27189 14176
rect 27125 14116 27129 14172
rect 27129 14116 27185 14172
rect 27185 14116 27189 14172
rect 27125 14112 27189 14116
rect 27205 14172 27269 14176
rect 27205 14116 27209 14172
rect 27209 14116 27265 14172
rect 27265 14116 27269 14172
rect 27205 14112 27269 14116
rect 5396 13908 5460 13972
rect 8892 13696 8956 13700
rect 8892 13640 8942 13696
rect 8942 13640 8956 13696
rect 8892 13636 8956 13640
rect 29684 13636 29748 13700
rect 7990 13628 8054 13632
rect 7990 13572 7994 13628
rect 7994 13572 8050 13628
rect 8050 13572 8054 13628
rect 7990 13568 8054 13572
rect 8070 13628 8134 13632
rect 8070 13572 8074 13628
rect 8074 13572 8130 13628
rect 8130 13572 8134 13628
rect 8070 13568 8134 13572
rect 8150 13628 8214 13632
rect 8150 13572 8154 13628
rect 8154 13572 8210 13628
rect 8210 13572 8214 13628
rect 8150 13568 8214 13572
rect 8230 13628 8294 13632
rect 8230 13572 8234 13628
rect 8234 13572 8290 13628
rect 8290 13572 8294 13628
rect 8230 13568 8294 13572
rect 15580 13628 15644 13632
rect 15580 13572 15584 13628
rect 15584 13572 15640 13628
rect 15640 13572 15644 13628
rect 15580 13568 15644 13572
rect 15660 13628 15724 13632
rect 15660 13572 15664 13628
rect 15664 13572 15720 13628
rect 15720 13572 15724 13628
rect 15660 13568 15724 13572
rect 15740 13628 15804 13632
rect 15740 13572 15744 13628
rect 15744 13572 15800 13628
rect 15800 13572 15804 13628
rect 15740 13568 15804 13572
rect 15820 13628 15884 13632
rect 15820 13572 15824 13628
rect 15824 13572 15880 13628
rect 15880 13572 15884 13628
rect 15820 13568 15884 13572
rect 23170 13628 23234 13632
rect 23170 13572 23174 13628
rect 23174 13572 23230 13628
rect 23230 13572 23234 13628
rect 23170 13568 23234 13572
rect 23250 13628 23314 13632
rect 23250 13572 23254 13628
rect 23254 13572 23310 13628
rect 23310 13572 23314 13628
rect 23250 13568 23314 13572
rect 23330 13628 23394 13632
rect 23330 13572 23334 13628
rect 23334 13572 23390 13628
rect 23390 13572 23394 13628
rect 23330 13568 23394 13572
rect 23410 13628 23474 13632
rect 23410 13572 23414 13628
rect 23414 13572 23470 13628
rect 23470 13572 23474 13628
rect 23410 13568 23474 13572
rect 30760 13628 30824 13632
rect 30760 13572 30764 13628
rect 30764 13572 30820 13628
rect 30820 13572 30824 13628
rect 30760 13568 30824 13572
rect 30840 13628 30904 13632
rect 30840 13572 30844 13628
rect 30844 13572 30900 13628
rect 30900 13572 30904 13628
rect 30840 13568 30904 13572
rect 30920 13628 30984 13632
rect 30920 13572 30924 13628
rect 30924 13572 30980 13628
rect 30980 13572 30984 13628
rect 30920 13568 30984 13572
rect 31000 13628 31064 13632
rect 31000 13572 31004 13628
rect 31004 13572 31060 13628
rect 31060 13572 31064 13628
rect 31000 13568 31064 13572
rect 23980 13500 24044 13564
rect 4195 13084 4259 13088
rect 4195 13028 4199 13084
rect 4199 13028 4255 13084
rect 4255 13028 4259 13084
rect 4195 13024 4259 13028
rect 4275 13084 4339 13088
rect 4275 13028 4279 13084
rect 4279 13028 4335 13084
rect 4335 13028 4339 13084
rect 4275 13024 4339 13028
rect 4355 13084 4419 13088
rect 4355 13028 4359 13084
rect 4359 13028 4415 13084
rect 4415 13028 4419 13084
rect 4355 13024 4419 13028
rect 4435 13084 4499 13088
rect 4435 13028 4439 13084
rect 4439 13028 4495 13084
rect 4495 13028 4499 13084
rect 4435 13024 4499 13028
rect 11785 13084 11849 13088
rect 11785 13028 11789 13084
rect 11789 13028 11845 13084
rect 11845 13028 11849 13084
rect 11785 13024 11849 13028
rect 11865 13084 11929 13088
rect 11865 13028 11869 13084
rect 11869 13028 11925 13084
rect 11925 13028 11929 13084
rect 11865 13024 11929 13028
rect 11945 13084 12009 13088
rect 11945 13028 11949 13084
rect 11949 13028 12005 13084
rect 12005 13028 12009 13084
rect 11945 13024 12009 13028
rect 12025 13084 12089 13088
rect 12025 13028 12029 13084
rect 12029 13028 12085 13084
rect 12085 13028 12089 13084
rect 12025 13024 12089 13028
rect 19375 13084 19439 13088
rect 19375 13028 19379 13084
rect 19379 13028 19435 13084
rect 19435 13028 19439 13084
rect 19375 13024 19439 13028
rect 19455 13084 19519 13088
rect 19455 13028 19459 13084
rect 19459 13028 19515 13084
rect 19515 13028 19519 13084
rect 19455 13024 19519 13028
rect 19535 13084 19599 13088
rect 19535 13028 19539 13084
rect 19539 13028 19595 13084
rect 19595 13028 19599 13084
rect 19535 13024 19599 13028
rect 19615 13084 19679 13088
rect 19615 13028 19619 13084
rect 19619 13028 19675 13084
rect 19675 13028 19679 13084
rect 19615 13024 19679 13028
rect 26965 13084 27029 13088
rect 26965 13028 26969 13084
rect 26969 13028 27025 13084
rect 27025 13028 27029 13084
rect 26965 13024 27029 13028
rect 27045 13084 27109 13088
rect 27045 13028 27049 13084
rect 27049 13028 27105 13084
rect 27105 13028 27109 13084
rect 27045 13024 27109 13028
rect 27125 13084 27189 13088
rect 27125 13028 27129 13084
rect 27129 13028 27185 13084
rect 27185 13028 27189 13084
rect 27125 13024 27189 13028
rect 27205 13084 27269 13088
rect 27205 13028 27209 13084
rect 27209 13028 27265 13084
rect 27265 13028 27269 13084
rect 27205 13024 27269 13028
rect 10548 12956 10612 13020
rect 29132 13016 29196 13020
rect 29132 12960 29146 13016
rect 29146 12960 29196 13016
rect 29132 12956 29196 12960
rect 6316 12684 6380 12748
rect 7788 12684 7852 12748
rect 2820 12412 2884 12476
rect 7990 12540 8054 12544
rect 7990 12484 7994 12540
rect 7994 12484 8050 12540
rect 8050 12484 8054 12540
rect 7990 12480 8054 12484
rect 8070 12540 8134 12544
rect 8070 12484 8074 12540
rect 8074 12484 8130 12540
rect 8130 12484 8134 12540
rect 8070 12480 8134 12484
rect 8150 12540 8214 12544
rect 8150 12484 8154 12540
rect 8154 12484 8210 12540
rect 8210 12484 8214 12540
rect 8150 12480 8214 12484
rect 8230 12540 8294 12544
rect 8230 12484 8234 12540
rect 8234 12484 8290 12540
rect 8290 12484 8294 12540
rect 8230 12480 8294 12484
rect 15580 12540 15644 12544
rect 15580 12484 15584 12540
rect 15584 12484 15640 12540
rect 15640 12484 15644 12540
rect 15580 12480 15644 12484
rect 15660 12540 15724 12544
rect 15660 12484 15664 12540
rect 15664 12484 15720 12540
rect 15720 12484 15724 12540
rect 15660 12480 15724 12484
rect 15740 12540 15804 12544
rect 15740 12484 15744 12540
rect 15744 12484 15800 12540
rect 15800 12484 15804 12540
rect 15740 12480 15804 12484
rect 15820 12540 15884 12544
rect 15820 12484 15824 12540
rect 15824 12484 15880 12540
rect 15880 12484 15884 12540
rect 15820 12480 15884 12484
rect 23170 12540 23234 12544
rect 23170 12484 23174 12540
rect 23174 12484 23230 12540
rect 23230 12484 23234 12540
rect 23170 12480 23234 12484
rect 23250 12540 23314 12544
rect 23250 12484 23254 12540
rect 23254 12484 23310 12540
rect 23310 12484 23314 12540
rect 23250 12480 23314 12484
rect 23330 12540 23394 12544
rect 23330 12484 23334 12540
rect 23334 12484 23390 12540
rect 23390 12484 23394 12540
rect 23330 12480 23394 12484
rect 23410 12540 23474 12544
rect 23410 12484 23414 12540
rect 23414 12484 23470 12540
rect 23470 12484 23474 12540
rect 23410 12480 23474 12484
rect 30760 12540 30824 12544
rect 30760 12484 30764 12540
rect 30764 12484 30820 12540
rect 30820 12484 30824 12540
rect 30760 12480 30824 12484
rect 30840 12540 30904 12544
rect 30840 12484 30844 12540
rect 30844 12484 30900 12540
rect 30900 12484 30904 12540
rect 30840 12480 30904 12484
rect 30920 12540 30984 12544
rect 30920 12484 30924 12540
rect 30924 12484 30980 12540
rect 30980 12484 30984 12540
rect 30920 12480 30984 12484
rect 31000 12540 31064 12544
rect 31000 12484 31004 12540
rect 31004 12484 31060 12540
rect 31060 12484 31064 12540
rect 31000 12480 31064 12484
rect 27660 12412 27724 12476
rect 28764 12276 28828 12340
rect 12572 12140 12636 12204
rect 11468 12004 11532 12068
rect 4195 11996 4259 12000
rect 4195 11940 4199 11996
rect 4199 11940 4255 11996
rect 4255 11940 4259 11996
rect 4195 11936 4259 11940
rect 4275 11996 4339 12000
rect 4275 11940 4279 11996
rect 4279 11940 4335 11996
rect 4335 11940 4339 11996
rect 4275 11936 4339 11940
rect 4355 11996 4419 12000
rect 4355 11940 4359 11996
rect 4359 11940 4415 11996
rect 4415 11940 4419 11996
rect 4355 11936 4419 11940
rect 4435 11996 4499 12000
rect 4435 11940 4439 11996
rect 4439 11940 4495 11996
rect 4495 11940 4499 11996
rect 4435 11936 4499 11940
rect 11785 11996 11849 12000
rect 11785 11940 11789 11996
rect 11789 11940 11845 11996
rect 11845 11940 11849 11996
rect 11785 11936 11849 11940
rect 11865 11996 11929 12000
rect 11865 11940 11869 11996
rect 11869 11940 11925 11996
rect 11925 11940 11929 11996
rect 11865 11936 11929 11940
rect 11945 11996 12009 12000
rect 11945 11940 11949 11996
rect 11949 11940 12005 11996
rect 12005 11940 12009 11996
rect 11945 11936 12009 11940
rect 12025 11996 12089 12000
rect 12025 11940 12029 11996
rect 12029 11940 12085 11996
rect 12085 11940 12089 11996
rect 12025 11936 12089 11940
rect 19375 11996 19439 12000
rect 19375 11940 19379 11996
rect 19379 11940 19435 11996
rect 19435 11940 19439 11996
rect 19375 11936 19439 11940
rect 19455 11996 19519 12000
rect 19455 11940 19459 11996
rect 19459 11940 19515 11996
rect 19515 11940 19519 11996
rect 19455 11936 19519 11940
rect 19535 11996 19599 12000
rect 19535 11940 19539 11996
rect 19539 11940 19595 11996
rect 19595 11940 19599 11996
rect 19535 11936 19599 11940
rect 19615 11996 19679 12000
rect 19615 11940 19619 11996
rect 19619 11940 19675 11996
rect 19675 11940 19679 11996
rect 19615 11936 19679 11940
rect 26965 11996 27029 12000
rect 26965 11940 26969 11996
rect 26969 11940 27025 11996
rect 27025 11940 27029 11996
rect 26965 11936 27029 11940
rect 27045 11996 27109 12000
rect 27045 11940 27049 11996
rect 27049 11940 27105 11996
rect 27105 11940 27109 11996
rect 27045 11936 27109 11940
rect 27125 11996 27189 12000
rect 27125 11940 27129 11996
rect 27129 11940 27185 11996
rect 27185 11940 27189 11996
rect 27125 11936 27189 11940
rect 27205 11996 27269 12000
rect 27205 11940 27209 11996
rect 27209 11940 27265 11996
rect 27265 11940 27269 11996
rect 27205 11936 27269 11940
rect 11284 11732 11348 11796
rect 6684 11596 6748 11660
rect 7990 11452 8054 11456
rect 7990 11396 7994 11452
rect 7994 11396 8050 11452
rect 8050 11396 8054 11452
rect 7990 11392 8054 11396
rect 8070 11452 8134 11456
rect 8070 11396 8074 11452
rect 8074 11396 8130 11452
rect 8130 11396 8134 11452
rect 8070 11392 8134 11396
rect 8150 11452 8214 11456
rect 8150 11396 8154 11452
rect 8154 11396 8210 11452
rect 8210 11396 8214 11452
rect 8150 11392 8214 11396
rect 8230 11452 8294 11456
rect 8230 11396 8234 11452
rect 8234 11396 8290 11452
rect 8290 11396 8294 11452
rect 8230 11392 8294 11396
rect 15580 11452 15644 11456
rect 15580 11396 15584 11452
rect 15584 11396 15640 11452
rect 15640 11396 15644 11452
rect 15580 11392 15644 11396
rect 15660 11452 15724 11456
rect 15660 11396 15664 11452
rect 15664 11396 15720 11452
rect 15720 11396 15724 11452
rect 15660 11392 15724 11396
rect 15740 11452 15804 11456
rect 15740 11396 15744 11452
rect 15744 11396 15800 11452
rect 15800 11396 15804 11452
rect 15740 11392 15804 11396
rect 15820 11452 15884 11456
rect 15820 11396 15824 11452
rect 15824 11396 15880 11452
rect 15880 11396 15884 11452
rect 15820 11392 15884 11396
rect 23170 11452 23234 11456
rect 23170 11396 23174 11452
rect 23174 11396 23230 11452
rect 23230 11396 23234 11452
rect 23170 11392 23234 11396
rect 23250 11452 23314 11456
rect 23250 11396 23254 11452
rect 23254 11396 23310 11452
rect 23310 11396 23314 11452
rect 23250 11392 23314 11396
rect 23330 11452 23394 11456
rect 23330 11396 23334 11452
rect 23334 11396 23390 11452
rect 23390 11396 23394 11452
rect 23330 11392 23394 11396
rect 23410 11452 23474 11456
rect 23410 11396 23414 11452
rect 23414 11396 23470 11452
rect 23470 11396 23474 11452
rect 23410 11392 23474 11396
rect 30760 11452 30824 11456
rect 30760 11396 30764 11452
rect 30764 11396 30820 11452
rect 30820 11396 30824 11452
rect 30760 11392 30824 11396
rect 30840 11452 30904 11456
rect 30840 11396 30844 11452
rect 30844 11396 30900 11452
rect 30900 11396 30904 11452
rect 30840 11392 30904 11396
rect 30920 11452 30984 11456
rect 30920 11396 30924 11452
rect 30924 11396 30980 11452
rect 30980 11396 30984 11452
rect 30920 11392 30984 11396
rect 31000 11452 31064 11456
rect 31000 11396 31004 11452
rect 31004 11396 31060 11452
rect 31060 11396 31064 11452
rect 31000 11392 31064 11396
rect 8708 11384 8772 11388
rect 8708 11328 8722 11384
rect 8722 11328 8772 11384
rect 8708 11324 8772 11328
rect 7052 11052 7116 11116
rect 3004 10916 3068 10980
rect 4195 10908 4259 10912
rect 4195 10852 4199 10908
rect 4199 10852 4255 10908
rect 4255 10852 4259 10908
rect 4195 10848 4259 10852
rect 4275 10908 4339 10912
rect 4275 10852 4279 10908
rect 4279 10852 4335 10908
rect 4335 10852 4339 10908
rect 4275 10848 4339 10852
rect 4355 10908 4419 10912
rect 4355 10852 4359 10908
rect 4359 10852 4415 10908
rect 4415 10852 4419 10908
rect 4355 10848 4419 10852
rect 4435 10908 4499 10912
rect 4435 10852 4439 10908
rect 4439 10852 4495 10908
rect 4495 10852 4499 10908
rect 4435 10848 4499 10852
rect 11785 10908 11849 10912
rect 11785 10852 11789 10908
rect 11789 10852 11845 10908
rect 11845 10852 11849 10908
rect 11785 10848 11849 10852
rect 11865 10908 11929 10912
rect 11865 10852 11869 10908
rect 11869 10852 11925 10908
rect 11925 10852 11929 10908
rect 11865 10848 11929 10852
rect 11945 10908 12009 10912
rect 11945 10852 11949 10908
rect 11949 10852 12005 10908
rect 12005 10852 12009 10908
rect 11945 10848 12009 10852
rect 12025 10908 12089 10912
rect 12025 10852 12029 10908
rect 12029 10852 12085 10908
rect 12085 10852 12089 10908
rect 12025 10848 12089 10852
rect 19375 10908 19439 10912
rect 19375 10852 19379 10908
rect 19379 10852 19435 10908
rect 19435 10852 19439 10908
rect 19375 10848 19439 10852
rect 19455 10908 19519 10912
rect 19455 10852 19459 10908
rect 19459 10852 19515 10908
rect 19515 10852 19519 10908
rect 19455 10848 19519 10852
rect 19535 10908 19599 10912
rect 19535 10852 19539 10908
rect 19539 10852 19595 10908
rect 19595 10852 19599 10908
rect 19535 10848 19599 10852
rect 19615 10908 19679 10912
rect 19615 10852 19619 10908
rect 19619 10852 19675 10908
rect 19675 10852 19679 10908
rect 19615 10848 19679 10852
rect 26965 10908 27029 10912
rect 26965 10852 26969 10908
rect 26969 10852 27025 10908
rect 27025 10852 27029 10908
rect 26965 10848 27029 10852
rect 27045 10908 27109 10912
rect 27045 10852 27049 10908
rect 27049 10852 27105 10908
rect 27105 10852 27109 10908
rect 27045 10848 27109 10852
rect 27125 10908 27189 10912
rect 27125 10852 27129 10908
rect 27129 10852 27185 10908
rect 27185 10852 27189 10908
rect 27125 10848 27189 10852
rect 27205 10908 27269 10912
rect 27205 10852 27209 10908
rect 27209 10852 27265 10908
rect 27265 10852 27269 10908
rect 27205 10848 27269 10852
rect 6684 10644 6748 10708
rect 7990 10364 8054 10368
rect 7990 10308 7994 10364
rect 7994 10308 8050 10364
rect 8050 10308 8054 10364
rect 7990 10304 8054 10308
rect 8070 10364 8134 10368
rect 8070 10308 8074 10364
rect 8074 10308 8130 10364
rect 8130 10308 8134 10364
rect 8070 10304 8134 10308
rect 8150 10364 8214 10368
rect 8150 10308 8154 10364
rect 8154 10308 8210 10364
rect 8210 10308 8214 10364
rect 8150 10304 8214 10308
rect 8230 10364 8294 10368
rect 8230 10308 8234 10364
rect 8234 10308 8290 10364
rect 8290 10308 8294 10364
rect 8230 10304 8294 10308
rect 15580 10364 15644 10368
rect 15580 10308 15584 10364
rect 15584 10308 15640 10364
rect 15640 10308 15644 10364
rect 15580 10304 15644 10308
rect 15660 10364 15724 10368
rect 15660 10308 15664 10364
rect 15664 10308 15720 10364
rect 15720 10308 15724 10364
rect 15660 10304 15724 10308
rect 15740 10364 15804 10368
rect 15740 10308 15744 10364
rect 15744 10308 15800 10364
rect 15800 10308 15804 10364
rect 15740 10304 15804 10308
rect 15820 10364 15884 10368
rect 15820 10308 15824 10364
rect 15824 10308 15880 10364
rect 15880 10308 15884 10364
rect 15820 10304 15884 10308
rect 23170 10364 23234 10368
rect 23170 10308 23174 10364
rect 23174 10308 23230 10364
rect 23230 10308 23234 10364
rect 23170 10304 23234 10308
rect 23250 10364 23314 10368
rect 23250 10308 23254 10364
rect 23254 10308 23310 10364
rect 23310 10308 23314 10364
rect 23250 10304 23314 10308
rect 23330 10364 23394 10368
rect 23330 10308 23334 10364
rect 23334 10308 23390 10364
rect 23390 10308 23394 10364
rect 23330 10304 23394 10308
rect 23410 10364 23474 10368
rect 23410 10308 23414 10364
rect 23414 10308 23470 10364
rect 23470 10308 23474 10364
rect 23410 10304 23474 10308
rect 30760 10364 30824 10368
rect 30760 10308 30764 10364
rect 30764 10308 30820 10364
rect 30820 10308 30824 10364
rect 30760 10304 30824 10308
rect 30840 10364 30904 10368
rect 30840 10308 30844 10364
rect 30844 10308 30900 10364
rect 30900 10308 30904 10364
rect 30840 10304 30904 10308
rect 30920 10364 30984 10368
rect 30920 10308 30924 10364
rect 30924 10308 30980 10364
rect 30980 10308 30984 10364
rect 30920 10304 30984 10308
rect 31000 10364 31064 10368
rect 31000 10308 31004 10364
rect 31004 10308 31060 10364
rect 31060 10308 31064 10364
rect 31000 10304 31064 10308
rect 17908 10236 17972 10300
rect 4195 9820 4259 9824
rect 4195 9764 4199 9820
rect 4199 9764 4255 9820
rect 4255 9764 4259 9820
rect 4195 9760 4259 9764
rect 4275 9820 4339 9824
rect 4275 9764 4279 9820
rect 4279 9764 4335 9820
rect 4335 9764 4339 9820
rect 4275 9760 4339 9764
rect 4355 9820 4419 9824
rect 4355 9764 4359 9820
rect 4359 9764 4415 9820
rect 4415 9764 4419 9820
rect 4355 9760 4419 9764
rect 4435 9820 4499 9824
rect 4435 9764 4439 9820
rect 4439 9764 4495 9820
rect 4495 9764 4499 9820
rect 4435 9760 4499 9764
rect 11785 9820 11849 9824
rect 11785 9764 11789 9820
rect 11789 9764 11845 9820
rect 11845 9764 11849 9820
rect 11785 9760 11849 9764
rect 11865 9820 11929 9824
rect 11865 9764 11869 9820
rect 11869 9764 11925 9820
rect 11925 9764 11929 9820
rect 11865 9760 11929 9764
rect 11945 9820 12009 9824
rect 11945 9764 11949 9820
rect 11949 9764 12005 9820
rect 12005 9764 12009 9820
rect 11945 9760 12009 9764
rect 12025 9820 12089 9824
rect 12025 9764 12029 9820
rect 12029 9764 12085 9820
rect 12085 9764 12089 9820
rect 12025 9760 12089 9764
rect 19375 9820 19439 9824
rect 19375 9764 19379 9820
rect 19379 9764 19435 9820
rect 19435 9764 19439 9820
rect 19375 9760 19439 9764
rect 19455 9820 19519 9824
rect 19455 9764 19459 9820
rect 19459 9764 19515 9820
rect 19515 9764 19519 9820
rect 19455 9760 19519 9764
rect 19535 9820 19599 9824
rect 19535 9764 19539 9820
rect 19539 9764 19595 9820
rect 19595 9764 19599 9820
rect 19535 9760 19599 9764
rect 19615 9820 19679 9824
rect 19615 9764 19619 9820
rect 19619 9764 19675 9820
rect 19675 9764 19679 9820
rect 19615 9760 19679 9764
rect 26965 9820 27029 9824
rect 26965 9764 26969 9820
rect 26969 9764 27025 9820
rect 27025 9764 27029 9820
rect 26965 9760 27029 9764
rect 27045 9820 27109 9824
rect 27045 9764 27049 9820
rect 27049 9764 27105 9820
rect 27105 9764 27109 9820
rect 27045 9760 27109 9764
rect 27125 9820 27189 9824
rect 27125 9764 27129 9820
rect 27129 9764 27185 9820
rect 27185 9764 27189 9820
rect 27125 9760 27189 9764
rect 27205 9820 27269 9824
rect 27205 9764 27209 9820
rect 27209 9764 27265 9820
rect 27265 9764 27269 9820
rect 27205 9760 27269 9764
rect 6132 9692 6196 9756
rect 6868 9692 6932 9756
rect 6316 9556 6380 9620
rect 7236 9556 7300 9620
rect 5028 9420 5092 9484
rect 7990 9276 8054 9280
rect 7990 9220 7994 9276
rect 7994 9220 8050 9276
rect 8050 9220 8054 9276
rect 7990 9216 8054 9220
rect 8070 9276 8134 9280
rect 8070 9220 8074 9276
rect 8074 9220 8130 9276
rect 8130 9220 8134 9276
rect 8070 9216 8134 9220
rect 8150 9276 8214 9280
rect 8150 9220 8154 9276
rect 8154 9220 8210 9276
rect 8210 9220 8214 9276
rect 8150 9216 8214 9220
rect 8230 9276 8294 9280
rect 8230 9220 8234 9276
rect 8234 9220 8290 9276
rect 8290 9220 8294 9276
rect 8230 9216 8294 9220
rect 15580 9276 15644 9280
rect 15580 9220 15584 9276
rect 15584 9220 15640 9276
rect 15640 9220 15644 9276
rect 15580 9216 15644 9220
rect 15660 9276 15724 9280
rect 15660 9220 15664 9276
rect 15664 9220 15720 9276
rect 15720 9220 15724 9276
rect 15660 9216 15724 9220
rect 15740 9276 15804 9280
rect 15740 9220 15744 9276
rect 15744 9220 15800 9276
rect 15800 9220 15804 9276
rect 15740 9216 15804 9220
rect 15820 9276 15884 9280
rect 15820 9220 15824 9276
rect 15824 9220 15880 9276
rect 15880 9220 15884 9276
rect 15820 9216 15884 9220
rect 23170 9276 23234 9280
rect 23170 9220 23174 9276
rect 23174 9220 23230 9276
rect 23230 9220 23234 9276
rect 23170 9216 23234 9220
rect 23250 9276 23314 9280
rect 23250 9220 23254 9276
rect 23254 9220 23310 9276
rect 23310 9220 23314 9276
rect 23250 9216 23314 9220
rect 23330 9276 23394 9280
rect 23330 9220 23334 9276
rect 23334 9220 23390 9276
rect 23390 9220 23394 9276
rect 23330 9216 23394 9220
rect 23410 9276 23474 9280
rect 23410 9220 23414 9276
rect 23414 9220 23470 9276
rect 23470 9220 23474 9276
rect 23410 9216 23474 9220
rect 30760 9276 30824 9280
rect 30760 9220 30764 9276
rect 30764 9220 30820 9276
rect 30820 9220 30824 9276
rect 30760 9216 30824 9220
rect 30840 9276 30904 9280
rect 30840 9220 30844 9276
rect 30844 9220 30900 9276
rect 30900 9220 30904 9276
rect 30840 9216 30904 9220
rect 30920 9276 30984 9280
rect 30920 9220 30924 9276
rect 30924 9220 30980 9276
rect 30980 9220 30984 9276
rect 30920 9216 30984 9220
rect 31000 9276 31064 9280
rect 31000 9220 31004 9276
rect 31004 9220 31060 9276
rect 31060 9220 31064 9276
rect 31000 9216 31064 9220
rect 24716 8876 24780 8940
rect 4195 8732 4259 8736
rect 4195 8676 4199 8732
rect 4199 8676 4255 8732
rect 4255 8676 4259 8732
rect 4195 8672 4259 8676
rect 4275 8732 4339 8736
rect 4275 8676 4279 8732
rect 4279 8676 4335 8732
rect 4335 8676 4339 8732
rect 4275 8672 4339 8676
rect 4355 8732 4419 8736
rect 4355 8676 4359 8732
rect 4359 8676 4415 8732
rect 4415 8676 4419 8732
rect 4355 8672 4419 8676
rect 4435 8732 4499 8736
rect 4435 8676 4439 8732
rect 4439 8676 4495 8732
rect 4495 8676 4499 8732
rect 4435 8672 4499 8676
rect 11785 8732 11849 8736
rect 11785 8676 11789 8732
rect 11789 8676 11845 8732
rect 11845 8676 11849 8732
rect 11785 8672 11849 8676
rect 11865 8732 11929 8736
rect 11865 8676 11869 8732
rect 11869 8676 11925 8732
rect 11925 8676 11929 8732
rect 11865 8672 11929 8676
rect 11945 8732 12009 8736
rect 11945 8676 11949 8732
rect 11949 8676 12005 8732
rect 12005 8676 12009 8732
rect 11945 8672 12009 8676
rect 12025 8732 12089 8736
rect 12025 8676 12029 8732
rect 12029 8676 12085 8732
rect 12085 8676 12089 8732
rect 12025 8672 12089 8676
rect 19375 8732 19439 8736
rect 19375 8676 19379 8732
rect 19379 8676 19435 8732
rect 19435 8676 19439 8732
rect 19375 8672 19439 8676
rect 19455 8732 19519 8736
rect 19455 8676 19459 8732
rect 19459 8676 19515 8732
rect 19515 8676 19519 8732
rect 19455 8672 19519 8676
rect 19535 8732 19599 8736
rect 19535 8676 19539 8732
rect 19539 8676 19595 8732
rect 19595 8676 19599 8732
rect 19535 8672 19599 8676
rect 19615 8732 19679 8736
rect 19615 8676 19619 8732
rect 19619 8676 19675 8732
rect 19675 8676 19679 8732
rect 19615 8672 19679 8676
rect 26965 8732 27029 8736
rect 26965 8676 26969 8732
rect 26969 8676 27025 8732
rect 27025 8676 27029 8732
rect 26965 8672 27029 8676
rect 27045 8732 27109 8736
rect 27045 8676 27049 8732
rect 27049 8676 27105 8732
rect 27105 8676 27109 8732
rect 27045 8672 27109 8676
rect 27125 8732 27189 8736
rect 27125 8676 27129 8732
rect 27129 8676 27185 8732
rect 27185 8676 27189 8732
rect 27125 8672 27189 8676
rect 27205 8732 27269 8736
rect 27205 8676 27209 8732
rect 27209 8676 27265 8732
rect 27265 8676 27269 8732
rect 27205 8672 27269 8676
rect 5948 8196 6012 8260
rect 7052 8196 7116 8260
rect 10180 8196 10244 8260
rect 7990 8188 8054 8192
rect 7990 8132 7994 8188
rect 7994 8132 8050 8188
rect 8050 8132 8054 8188
rect 7990 8128 8054 8132
rect 8070 8188 8134 8192
rect 8070 8132 8074 8188
rect 8074 8132 8130 8188
rect 8130 8132 8134 8188
rect 8070 8128 8134 8132
rect 8150 8188 8214 8192
rect 8150 8132 8154 8188
rect 8154 8132 8210 8188
rect 8210 8132 8214 8188
rect 8150 8128 8214 8132
rect 8230 8188 8294 8192
rect 8230 8132 8234 8188
rect 8234 8132 8290 8188
rect 8290 8132 8294 8188
rect 8230 8128 8294 8132
rect 15580 8188 15644 8192
rect 15580 8132 15584 8188
rect 15584 8132 15640 8188
rect 15640 8132 15644 8188
rect 15580 8128 15644 8132
rect 15660 8188 15724 8192
rect 15660 8132 15664 8188
rect 15664 8132 15720 8188
rect 15720 8132 15724 8188
rect 15660 8128 15724 8132
rect 15740 8188 15804 8192
rect 15740 8132 15744 8188
rect 15744 8132 15800 8188
rect 15800 8132 15804 8188
rect 15740 8128 15804 8132
rect 15820 8188 15884 8192
rect 15820 8132 15824 8188
rect 15824 8132 15880 8188
rect 15880 8132 15884 8188
rect 15820 8128 15884 8132
rect 23170 8188 23234 8192
rect 23170 8132 23174 8188
rect 23174 8132 23230 8188
rect 23230 8132 23234 8188
rect 23170 8128 23234 8132
rect 23250 8188 23314 8192
rect 23250 8132 23254 8188
rect 23254 8132 23310 8188
rect 23310 8132 23314 8188
rect 23250 8128 23314 8132
rect 23330 8188 23394 8192
rect 23330 8132 23334 8188
rect 23334 8132 23390 8188
rect 23390 8132 23394 8188
rect 23330 8128 23394 8132
rect 23410 8188 23474 8192
rect 23410 8132 23414 8188
rect 23414 8132 23470 8188
rect 23470 8132 23474 8188
rect 23410 8128 23474 8132
rect 30760 8188 30824 8192
rect 30760 8132 30764 8188
rect 30764 8132 30820 8188
rect 30820 8132 30824 8188
rect 30760 8128 30824 8132
rect 30840 8188 30904 8192
rect 30840 8132 30844 8188
rect 30844 8132 30900 8188
rect 30900 8132 30904 8188
rect 30840 8128 30904 8132
rect 30920 8188 30984 8192
rect 30920 8132 30924 8188
rect 30924 8132 30980 8188
rect 30980 8132 30984 8188
rect 30920 8128 30984 8132
rect 31000 8188 31064 8192
rect 31000 8132 31004 8188
rect 31004 8132 31060 8188
rect 31060 8132 31064 8188
rect 31000 8128 31064 8132
rect 26188 7924 26252 7988
rect 4195 7644 4259 7648
rect 4195 7588 4199 7644
rect 4199 7588 4255 7644
rect 4255 7588 4259 7644
rect 4195 7584 4259 7588
rect 4275 7644 4339 7648
rect 4275 7588 4279 7644
rect 4279 7588 4335 7644
rect 4335 7588 4339 7644
rect 4275 7584 4339 7588
rect 4355 7644 4419 7648
rect 4355 7588 4359 7644
rect 4359 7588 4415 7644
rect 4415 7588 4419 7644
rect 4355 7584 4419 7588
rect 4435 7644 4499 7648
rect 4435 7588 4439 7644
rect 4439 7588 4495 7644
rect 4495 7588 4499 7644
rect 4435 7584 4499 7588
rect 6868 7380 6932 7444
rect 11785 7644 11849 7648
rect 11785 7588 11789 7644
rect 11789 7588 11845 7644
rect 11845 7588 11849 7644
rect 11785 7584 11849 7588
rect 11865 7644 11929 7648
rect 11865 7588 11869 7644
rect 11869 7588 11925 7644
rect 11925 7588 11929 7644
rect 11865 7584 11929 7588
rect 11945 7644 12009 7648
rect 11945 7588 11949 7644
rect 11949 7588 12005 7644
rect 12005 7588 12009 7644
rect 11945 7584 12009 7588
rect 12025 7644 12089 7648
rect 12025 7588 12029 7644
rect 12029 7588 12085 7644
rect 12085 7588 12089 7644
rect 12025 7584 12089 7588
rect 19375 7644 19439 7648
rect 19375 7588 19379 7644
rect 19379 7588 19435 7644
rect 19435 7588 19439 7644
rect 19375 7584 19439 7588
rect 19455 7644 19519 7648
rect 19455 7588 19459 7644
rect 19459 7588 19515 7644
rect 19515 7588 19519 7644
rect 19455 7584 19519 7588
rect 19535 7644 19599 7648
rect 19535 7588 19539 7644
rect 19539 7588 19595 7644
rect 19595 7588 19599 7644
rect 19535 7584 19599 7588
rect 19615 7644 19679 7648
rect 19615 7588 19619 7644
rect 19619 7588 19675 7644
rect 19675 7588 19679 7644
rect 19615 7584 19679 7588
rect 26965 7644 27029 7648
rect 26965 7588 26969 7644
rect 26969 7588 27025 7644
rect 27025 7588 27029 7644
rect 26965 7584 27029 7588
rect 27045 7644 27109 7648
rect 27045 7588 27049 7644
rect 27049 7588 27105 7644
rect 27105 7588 27109 7644
rect 27045 7584 27109 7588
rect 27125 7644 27189 7648
rect 27125 7588 27129 7644
rect 27129 7588 27185 7644
rect 27185 7588 27189 7644
rect 27125 7584 27189 7588
rect 27205 7644 27269 7648
rect 27205 7588 27209 7644
rect 27209 7588 27265 7644
rect 27265 7588 27269 7644
rect 27205 7584 27269 7588
rect 16804 7108 16868 7172
rect 7990 7100 8054 7104
rect 7990 7044 7994 7100
rect 7994 7044 8050 7100
rect 8050 7044 8054 7100
rect 7990 7040 8054 7044
rect 8070 7100 8134 7104
rect 8070 7044 8074 7100
rect 8074 7044 8130 7100
rect 8130 7044 8134 7100
rect 8070 7040 8134 7044
rect 8150 7100 8214 7104
rect 8150 7044 8154 7100
rect 8154 7044 8210 7100
rect 8210 7044 8214 7100
rect 8150 7040 8214 7044
rect 8230 7100 8294 7104
rect 8230 7044 8234 7100
rect 8234 7044 8290 7100
rect 8290 7044 8294 7100
rect 8230 7040 8294 7044
rect 15580 7100 15644 7104
rect 15580 7044 15584 7100
rect 15584 7044 15640 7100
rect 15640 7044 15644 7100
rect 15580 7040 15644 7044
rect 15660 7100 15724 7104
rect 15660 7044 15664 7100
rect 15664 7044 15720 7100
rect 15720 7044 15724 7100
rect 15660 7040 15724 7044
rect 15740 7100 15804 7104
rect 15740 7044 15744 7100
rect 15744 7044 15800 7100
rect 15800 7044 15804 7100
rect 15740 7040 15804 7044
rect 15820 7100 15884 7104
rect 15820 7044 15824 7100
rect 15824 7044 15880 7100
rect 15880 7044 15884 7100
rect 15820 7040 15884 7044
rect 23170 7100 23234 7104
rect 23170 7044 23174 7100
rect 23174 7044 23230 7100
rect 23230 7044 23234 7100
rect 23170 7040 23234 7044
rect 23250 7100 23314 7104
rect 23250 7044 23254 7100
rect 23254 7044 23310 7100
rect 23310 7044 23314 7100
rect 23250 7040 23314 7044
rect 23330 7100 23394 7104
rect 23330 7044 23334 7100
rect 23334 7044 23390 7100
rect 23390 7044 23394 7100
rect 23330 7040 23394 7044
rect 23410 7100 23474 7104
rect 23410 7044 23414 7100
rect 23414 7044 23470 7100
rect 23470 7044 23474 7100
rect 23410 7040 23474 7044
rect 30760 7100 30824 7104
rect 30760 7044 30764 7100
rect 30764 7044 30820 7100
rect 30820 7044 30824 7100
rect 30760 7040 30824 7044
rect 30840 7100 30904 7104
rect 30840 7044 30844 7100
rect 30844 7044 30900 7100
rect 30900 7044 30904 7100
rect 30840 7040 30904 7044
rect 30920 7100 30984 7104
rect 30920 7044 30924 7100
rect 30924 7044 30980 7100
rect 30980 7044 30984 7100
rect 30920 7040 30984 7044
rect 31000 7100 31064 7104
rect 31000 7044 31004 7100
rect 31004 7044 31060 7100
rect 31060 7044 31064 7100
rect 31000 7040 31064 7044
rect 6132 6972 6196 7036
rect 16620 6972 16684 7036
rect 6684 6700 6748 6764
rect 4195 6556 4259 6560
rect 4195 6500 4199 6556
rect 4199 6500 4255 6556
rect 4255 6500 4259 6556
rect 4195 6496 4259 6500
rect 4275 6556 4339 6560
rect 4275 6500 4279 6556
rect 4279 6500 4335 6556
rect 4335 6500 4339 6556
rect 4275 6496 4339 6500
rect 4355 6556 4419 6560
rect 4355 6500 4359 6556
rect 4359 6500 4415 6556
rect 4415 6500 4419 6556
rect 4355 6496 4419 6500
rect 4435 6556 4499 6560
rect 4435 6500 4439 6556
rect 4439 6500 4495 6556
rect 4495 6500 4499 6556
rect 4435 6496 4499 6500
rect 11785 6556 11849 6560
rect 11785 6500 11789 6556
rect 11789 6500 11845 6556
rect 11845 6500 11849 6556
rect 11785 6496 11849 6500
rect 11865 6556 11929 6560
rect 11865 6500 11869 6556
rect 11869 6500 11925 6556
rect 11925 6500 11929 6556
rect 11865 6496 11929 6500
rect 11945 6556 12009 6560
rect 11945 6500 11949 6556
rect 11949 6500 12005 6556
rect 12005 6500 12009 6556
rect 11945 6496 12009 6500
rect 12025 6556 12089 6560
rect 12025 6500 12029 6556
rect 12029 6500 12085 6556
rect 12085 6500 12089 6556
rect 12025 6496 12089 6500
rect 19375 6556 19439 6560
rect 19375 6500 19379 6556
rect 19379 6500 19435 6556
rect 19435 6500 19439 6556
rect 19375 6496 19439 6500
rect 19455 6556 19519 6560
rect 19455 6500 19459 6556
rect 19459 6500 19515 6556
rect 19515 6500 19519 6556
rect 19455 6496 19519 6500
rect 19535 6556 19599 6560
rect 19535 6500 19539 6556
rect 19539 6500 19595 6556
rect 19595 6500 19599 6556
rect 19535 6496 19599 6500
rect 19615 6556 19679 6560
rect 19615 6500 19619 6556
rect 19619 6500 19675 6556
rect 19675 6500 19679 6556
rect 19615 6496 19679 6500
rect 26965 6556 27029 6560
rect 26965 6500 26969 6556
rect 26969 6500 27025 6556
rect 27025 6500 27029 6556
rect 26965 6496 27029 6500
rect 27045 6556 27109 6560
rect 27045 6500 27049 6556
rect 27049 6500 27105 6556
rect 27105 6500 27109 6556
rect 27045 6496 27109 6500
rect 27125 6556 27189 6560
rect 27125 6500 27129 6556
rect 27129 6500 27185 6556
rect 27185 6500 27189 6556
rect 27125 6496 27189 6500
rect 27205 6556 27269 6560
rect 27205 6500 27209 6556
rect 27209 6500 27265 6556
rect 27265 6500 27269 6556
rect 27205 6496 27269 6500
rect 7990 6012 8054 6016
rect 7990 5956 7994 6012
rect 7994 5956 8050 6012
rect 8050 5956 8054 6012
rect 7990 5952 8054 5956
rect 8070 6012 8134 6016
rect 8070 5956 8074 6012
rect 8074 5956 8130 6012
rect 8130 5956 8134 6012
rect 8070 5952 8134 5956
rect 8150 6012 8214 6016
rect 8150 5956 8154 6012
rect 8154 5956 8210 6012
rect 8210 5956 8214 6012
rect 8150 5952 8214 5956
rect 8230 6012 8294 6016
rect 8230 5956 8234 6012
rect 8234 5956 8290 6012
rect 8290 5956 8294 6012
rect 8230 5952 8294 5956
rect 15580 6012 15644 6016
rect 15580 5956 15584 6012
rect 15584 5956 15640 6012
rect 15640 5956 15644 6012
rect 15580 5952 15644 5956
rect 15660 6012 15724 6016
rect 15660 5956 15664 6012
rect 15664 5956 15720 6012
rect 15720 5956 15724 6012
rect 15660 5952 15724 5956
rect 15740 6012 15804 6016
rect 15740 5956 15744 6012
rect 15744 5956 15800 6012
rect 15800 5956 15804 6012
rect 15740 5952 15804 5956
rect 15820 6012 15884 6016
rect 15820 5956 15824 6012
rect 15824 5956 15880 6012
rect 15880 5956 15884 6012
rect 15820 5952 15884 5956
rect 23170 6012 23234 6016
rect 23170 5956 23174 6012
rect 23174 5956 23230 6012
rect 23230 5956 23234 6012
rect 23170 5952 23234 5956
rect 23250 6012 23314 6016
rect 23250 5956 23254 6012
rect 23254 5956 23310 6012
rect 23310 5956 23314 6012
rect 23250 5952 23314 5956
rect 23330 6012 23394 6016
rect 23330 5956 23334 6012
rect 23334 5956 23390 6012
rect 23390 5956 23394 6012
rect 23330 5952 23394 5956
rect 23410 6012 23474 6016
rect 23410 5956 23414 6012
rect 23414 5956 23470 6012
rect 23470 5956 23474 6012
rect 23410 5952 23474 5956
rect 30760 6012 30824 6016
rect 30760 5956 30764 6012
rect 30764 5956 30820 6012
rect 30820 5956 30824 6012
rect 30760 5952 30824 5956
rect 30840 6012 30904 6016
rect 30840 5956 30844 6012
rect 30844 5956 30900 6012
rect 30900 5956 30904 6012
rect 30840 5952 30904 5956
rect 30920 6012 30984 6016
rect 30920 5956 30924 6012
rect 30924 5956 30980 6012
rect 30980 5956 30984 6012
rect 30920 5952 30984 5956
rect 31000 6012 31064 6016
rect 31000 5956 31004 6012
rect 31004 5956 31060 6012
rect 31060 5956 31064 6012
rect 31000 5952 31064 5956
rect 3004 5476 3068 5540
rect 8524 5476 8588 5540
rect 26188 5476 26252 5540
rect 4195 5468 4259 5472
rect 4195 5412 4199 5468
rect 4199 5412 4255 5468
rect 4255 5412 4259 5468
rect 4195 5408 4259 5412
rect 4275 5468 4339 5472
rect 4275 5412 4279 5468
rect 4279 5412 4335 5468
rect 4335 5412 4339 5468
rect 4275 5408 4339 5412
rect 4355 5468 4419 5472
rect 4355 5412 4359 5468
rect 4359 5412 4415 5468
rect 4415 5412 4419 5468
rect 4355 5408 4419 5412
rect 4435 5468 4499 5472
rect 4435 5412 4439 5468
rect 4439 5412 4495 5468
rect 4495 5412 4499 5468
rect 4435 5408 4499 5412
rect 11785 5468 11849 5472
rect 11785 5412 11789 5468
rect 11789 5412 11845 5468
rect 11845 5412 11849 5468
rect 11785 5408 11849 5412
rect 11865 5468 11929 5472
rect 11865 5412 11869 5468
rect 11869 5412 11925 5468
rect 11925 5412 11929 5468
rect 11865 5408 11929 5412
rect 11945 5468 12009 5472
rect 11945 5412 11949 5468
rect 11949 5412 12005 5468
rect 12005 5412 12009 5468
rect 11945 5408 12009 5412
rect 12025 5468 12089 5472
rect 12025 5412 12029 5468
rect 12029 5412 12085 5468
rect 12085 5412 12089 5468
rect 12025 5408 12089 5412
rect 19375 5468 19439 5472
rect 19375 5412 19379 5468
rect 19379 5412 19435 5468
rect 19435 5412 19439 5468
rect 19375 5408 19439 5412
rect 19455 5468 19519 5472
rect 19455 5412 19459 5468
rect 19459 5412 19515 5468
rect 19515 5412 19519 5468
rect 19455 5408 19519 5412
rect 19535 5468 19599 5472
rect 19535 5412 19539 5468
rect 19539 5412 19595 5468
rect 19595 5412 19599 5468
rect 19535 5408 19599 5412
rect 19615 5468 19679 5472
rect 19615 5412 19619 5468
rect 19619 5412 19675 5468
rect 19675 5412 19679 5468
rect 19615 5408 19679 5412
rect 26965 5468 27029 5472
rect 26965 5412 26969 5468
rect 26969 5412 27025 5468
rect 27025 5412 27029 5468
rect 26965 5408 27029 5412
rect 27045 5468 27109 5472
rect 27045 5412 27049 5468
rect 27049 5412 27105 5468
rect 27105 5412 27109 5468
rect 27045 5408 27109 5412
rect 27125 5468 27189 5472
rect 27125 5412 27129 5468
rect 27129 5412 27185 5468
rect 27185 5412 27189 5468
rect 27125 5408 27189 5412
rect 27205 5468 27269 5472
rect 27205 5412 27209 5468
rect 27209 5412 27265 5468
rect 27265 5412 27269 5468
rect 27205 5408 27269 5412
rect 7990 4924 8054 4928
rect 7990 4868 7994 4924
rect 7994 4868 8050 4924
rect 8050 4868 8054 4924
rect 7990 4864 8054 4868
rect 8070 4924 8134 4928
rect 8070 4868 8074 4924
rect 8074 4868 8130 4924
rect 8130 4868 8134 4924
rect 8070 4864 8134 4868
rect 8150 4924 8214 4928
rect 8150 4868 8154 4924
rect 8154 4868 8210 4924
rect 8210 4868 8214 4924
rect 8150 4864 8214 4868
rect 8230 4924 8294 4928
rect 8230 4868 8234 4924
rect 8234 4868 8290 4924
rect 8290 4868 8294 4924
rect 8230 4864 8294 4868
rect 15580 4924 15644 4928
rect 15580 4868 15584 4924
rect 15584 4868 15640 4924
rect 15640 4868 15644 4924
rect 15580 4864 15644 4868
rect 15660 4924 15724 4928
rect 15660 4868 15664 4924
rect 15664 4868 15720 4924
rect 15720 4868 15724 4924
rect 15660 4864 15724 4868
rect 15740 4924 15804 4928
rect 15740 4868 15744 4924
rect 15744 4868 15800 4924
rect 15800 4868 15804 4924
rect 15740 4864 15804 4868
rect 15820 4924 15884 4928
rect 15820 4868 15824 4924
rect 15824 4868 15880 4924
rect 15880 4868 15884 4924
rect 15820 4864 15884 4868
rect 23170 4924 23234 4928
rect 23170 4868 23174 4924
rect 23174 4868 23230 4924
rect 23230 4868 23234 4924
rect 23170 4864 23234 4868
rect 23250 4924 23314 4928
rect 23250 4868 23254 4924
rect 23254 4868 23310 4924
rect 23310 4868 23314 4924
rect 23250 4864 23314 4868
rect 23330 4924 23394 4928
rect 23330 4868 23334 4924
rect 23334 4868 23390 4924
rect 23390 4868 23394 4924
rect 23330 4864 23394 4868
rect 23410 4924 23474 4928
rect 23410 4868 23414 4924
rect 23414 4868 23470 4924
rect 23470 4868 23474 4924
rect 23410 4864 23474 4868
rect 30760 4924 30824 4928
rect 30760 4868 30764 4924
rect 30764 4868 30820 4924
rect 30820 4868 30824 4924
rect 30760 4864 30824 4868
rect 30840 4924 30904 4928
rect 30840 4868 30844 4924
rect 30844 4868 30900 4924
rect 30900 4868 30904 4924
rect 30840 4864 30904 4868
rect 30920 4924 30984 4928
rect 30920 4868 30924 4924
rect 30924 4868 30980 4924
rect 30980 4868 30984 4924
rect 30920 4864 30984 4868
rect 31000 4924 31064 4928
rect 31000 4868 31004 4924
rect 31004 4868 31060 4924
rect 31060 4868 31064 4924
rect 31000 4864 31064 4868
rect 16620 4660 16684 4724
rect 16804 4524 16868 4588
rect 4195 4380 4259 4384
rect 4195 4324 4199 4380
rect 4199 4324 4255 4380
rect 4255 4324 4259 4380
rect 4195 4320 4259 4324
rect 4275 4380 4339 4384
rect 4275 4324 4279 4380
rect 4279 4324 4335 4380
rect 4335 4324 4339 4380
rect 4275 4320 4339 4324
rect 4355 4380 4419 4384
rect 4355 4324 4359 4380
rect 4359 4324 4415 4380
rect 4415 4324 4419 4380
rect 4355 4320 4419 4324
rect 4435 4380 4499 4384
rect 4435 4324 4439 4380
rect 4439 4324 4495 4380
rect 4495 4324 4499 4380
rect 4435 4320 4499 4324
rect 11785 4380 11849 4384
rect 11785 4324 11789 4380
rect 11789 4324 11845 4380
rect 11845 4324 11849 4380
rect 11785 4320 11849 4324
rect 11865 4380 11929 4384
rect 11865 4324 11869 4380
rect 11869 4324 11925 4380
rect 11925 4324 11929 4380
rect 11865 4320 11929 4324
rect 11945 4380 12009 4384
rect 11945 4324 11949 4380
rect 11949 4324 12005 4380
rect 12005 4324 12009 4380
rect 11945 4320 12009 4324
rect 12025 4380 12089 4384
rect 12025 4324 12029 4380
rect 12029 4324 12085 4380
rect 12085 4324 12089 4380
rect 12025 4320 12089 4324
rect 19375 4380 19439 4384
rect 19375 4324 19379 4380
rect 19379 4324 19435 4380
rect 19435 4324 19439 4380
rect 19375 4320 19439 4324
rect 19455 4380 19519 4384
rect 19455 4324 19459 4380
rect 19459 4324 19515 4380
rect 19515 4324 19519 4380
rect 19455 4320 19519 4324
rect 19535 4380 19599 4384
rect 19535 4324 19539 4380
rect 19539 4324 19595 4380
rect 19595 4324 19599 4380
rect 19535 4320 19599 4324
rect 19615 4380 19679 4384
rect 19615 4324 19619 4380
rect 19619 4324 19675 4380
rect 19675 4324 19679 4380
rect 19615 4320 19679 4324
rect 26965 4380 27029 4384
rect 26965 4324 26969 4380
rect 26969 4324 27025 4380
rect 27025 4324 27029 4380
rect 26965 4320 27029 4324
rect 27045 4380 27109 4384
rect 27045 4324 27049 4380
rect 27049 4324 27105 4380
rect 27105 4324 27109 4380
rect 27045 4320 27109 4324
rect 27125 4380 27189 4384
rect 27125 4324 27129 4380
rect 27129 4324 27185 4380
rect 27185 4324 27189 4380
rect 27125 4320 27189 4324
rect 27205 4380 27269 4384
rect 27205 4324 27209 4380
rect 27209 4324 27265 4380
rect 27265 4324 27269 4380
rect 27205 4320 27269 4324
rect 2820 4040 2884 4044
rect 17908 4116 17972 4180
rect 2820 3984 2834 4040
rect 2834 3984 2884 4040
rect 2820 3980 2884 3984
rect 7236 3844 7300 3908
rect 7990 3836 8054 3840
rect 7990 3780 7994 3836
rect 7994 3780 8050 3836
rect 8050 3780 8054 3836
rect 7990 3776 8054 3780
rect 8070 3836 8134 3840
rect 8070 3780 8074 3836
rect 8074 3780 8130 3836
rect 8130 3780 8134 3836
rect 8070 3776 8134 3780
rect 8150 3836 8214 3840
rect 8150 3780 8154 3836
rect 8154 3780 8210 3836
rect 8210 3780 8214 3836
rect 8150 3776 8214 3780
rect 8230 3836 8294 3840
rect 8230 3780 8234 3836
rect 8234 3780 8290 3836
rect 8290 3780 8294 3836
rect 8230 3776 8294 3780
rect 15580 3836 15644 3840
rect 15580 3780 15584 3836
rect 15584 3780 15640 3836
rect 15640 3780 15644 3836
rect 15580 3776 15644 3780
rect 15660 3836 15724 3840
rect 15660 3780 15664 3836
rect 15664 3780 15720 3836
rect 15720 3780 15724 3836
rect 15660 3776 15724 3780
rect 15740 3836 15804 3840
rect 15740 3780 15744 3836
rect 15744 3780 15800 3836
rect 15800 3780 15804 3836
rect 15740 3776 15804 3780
rect 15820 3836 15884 3840
rect 15820 3780 15824 3836
rect 15824 3780 15880 3836
rect 15880 3780 15884 3836
rect 15820 3776 15884 3780
rect 24716 3980 24780 4044
rect 23170 3836 23234 3840
rect 23170 3780 23174 3836
rect 23174 3780 23230 3836
rect 23230 3780 23234 3836
rect 23170 3776 23234 3780
rect 23250 3836 23314 3840
rect 23250 3780 23254 3836
rect 23254 3780 23310 3836
rect 23310 3780 23314 3836
rect 23250 3776 23314 3780
rect 23330 3836 23394 3840
rect 23330 3780 23334 3836
rect 23334 3780 23390 3836
rect 23390 3780 23394 3836
rect 23330 3776 23394 3780
rect 23410 3836 23474 3840
rect 23410 3780 23414 3836
rect 23414 3780 23470 3836
rect 23470 3780 23474 3836
rect 23410 3776 23474 3780
rect 30760 3836 30824 3840
rect 30760 3780 30764 3836
rect 30764 3780 30820 3836
rect 30820 3780 30824 3836
rect 30760 3776 30824 3780
rect 30840 3836 30904 3840
rect 30840 3780 30844 3836
rect 30844 3780 30900 3836
rect 30900 3780 30904 3836
rect 30840 3776 30904 3780
rect 30920 3836 30984 3840
rect 30920 3780 30924 3836
rect 30924 3780 30980 3836
rect 30980 3780 30984 3836
rect 30920 3776 30984 3780
rect 31000 3836 31064 3840
rect 31000 3780 31004 3836
rect 31004 3780 31060 3836
rect 31060 3780 31064 3836
rect 31000 3776 31064 3780
rect 4195 3292 4259 3296
rect 4195 3236 4199 3292
rect 4199 3236 4255 3292
rect 4255 3236 4259 3292
rect 4195 3232 4259 3236
rect 4275 3292 4339 3296
rect 4275 3236 4279 3292
rect 4279 3236 4335 3292
rect 4335 3236 4339 3292
rect 4275 3232 4339 3236
rect 4355 3292 4419 3296
rect 4355 3236 4359 3292
rect 4359 3236 4415 3292
rect 4415 3236 4419 3292
rect 4355 3232 4419 3236
rect 4435 3292 4499 3296
rect 4435 3236 4439 3292
rect 4439 3236 4495 3292
rect 4495 3236 4499 3292
rect 4435 3232 4499 3236
rect 11785 3292 11849 3296
rect 11785 3236 11789 3292
rect 11789 3236 11845 3292
rect 11845 3236 11849 3292
rect 11785 3232 11849 3236
rect 11865 3292 11929 3296
rect 11865 3236 11869 3292
rect 11869 3236 11925 3292
rect 11925 3236 11929 3292
rect 11865 3232 11929 3236
rect 11945 3292 12009 3296
rect 11945 3236 11949 3292
rect 11949 3236 12005 3292
rect 12005 3236 12009 3292
rect 11945 3232 12009 3236
rect 12025 3292 12089 3296
rect 12025 3236 12029 3292
rect 12029 3236 12085 3292
rect 12085 3236 12089 3292
rect 12025 3232 12089 3236
rect 8524 3028 8588 3092
rect 19375 3292 19439 3296
rect 19375 3236 19379 3292
rect 19379 3236 19435 3292
rect 19435 3236 19439 3292
rect 19375 3232 19439 3236
rect 19455 3292 19519 3296
rect 19455 3236 19459 3292
rect 19459 3236 19515 3292
rect 19515 3236 19519 3292
rect 19455 3232 19519 3236
rect 19535 3292 19599 3296
rect 19535 3236 19539 3292
rect 19539 3236 19595 3292
rect 19595 3236 19599 3292
rect 19535 3232 19599 3236
rect 19615 3292 19679 3296
rect 19615 3236 19619 3292
rect 19619 3236 19675 3292
rect 19675 3236 19679 3292
rect 19615 3232 19679 3236
rect 26965 3292 27029 3296
rect 26965 3236 26969 3292
rect 26969 3236 27025 3292
rect 27025 3236 27029 3292
rect 26965 3232 27029 3236
rect 27045 3292 27109 3296
rect 27045 3236 27049 3292
rect 27049 3236 27105 3292
rect 27105 3236 27109 3292
rect 27045 3232 27109 3236
rect 27125 3292 27189 3296
rect 27125 3236 27129 3292
rect 27129 3236 27185 3292
rect 27185 3236 27189 3292
rect 27125 3232 27189 3236
rect 27205 3292 27269 3296
rect 27205 3236 27209 3292
rect 27209 3236 27265 3292
rect 27265 3236 27269 3292
rect 27205 3232 27269 3236
rect 7990 2748 8054 2752
rect 7990 2692 7994 2748
rect 7994 2692 8050 2748
rect 8050 2692 8054 2748
rect 7990 2688 8054 2692
rect 8070 2748 8134 2752
rect 8070 2692 8074 2748
rect 8074 2692 8130 2748
rect 8130 2692 8134 2748
rect 8070 2688 8134 2692
rect 8150 2748 8214 2752
rect 8150 2692 8154 2748
rect 8154 2692 8210 2748
rect 8210 2692 8214 2748
rect 8150 2688 8214 2692
rect 8230 2748 8294 2752
rect 8230 2692 8234 2748
rect 8234 2692 8290 2748
rect 8290 2692 8294 2748
rect 8230 2688 8294 2692
rect 15580 2748 15644 2752
rect 15580 2692 15584 2748
rect 15584 2692 15640 2748
rect 15640 2692 15644 2748
rect 15580 2688 15644 2692
rect 15660 2748 15724 2752
rect 15660 2692 15664 2748
rect 15664 2692 15720 2748
rect 15720 2692 15724 2748
rect 15660 2688 15724 2692
rect 15740 2748 15804 2752
rect 15740 2692 15744 2748
rect 15744 2692 15800 2748
rect 15800 2692 15804 2748
rect 15740 2688 15804 2692
rect 15820 2748 15884 2752
rect 15820 2692 15824 2748
rect 15824 2692 15880 2748
rect 15880 2692 15884 2748
rect 15820 2688 15884 2692
rect 23170 2748 23234 2752
rect 23170 2692 23174 2748
rect 23174 2692 23230 2748
rect 23230 2692 23234 2748
rect 23170 2688 23234 2692
rect 23250 2748 23314 2752
rect 23250 2692 23254 2748
rect 23254 2692 23310 2748
rect 23310 2692 23314 2748
rect 23250 2688 23314 2692
rect 23330 2748 23394 2752
rect 23330 2692 23334 2748
rect 23334 2692 23390 2748
rect 23390 2692 23394 2748
rect 23330 2688 23394 2692
rect 23410 2748 23474 2752
rect 23410 2692 23414 2748
rect 23414 2692 23470 2748
rect 23470 2692 23474 2748
rect 23410 2688 23474 2692
rect 30760 2748 30824 2752
rect 30760 2692 30764 2748
rect 30764 2692 30820 2748
rect 30820 2692 30824 2748
rect 30760 2688 30824 2692
rect 30840 2748 30904 2752
rect 30840 2692 30844 2748
rect 30844 2692 30900 2748
rect 30900 2692 30904 2748
rect 30840 2688 30904 2692
rect 30920 2748 30984 2752
rect 30920 2692 30924 2748
rect 30924 2692 30980 2748
rect 30980 2692 30984 2748
rect 30920 2688 30984 2692
rect 31000 2748 31064 2752
rect 31000 2692 31004 2748
rect 31004 2692 31060 2748
rect 31060 2692 31064 2748
rect 31000 2688 31064 2692
rect 5028 2484 5092 2548
rect 3924 2408 3988 2412
rect 3924 2352 3974 2408
rect 3974 2352 3988 2408
rect 3924 2348 3988 2352
rect 4195 2204 4259 2208
rect 4195 2148 4199 2204
rect 4199 2148 4255 2204
rect 4255 2148 4259 2204
rect 4195 2144 4259 2148
rect 4275 2204 4339 2208
rect 4275 2148 4279 2204
rect 4279 2148 4335 2204
rect 4335 2148 4339 2204
rect 4275 2144 4339 2148
rect 4355 2204 4419 2208
rect 4355 2148 4359 2204
rect 4359 2148 4415 2204
rect 4415 2148 4419 2204
rect 4355 2144 4419 2148
rect 4435 2204 4499 2208
rect 4435 2148 4439 2204
rect 4439 2148 4495 2204
rect 4495 2148 4499 2204
rect 4435 2144 4499 2148
rect 11785 2204 11849 2208
rect 11785 2148 11789 2204
rect 11789 2148 11845 2204
rect 11845 2148 11849 2204
rect 11785 2144 11849 2148
rect 11865 2204 11929 2208
rect 11865 2148 11869 2204
rect 11869 2148 11925 2204
rect 11925 2148 11929 2204
rect 11865 2144 11929 2148
rect 11945 2204 12009 2208
rect 11945 2148 11949 2204
rect 11949 2148 12005 2204
rect 12005 2148 12009 2204
rect 11945 2144 12009 2148
rect 12025 2204 12089 2208
rect 12025 2148 12029 2204
rect 12029 2148 12085 2204
rect 12085 2148 12089 2204
rect 12025 2144 12089 2148
rect 19375 2204 19439 2208
rect 19375 2148 19379 2204
rect 19379 2148 19435 2204
rect 19435 2148 19439 2204
rect 19375 2144 19439 2148
rect 19455 2204 19519 2208
rect 19455 2148 19459 2204
rect 19459 2148 19515 2204
rect 19515 2148 19519 2204
rect 19455 2144 19519 2148
rect 19535 2204 19599 2208
rect 19535 2148 19539 2204
rect 19539 2148 19595 2204
rect 19595 2148 19599 2204
rect 19535 2144 19599 2148
rect 19615 2204 19679 2208
rect 19615 2148 19619 2204
rect 19619 2148 19675 2204
rect 19675 2148 19679 2204
rect 19615 2144 19679 2148
rect 26965 2204 27029 2208
rect 26965 2148 26969 2204
rect 26969 2148 27025 2204
rect 27025 2148 27029 2204
rect 26965 2144 27029 2148
rect 27045 2204 27109 2208
rect 27045 2148 27049 2204
rect 27049 2148 27105 2204
rect 27105 2148 27109 2204
rect 27045 2144 27109 2148
rect 27125 2204 27189 2208
rect 27125 2148 27129 2204
rect 27129 2148 27185 2204
rect 27185 2148 27189 2204
rect 27125 2144 27189 2148
rect 27205 2204 27269 2208
rect 27205 2148 27209 2204
rect 27209 2148 27265 2204
rect 27265 2148 27269 2204
rect 27205 2144 27269 2148
rect 7990 1660 8054 1664
rect 7990 1604 7994 1660
rect 7994 1604 8050 1660
rect 8050 1604 8054 1660
rect 7990 1600 8054 1604
rect 8070 1660 8134 1664
rect 8070 1604 8074 1660
rect 8074 1604 8130 1660
rect 8130 1604 8134 1660
rect 8070 1600 8134 1604
rect 8150 1660 8214 1664
rect 8150 1604 8154 1660
rect 8154 1604 8210 1660
rect 8210 1604 8214 1660
rect 8150 1600 8214 1604
rect 8230 1660 8294 1664
rect 8230 1604 8234 1660
rect 8234 1604 8290 1660
rect 8290 1604 8294 1660
rect 8230 1600 8294 1604
rect 15580 1660 15644 1664
rect 15580 1604 15584 1660
rect 15584 1604 15640 1660
rect 15640 1604 15644 1660
rect 15580 1600 15644 1604
rect 15660 1660 15724 1664
rect 15660 1604 15664 1660
rect 15664 1604 15720 1660
rect 15720 1604 15724 1660
rect 15660 1600 15724 1604
rect 15740 1660 15804 1664
rect 15740 1604 15744 1660
rect 15744 1604 15800 1660
rect 15800 1604 15804 1660
rect 15740 1600 15804 1604
rect 15820 1660 15884 1664
rect 15820 1604 15824 1660
rect 15824 1604 15880 1660
rect 15880 1604 15884 1660
rect 15820 1600 15884 1604
rect 23170 1660 23234 1664
rect 23170 1604 23174 1660
rect 23174 1604 23230 1660
rect 23230 1604 23234 1660
rect 23170 1600 23234 1604
rect 23250 1660 23314 1664
rect 23250 1604 23254 1660
rect 23254 1604 23310 1660
rect 23310 1604 23314 1660
rect 23250 1600 23314 1604
rect 23330 1660 23394 1664
rect 23330 1604 23334 1660
rect 23334 1604 23390 1660
rect 23390 1604 23394 1660
rect 23330 1600 23394 1604
rect 23410 1660 23474 1664
rect 23410 1604 23414 1660
rect 23414 1604 23470 1660
rect 23470 1604 23474 1660
rect 23410 1600 23474 1604
rect 30760 1660 30824 1664
rect 30760 1604 30764 1660
rect 30764 1604 30820 1660
rect 30820 1604 30824 1660
rect 30760 1600 30824 1604
rect 30840 1660 30904 1664
rect 30840 1604 30844 1660
rect 30844 1604 30900 1660
rect 30900 1604 30904 1660
rect 30840 1600 30904 1604
rect 30920 1660 30984 1664
rect 30920 1604 30924 1660
rect 30924 1604 30980 1660
rect 30980 1604 30984 1660
rect 30920 1600 30984 1604
rect 31000 1660 31064 1664
rect 31000 1604 31004 1660
rect 31004 1604 31060 1660
rect 31060 1604 31064 1660
rect 31000 1600 31064 1604
rect 4195 1116 4259 1120
rect 4195 1060 4199 1116
rect 4199 1060 4255 1116
rect 4255 1060 4259 1116
rect 4195 1056 4259 1060
rect 4275 1116 4339 1120
rect 4275 1060 4279 1116
rect 4279 1060 4335 1116
rect 4335 1060 4339 1116
rect 4275 1056 4339 1060
rect 4355 1116 4419 1120
rect 4355 1060 4359 1116
rect 4359 1060 4415 1116
rect 4415 1060 4419 1116
rect 4355 1056 4419 1060
rect 4435 1116 4499 1120
rect 4435 1060 4439 1116
rect 4439 1060 4495 1116
rect 4495 1060 4499 1116
rect 4435 1056 4499 1060
rect 11785 1116 11849 1120
rect 11785 1060 11789 1116
rect 11789 1060 11845 1116
rect 11845 1060 11849 1116
rect 11785 1056 11849 1060
rect 11865 1116 11929 1120
rect 11865 1060 11869 1116
rect 11869 1060 11925 1116
rect 11925 1060 11929 1116
rect 11865 1056 11929 1060
rect 11945 1116 12009 1120
rect 11945 1060 11949 1116
rect 11949 1060 12005 1116
rect 12005 1060 12009 1116
rect 11945 1056 12009 1060
rect 12025 1116 12089 1120
rect 12025 1060 12029 1116
rect 12029 1060 12085 1116
rect 12085 1060 12089 1116
rect 12025 1056 12089 1060
rect 19375 1116 19439 1120
rect 19375 1060 19379 1116
rect 19379 1060 19435 1116
rect 19435 1060 19439 1116
rect 19375 1056 19439 1060
rect 19455 1116 19519 1120
rect 19455 1060 19459 1116
rect 19459 1060 19515 1116
rect 19515 1060 19519 1116
rect 19455 1056 19519 1060
rect 19535 1116 19599 1120
rect 19535 1060 19539 1116
rect 19539 1060 19595 1116
rect 19595 1060 19599 1116
rect 19535 1056 19599 1060
rect 19615 1116 19679 1120
rect 19615 1060 19619 1116
rect 19619 1060 19675 1116
rect 19675 1060 19679 1116
rect 19615 1056 19679 1060
rect 26965 1116 27029 1120
rect 26965 1060 26969 1116
rect 26969 1060 27025 1116
rect 27025 1060 27029 1116
rect 26965 1056 27029 1060
rect 27045 1116 27109 1120
rect 27045 1060 27049 1116
rect 27049 1060 27105 1116
rect 27105 1060 27109 1116
rect 27045 1056 27109 1060
rect 27125 1116 27189 1120
rect 27125 1060 27129 1116
rect 27129 1060 27185 1116
rect 27185 1060 27189 1116
rect 27125 1056 27189 1060
rect 27205 1116 27269 1120
rect 27205 1060 27209 1116
rect 27209 1060 27265 1116
rect 27265 1060 27269 1116
rect 27205 1056 27269 1060
rect 7990 572 8054 576
rect 7990 516 7994 572
rect 7994 516 8050 572
rect 8050 516 8054 572
rect 7990 512 8054 516
rect 8070 572 8134 576
rect 8070 516 8074 572
rect 8074 516 8130 572
rect 8130 516 8134 572
rect 8070 512 8134 516
rect 8150 572 8214 576
rect 8150 516 8154 572
rect 8154 516 8210 572
rect 8210 516 8214 572
rect 8150 512 8214 516
rect 8230 572 8294 576
rect 8230 516 8234 572
rect 8234 516 8290 572
rect 8290 516 8294 572
rect 8230 512 8294 516
rect 15580 572 15644 576
rect 15580 516 15584 572
rect 15584 516 15640 572
rect 15640 516 15644 572
rect 15580 512 15644 516
rect 15660 572 15724 576
rect 15660 516 15664 572
rect 15664 516 15720 572
rect 15720 516 15724 572
rect 15660 512 15724 516
rect 15740 572 15804 576
rect 15740 516 15744 572
rect 15744 516 15800 572
rect 15800 516 15804 572
rect 15740 512 15804 516
rect 15820 572 15884 576
rect 15820 516 15824 572
rect 15824 516 15880 572
rect 15880 516 15884 572
rect 15820 512 15884 516
rect 23170 572 23234 576
rect 23170 516 23174 572
rect 23174 516 23230 572
rect 23230 516 23234 572
rect 23170 512 23234 516
rect 23250 572 23314 576
rect 23250 516 23254 572
rect 23254 516 23310 572
rect 23310 516 23314 572
rect 23250 512 23314 516
rect 23330 572 23394 576
rect 23330 516 23334 572
rect 23334 516 23390 572
rect 23390 516 23394 572
rect 23330 512 23394 516
rect 23410 572 23474 576
rect 23410 516 23414 572
rect 23414 516 23470 572
rect 23470 516 23474 572
rect 23410 512 23474 516
rect 30760 572 30824 576
rect 30760 516 30764 572
rect 30764 516 30820 572
rect 30820 516 30824 572
rect 30760 512 30824 516
rect 30840 572 30904 576
rect 30840 516 30844 572
rect 30844 516 30900 572
rect 30900 516 30904 572
rect 30840 512 30904 516
rect 30920 572 30984 576
rect 30920 516 30924 572
rect 30924 516 30980 572
rect 30980 516 30984 572
rect 30920 512 30984 516
rect 31000 572 31064 576
rect 31000 516 31004 572
rect 31004 516 31060 572
rect 31060 516 31064 572
rect 31000 512 31064 516
<< metal4 >>
rect 4294 22130 4354 22304
rect 4478 22174 4722 22234
rect 4478 22130 4538 22174
rect 4294 22070 4538 22130
rect 4187 21792 4507 21808
rect 4187 21728 4195 21792
rect 4259 21728 4275 21792
rect 4339 21728 4355 21792
rect 4419 21728 4435 21792
rect 4499 21728 4507 21792
rect 3923 20772 3989 20773
rect 3923 20708 3924 20772
rect 3988 20708 3989 20772
rect 3923 20707 3989 20708
rect 2819 12476 2885 12477
rect 2819 12412 2820 12476
rect 2884 12412 2885 12476
rect 2819 12411 2885 12412
rect 2822 4045 2882 12411
rect 3003 10980 3069 10981
rect 3003 10916 3004 10980
rect 3068 10916 3069 10980
rect 3003 10915 3069 10916
rect 3006 5541 3066 10915
rect 3003 5540 3069 5541
rect 3003 5476 3004 5540
rect 3068 5476 3069 5540
rect 3003 5475 3069 5476
rect 2819 4044 2885 4045
rect 2819 3980 2820 4044
rect 2884 3980 2885 4044
rect 2819 3979 2885 3980
rect 3926 2413 3986 20707
rect 4187 20704 4507 21728
rect 4187 20640 4195 20704
rect 4259 20640 4275 20704
rect 4339 20640 4355 20704
rect 4419 20640 4435 20704
rect 4499 20640 4507 20704
rect 4187 19616 4507 20640
rect 4187 19552 4195 19616
rect 4259 19552 4275 19616
rect 4339 19552 4355 19616
rect 4419 19552 4435 19616
rect 4499 19552 4507 19616
rect 4187 18528 4507 19552
rect 4187 18464 4195 18528
rect 4259 18464 4275 18528
rect 4339 18464 4355 18528
rect 4419 18464 4435 18528
rect 4499 18464 4507 18528
rect 4187 17440 4507 18464
rect 4662 18461 4722 22174
rect 4846 22130 4906 22304
rect 5030 22174 5274 22234
rect 5030 22130 5090 22174
rect 4846 22070 5090 22130
rect 5214 18461 5274 22174
rect 5398 18733 5458 22304
rect 5395 18732 5461 18733
rect 5395 18668 5396 18732
rect 5460 18668 5461 18732
rect 5395 18667 5461 18668
rect 4659 18460 4725 18461
rect 4659 18396 4660 18460
rect 4724 18396 4725 18460
rect 4659 18395 4725 18396
rect 5211 18460 5277 18461
rect 5211 18396 5212 18460
rect 5276 18396 5277 18460
rect 5211 18395 5277 18396
rect 5395 18052 5461 18053
rect 5395 17988 5396 18052
rect 5460 17988 5461 18052
rect 5395 17987 5461 17988
rect 4187 17376 4195 17440
rect 4259 17376 4275 17440
rect 4339 17376 4355 17440
rect 4419 17376 4435 17440
rect 4499 17376 4507 17440
rect 4187 16352 4507 17376
rect 4187 16288 4195 16352
rect 4259 16288 4275 16352
rect 4339 16288 4355 16352
rect 4419 16288 4435 16352
rect 4499 16288 4507 16352
rect 4187 15264 4507 16288
rect 4187 15200 4195 15264
rect 4259 15200 4275 15264
rect 4339 15200 4355 15264
rect 4419 15200 4435 15264
rect 4499 15200 4507 15264
rect 4187 14176 4507 15200
rect 4187 14112 4195 14176
rect 4259 14112 4275 14176
rect 4339 14112 4355 14176
rect 4419 14112 4435 14176
rect 4499 14112 4507 14176
rect 4187 13088 4507 14112
rect 5398 13973 5458 17987
rect 5950 17373 6010 22304
rect 6502 18189 6562 22304
rect 7054 18325 7114 22304
rect 7606 20637 7666 22304
rect 7790 22174 8034 22234
rect 7603 20636 7669 20637
rect 7603 20572 7604 20636
rect 7668 20572 7669 20636
rect 7603 20571 7669 20572
rect 7051 18324 7117 18325
rect 7051 18260 7052 18324
rect 7116 18260 7117 18324
rect 7051 18259 7117 18260
rect 6499 18188 6565 18189
rect 6499 18124 6500 18188
rect 6564 18124 6565 18188
rect 6499 18123 6565 18124
rect 6683 18052 6749 18053
rect 6683 17988 6684 18052
rect 6748 17988 6749 18052
rect 6683 17987 6749 17988
rect 5947 17372 6013 17373
rect 5947 17308 5948 17372
rect 6012 17308 6013 17372
rect 5947 17307 6013 17308
rect 5947 16692 6013 16693
rect 5947 16628 5948 16692
rect 6012 16628 6013 16692
rect 5947 16627 6013 16628
rect 5395 13972 5461 13973
rect 5395 13908 5396 13972
rect 5460 13908 5461 13972
rect 5395 13907 5461 13908
rect 4187 13024 4195 13088
rect 4259 13024 4275 13088
rect 4339 13024 4355 13088
rect 4419 13024 4435 13088
rect 4499 13024 4507 13088
rect 4187 12000 4507 13024
rect 4187 11936 4195 12000
rect 4259 11936 4275 12000
rect 4339 11936 4355 12000
rect 4419 11936 4435 12000
rect 4499 11936 4507 12000
rect 4187 10912 4507 11936
rect 4187 10848 4195 10912
rect 4259 10848 4275 10912
rect 4339 10848 4355 10912
rect 4419 10848 4435 10912
rect 4499 10848 4507 10912
rect 4187 9824 4507 10848
rect 4187 9760 4195 9824
rect 4259 9760 4275 9824
rect 4339 9760 4355 9824
rect 4419 9760 4435 9824
rect 4499 9760 4507 9824
rect 4187 8736 4507 9760
rect 5027 9484 5093 9485
rect 5027 9420 5028 9484
rect 5092 9420 5093 9484
rect 5027 9419 5093 9420
rect 4187 8672 4195 8736
rect 4259 8672 4275 8736
rect 4339 8672 4355 8736
rect 4419 8672 4435 8736
rect 4499 8672 4507 8736
rect 4187 7648 4507 8672
rect 4187 7584 4195 7648
rect 4259 7584 4275 7648
rect 4339 7584 4355 7648
rect 4419 7584 4435 7648
rect 4499 7584 4507 7648
rect 4187 6560 4507 7584
rect 4187 6496 4195 6560
rect 4259 6496 4275 6560
rect 4339 6496 4355 6560
rect 4419 6496 4435 6560
rect 4499 6496 4507 6560
rect 4187 5472 4507 6496
rect 4187 5408 4195 5472
rect 4259 5408 4275 5472
rect 4339 5408 4355 5472
rect 4419 5408 4435 5472
rect 4499 5408 4507 5472
rect 4187 4384 4507 5408
rect 4187 4320 4195 4384
rect 4259 4320 4275 4384
rect 4339 4320 4355 4384
rect 4419 4320 4435 4384
rect 4499 4320 4507 4384
rect 4187 3296 4507 4320
rect 4187 3232 4195 3296
rect 4259 3232 4275 3296
rect 4339 3232 4355 3296
rect 4419 3232 4435 3296
rect 4499 3232 4507 3296
rect 3923 2412 3989 2413
rect 3923 2348 3924 2412
rect 3988 2348 3989 2412
rect 3923 2347 3989 2348
rect 4187 2208 4507 3232
rect 5030 2549 5090 9419
rect 5950 8261 6010 16627
rect 6315 12748 6381 12749
rect 6315 12684 6316 12748
rect 6380 12684 6381 12748
rect 6315 12683 6381 12684
rect 6131 9756 6197 9757
rect 6131 9692 6132 9756
rect 6196 9692 6197 9756
rect 6131 9691 6197 9692
rect 5947 8260 6013 8261
rect 5947 8196 5948 8260
rect 6012 8196 6013 8260
rect 5947 8195 6013 8196
rect 6134 7037 6194 9691
rect 6318 9621 6378 12683
rect 6686 11661 6746 17987
rect 7790 12749 7850 22174
rect 7974 22130 8034 22174
rect 8158 22130 8218 22304
rect 7974 22070 8218 22130
rect 7982 21248 8302 21808
rect 7982 21184 7990 21248
rect 8054 21184 8070 21248
rect 8134 21184 8150 21248
rect 8214 21184 8230 21248
rect 8294 21184 8302 21248
rect 7982 20160 8302 21184
rect 7982 20096 7990 20160
rect 8054 20096 8070 20160
rect 8134 20096 8150 20160
rect 8214 20096 8230 20160
rect 8294 20096 8302 20160
rect 7982 19072 8302 20096
rect 8710 19141 8770 22304
rect 8891 20772 8957 20773
rect 8891 20708 8892 20772
rect 8956 20708 8957 20772
rect 8891 20707 8957 20708
rect 8707 19140 8773 19141
rect 8707 19076 8708 19140
rect 8772 19076 8773 19140
rect 8707 19075 8773 19076
rect 7982 19008 7990 19072
rect 8054 19008 8070 19072
rect 8134 19008 8150 19072
rect 8214 19008 8230 19072
rect 8294 19008 8302 19072
rect 7982 17984 8302 19008
rect 8707 18732 8773 18733
rect 8707 18668 8708 18732
rect 8772 18668 8773 18732
rect 8707 18667 8773 18668
rect 7982 17920 7990 17984
rect 8054 17920 8070 17984
rect 8134 17920 8150 17984
rect 8214 17920 8230 17984
rect 8294 17920 8302 17984
rect 7982 16896 8302 17920
rect 7982 16832 7990 16896
rect 8054 16832 8070 16896
rect 8134 16832 8150 16896
rect 8214 16832 8230 16896
rect 8294 16832 8302 16896
rect 7982 15808 8302 16832
rect 8523 16828 8589 16829
rect 8523 16764 8524 16828
rect 8588 16764 8589 16828
rect 8523 16763 8589 16764
rect 7982 15744 7990 15808
rect 8054 15744 8070 15808
rect 8134 15744 8150 15808
rect 8214 15744 8230 15808
rect 8294 15744 8302 15808
rect 7982 14720 8302 15744
rect 8526 15197 8586 16763
rect 8523 15196 8589 15197
rect 8523 15132 8524 15196
rect 8588 15132 8589 15196
rect 8523 15131 8589 15132
rect 7982 14656 7990 14720
rect 8054 14656 8070 14720
rect 8134 14656 8150 14720
rect 8214 14656 8230 14720
rect 8294 14656 8302 14720
rect 7982 13632 8302 14656
rect 7982 13568 7990 13632
rect 8054 13568 8070 13632
rect 8134 13568 8150 13632
rect 8214 13568 8230 13632
rect 8294 13568 8302 13632
rect 7787 12748 7853 12749
rect 7787 12684 7788 12748
rect 7852 12684 7853 12748
rect 7787 12683 7853 12684
rect 7982 12544 8302 13568
rect 7982 12480 7990 12544
rect 8054 12480 8070 12544
rect 8134 12480 8150 12544
rect 8214 12480 8230 12544
rect 8294 12480 8302 12544
rect 6683 11660 6749 11661
rect 6683 11596 6684 11660
rect 6748 11596 6749 11660
rect 6683 11595 6749 11596
rect 7982 11456 8302 12480
rect 7982 11392 7990 11456
rect 8054 11392 8070 11456
rect 8134 11392 8150 11456
rect 8214 11392 8230 11456
rect 8294 11392 8302 11456
rect 7051 11116 7117 11117
rect 7051 11052 7052 11116
rect 7116 11052 7117 11116
rect 7051 11051 7117 11052
rect 6683 10708 6749 10709
rect 6683 10644 6684 10708
rect 6748 10644 6749 10708
rect 6683 10643 6749 10644
rect 6315 9620 6381 9621
rect 6315 9556 6316 9620
rect 6380 9556 6381 9620
rect 6315 9555 6381 9556
rect 6131 7036 6197 7037
rect 6131 6972 6132 7036
rect 6196 6972 6197 7036
rect 6131 6971 6197 6972
rect 6686 6765 6746 10643
rect 6867 9756 6933 9757
rect 6867 9692 6868 9756
rect 6932 9692 6933 9756
rect 6867 9691 6933 9692
rect 6870 7445 6930 9691
rect 7054 8261 7114 11051
rect 7982 10368 8302 11392
rect 8710 11389 8770 18667
rect 8894 13701 8954 20707
rect 9262 18869 9322 22304
rect 9814 19141 9874 22304
rect 10366 22130 10426 22304
rect 10731 22268 10797 22269
rect 10731 22234 10732 22268
rect 10550 22204 10732 22234
rect 10796 22204 10797 22268
rect 10550 22203 10797 22204
rect 10550 22174 10794 22203
rect 10550 22130 10610 22174
rect 10366 22070 10610 22130
rect 10179 20772 10245 20773
rect 10179 20708 10180 20772
rect 10244 20708 10245 20772
rect 10179 20707 10245 20708
rect 9811 19140 9877 19141
rect 9811 19076 9812 19140
rect 9876 19076 9877 19140
rect 9811 19075 9877 19076
rect 9259 18868 9325 18869
rect 9259 18804 9260 18868
rect 9324 18804 9325 18868
rect 9259 18803 9325 18804
rect 8891 13700 8957 13701
rect 8891 13636 8892 13700
rect 8956 13636 8957 13700
rect 8891 13635 8957 13636
rect 8707 11388 8773 11389
rect 8707 11324 8708 11388
rect 8772 11324 8773 11388
rect 8707 11323 8773 11324
rect 7982 10304 7990 10368
rect 8054 10304 8070 10368
rect 8134 10304 8150 10368
rect 8214 10304 8230 10368
rect 8294 10304 8302 10368
rect 7235 9620 7301 9621
rect 7235 9556 7236 9620
rect 7300 9556 7301 9620
rect 7235 9555 7301 9556
rect 7051 8260 7117 8261
rect 7051 8196 7052 8260
rect 7116 8196 7117 8260
rect 7051 8195 7117 8196
rect 6867 7444 6933 7445
rect 6867 7380 6868 7444
rect 6932 7380 6933 7444
rect 6867 7379 6933 7380
rect 6683 6764 6749 6765
rect 6683 6700 6684 6764
rect 6748 6700 6749 6764
rect 6683 6699 6749 6700
rect 7238 3909 7298 9555
rect 7982 9280 8302 10304
rect 7982 9216 7990 9280
rect 8054 9216 8070 9280
rect 8134 9216 8150 9280
rect 8214 9216 8230 9280
rect 8294 9216 8302 9280
rect 7982 8192 8302 9216
rect 10182 8261 10242 20707
rect 10918 19277 10978 22304
rect 11283 21044 11349 21045
rect 11283 20980 11284 21044
rect 11348 20980 11349 21044
rect 11283 20979 11349 20980
rect 10915 19276 10981 19277
rect 10915 19212 10916 19276
rect 10980 19212 10981 19276
rect 10915 19211 10981 19212
rect 10547 18460 10613 18461
rect 10547 18396 10548 18460
rect 10612 18396 10613 18460
rect 10547 18395 10613 18396
rect 10550 13021 10610 18395
rect 10547 13020 10613 13021
rect 10547 12956 10548 13020
rect 10612 12956 10613 13020
rect 10547 12955 10613 12956
rect 11286 11797 11346 20979
rect 11470 20909 11530 22304
rect 12022 22130 12082 22304
rect 12022 22070 12266 22130
rect 12206 21861 12266 22070
rect 12203 21860 12269 21861
rect 11777 21792 12097 21808
rect 12203 21796 12204 21860
rect 12268 21796 12269 21860
rect 12203 21795 12269 21796
rect 11777 21728 11785 21792
rect 11849 21728 11865 21792
rect 11929 21728 11945 21792
rect 12009 21728 12025 21792
rect 12089 21728 12097 21792
rect 11467 20908 11533 20909
rect 11467 20844 11468 20908
rect 11532 20844 11533 20908
rect 11467 20843 11533 20844
rect 11777 20704 12097 21728
rect 11777 20640 11785 20704
rect 11849 20640 11865 20704
rect 11929 20640 11945 20704
rect 12009 20640 12025 20704
rect 12089 20640 12097 20704
rect 11777 19616 12097 20640
rect 11777 19552 11785 19616
rect 11849 19552 11865 19616
rect 11929 19552 11945 19616
rect 12009 19552 12025 19616
rect 12089 19552 12097 19616
rect 11467 19412 11533 19413
rect 11467 19348 11468 19412
rect 11532 19348 11533 19412
rect 11467 19347 11533 19348
rect 11470 12069 11530 19347
rect 11777 18528 12097 19552
rect 12574 19277 12634 22304
rect 13126 22130 13186 22304
rect 13310 22174 13554 22234
rect 13310 22130 13370 22174
rect 13126 22070 13370 22130
rect 13494 21450 13554 22174
rect 13678 21589 13738 22304
rect 13675 21588 13741 21589
rect 13675 21524 13676 21588
rect 13740 21524 13741 21588
rect 13675 21523 13741 21524
rect 13675 21452 13741 21453
rect 13675 21450 13676 21452
rect 13494 21390 13676 21450
rect 13675 21388 13676 21390
rect 13740 21388 13741 21452
rect 13675 21387 13741 21388
rect 12571 19276 12637 19277
rect 12571 19212 12572 19276
rect 12636 19212 12637 19276
rect 12571 19211 12637 19212
rect 11777 18464 11785 18528
rect 11849 18464 11865 18528
rect 11929 18464 11945 18528
rect 12009 18464 12025 18528
rect 12089 18464 12097 18528
rect 11777 17440 12097 18464
rect 11777 17376 11785 17440
rect 11849 17376 11865 17440
rect 11929 17376 11945 17440
rect 12009 17376 12025 17440
rect 12089 17376 12097 17440
rect 11777 16352 12097 17376
rect 14230 16421 14290 22304
rect 14782 19277 14842 22304
rect 15334 20770 15394 22304
rect 15886 22130 15946 22304
rect 15886 22070 16130 22130
rect 15150 20710 15394 20770
rect 15572 21248 15892 21808
rect 15572 21184 15580 21248
rect 15644 21184 15660 21248
rect 15724 21184 15740 21248
rect 15804 21184 15820 21248
rect 15884 21184 15892 21248
rect 15150 20637 15210 20710
rect 15147 20636 15213 20637
rect 15147 20572 15148 20636
rect 15212 20572 15213 20636
rect 15147 20571 15213 20572
rect 15572 20160 15892 21184
rect 15572 20096 15580 20160
rect 15644 20096 15660 20160
rect 15724 20096 15740 20160
rect 15804 20096 15820 20160
rect 15884 20096 15892 20160
rect 14779 19276 14845 19277
rect 14779 19212 14780 19276
rect 14844 19212 14845 19276
rect 14779 19211 14845 19212
rect 15572 19072 15892 20096
rect 16070 19277 16130 22070
rect 16438 19277 16498 22304
rect 16990 21589 17050 22304
rect 17542 22104 17602 22304
rect 18094 22104 18154 22304
rect 18646 22104 18706 22304
rect 19198 22104 19258 22304
rect 19750 22104 19810 22304
rect 20302 22104 20362 22304
rect 20854 22104 20914 22304
rect 21406 22104 21466 22304
rect 19367 21792 19687 21808
rect 19367 21728 19375 21792
rect 19439 21728 19455 21792
rect 19519 21728 19535 21792
rect 19599 21728 19615 21792
rect 19679 21728 19687 21792
rect 16987 21588 17053 21589
rect 16987 21524 16988 21588
rect 17052 21524 17053 21588
rect 16987 21523 17053 21524
rect 19367 20704 19687 21728
rect 19367 20640 19375 20704
rect 19439 20640 19455 20704
rect 19519 20640 19535 20704
rect 19599 20640 19615 20704
rect 19679 20640 19687 20704
rect 19367 19616 19687 20640
rect 21958 19957 22018 22304
rect 21955 19956 22021 19957
rect 21955 19892 21956 19956
rect 22020 19892 22021 19956
rect 21955 19891 22021 19892
rect 19367 19552 19375 19616
rect 19439 19552 19455 19616
rect 19519 19552 19535 19616
rect 19599 19552 19615 19616
rect 19679 19552 19687 19616
rect 16067 19276 16133 19277
rect 16067 19212 16068 19276
rect 16132 19212 16133 19276
rect 16067 19211 16133 19212
rect 16435 19276 16501 19277
rect 16435 19212 16436 19276
rect 16500 19212 16501 19276
rect 16435 19211 16501 19212
rect 15572 19008 15580 19072
rect 15644 19008 15660 19072
rect 15724 19008 15740 19072
rect 15804 19008 15820 19072
rect 15884 19008 15892 19072
rect 15572 17984 15892 19008
rect 15572 17920 15580 17984
rect 15644 17920 15660 17984
rect 15724 17920 15740 17984
rect 15804 17920 15820 17984
rect 15884 17920 15892 17984
rect 15572 16896 15892 17920
rect 15572 16832 15580 16896
rect 15644 16832 15660 16896
rect 15724 16832 15740 16896
rect 15804 16832 15820 16896
rect 15884 16832 15892 16896
rect 14227 16420 14293 16421
rect 14227 16356 14228 16420
rect 14292 16356 14293 16420
rect 14227 16355 14293 16356
rect 11777 16288 11785 16352
rect 11849 16288 11865 16352
rect 11929 16288 11945 16352
rect 12009 16288 12025 16352
rect 12089 16288 12097 16352
rect 11777 15264 12097 16288
rect 15572 15808 15892 16832
rect 15572 15744 15580 15808
rect 15644 15744 15660 15808
rect 15724 15744 15740 15808
rect 15804 15744 15820 15808
rect 15884 15744 15892 15808
rect 12571 15740 12637 15741
rect 12571 15676 12572 15740
rect 12636 15676 12637 15740
rect 12571 15675 12637 15676
rect 11777 15200 11785 15264
rect 11849 15200 11865 15264
rect 11929 15200 11945 15264
rect 12009 15200 12025 15264
rect 12089 15200 12097 15264
rect 11777 14176 12097 15200
rect 11777 14112 11785 14176
rect 11849 14112 11865 14176
rect 11929 14112 11945 14176
rect 12009 14112 12025 14176
rect 12089 14112 12097 14176
rect 11777 13088 12097 14112
rect 11777 13024 11785 13088
rect 11849 13024 11865 13088
rect 11929 13024 11945 13088
rect 12009 13024 12025 13088
rect 12089 13024 12097 13088
rect 11467 12068 11533 12069
rect 11467 12004 11468 12068
rect 11532 12004 11533 12068
rect 11467 12003 11533 12004
rect 11777 12000 12097 13024
rect 12574 12205 12634 15675
rect 15572 14720 15892 15744
rect 15572 14656 15580 14720
rect 15644 14656 15660 14720
rect 15724 14656 15740 14720
rect 15804 14656 15820 14720
rect 15884 14656 15892 14720
rect 15572 13632 15892 14656
rect 15572 13568 15580 13632
rect 15644 13568 15660 13632
rect 15724 13568 15740 13632
rect 15804 13568 15820 13632
rect 15884 13568 15892 13632
rect 15572 12544 15892 13568
rect 15572 12480 15580 12544
rect 15644 12480 15660 12544
rect 15724 12480 15740 12544
rect 15804 12480 15820 12544
rect 15884 12480 15892 12544
rect 12571 12204 12637 12205
rect 12571 12140 12572 12204
rect 12636 12140 12637 12204
rect 12571 12139 12637 12140
rect 11777 11936 11785 12000
rect 11849 11936 11865 12000
rect 11929 11936 11945 12000
rect 12009 11936 12025 12000
rect 12089 11936 12097 12000
rect 11283 11796 11349 11797
rect 11283 11732 11284 11796
rect 11348 11732 11349 11796
rect 11283 11731 11349 11732
rect 11777 10912 12097 11936
rect 11777 10848 11785 10912
rect 11849 10848 11865 10912
rect 11929 10848 11945 10912
rect 12009 10848 12025 10912
rect 12089 10848 12097 10912
rect 11777 9824 12097 10848
rect 11777 9760 11785 9824
rect 11849 9760 11865 9824
rect 11929 9760 11945 9824
rect 12009 9760 12025 9824
rect 12089 9760 12097 9824
rect 11777 8736 12097 9760
rect 11777 8672 11785 8736
rect 11849 8672 11865 8736
rect 11929 8672 11945 8736
rect 12009 8672 12025 8736
rect 12089 8672 12097 8736
rect 10179 8260 10245 8261
rect 10179 8196 10180 8260
rect 10244 8196 10245 8260
rect 10179 8195 10245 8196
rect 7982 8128 7990 8192
rect 8054 8128 8070 8192
rect 8134 8128 8150 8192
rect 8214 8128 8230 8192
rect 8294 8128 8302 8192
rect 7982 7104 8302 8128
rect 7982 7040 7990 7104
rect 8054 7040 8070 7104
rect 8134 7040 8150 7104
rect 8214 7040 8230 7104
rect 8294 7040 8302 7104
rect 7982 6016 8302 7040
rect 7982 5952 7990 6016
rect 8054 5952 8070 6016
rect 8134 5952 8150 6016
rect 8214 5952 8230 6016
rect 8294 5952 8302 6016
rect 7982 4928 8302 5952
rect 11777 7648 12097 8672
rect 11777 7584 11785 7648
rect 11849 7584 11865 7648
rect 11929 7584 11945 7648
rect 12009 7584 12025 7648
rect 12089 7584 12097 7648
rect 11777 6560 12097 7584
rect 11777 6496 11785 6560
rect 11849 6496 11865 6560
rect 11929 6496 11945 6560
rect 12009 6496 12025 6560
rect 12089 6496 12097 6560
rect 8523 5540 8589 5541
rect 8523 5476 8524 5540
rect 8588 5476 8589 5540
rect 8523 5475 8589 5476
rect 7982 4864 7990 4928
rect 8054 4864 8070 4928
rect 8134 4864 8150 4928
rect 8214 4864 8230 4928
rect 8294 4864 8302 4928
rect 7235 3908 7301 3909
rect 7235 3844 7236 3908
rect 7300 3844 7301 3908
rect 7235 3843 7301 3844
rect 7982 3840 8302 4864
rect 7982 3776 7990 3840
rect 8054 3776 8070 3840
rect 8134 3776 8150 3840
rect 8214 3776 8230 3840
rect 8294 3776 8302 3840
rect 7982 2752 8302 3776
rect 8526 3093 8586 5475
rect 11777 5472 12097 6496
rect 11777 5408 11785 5472
rect 11849 5408 11865 5472
rect 11929 5408 11945 5472
rect 12009 5408 12025 5472
rect 12089 5408 12097 5472
rect 11777 4384 12097 5408
rect 11777 4320 11785 4384
rect 11849 4320 11865 4384
rect 11929 4320 11945 4384
rect 12009 4320 12025 4384
rect 12089 4320 12097 4384
rect 11777 3296 12097 4320
rect 11777 3232 11785 3296
rect 11849 3232 11865 3296
rect 11929 3232 11945 3296
rect 12009 3232 12025 3296
rect 12089 3232 12097 3296
rect 8523 3092 8589 3093
rect 8523 3028 8524 3092
rect 8588 3028 8589 3092
rect 8523 3027 8589 3028
rect 7982 2688 7990 2752
rect 8054 2688 8070 2752
rect 8134 2688 8150 2752
rect 8214 2688 8230 2752
rect 8294 2688 8302 2752
rect 5027 2548 5093 2549
rect 5027 2484 5028 2548
rect 5092 2484 5093 2548
rect 5027 2483 5093 2484
rect 4187 2144 4195 2208
rect 4259 2144 4275 2208
rect 4339 2144 4355 2208
rect 4419 2144 4435 2208
rect 4499 2144 4507 2208
rect 4187 1120 4507 2144
rect 4187 1056 4195 1120
rect 4259 1056 4275 1120
rect 4339 1056 4355 1120
rect 4419 1056 4435 1120
rect 4499 1056 4507 1120
rect 4187 496 4507 1056
rect 7982 1664 8302 2688
rect 7982 1600 7990 1664
rect 8054 1600 8070 1664
rect 8134 1600 8150 1664
rect 8214 1600 8230 1664
rect 8294 1600 8302 1664
rect 7982 576 8302 1600
rect 7982 512 7990 576
rect 8054 512 8070 576
rect 8134 512 8150 576
rect 8214 512 8230 576
rect 8294 512 8302 576
rect 7982 496 8302 512
rect 11777 2208 12097 3232
rect 11777 2144 11785 2208
rect 11849 2144 11865 2208
rect 11929 2144 11945 2208
rect 12009 2144 12025 2208
rect 12089 2144 12097 2208
rect 11777 1120 12097 2144
rect 11777 1056 11785 1120
rect 11849 1056 11865 1120
rect 11929 1056 11945 1120
rect 12009 1056 12025 1120
rect 12089 1056 12097 1120
rect 11777 496 12097 1056
rect 15572 11456 15892 12480
rect 15572 11392 15580 11456
rect 15644 11392 15660 11456
rect 15724 11392 15740 11456
rect 15804 11392 15820 11456
rect 15884 11392 15892 11456
rect 15572 10368 15892 11392
rect 15572 10304 15580 10368
rect 15644 10304 15660 10368
rect 15724 10304 15740 10368
rect 15804 10304 15820 10368
rect 15884 10304 15892 10368
rect 15572 9280 15892 10304
rect 19367 18528 19687 19552
rect 19367 18464 19375 18528
rect 19439 18464 19455 18528
rect 19519 18464 19535 18528
rect 19599 18464 19615 18528
rect 19679 18464 19687 18528
rect 19367 17440 19687 18464
rect 22510 18053 22570 22304
rect 23062 22130 23122 22304
rect 22878 22070 23122 22130
rect 22878 18053 22938 22070
rect 23162 21248 23482 21808
rect 23162 21184 23170 21248
rect 23234 21184 23250 21248
rect 23314 21184 23330 21248
rect 23394 21184 23410 21248
rect 23474 21184 23482 21248
rect 23162 20160 23482 21184
rect 23614 20637 23674 22304
rect 23611 20636 23677 20637
rect 23611 20572 23612 20636
rect 23676 20572 23677 20636
rect 23611 20571 23677 20572
rect 23162 20096 23170 20160
rect 23234 20096 23250 20160
rect 23314 20096 23330 20160
rect 23394 20096 23410 20160
rect 23474 20096 23482 20160
rect 23162 19072 23482 20096
rect 23162 19008 23170 19072
rect 23234 19008 23250 19072
rect 23314 19008 23330 19072
rect 23394 19008 23410 19072
rect 23474 19008 23482 19072
rect 22507 18052 22573 18053
rect 22507 17988 22508 18052
rect 22572 17988 22573 18052
rect 22507 17987 22573 17988
rect 22875 18052 22941 18053
rect 22875 17988 22876 18052
rect 22940 17988 22941 18052
rect 22875 17987 22941 17988
rect 19367 17376 19375 17440
rect 19439 17376 19455 17440
rect 19519 17376 19535 17440
rect 19599 17376 19615 17440
rect 19679 17376 19687 17440
rect 19367 16352 19687 17376
rect 19367 16288 19375 16352
rect 19439 16288 19455 16352
rect 19519 16288 19535 16352
rect 19599 16288 19615 16352
rect 19679 16288 19687 16352
rect 19367 15264 19687 16288
rect 19367 15200 19375 15264
rect 19439 15200 19455 15264
rect 19519 15200 19535 15264
rect 19599 15200 19615 15264
rect 19679 15200 19687 15264
rect 19367 14176 19687 15200
rect 19367 14112 19375 14176
rect 19439 14112 19455 14176
rect 19519 14112 19535 14176
rect 19599 14112 19615 14176
rect 19679 14112 19687 14176
rect 19367 13088 19687 14112
rect 19367 13024 19375 13088
rect 19439 13024 19455 13088
rect 19519 13024 19535 13088
rect 19599 13024 19615 13088
rect 19679 13024 19687 13088
rect 19367 12000 19687 13024
rect 19367 11936 19375 12000
rect 19439 11936 19455 12000
rect 19519 11936 19535 12000
rect 19599 11936 19615 12000
rect 19679 11936 19687 12000
rect 19367 10912 19687 11936
rect 19367 10848 19375 10912
rect 19439 10848 19455 10912
rect 19519 10848 19535 10912
rect 19599 10848 19615 10912
rect 19679 10848 19687 10912
rect 17907 10300 17973 10301
rect 17907 10236 17908 10300
rect 17972 10236 17973 10300
rect 17907 10235 17973 10236
rect 15572 9216 15580 9280
rect 15644 9216 15660 9280
rect 15724 9216 15740 9280
rect 15804 9216 15820 9280
rect 15884 9216 15892 9280
rect 15572 8192 15892 9216
rect 15572 8128 15580 8192
rect 15644 8128 15660 8192
rect 15724 8128 15740 8192
rect 15804 8128 15820 8192
rect 15884 8128 15892 8192
rect 15572 7104 15892 8128
rect 16803 7172 16869 7173
rect 16803 7108 16804 7172
rect 16868 7108 16869 7172
rect 16803 7107 16869 7108
rect 15572 7040 15580 7104
rect 15644 7040 15660 7104
rect 15724 7040 15740 7104
rect 15804 7040 15820 7104
rect 15884 7040 15892 7104
rect 15572 6016 15892 7040
rect 16619 7036 16685 7037
rect 16619 6972 16620 7036
rect 16684 6972 16685 7036
rect 16619 6971 16685 6972
rect 15572 5952 15580 6016
rect 15644 5952 15660 6016
rect 15724 5952 15740 6016
rect 15804 5952 15820 6016
rect 15884 5952 15892 6016
rect 15572 4928 15892 5952
rect 15572 4864 15580 4928
rect 15644 4864 15660 4928
rect 15724 4864 15740 4928
rect 15804 4864 15820 4928
rect 15884 4864 15892 4928
rect 15572 3840 15892 4864
rect 16622 4725 16682 6971
rect 16619 4724 16685 4725
rect 16619 4660 16620 4724
rect 16684 4660 16685 4724
rect 16619 4659 16685 4660
rect 16806 4589 16866 7107
rect 16803 4588 16869 4589
rect 16803 4524 16804 4588
rect 16868 4524 16869 4588
rect 16803 4523 16869 4524
rect 17910 4181 17970 10235
rect 19367 9824 19687 10848
rect 19367 9760 19375 9824
rect 19439 9760 19455 9824
rect 19519 9760 19535 9824
rect 19599 9760 19615 9824
rect 19679 9760 19687 9824
rect 19367 8736 19687 9760
rect 19367 8672 19375 8736
rect 19439 8672 19455 8736
rect 19519 8672 19535 8736
rect 19599 8672 19615 8736
rect 19679 8672 19687 8736
rect 19367 7648 19687 8672
rect 19367 7584 19375 7648
rect 19439 7584 19455 7648
rect 19519 7584 19535 7648
rect 19599 7584 19615 7648
rect 19679 7584 19687 7648
rect 19367 6560 19687 7584
rect 19367 6496 19375 6560
rect 19439 6496 19455 6560
rect 19519 6496 19535 6560
rect 19599 6496 19615 6560
rect 19679 6496 19687 6560
rect 19367 5472 19687 6496
rect 19367 5408 19375 5472
rect 19439 5408 19455 5472
rect 19519 5408 19535 5472
rect 19599 5408 19615 5472
rect 19679 5408 19687 5472
rect 19367 4384 19687 5408
rect 19367 4320 19375 4384
rect 19439 4320 19455 4384
rect 19519 4320 19535 4384
rect 19599 4320 19615 4384
rect 19679 4320 19687 4384
rect 17907 4180 17973 4181
rect 17907 4116 17908 4180
rect 17972 4116 17973 4180
rect 17907 4115 17973 4116
rect 15572 3776 15580 3840
rect 15644 3776 15660 3840
rect 15724 3776 15740 3840
rect 15804 3776 15820 3840
rect 15884 3776 15892 3840
rect 15572 2752 15892 3776
rect 15572 2688 15580 2752
rect 15644 2688 15660 2752
rect 15724 2688 15740 2752
rect 15804 2688 15820 2752
rect 15884 2688 15892 2752
rect 15572 1664 15892 2688
rect 15572 1600 15580 1664
rect 15644 1600 15660 1664
rect 15724 1600 15740 1664
rect 15804 1600 15820 1664
rect 15884 1600 15892 1664
rect 15572 576 15892 1600
rect 15572 512 15580 576
rect 15644 512 15660 576
rect 15724 512 15740 576
rect 15804 512 15820 576
rect 15884 512 15892 576
rect 15572 496 15892 512
rect 19367 3296 19687 4320
rect 19367 3232 19375 3296
rect 19439 3232 19455 3296
rect 19519 3232 19535 3296
rect 19599 3232 19615 3296
rect 19679 3232 19687 3296
rect 19367 2208 19687 3232
rect 19367 2144 19375 2208
rect 19439 2144 19455 2208
rect 19519 2144 19535 2208
rect 19599 2144 19615 2208
rect 19679 2144 19687 2208
rect 19367 1120 19687 2144
rect 19367 1056 19375 1120
rect 19439 1056 19455 1120
rect 19519 1056 19535 1120
rect 19599 1056 19615 1120
rect 19679 1056 19687 1120
rect 19367 496 19687 1056
rect 23162 17984 23482 19008
rect 23979 18868 24045 18869
rect 23979 18804 23980 18868
rect 24044 18804 24045 18868
rect 23979 18803 24045 18804
rect 23162 17920 23170 17984
rect 23234 17920 23250 17984
rect 23314 17920 23330 17984
rect 23394 17920 23410 17984
rect 23474 17920 23482 17984
rect 23162 16896 23482 17920
rect 23162 16832 23170 16896
rect 23234 16832 23250 16896
rect 23314 16832 23330 16896
rect 23394 16832 23410 16896
rect 23474 16832 23482 16896
rect 23162 15808 23482 16832
rect 23162 15744 23170 15808
rect 23234 15744 23250 15808
rect 23314 15744 23330 15808
rect 23394 15744 23410 15808
rect 23474 15744 23482 15808
rect 23162 14720 23482 15744
rect 23162 14656 23170 14720
rect 23234 14656 23250 14720
rect 23314 14656 23330 14720
rect 23394 14656 23410 14720
rect 23474 14656 23482 14720
rect 23162 13632 23482 14656
rect 23162 13568 23170 13632
rect 23234 13568 23250 13632
rect 23314 13568 23330 13632
rect 23394 13568 23410 13632
rect 23474 13568 23482 13632
rect 23162 12544 23482 13568
rect 23982 13565 24042 18803
rect 24166 18189 24226 22304
rect 24718 19277 24778 22304
rect 24902 22174 25146 22234
rect 24902 21045 24962 22174
rect 25086 22130 25146 22174
rect 25270 22130 25330 22304
rect 25086 22070 25330 22130
rect 25454 22174 25698 22234
rect 25454 21589 25514 22174
rect 25638 22130 25698 22174
rect 25822 22130 25882 22304
rect 25638 22070 25882 22130
rect 25451 21588 25517 21589
rect 25451 21524 25452 21588
rect 25516 21524 25517 21588
rect 25451 21523 25517 21524
rect 26374 21181 26434 22304
rect 26926 22104 26986 22304
rect 27478 22104 27538 22304
rect 26957 21792 27277 21808
rect 26957 21728 26965 21792
rect 27029 21728 27045 21792
rect 27109 21728 27125 21792
rect 27189 21728 27205 21792
rect 27269 21728 27277 21792
rect 26371 21180 26437 21181
rect 26371 21116 26372 21180
rect 26436 21116 26437 21180
rect 26371 21115 26437 21116
rect 24899 21044 24965 21045
rect 24899 20980 24900 21044
rect 24964 20980 24965 21044
rect 24899 20979 24965 20980
rect 26957 20704 27277 21728
rect 28763 21452 28829 21453
rect 28763 21388 28764 21452
rect 28828 21388 28829 21452
rect 28763 21387 28829 21388
rect 26957 20640 26965 20704
rect 27029 20640 27045 20704
rect 27109 20640 27125 20704
rect 27189 20640 27205 20704
rect 27269 20640 27277 20704
rect 26957 19616 27277 20640
rect 27659 20500 27725 20501
rect 27659 20436 27660 20500
rect 27724 20436 27725 20500
rect 27659 20435 27725 20436
rect 26957 19552 26965 19616
rect 27029 19552 27045 19616
rect 27109 19552 27125 19616
rect 27189 19552 27205 19616
rect 27269 19552 27277 19616
rect 26555 19412 26621 19413
rect 26555 19348 26556 19412
rect 26620 19348 26621 19412
rect 26555 19347 26621 19348
rect 24715 19276 24781 19277
rect 24715 19212 24716 19276
rect 24780 19212 24781 19276
rect 24715 19211 24781 19212
rect 24163 18188 24229 18189
rect 24163 18124 24164 18188
rect 24228 18124 24229 18188
rect 24163 18123 24229 18124
rect 26558 15197 26618 19347
rect 26957 18528 27277 19552
rect 26957 18464 26965 18528
rect 27029 18464 27045 18528
rect 27109 18464 27125 18528
rect 27189 18464 27205 18528
rect 27269 18464 27277 18528
rect 26957 17440 27277 18464
rect 26957 17376 26965 17440
rect 27029 17376 27045 17440
rect 27109 17376 27125 17440
rect 27189 17376 27205 17440
rect 27269 17376 27277 17440
rect 26957 16352 27277 17376
rect 26957 16288 26965 16352
rect 27029 16288 27045 16352
rect 27109 16288 27125 16352
rect 27189 16288 27205 16352
rect 27269 16288 27277 16352
rect 26957 15264 27277 16288
rect 26957 15200 26965 15264
rect 27029 15200 27045 15264
rect 27109 15200 27125 15264
rect 27189 15200 27205 15264
rect 27269 15200 27277 15264
rect 26555 15196 26621 15197
rect 26555 15132 26556 15196
rect 26620 15132 26621 15196
rect 26555 15131 26621 15132
rect 26957 14176 27277 15200
rect 26957 14112 26965 14176
rect 27029 14112 27045 14176
rect 27109 14112 27125 14176
rect 27189 14112 27205 14176
rect 27269 14112 27277 14176
rect 23979 13564 24045 13565
rect 23979 13500 23980 13564
rect 24044 13500 24045 13564
rect 23979 13499 24045 13500
rect 23162 12480 23170 12544
rect 23234 12480 23250 12544
rect 23314 12480 23330 12544
rect 23394 12480 23410 12544
rect 23474 12480 23482 12544
rect 23162 11456 23482 12480
rect 23162 11392 23170 11456
rect 23234 11392 23250 11456
rect 23314 11392 23330 11456
rect 23394 11392 23410 11456
rect 23474 11392 23482 11456
rect 23162 10368 23482 11392
rect 23162 10304 23170 10368
rect 23234 10304 23250 10368
rect 23314 10304 23330 10368
rect 23394 10304 23410 10368
rect 23474 10304 23482 10368
rect 23162 9280 23482 10304
rect 23162 9216 23170 9280
rect 23234 9216 23250 9280
rect 23314 9216 23330 9280
rect 23394 9216 23410 9280
rect 23474 9216 23482 9280
rect 23162 8192 23482 9216
rect 26957 13088 27277 14112
rect 26957 13024 26965 13088
rect 27029 13024 27045 13088
rect 27109 13024 27125 13088
rect 27189 13024 27205 13088
rect 27269 13024 27277 13088
rect 26957 12000 27277 13024
rect 27662 12477 27722 20435
rect 27659 12476 27725 12477
rect 27659 12412 27660 12476
rect 27724 12412 27725 12476
rect 27659 12411 27725 12412
rect 28766 12341 28826 21387
rect 30752 21248 31072 21808
rect 30752 21184 30760 21248
rect 30824 21184 30840 21248
rect 30904 21184 30920 21248
rect 30984 21184 31000 21248
rect 31064 21184 31072 21248
rect 30752 20160 31072 21184
rect 30752 20096 30760 20160
rect 30824 20096 30840 20160
rect 30904 20096 30920 20160
rect 30984 20096 31000 20160
rect 31064 20096 31072 20160
rect 30752 19072 31072 20096
rect 30752 19008 30760 19072
rect 30824 19008 30840 19072
rect 30904 19008 30920 19072
rect 30984 19008 31000 19072
rect 31064 19008 31072 19072
rect 30752 17984 31072 19008
rect 30752 17920 30760 17984
rect 30824 17920 30840 17984
rect 30904 17920 30920 17984
rect 30984 17920 31000 17984
rect 31064 17920 31072 17984
rect 29499 17100 29565 17101
rect 29499 17036 29500 17100
rect 29564 17036 29565 17100
rect 29499 17035 29565 17036
rect 29315 16828 29381 16829
rect 29315 16764 29316 16828
rect 29380 16764 29381 16828
rect 29315 16763 29381 16764
rect 29131 16556 29197 16557
rect 29131 16492 29132 16556
rect 29196 16492 29197 16556
rect 29131 16491 29197 16492
rect 29134 13021 29194 16491
rect 29318 15741 29378 16763
rect 29502 16149 29562 17035
rect 30752 16896 31072 17920
rect 30752 16832 30760 16896
rect 30824 16832 30840 16896
rect 30904 16832 30920 16896
rect 30984 16832 31000 16896
rect 31064 16832 31072 16896
rect 29683 16420 29749 16421
rect 29683 16356 29684 16420
rect 29748 16356 29749 16420
rect 29683 16355 29749 16356
rect 29499 16148 29565 16149
rect 29499 16084 29500 16148
rect 29564 16084 29565 16148
rect 29499 16083 29565 16084
rect 29315 15740 29381 15741
rect 29315 15676 29316 15740
rect 29380 15676 29381 15740
rect 29315 15675 29381 15676
rect 29686 13701 29746 16355
rect 30752 15808 31072 16832
rect 30752 15744 30760 15808
rect 30824 15744 30840 15808
rect 30904 15744 30920 15808
rect 30984 15744 31000 15808
rect 31064 15744 31072 15808
rect 30752 14720 31072 15744
rect 30752 14656 30760 14720
rect 30824 14656 30840 14720
rect 30904 14656 30920 14720
rect 30984 14656 31000 14720
rect 31064 14656 31072 14720
rect 29683 13700 29749 13701
rect 29683 13636 29684 13700
rect 29748 13636 29749 13700
rect 29683 13635 29749 13636
rect 30752 13632 31072 14656
rect 30752 13568 30760 13632
rect 30824 13568 30840 13632
rect 30904 13568 30920 13632
rect 30984 13568 31000 13632
rect 31064 13568 31072 13632
rect 29131 13020 29197 13021
rect 29131 12956 29132 13020
rect 29196 12956 29197 13020
rect 29131 12955 29197 12956
rect 30752 12544 31072 13568
rect 30752 12480 30760 12544
rect 30824 12480 30840 12544
rect 30904 12480 30920 12544
rect 30984 12480 31000 12544
rect 31064 12480 31072 12544
rect 28763 12340 28829 12341
rect 28763 12276 28764 12340
rect 28828 12276 28829 12340
rect 28763 12275 28829 12276
rect 26957 11936 26965 12000
rect 27029 11936 27045 12000
rect 27109 11936 27125 12000
rect 27189 11936 27205 12000
rect 27269 11936 27277 12000
rect 26957 10912 27277 11936
rect 26957 10848 26965 10912
rect 27029 10848 27045 10912
rect 27109 10848 27125 10912
rect 27189 10848 27205 10912
rect 27269 10848 27277 10912
rect 26957 9824 27277 10848
rect 26957 9760 26965 9824
rect 27029 9760 27045 9824
rect 27109 9760 27125 9824
rect 27189 9760 27205 9824
rect 27269 9760 27277 9824
rect 24715 8940 24781 8941
rect 24715 8876 24716 8940
rect 24780 8876 24781 8940
rect 24715 8875 24781 8876
rect 23162 8128 23170 8192
rect 23234 8128 23250 8192
rect 23314 8128 23330 8192
rect 23394 8128 23410 8192
rect 23474 8128 23482 8192
rect 23162 7104 23482 8128
rect 23162 7040 23170 7104
rect 23234 7040 23250 7104
rect 23314 7040 23330 7104
rect 23394 7040 23410 7104
rect 23474 7040 23482 7104
rect 23162 6016 23482 7040
rect 23162 5952 23170 6016
rect 23234 5952 23250 6016
rect 23314 5952 23330 6016
rect 23394 5952 23410 6016
rect 23474 5952 23482 6016
rect 23162 4928 23482 5952
rect 23162 4864 23170 4928
rect 23234 4864 23250 4928
rect 23314 4864 23330 4928
rect 23394 4864 23410 4928
rect 23474 4864 23482 4928
rect 23162 3840 23482 4864
rect 24718 4045 24778 8875
rect 26957 8736 27277 9760
rect 26957 8672 26965 8736
rect 27029 8672 27045 8736
rect 27109 8672 27125 8736
rect 27189 8672 27205 8736
rect 27269 8672 27277 8736
rect 26187 7988 26253 7989
rect 26187 7924 26188 7988
rect 26252 7924 26253 7988
rect 26187 7923 26253 7924
rect 26190 5541 26250 7923
rect 26957 7648 27277 8672
rect 26957 7584 26965 7648
rect 27029 7584 27045 7648
rect 27109 7584 27125 7648
rect 27189 7584 27205 7648
rect 27269 7584 27277 7648
rect 26957 6560 27277 7584
rect 26957 6496 26965 6560
rect 27029 6496 27045 6560
rect 27109 6496 27125 6560
rect 27189 6496 27205 6560
rect 27269 6496 27277 6560
rect 26187 5540 26253 5541
rect 26187 5476 26188 5540
rect 26252 5476 26253 5540
rect 26187 5475 26253 5476
rect 26957 5472 27277 6496
rect 26957 5408 26965 5472
rect 27029 5408 27045 5472
rect 27109 5408 27125 5472
rect 27189 5408 27205 5472
rect 27269 5408 27277 5472
rect 26957 4384 27277 5408
rect 26957 4320 26965 4384
rect 27029 4320 27045 4384
rect 27109 4320 27125 4384
rect 27189 4320 27205 4384
rect 27269 4320 27277 4384
rect 24715 4044 24781 4045
rect 24715 3980 24716 4044
rect 24780 3980 24781 4044
rect 24715 3979 24781 3980
rect 23162 3776 23170 3840
rect 23234 3776 23250 3840
rect 23314 3776 23330 3840
rect 23394 3776 23410 3840
rect 23474 3776 23482 3840
rect 23162 2752 23482 3776
rect 23162 2688 23170 2752
rect 23234 2688 23250 2752
rect 23314 2688 23330 2752
rect 23394 2688 23410 2752
rect 23474 2688 23482 2752
rect 23162 1664 23482 2688
rect 23162 1600 23170 1664
rect 23234 1600 23250 1664
rect 23314 1600 23330 1664
rect 23394 1600 23410 1664
rect 23474 1600 23482 1664
rect 23162 576 23482 1600
rect 23162 512 23170 576
rect 23234 512 23250 576
rect 23314 512 23330 576
rect 23394 512 23410 576
rect 23474 512 23482 576
rect 23162 496 23482 512
rect 26957 3296 27277 4320
rect 26957 3232 26965 3296
rect 27029 3232 27045 3296
rect 27109 3232 27125 3296
rect 27189 3232 27205 3296
rect 27269 3232 27277 3296
rect 26957 2208 27277 3232
rect 26957 2144 26965 2208
rect 27029 2144 27045 2208
rect 27109 2144 27125 2208
rect 27189 2144 27205 2208
rect 27269 2144 27277 2208
rect 26957 1120 27277 2144
rect 26957 1056 26965 1120
rect 27029 1056 27045 1120
rect 27109 1056 27125 1120
rect 27189 1056 27205 1120
rect 27269 1056 27277 1120
rect 26957 496 27277 1056
rect 30752 11456 31072 12480
rect 30752 11392 30760 11456
rect 30824 11392 30840 11456
rect 30904 11392 30920 11456
rect 30984 11392 31000 11456
rect 31064 11392 31072 11456
rect 30752 10368 31072 11392
rect 30752 10304 30760 10368
rect 30824 10304 30840 10368
rect 30904 10304 30920 10368
rect 30984 10304 31000 10368
rect 31064 10304 31072 10368
rect 30752 9280 31072 10304
rect 30752 9216 30760 9280
rect 30824 9216 30840 9280
rect 30904 9216 30920 9280
rect 30984 9216 31000 9280
rect 31064 9216 31072 9280
rect 30752 8192 31072 9216
rect 30752 8128 30760 8192
rect 30824 8128 30840 8192
rect 30904 8128 30920 8192
rect 30984 8128 31000 8192
rect 31064 8128 31072 8192
rect 30752 7104 31072 8128
rect 30752 7040 30760 7104
rect 30824 7040 30840 7104
rect 30904 7040 30920 7104
rect 30984 7040 31000 7104
rect 31064 7040 31072 7104
rect 30752 6016 31072 7040
rect 30752 5952 30760 6016
rect 30824 5952 30840 6016
rect 30904 5952 30920 6016
rect 30984 5952 31000 6016
rect 31064 5952 31072 6016
rect 30752 4928 31072 5952
rect 30752 4864 30760 4928
rect 30824 4864 30840 4928
rect 30904 4864 30920 4928
rect 30984 4864 31000 4928
rect 31064 4864 31072 4928
rect 30752 3840 31072 4864
rect 30752 3776 30760 3840
rect 30824 3776 30840 3840
rect 30904 3776 30920 3840
rect 30984 3776 31000 3840
rect 31064 3776 31072 3840
rect 30752 2752 31072 3776
rect 30752 2688 30760 2752
rect 30824 2688 30840 2752
rect 30904 2688 30920 2752
rect 30984 2688 31000 2752
rect 31064 2688 31072 2752
rect 30752 1664 31072 2688
rect 30752 1600 30760 1664
rect 30824 1600 30840 1664
rect 30904 1600 30920 1664
rect 30984 1600 31000 1664
rect 31064 1600 31072 1664
rect 30752 576 31072 1600
rect 30752 512 30760 576
rect 30824 512 30840 576
rect 30904 512 30920 576
rect 30984 512 31000 576
rect 31064 512 31072 576
rect 30752 496 31072 512
use sky130_fd_sc_hd__inv_2  _05_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 30360 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _06_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 21344 0 1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _07_
timestamp 1693170804
transform 1 0 23828 0 1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _08_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 22908 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _09_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 25668 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _10_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 18676 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _11_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 21804 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 13892 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _21_
timestamp 1693170804
transform 1 0 13524 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _22_
timestamp 1693170804
transform 1 0 10672 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _23_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8096 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _24_
timestamp 1693170804
transform 1 0 18676 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _25_
timestamp 1693170804
transform 1 0 5796 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _26_
timestamp 1693170804
transform 1 0 4600 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _27_
timestamp 1693170804
transform 1 0 5152 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1693170804
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1693170804
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1693170804
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1693170804
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1693170804
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1693170804
transform 1 0 21436 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1693170804
transform 1 0 23276 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1693170804
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1693170804
transform 1 0 4692 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1693170804
transform 1 0 5520 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1693170804
transform 1 0 3680 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1693170804
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1693170804
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1693170804
transform 1 0 3404 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1693170804
transform 1 0 4048 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1693170804
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1693170804
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1693170804
transform 1 0 3680 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1693170804
transform 1 0 11776 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1693170804
transform 1 0 3680 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2i_2  ct.cw.cc_test_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28980 0 1 20128
box -38 -48 1050 592
use sky130_ht_sc_tt05__mux2i_2  ct.cw.cc_test_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698685089
transform 1 0 28980 0 1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__maj3_2  ct.cw.cc_test_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28980 0 1 21216
box -38 -48 866 592
use sky130_ht_sc_tt05__maj3_2  ct.cw.cc_test_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698685089
transform 1 0 28980 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dlrtp_1  ct.cw.cc_test_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28980 0 1 19040
box -38 -48 1234 592
use sky130_ht_sc_tt05__dlrtp_1  ct.cw.cc_test_5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698685089
transform 1 0 28980 0 1 17952
box -38 -48 1418 592
use sky130_fd_sc_hd__dfrtp_1  ct.cw.cc_test_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 26588 0 -1 19040
box -38 -48 1878 592
use sky130_ht_sc_tt05__dfrtp_1  ct.cw.cc_test_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698685089
transform 1 0 24564 0 1 19040
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[0\].bits\[0\].cc_flop $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 19412 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[0\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 21988 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[0\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 28704 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[0\].cc_clkbuf
timestamp 1693170804
transform 1 0 29808 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[1\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[1\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 14260 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[1\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[1\].cc_clkbuf
timestamp 1693170804
transform 1 0 24288 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[2\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 16836 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[2\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[2\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 14260 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[2\].cc_clkbuf
timestamp 1693170804
transform 1 0 29992 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[3\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[3\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[3\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 17204 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[3\].cc_clkbuf
timestamp 1693170804
transform 1 0 28152 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[4\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 26404 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[4\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 27048 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[4\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[4\].cc_clkbuf
timestamp 1693170804
transform 1 0 24012 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[5\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 26404 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[5\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 27048 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[5\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 26404 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[5\].cc_clkbuf
timestamp 1693170804
transform 1 0 23552 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[6\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 24380 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[6\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[6\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 26404 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[6\].cc_clkbuf
timestamp 1693170804
transform 1 0 22172 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[7\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 20424 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[7\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 21252 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[7\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[7\].cc_clkbuf
timestamp 1693170804
transform 1 0 21252 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[8\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 18676 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[8\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 18676 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[8\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 16836 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[8\].cc_clkbuf
timestamp 1693170804
transform 1 0 20424 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[9\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 17848 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[9\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 17848 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[9\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 18676 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[9\].cc_clkbuf
timestamp 1693170804
transform 1 0 17848 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[10\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 16100 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[10\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 16100 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[10\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 15916 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[10\].cc_clkbuf
timestamp 1693170804
transform 1 0 13616 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[11\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 16100 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[11\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 14168 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[11\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 14260 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[11\].cc_clkbuf
timestamp 1693170804
transform 1 0 13708 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[0\].cc_scanflop $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 12052 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 11868 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 12972 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 11132 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 5520 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 8464 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8096 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 11500 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 15732 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[0\].cc_clkbuf
timestamp 1693170804
transform 1 0 10304 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[0\].rs_mbuf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 16100 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 10948 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 3404 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 10764 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 8464 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 14076 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 8924 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 5336 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10856 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[1\].cc_clkbuf
timestamp 1693170804
transform 1 0 4784 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[1\].rs_mbuf
timestamp 1693170804
transform 1 0 10948 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 9476 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 9200 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 9752 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3128 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[2\].bits\[4\].rs_cbuf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 11500 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 4232 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[2\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 6440 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[2\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[2\].cc_clkbuf
timestamp 1693170804
transform 1 0 4232 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[2\].rs_mbuf
timestamp 1693170804
transform 1 0 3680 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 13432 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 14076 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 5980 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 12328 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 12328 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 11132 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 16928 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[3\].cc_clkbuf
timestamp 1693170804
transform 1 0 3220 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[3\].rs_mbuf
timestamp 1693170804
transform 1 0 3864 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 4416 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 4692 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[4\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[4\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 11684 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[4\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 16928 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[4\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[4\].cc_clkbuf
timestamp 1693170804
transform 1 0 3220 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[4\].rs_mbuf
timestamp 1693170804
transform 1 0 3220 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 4416 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3772 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 4692 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3772 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 4968 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 15548 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 1196 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[5\].cc_clkbuf
timestamp 1693170804
transform 1 0 3220 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[5\].rs_mbuf
timestamp 1693170804
transform 1 0 3220 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6348 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 6072 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 6348 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 9384 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 8280 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 9936 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[6\].cc_clkbuf
timestamp 1693170804
transform 1 0 5796 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[6\].rs_mbuf
timestamp 1693170804
transform 1 0 8832 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 10304 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 12236 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 11960 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[7\].cc_clkbuf
timestamp 1693170804
transform 1 0 10948 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[7\].rs_mbuf
timestamp 1693170804
transform 1 0 11040 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 14168 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 13616 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 14720 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 14168 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 13892 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 14720 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 15640 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 14444 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 14444 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 15916 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[8\].cc_clkbuf
timestamp 1693170804
transform 1 0 13524 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[8\].rs_mbuf
timestamp 1693170804
transform 1 0 14996 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 18676 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 18952 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 17204 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 18216 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 17112 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 19320 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 17480 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 17204 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 17112 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 17756 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 17112 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 19228 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[9\].cc_clkbuf
timestamp 1693170804
transform 1 0 16100 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[9\].rs_mbuf
timestamp 1693170804
transform 1 0 18676 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 19504 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 19780 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 19596 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 19872 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 20240 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 20608 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 22816 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 20608 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 23368 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[10\].cc_clkbuf
timestamp 1693170804
transform 1 0 18032 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[10\].rs_mbuf
timestamp 1693170804
transform 1 0 20884 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 22448 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 22172 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 22724 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 23000 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 24840 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24840 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[11\].cc_clkbuf
timestamp 1693170804
transform 1 0 22816 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[11\].rs_mbuf
timestamp 1693170804
transform 1 0 24288 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 26036 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 26036 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 28336 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 29900 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 30176 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[12\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[12\].cc_clkbuf
timestamp 1693170804
transform 1 0 25668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[12\].rs_mbuf
timestamp 1693170804
transform 1 0 29808 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 24012 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 23736 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 24012 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 27140 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 28336 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 28428 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 29348 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 30268 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 28428 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 29624 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[13\].cc_clkbuf
timestamp 1693170804
transform 1 0 28980 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[13\].rs_mbuf
timestamp 1693170804
transform 1 0 26588 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 21896 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 23092 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 23368 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 24196 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 28060 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 28612 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 29348 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 27784 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 28060 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 29624 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[14\].cc_clkbuf
timestamp 1693170804
transform 1 0 27416 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[14\].rs_mbuf
timestamp 1693170804
transform 1 0 26036 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 20332 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 20608 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 23000 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 29992 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 27692 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 29716 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 27508 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 27692 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 28428 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[15\].cc_clkbuf
timestamp 1693170804
transform 1 0 25668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[15\].rs_mbuf
timestamp 1693170804
transform 1 0 26404 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 19136 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 19412 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 19688 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 22356 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26312 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 28244 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26220 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 27968 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 23184 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 27692 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[16\].cc_clkbuf
timestamp 1693170804
transform 1 0 26956 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[16\].rs_mbuf
timestamp 1693170804
transform 1 0 19044 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16836 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 16928 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 17940 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 20148 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 20608 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 25944 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 27416 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 20332 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24564 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 25668 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[17\].cc_clkbuf
timestamp 1693170804
transform 1 0 18676 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[17\].rs_mbuf
timestamp 1693170804
transform 1 0 16836 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 17388 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 18124 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 19596 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 17388 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 20148 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 24104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[18\].cc_clkbuf
timestamp 1693170804
transform 1 0 20608 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[18\].rs_mbuf
timestamp 1693170804
transform 1 0 16836 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 17756 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 19688 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 21804 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 22264 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[19\].cc_clkbuf
timestamp 1693170804
transform 1 0 19596 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[19\].rs_mbuf
timestamp 1693170804
transform 1 0 19136 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 27876 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 29900 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 27508 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 28520 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 25668 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 27508 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 26496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 24472 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 25944 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 28152 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 26772 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[20\].cc_clkbuf
timestamp 1693170804
transform 1 0 23092 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[20\].rs_mbuf
timestamp 1693170804
transform 1 0 26036 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 27876 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 28520 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 28428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 18952 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[21\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 27508 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[21\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 27232 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[21\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 16744 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[21\].cc_clkbuf
timestamp 1693170804
transform 1 0 27140 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[21\].rs_mbuf
timestamp 1693170804
transform 1 0 27324 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 26956 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 27232 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18952 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 26588 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26312 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 26956 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26220 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26220 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 26680 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 26680 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[22\].cc_clkbuf
timestamp 1693170804
transform 1 0 27140 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[22\].rs_mbuf
timestamp 1693170804
transform 1 0 26680 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 11500 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[23\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 25944 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 25668 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 24012 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 26036 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 24012 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 24196 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 23920 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 13616 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[23\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[23\].cc_clkbuf
timestamp 1693170804
transform 1 0 26404 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[23\].rs_mbuf
timestamp 1693170804
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 23736 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 23092 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 22816 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 21804 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 21896 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 22540 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 22816 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[24\].cc_clkbuf
timestamp 1693170804
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[24\].rs_mbuf
timestamp 1693170804
transform 1 0 22264 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 23092 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 19964 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 19872 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 20792 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 23368 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 20792 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[25\].cc_clkbuf
timestamp 1693170804
transform 1 0 20608 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[25\].rs_mbuf
timestamp 1693170804
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 20516 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 19320 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 17940 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 18216 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 18676 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 20792 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 19596 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[26\].cc_clkbuf
timestamp 1693170804
transform 1 0 18768 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[26\].rs_mbuf
timestamp 1693170804
transform 1 0 18032 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 17664 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 16284 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 15824 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 17388 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 15824 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 18032 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 15824 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[27\].cc_clkbuf
timestamp 1693170804
transform 1 0 18032 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[27\].rs_mbuf
timestamp 1693170804
transform 1 0 16836 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13708 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 13708 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 8464 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 12880 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13616 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 13800 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 13616 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10028 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[28\].cc_clkbuf
timestamp 1693170804
transform 1 0 12328 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[28\].rs_mbuf
timestamp 1693170804
transform 1 0 12880 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 11500 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 8740 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 11040 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 12604 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 12328 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10304 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[29\].cc_clkbuf
timestamp 1693170804
transform 1 0 11040 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[29\].rs_mbuf
timestamp 1693170804
transform 1 0 11040 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 4876 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 8740 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 10028 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 9844 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10304 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 3588 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 9016 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[30\].cc_clkbuf
timestamp 1693170804
transform 1 0 10948 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[30\].rs_mbuf
timestamp 1693170804
transform 1 0 9292 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 7452 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 8648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 7820 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 3956 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 7728 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 5980 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[31\].cc_clkbuf
timestamp 1693170804
transform 1 0 8372 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[31\].rs_mbuf
timestamp 1693170804
transform 1 0 8096 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[32\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 8924 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 15732 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[32\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 9200 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 5888 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 6624 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 6900 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 5888 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[32\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 8648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 7176 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[32\].cc_clkbuf
timestamp 1693170804
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[32\].rs_mbuf
timestamp 1693170804
transform 1 0 5796 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 13616 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 11316 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3680 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 5152 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 1288 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 1012 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 17204 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[33\].cc_clkbuf
timestamp 1693170804
transform 1 0 2392 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[33\].rs_mbuf
timestamp 1693170804
transform 1 0 6808 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 11500 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 18676 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 7452 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[34\].cc_clkbuf
timestamp 1693170804
transform 1 0 5796 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[34\].rs_mbuf
timestamp 1693170804
transform 1 0 5796 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 1196 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 5520 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 6348 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 1104 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 5520 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[35\].cc_clkbuf
timestamp 1693170804
transform 1 0 3864 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[35\].rs_mbuf
timestamp 1693170804
transform 1 0 5796 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 9384 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 8648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 8924 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 6716 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 9476 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 8464 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 8740 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[36\].cc_clkbuf
timestamp 1693170804
transform 1 0 5796 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[36\].rs_mbuf
timestamp 1693170804
transform 1 0 7728 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16928 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 14720 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 15640 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 15916 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 14536 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 14628 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 13892 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 14812 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 12788 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 12144 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 13064 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[37\].cc_clkbuf
timestamp 1693170804
transform 1 0 10948 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[37\].rs_mbuf
timestamp 1693170804
transform 1 0 14168 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13892 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 14720 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13708 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 13432 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13708 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 14996 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11132 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10304 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11132 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 11132 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[38\].cc_clkbuf
timestamp 1693170804
transform 1 0 12236 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[38\].rs_mbuf
timestamp 1693170804
transform 1 0 12880 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 12512 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 12512 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 12236 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 12604 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 12788 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 12512 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 12880 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8924 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10028 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 9660 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[39\].cc_clkbuf
timestamp 1693170804
transform 1 0 11776 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[39\].rs_mbuf
timestamp 1693170804
transform 1 0 14720 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 9568 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 10304 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 9568 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 9292 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 9568 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 10028 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 7636 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 7360 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[40\].cc_clkbuf
timestamp 1693170804
transform 1 0 9016 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[40\].rs_mbuf
timestamp 1693170804
transform 1 0 8464 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 6164 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6624 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 6164 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 9016 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6716 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 8740 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 6440 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 6072 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[41\].cc_clkbuf
timestamp 1693170804
transform 1 0 7728 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[41\].rs_mbuf
timestamp 1693170804
transform 1 0 5888 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3772 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3772 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 1196 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 3496 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 3496 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[42\].cc_clkbuf
timestamp 1693170804
transform 1 0 4508 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[42\].rs_mbuf
timestamp 1693170804
transform 1 0 3680 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 1472 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 1472 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 3496 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 1012 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 1564 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[43\].cc_clkbuf
timestamp 1693170804
transform 1 0 920 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[43\].rs_mbuf
timestamp 1693170804
transform 1 0 5060 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dlclkp_4  ct.ro.cc_clock_gate $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 19596 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_4  ct.ro.cc_clock_inv $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 23276 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  ct.ro.cc_ring_osc_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 19596 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  ct.ro.cc_ring_osc_1
timestamp 1693170804
transform 1 0 23000 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  ct.ro.cc_ring_osc_2
timestamp 1693170804
transform 1 0 23276 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[1\].cc_div_flop $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 18952 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[2\].cc_div_flop
timestamp 1693170804
transform 1 0 19320 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[3\].cc_div_flop
timestamp 1693170804
transform 1 0 21252 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[4\].cc_div_flop
timestamp 1693170804
transform 1 0 23460 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[5\].cc_div_flop
timestamp 1693170804
transform 1 0 22172 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[6\].cc_div_flop
timestamp 1693170804
transform 1 0 21528 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[7\].cc_div_flop
timestamp 1693170804
transform 1 0 23828 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2i_2  cw.cc_test_0
timestamp 1693170804
transform 1 0 16192 0 -1 21216
box -38 -48 1050 592
use sky130_ht_sc_tt05__mux2i_2  cw.cc_test_1
timestamp 1698685089
transform 1 0 16100 0 -1 17952
box -38 -48 1050 592
use sky130_fd_sc_hd__maj3_2  cw.cc_test_2
timestamp 1693170804
transform 1 0 17664 0 1 19040
box -38 -48 866 592
use sky130_ht_sc_tt05__maj3_2  cw.cc_test_3
timestamp 1698685089
transform 1 0 11224 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dlrtp_1  cw.cc_test_4
timestamp 1693170804
transform 1 0 14444 0 1 16864
box -38 -48 1234 592
use sky130_ht_sc_tt05__dlrtp_1  cw.cc_test_5
timestamp 1698685089
transform 1 0 12052 0 -1 16864
box -38 -48 1418 592
use sky130_fd_sc_hd__dfrtp_1  cw.cc_test_6
timestamp 1693170804
transform 1 0 14260 0 1 20128
box -38 -48 1878 592
use sky130_ht_sc_tt05__dfrtp_1  cw.cc_test_7
timestamp 1698685089
transform 1 0 13892 0 -1 21216
box -38 -48 2154 592
use sky130_fd_sc_hd__buf_2  fanout5
timestamp 1693170804
transform 1 0 9016 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 13524 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout7
timestamp 1693170804
transform 1 0 13524 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout8
timestamp 1693170804
transform 1 0 26864 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout9
timestamp 1693170804
transform 1 0 29716 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout10
timestamp 1693170804
transform 1 0 8188 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout11
timestamp 1693170804
transform 1 0 11776 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout12
timestamp 1693170804
transform 1 0 11040 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 1693170804
transform 1 0 28980 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1693170804
transform 1 0 29992 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout15
timestamp 1693170804
transform 1 0 8372 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 1693170804
transform 1 0 12144 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout17
timestamp 1693170804
transform 1 0 13524 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 1693170804
transform 1 0 28980 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout19
timestamp 1693170804
transform 1 0 28980 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout20
timestamp 1693170804
transform 1 0 29348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1693170804
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout22
timestamp 1693170804
transform 1 0 13064 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1693170804
transform 1 0 16100 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 1693170804
transform 1 0 29348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1693170804
transform 1 0 28980 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout26
timestamp 1693170804
transform 1 0 30176 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout27
timestamp 1693170804
transform 1 0 15088 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1693170804
transform 1 0 16652 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout29
timestamp 1693170804
transform 1 0 10856 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout30
timestamp 1693170804
transform 1 0 23828 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 1693170804
transform 1 0 30084 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout32
timestamp 1693170804
transform 1 0 28980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 1693170804
transform 1 0 5336 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout34
timestamp 1693170804
transform 1 0 12328 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout35
timestamp 1693170804
transform 1 0 10856 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout36
timestamp 1693170804
transform 1 0 27140 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout37
timestamp 1693170804
transform 1 0 28244 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp 1693170804
transform 1 0 30268 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 1693170804
transform 1 0 13432 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout40
timestamp 1693170804
transform 1 0 16100 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout41
timestamp 1693170804
transform 1 0 8280 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1693170804
transform 1 0 29532 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 1693170804
transform 1 0 28244 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 1693170804
transform 1 0 29532 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 1693170804
transform 1 0 11500 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout46
timestamp 1693170804
transform 1 0 13524 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 1693170804
transform 1 0 13156 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout48
timestamp 1693170804
transform 1 0 30084 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1693170804
transform 1 0 25760 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp 1693170804
transform 1 0 26312 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 1693170804
transform 1 0 14076 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout52
timestamp 1693170804
transform 1 0 7728 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout53
timestamp 1693170804
transform 1 0 25668 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout54
timestamp 1693170804
transform 1 0 25760 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout55
timestamp 1693170804
transform 1 0 26036 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 828 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3220 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_36
timestamp 1693170804
transform 1 0 3864 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4232 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_44
timestamp 1693170804
transform 1 0 4600 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28980 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_321 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 30084 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_6
timestamp 1693170804
transform 1 0 1104 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_63
timestamp 1693170804
transform 1 0 6348 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1693170804
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1693170804
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1693170804
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_317 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 29716 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_325
timestamp 1693170804
transform 1 0 30452 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 1693170804
transform 1 0 828 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_56
timestamp 1693170804
transform 1 0 5704 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 1693170804
transform 1 0 8372 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 1693170804
transform 1 0 13524 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1693170804
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_277 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 26036 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1693170804
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_312
timestamp 1693170804
transform 1 0 29256 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_324
timestamp 1693170804
transform 1 0 30360 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_3
timestamp 1693170804
transform 1 0 828 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_7
timestamp 1693170804
transform 1 0 1196 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_32
timestamp 1693170804
transform 1 0 3496 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_36
timestamp 1693170804
transform 1 0 3864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_48
timestamp 1693170804
transform 1 0 4968 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 1693170804
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_74
timestamp 1693170804
transform 1 0 7360 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_102
timestamp 1693170804
transform 1 0 9936 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1693170804
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_217
timestamp 1693170804
transform 1 0 20516 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_255
timestamp 1693170804
transform 1 0 24012 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_287
timestamp 1693170804
transform 1 0 26956 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_295
timestamp 1693170804
transform 1 0 27692 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_324
timestamp 1693170804
transform 1 0 30360 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_3
timestamp 1693170804
transform 1 0 828 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29
timestamp 1693170804
transform 1 0 3220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_33
timestamp 1693170804
transform 1 0 3588 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_58
timestamp 1693170804
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_91
timestamp 1693170804
transform 1 0 8924 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_141
timestamp 1693170804
transform 1 0 13524 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1693170804
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_277
timestamp 1693170804
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_306
timestamp 1693170804
transform 1 0 28704 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1693170804
transform 1 0 28980 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_321
timestamp 1693170804
transform 1 0 30084 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_3
timestamp 1693170804
transform 1 0 828 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_14
timestamp 1693170804
transform 1 0 1840 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_26
timestamp 1693170804
transform 1 0 2944 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_30
timestamp 1693170804
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1693170804
transform 1 0 5796 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp 1693170804
transform 1 0 10948 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1693170804
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1693170804
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_290
timestamp 1693170804
transform 1 0 27232 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_321
timestamp 1693170804
transform 1 0 30084 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 1693170804
transform 1 0 828 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_56
timestamp 1693170804
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1693170804
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_88
timestamp 1693170804
transform 1 0 8648 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_168
timestamp 1693170804
transform 1 0 16008 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_197
timestamp 1693170804
transform 1 0 18676 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_234
timestamp 1693170804
transform 1 0 22080 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_248
timestamp 1693170804
transform 1 0 23368 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1693170804
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_303
timestamp 1693170804
transform 1 0 28428 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1693170804
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1693170804
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_321
timestamp 1693170804
transform 1 0 30084 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 1693170804
transform 1 0 828 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_7
timestamp 1693170804
transform 1 0 1196 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_63
timestamp 1693170804
transform 1 0 6348 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1693170804
transform 1 0 10948 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1693170804
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_228
timestamp 1693170804
transform 1 0 21528 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1693170804
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_281
timestamp 1693170804
transform 1 0 26404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_289
timestamp 1693170804
transform 1 0 27140 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_317
timestamp 1693170804
transform 1 0 29716 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_325
timestamp 1693170804
transform 1 0 30452 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1693170804
transform 1 0 828 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_56
timestamp 1693170804
transform 1 0 5704 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_91
timestamp 1693170804
transform 1 0 8924 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_141
timestamp 1693170804
transform 1 0 13524 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_245
timestamp 1693170804
transform 1 0 23092 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_249
timestamp 1693170804
transform 1 0 23460 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_280
timestamp 1693170804
transform 1 0 26312 0 1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_315
timestamp 1693170804
transform 1 0 29532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_6
timestamp 1693170804
transform 1 0 1104 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_32
timestamp 1693170804
transform 1 0 3496 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_48
timestamp 1693170804
transform 1 0 4968 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_52
timestamp 1693170804
transform 1 0 5336 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_78
timestamp 1693170804
transform 1 0 7728 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 1693170804
transform 1 0 10948 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1693170804
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_228
timestamp 1693170804
transform 1 0 21528 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_317
timestamp 1693170804
transform 1 0 29716 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_325
timestamp 1693170804
transform 1 0 30452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 1693170804
transform 1 0 828 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 1693170804
transform 1 0 3220 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_121
timestamp 1693170804
transform 1 0 11684 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1693170804
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_200
timestamp 1693170804
transform 1 0 18952 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_235
timestamp 1693170804
transform 1 0 22172 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1693170804
transform 1 0 23092 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1693170804
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_253
timestamp 1693170804
transform 1 0 23828 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_312
timestamp 1693170804
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_324
timestamp 1693170804
transform 1 0 30360 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_30
timestamp 1693170804
transform 1 0 3312 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_63
timestamp 1693170804
transform 1 0 6348 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_125
timestamp 1693170804
transform 1 0 12052 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_150
timestamp 1693170804
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1693170804
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_169
timestamp 1693170804
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_174
timestamp 1693170804
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_225
timestamp 1693170804
transform 1 0 21252 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_229
timestamp 1693170804
transform 1 0 21620 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_255
timestamp 1693170804
transform 1 0 24012 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_281
timestamp 1693170804
transform 1 0 26404 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_319
timestamp 1693170804
transform 1 0 29900 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 1693170804
transform 1 0 828 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1693170804
transform 1 0 3220 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1693170804
transform 1 0 8372 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_141
timestamp 1693170804
transform 1 0 13524 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1693170804
transform 1 0 23644 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_283
timestamp 1693170804
transform 1 0 26588 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_315
timestamp 1693170804
transform 1 0 29532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_3
timestamp 1693170804
transform 1 0 828 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_31
timestamp 1693170804
transform 1 0 3404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_63
timestamp 1693170804
transform 1 0 6348 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_119
timestamp 1693170804
transform 1 0 11500 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_220
timestamp 1693170804
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1693170804
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_281
timestamp 1693170804
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_288
timestamp 1693170804
transform 1 0 27048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_322
timestamp 1693170804
transform 1 0 30176 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_326
timestamp 1693170804
transform 1 0 30544 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 1693170804
transform 1 0 828 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_53
timestamp 1693170804
transform 1 0 5428 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_94
timestamp 1693170804
transform 1 0 9200 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_126
timestamp 1693170804
transform 1 0 12144 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1693170804
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 1693170804
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1693170804
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_221
timestamp 1693170804
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_277
timestamp 1693170804
transform 1 0 26036 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1693170804
transform 1 0 28796 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 1693170804
transform 1 0 828 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_63
timestamp 1693170804
transform 1 0 6348 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_73
timestamp 1693170804
transform 1 0 7268 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_101
timestamp 1693170804
transform 1 0 9844 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1693170804
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_139
timestamp 1693170804
transform 1 0 13340 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1693170804
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1693170804
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_173
timestamp 1693170804
transform 1 0 16468 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_216
timestamp 1693170804
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1693170804
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_305
timestamp 1693170804
transform 1 0 28612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_325
timestamp 1693170804
transform 1 0 30452 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 1693170804
transform 1 0 828 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_29
timestamp 1693170804
transform 1 0 3220 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_89
timestamp 1693170804
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1693170804
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_168
timestamp 1693170804
transform 1 0 16008 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_245
timestamp 1693170804
transform 1 0 23092 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_259
timestamp 1693170804
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_285
timestamp 1693170804
transform 1 0 26772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_304
timestamp 1693170804
transform 1 0 28520 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1693170804
transform 1 0 28980 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_321
timestamp 1693170804
transform 1 0 30084 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 1693170804
transform 1 0 828 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1693170804
transform 1 0 5796 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 1693170804
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_139
timestamp 1693170804
transform 1 0 13340 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_175
timestamp 1693170804
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_210
timestamp 1693170804
transform 1 0 19872 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_214
timestamp 1693170804
transform 1 0 20240 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_249
timestamp 1693170804
transform 1 0 23460 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_255
timestamp 1693170804
transform 1 0 24012 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_3
timestamp 1693170804
transform 1 0 828 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_53
timestamp 1693170804
transform 1 0 5428 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_85
timestamp 1693170804
transform 1 0 8372 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_96
timestamp 1693170804
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_169
timestamp 1693170804
transform 1 0 16100 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_203
timestamp 1693170804
transform 1 0 19228 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_211
timestamp 1693170804
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_240
timestamp 1693170804
transform 1 0 22632 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_247
timestamp 1693170804
transform 1 0 23276 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1693170804
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_277
timestamp 1693170804
transform 1 0 26036 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_306
timestamp 1693170804
transform 1 0 28704 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_323
timestamp 1693170804
transform 1 0 30268 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_3
timestamp 1693170804
transform 1 0 828 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1693170804
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_81
timestamp 1693170804
transform 1 0 8004 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_87
timestamp 1693170804
transform 1 0 8556 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_160
timestamp 1693170804
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_164
timestamp 1693170804
transform 1 0 15640 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_169
timestamp 1693170804
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_173
timestamp 1693170804
transform 1 0 16468 0 -1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_207
timestamp 1693170804
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_219
timestamp 1693170804
transform 1 0 20700 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1693170804
transform 1 0 21068 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1693170804
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_326
timestamp 1693170804
transform 1 0 30544 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_3
timestamp 1693170804
transform 1 0 828 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_59
timestamp 1693170804
transform 1 0 5980 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_91
timestamp 1693170804
transform 1 0 8924 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_131
timestamp 1693170804
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_165
timestamp 1693170804
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_245
timestamp 1693170804
transform 1 0 23092 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_319
timestamp 1693170804
transform 1 0 29900 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1693170804
transform 1 0 828 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_60
timestamp 1693170804
transform 1 0 6072 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_125
timestamp 1693170804
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1693170804
transform 1 0 15824 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_172
timestamp 1693170804
transform 1 0 16376 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_211
timestamp 1693170804
transform 1 0 19964 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1693170804
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_3
timestamp 1693170804
transform 1 0 828 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_35
timestamp 1693170804
transform 1 0 3772 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1693170804
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1693170804
transform 1 0 23644 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_283
timestamp 1693170804
transform 1 0 26588 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_325
timestamp 1693170804
transform 1 0 30452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp 1693170804
transform 1 0 828 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_60
timestamp 1693170804
transform 1 0 6072 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_113
timestamp 1693170804
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_163
timestamp 1693170804
transform 1 0 15548 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1693170804
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1693170804
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_225
timestamp 1693170804
transform 1 0 21252 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_3
timestamp 1693170804
transform 1 0 828 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_59
timestamp 1693170804
transform 1 0 5980 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_115
timestamp 1693170804
transform 1 0 11132 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1693170804
transform 1 0 13524 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_203
timestamp 1693170804
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_207
timestamp 1693170804
transform 1 0 19596 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_253
timestamp 1693170804
transform 1 0 23828 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_279
timestamp 1693170804
transform 1 0 26220 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_326
timestamp 1693170804
transform 1 0 30544 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_3
timestamp 1693170804
transform 1 0 828 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_40
timestamp 1693170804
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_51
timestamp 1693170804
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_105
timestamp 1693170804
transform 1 0 10212 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_113
timestamp 1693170804
transform 1 0 10948 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_179
timestamp 1693170804
transform 1 0 17020 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_210
timestamp 1693170804
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_220
timestamp 1693170804
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1693170804
transform 1 0 26220 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_281
timestamp 1693170804
transform 1 0 26404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_298
timestamp 1693170804
transform 1 0 27968 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_3
timestamp 1693170804
transform 1 0 828 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_59
timestamp 1693170804
transform 1 0 5980 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_85
timestamp 1693170804
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_111
timestamp 1693170804
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_147
timestamp 1693170804
transform 1 0 14076 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_209
timestamp 1693170804
transform 1 0 19780 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_234
timestamp 1693170804
transform 1 0 22080 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_247
timestamp 1693170804
transform 1 0 23276 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1693170804
transform 1 0 28796 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_319
timestamp 1693170804
transform 1 0 29900 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_3
timestamp 1693170804
transform 1 0 828 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1693170804
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_119
timestamp 1693170804
transform 1 0 11500 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_273
timestamp 1693170804
transform 1 0 25668 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_3
timestamp 1693170804
transform 1 0 828 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_59
timestamp 1693170804
transform 1 0 5980 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_85
timestamp 1693170804
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_111
timestamp 1693170804
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_150
timestamp 1693170804
transform 1 0 14352 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_227
timestamp 1693170804
transform 1 0 21436 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1693170804
transform 1 0 28796 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_3
timestamp 1693170804
transform 1 0 828 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_31
timestamp 1693170804
transform 1 0 3404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1693170804
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_113
timestamp 1693170804
transform 1 0 10948 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_120
timestamp 1693170804
transform 1 0 11592 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_124
timestamp 1693170804
transform 1 0 11960 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_143
timestamp 1693170804
transform 1 0 13708 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_178
timestamp 1693170804
transform 1 0 16928 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_204
timestamp 1693170804
transform 1 0 19320 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1693170804
transform 1 0 26220 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_3
timestamp 1693170804
transform 1 0 828 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_35
timestamp 1693170804
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_150
timestamp 1693170804
transform 1 0 14352 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_170
timestamp 1693170804
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_216
timestamp 1693170804
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1693170804
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_256
timestamp 1693170804
transform 1 0 24104 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1693170804
transform 1 0 28796 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_326
timestamp 1693170804
transform 1 0 30544 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_3
timestamp 1693170804
transform 1 0 828 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_63
timestamp 1693170804
transform 1 0 6348 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_204
timestamp 1693170804
transform 1 0 19320 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_252
timestamp 1693170804
transform 1 0 23736 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_300
timestamp 1693170804
transform 1 0 28152 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_326
timestamp 1693170804
transform 1 0 30544 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_3
timestamp 1693170804
transform 1 0 828 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_35
timestamp 1693170804
transform 1 0 3772 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 1693170804
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_111
timestamp 1693170804
transform 1 0 10764 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_175
timestamp 1693170804
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_216
timestamp 1693170804
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_245
timestamp 1693170804
transform 1 0 23092 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_256
timestamp 1693170804
transform 1 0 24104 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1693170804
transform 1 0 28796 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_3
timestamp 1693170804
transform 1 0 828 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_32
timestamp 1693170804
transform 1 0 3496 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_42
timestamp 1693170804
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_57
timestamp 1693170804
transform 1 0 5796 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_83
timestamp 1693170804
transform 1 0 8188 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_147
timestamp 1693170804
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1693170804
transform 1 0 20976 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_249
timestamp 1693170804
transform 1 0 23460 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_281
timestamp 1693170804
transform 1 0 26404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_3
timestamp 1693170804
transform 1 0 828 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_29
timestamp 1693170804
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_76
timestamp 1693170804
transform 1 0 7544 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_109
timestamp 1693170804
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_138
timestamp 1693170804
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_141
timestamp 1693170804
transform 1 0 13524 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1693170804
transform 1 0 18492 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_241
timestamp 1693170804
transform 1 0 22724 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_253
timestamp 1693170804
transform 1 0 23828 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_326
timestamp 1693170804
transform 1 0 30544 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_3
timestamp 1693170804
transform 1 0 828 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_28
timestamp 1693170804
transform 1 0 3128 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_81
timestamp 1693170804
transform 1 0 8004 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_110
timestamp 1693170804
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_234
timestamp 1693170804
transform 1 0 22080 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_278
timestamp 1693170804
transform 1 0 26128 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_3
timestamp 1693170804
transform 1 0 828 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_35
timestamp 1693170804
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_85
timestamp 1693170804
transform 1 0 8372 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_141
timestamp 1693170804
transform 1 0 13524 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_194
timestamp 1693170804
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_202
timestamp 1693170804
transform 1 0 19136 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_283
timestamp 1693170804
transform 1 0 26588 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_326
timestamp 1693170804
transform 1 0 30544 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_3
timestamp 1693170804
transform 1 0 828 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_81
timestamp 1693170804
transform 1 0 8004 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_143
timestamp 1693170804
transform 1 0 13708 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_169
timestamp 1693170804
transform 1 0 16100 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1693170804
transform 1 0 26220 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_300
timestamp 1693170804
transform 1 0 28152 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_326
timestamp 1693170804
transform 1 0 30544 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_3
timestamp 1693170804
transform 1 0 828 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_113
timestamp 1693170804
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1693170804
transform 1 0 13340 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_147
timestamp 1693170804
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_175
timestamp 1693170804
transform 1 0 16652 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_203
timestamp 1693170804
transform 1 0 19228 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_225
timestamp 1693170804
transform 1 0 21252 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 1693170804
transform 1 0 28704 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1693170804
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1693170804
transform 1 0 30268 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1693170804
transform 1 0 30084 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1693170804
transform 1 0 28152 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_39
timestamp 1693170804
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1693170804
transform -1 0 30912 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_40
timestamp 1693170804
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1693170804
transform -1 0 30912 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_41
timestamp 1693170804
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1693170804
transform -1 0 30912 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_42
timestamp 1693170804
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1693170804
transform -1 0 30912 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_43
timestamp 1693170804
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1693170804
transform -1 0 30912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_44
timestamp 1693170804
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1693170804
transform -1 0 30912 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_45
timestamp 1693170804
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1693170804
transform -1 0 30912 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_46
timestamp 1693170804
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1693170804
transform -1 0 30912 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_47
timestamp 1693170804
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1693170804
transform -1 0 30912 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_48
timestamp 1693170804
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1693170804
transform -1 0 30912 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_49
timestamp 1693170804
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1693170804
transform -1 0 30912 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_50
timestamp 1693170804
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1693170804
transform -1 0 30912 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_51
timestamp 1693170804
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1693170804
transform -1 0 30912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_52
timestamp 1693170804
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1693170804
transform -1 0 30912 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_53
timestamp 1693170804
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1693170804
transform -1 0 30912 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_54
timestamp 1693170804
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1693170804
transform -1 0 30912 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_55
timestamp 1693170804
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1693170804
transform -1 0 30912 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_56
timestamp 1693170804
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1693170804
transform -1 0 30912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_57
timestamp 1693170804
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1693170804
transform -1 0 30912 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_58
timestamp 1693170804
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1693170804
transform -1 0 30912 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_59
timestamp 1693170804
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1693170804
transform -1 0 30912 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_60
timestamp 1693170804
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1693170804
transform -1 0 30912 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_61
timestamp 1693170804
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1693170804
transform -1 0 30912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_62
timestamp 1693170804
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1693170804
transform -1 0 30912 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_63
timestamp 1693170804
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1693170804
transform -1 0 30912 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_64
timestamp 1693170804
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1693170804
transform -1 0 30912 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_65
timestamp 1693170804
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1693170804
transform -1 0 30912 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_66
timestamp 1693170804
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1693170804
transform -1 0 30912 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_67
timestamp 1693170804
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1693170804
transform -1 0 30912 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_68
timestamp 1693170804
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1693170804
transform -1 0 30912 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_69
timestamp 1693170804
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1693170804
transform -1 0 30912 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_70
timestamp 1693170804
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1693170804
transform -1 0 30912 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_71
timestamp 1693170804
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1693170804
transform -1 0 30912 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_72
timestamp 1693170804
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1693170804
transform -1 0 30912 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_73
timestamp 1693170804
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1693170804
transform -1 0 30912 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_74
timestamp 1693170804
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1693170804
transform -1 0 30912 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_75
timestamp 1693170804
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1693170804
transform -1 0 30912 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_76
timestamp 1693170804
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1693170804
transform -1 0 30912 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_77
timestamp 1693170804
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1693170804
transform -1 0 30912 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp 1693170804
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp 1693170804
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_81
timestamp 1693170804
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82
timestamp 1693170804
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_83
timestamp 1693170804
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 1693170804
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1693170804
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1693170804
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1693170804
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1693170804
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_89
timestamp 1693170804
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_90
timestamp 1693170804
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_91
timestamp 1693170804
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1693170804
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1693170804
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_94
timestamp 1693170804
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_95
timestamp 1693170804
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1693170804
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1693170804
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1693170804
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1693170804
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1693170804
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1693170804
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1693170804
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1693170804
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_104
timestamp 1693170804
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1693170804
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1693170804
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1693170804
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_108
timestamp 1693170804
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_109
timestamp 1693170804
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_110
timestamp 1693170804
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1693170804
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_112
timestamp 1693170804
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_113
timestamp 1693170804
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_114
timestamp 1693170804
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_115
timestamp 1693170804
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_116
timestamp 1693170804
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_117
timestamp 1693170804
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_118
timestamp 1693170804
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_119
timestamp 1693170804
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_120
timestamp 1693170804
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_121
timestamp 1693170804
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_122
timestamp 1693170804
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_123
timestamp 1693170804
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_124
timestamp 1693170804
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_125
timestamp 1693170804
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_126
timestamp 1693170804
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_127
timestamp 1693170804
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_128
timestamp 1693170804
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_129
timestamp 1693170804
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_130
timestamp 1693170804
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_131
timestamp 1693170804
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_132
timestamp 1693170804
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_133
timestamp 1693170804
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_134
timestamp 1693170804
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_135
timestamp 1693170804
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_136
timestamp 1693170804
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_137
timestamp 1693170804
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_138
timestamp 1693170804
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_139
timestamp 1693170804
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_140
timestamp 1693170804
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 1693170804
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_142
timestamp 1693170804
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 1693170804
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp 1693170804
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp 1693170804
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp 1693170804
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp 1693170804
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp 1693170804
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_149
timestamp 1693170804
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_150
timestamp 1693170804
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_151
timestamp 1693170804
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_152
timestamp 1693170804
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_153
timestamp 1693170804
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_154
timestamp 1693170804
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_155
timestamp 1693170804
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_156
timestamp 1693170804
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_157
timestamp 1693170804
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_158
timestamp 1693170804
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_159
timestamp 1693170804
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_160
timestamp 1693170804
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_161
timestamp 1693170804
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_162
timestamp 1693170804
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp 1693170804
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_164
timestamp 1693170804
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_165
timestamp 1693170804
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_166
timestamp 1693170804
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_167
timestamp 1693170804
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_168
timestamp 1693170804
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_169
timestamp 1693170804
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_170
timestamp 1693170804
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_171
timestamp 1693170804
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_172
timestamp 1693170804
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_173
timestamp 1693170804
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_174
timestamp 1693170804
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_175
timestamp 1693170804
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_176
timestamp 1693170804
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_177
timestamp 1693170804
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_178
timestamp 1693170804
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_179
timestamp 1693170804
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_180
timestamp 1693170804
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_181
timestamp 1693170804
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_182
timestamp 1693170804
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_183
timestamp 1693170804
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_184
timestamp 1693170804
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 1693170804
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_186
timestamp 1693170804
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_187
timestamp 1693170804
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_188
timestamp 1693170804
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_189
timestamp 1693170804
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_190
timestamp 1693170804
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_191
timestamp 1693170804
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_192
timestamp 1693170804
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_193
timestamp 1693170804
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_194
timestamp 1693170804
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_195
timestamp 1693170804
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_196
timestamp 1693170804
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_197
timestamp 1693170804
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_198
timestamp 1693170804
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_199
timestamp 1693170804
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_200
timestamp 1693170804
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_201
timestamp 1693170804
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_202
timestamp 1693170804
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_203
timestamp 1693170804
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_204
timestamp 1693170804
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_205
timestamp 1693170804
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_206
timestamp 1693170804
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_207
timestamp 1693170804
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_208
timestamp 1693170804
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp 1693170804
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_210
timestamp 1693170804
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_211
timestamp 1693170804
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_212
timestamp 1693170804
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_213
timestamp 1693170804
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp 1693170804
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_215
timestamp 1693170804
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_216
timestamp 1693170804
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_217
timestamp 1693170804
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_218
timestamp 1693170804
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp 1693170804
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp 1693170804
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_221
timestamp 1693170804
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_222
timestamp 1693170804
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_223
timestamp 1693170804
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp 1693170804
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp 1693170804
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_226
timestamp 1693170804
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_227
timestamp 1693170804
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_228
timestamp 1693170804
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp 1693170804
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp 1693170804
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp 1693170804
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_232
timestamp 1693170804
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_233
timestamp 1693170804
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp 1693170804
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp 1693170804
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp 1693170804
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_237
timestamp 1693170804
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_238
timestamp 1693170804
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp 1693170804
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp 1693170804
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp 1693170804
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp 1693170804
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_243
timestamp 1693170804
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp 1693170804
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp 1693170804
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp 1693170804
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp 1693170804
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_248
timestamp 1693170804
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp 1693170804
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp 1693170804
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp 1693170804
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp 1693170804
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 1693170804
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp 1693170804
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp 1693170804
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp 1693170804
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp 1693170804
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 1693170804
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp 1693170804
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp 1693170804
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp 1693170804
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp 1693170804
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 1693170804
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 1693170804
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1693170804
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp 1693170804
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp 1693170804
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 1693170804
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 1693170804
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp 1693170804
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp 1693170804
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp 1693170804
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 1693170804
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 1693170804
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1693170804
transform 1 0 28888 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp 1693170804
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp 1693170804
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 1693170804
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 1693170804
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1693170804
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp 1693170804
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp 1693170804
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 1693170804
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 1693170804
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1693170804
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 1693170804
transform 1 0 28888 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp 1693170804
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 1693170804
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 1693170804
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1693170804
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 1693170804
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp 1693170804
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 1693170804
transform 1 0 5704 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 1693170804
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1693170804
transform 1 0 10856 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 1693170804
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 1693170804
transform 1 0 16008 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_298
timestamp 1693170804
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp 1693170804
transform 1 0 21160 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_300
timestamp 1693170804
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp 1693170804
transform 1 0 26312 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_302
timestamp 1693170804
transform 1 0 28888 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 11776 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_57
timestamp 1693170804
transform 1 0 10948 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_58
timestamp 1693170804
transform 1 0 10580 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_59
timestamp 1693170804
transform 1 0 8648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_60
timestamp 1693170804
transform 1 0 11408 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_61
timestamp 1693170804
transform 1 0 16376 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_62
timestamp 1693170804
transform 1 0 11224 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_63
timestamp 1693170804
transform 1 0 12052 0 1 12512
box -38 -48 314 592
<< labels >>
flabel metal4 s 7982 496 8302 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15572 496 15892 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 23162 496 23482 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 30752 496 31072 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4187 496 4507 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11777 496 12097 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19367 496 19687 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26957 496 27277 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26926 22104 26986 22304 0 FreeSans 480 90 0 0 clk
port 2 nsew signal input
flabel metal4 s 27478 22104 27538 22304 0 FreeSans 480 90 0 0 ena
port 3 nsew signal input
flabel metal4 s 26374 22104 26434 22304 0 FreeSans 480 90 0 0 rst_n
port 4 nsew signal input
flabel metal4 s 25822 22104 25882 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 5 nsew signal input
flabel metal4 s 25270 22104 25330 22304 0 FreeSans 480 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal4 s 24718 22104 24778 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal4 s 24166 22104 24226 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal4 s 23614 22104 23674 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal4 s 23062 22104 23122 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal4 s 22510 22104 22570 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal4 s 21958 22104 22018 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal4 s 21406 22104 21466 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal4 s 20854 22104 20914 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal4 s 20302 22104 20362 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal4 s 19750 22104 19810 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal4 s 19198 22104 19258 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal4 s 18646 22104 18706 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal4 s 18094 22104 18154 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal4 s 17542 22104 17602 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal4 s 8158 22104 8218 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 21 nsew signal tristate
flabel metal4 s 7606 22104 7666 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 22 nsew signal tristate
flabel metal4 s 7054 22104 7114 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 23 nsew signal tristate
flabel metal4 s 6502 22104 6562 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 24 nsew signal tristate
flabel metal4 s 5950 22104 6010 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 25 nsew signal tristate
flabel metal4 s 5398 22104 5458 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 26 nsew signal tristate
flabel metal4 s 4846 22104 4906 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 27 nsew signal tristate
flabel metal4 s 4294 22104 4354 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 28 nsew signal tristate
flabel metal4 s 12574 22104 12634 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 29 nsew signal tristate
flabel metal4 s 12022 22104 12082 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 30 nsew signal tristate
flabel metal4 s 11470 22104 11530 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 31 nsew signal tristate
flabel metal4 s 10918 22104 10978 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 32 nsew signal tristate
flabel metal4 s 10366 22104 10426 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 33 nsew signal tristate
flabel metal4 s 9814 22104 9874 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 34 nsew signal tristate
flabel metal4 s 9262 22104 9322 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 35 nsew signal tristate
flabel metal4 s 8710 22104 8770 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 36 nsew signal tristate
flabel metal4 s 16990 22104 17050 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 37 nsew signal tristate
flabel metal4 s 16438 22104 16498 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 38 nsew signal tristate
flabel metal4 s 15886 22104 15946 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 39 nsew signal tristate
flabel metal4 s 15334 22104 15394 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 40 nsew signal tristate
flabel metal4 s 14782 22104 14842 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 41 nsew signal tristate
flabel metal4 s 14230 22104 14290 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 42 nsew signal tristate
flabel metal4 s 13678 22104 13738 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 43 nsew signal tristate
flabel metal4 s 13126 22104 13186 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 44 nsew signal tristate
rlabel via1 15812 21216 15812 21216 0 VGND
rlabel metal1 15732 21760 15732 21760 0 VPWR
rlabel metal2 26174 16699 26174 16699 0 _00_
rlabel metal1 23184 19278 23184 19278 0 _01_
rlabel metal1 23966 19278 23966 19278 0 _02_
rlabel metal1 23598 19142 23598 19142 0 _03_
rlabel metal1 21988 19890 21988 19890 0 _04_
rlabel metal1 25070 19142 25070 19142 0 ct.cw.source\[0\]
rlabel metal1 25484 19142 25484 19142 0 ct.cw.source\[1\]
rlabel metal1 28343 18870 28343 18870 0 ct.cw.source\[2\]
rlabel metal2 1978 13345 1978 13345 0 ct.cw.target\[0\]
rlabel metal2 1978 11169 1978 11169 0 ct.cw.target\[1\]
rlabel metal2 2070 14433 2070 14433 0 ct.cw.target\[2\]
rlabel via2 2162 12835 2162 12835 0 ct.cw.target\[3\]
rlabel metal1 1794 9146 1794 9146 0 ct.cw.target\[4\]
rlabel metal1 14720 16014 14720 16014 0 ct.cw.target\[5\]
rlabel metal1 16146 17068 16146 17068 0 ct.cw.target\[6\]
rlabel metal1 13616 15946 13616 15946 0 ct.cw.target\[7\]
rlabel metal1 29486 13362 29486 13362 0 ct.ic.data_chain\[10\]
rlabel metal1 15318 21454 15318 21454 0 ct.ic.data_chain\[11\]
rlabel metal1 19734 21896 19734 21896 0 ct.ic.data_chain\[12\]
rlabel metal1 28842 15538 28842 15538 0 ct.ic.data_chain\[13\]
rlabel metal1 17526 21930 17526 21930 0 ct.ic.data_chain\[14\]
rlabel metal1 27048 21454 27048 21454 0 ct.ic.data_chain\[15\]
rlabel metal1 27922 17170 27922 17170 0 ct.ic.data_chain\[16\]
rlabel metal1 28612 16626 28612 16626 0 ct.ic.data_chain\[17\]
rlabel metal1 26634 19890 26634 19890 0 ct.ic.data_chain\[18\]
rlabel metal2 21114 17221 21114 17221 0 ct.ic.data_chain\[19\]
rlabel metal1 27094 20910 27094 20910 0 ct.ic.data_chain\[20\]
rlabel metal2 23506 19618 23506 19618 0 ct.ic.data_chain\[21\]
rlabel metal1 20930 18904 20930 18904 0 ct.ic.data_chain\[22\]
rlabel metal1 23598 17748 23598 17748 0 ct.ic.data_chain\[23\]
rlabel metal1 20424 18394 20424 18394 0 ct.ic.data_chain\[24\]
rlabel metal1 20930 17306 20930 17306 0 ct.ic.data_chain\[25\]
rlabel metal1 19550 17714 19550 17714 0 ct.ic.data_chain\[26\]
rlabel metal1 19044 18258 19044 18258 0 ct.ic.data_chain\[27\]
rlabel metal1 19090 17170 19090 17170 0 ct.ic.data_chain\[28\]
rlabel metal1 17894 18258 17894 18258 0 ct.ic.data_chain\[29\]
rlabel metal2 18170 19244 18170 19244 0 ct.ic.data_chain\[30\]
rlabel metal1 17848 18938 17848 18938 0 ct.ic.data_chain\[31\]
rlabel metal1 18906 19278 18906 19278 0 ct.ic.data_chain\[32\]
rlabel metal1 16974 19890 16974 19890 0 ct.ic.data_chain\[33\]
rlabel metal1 16238 18802 16238 18802 0 ct.ic.data_chain\[34\]
rlabel metal1 16054 19346 16054 19346 0 ct.ic.data_chain\[35\]
rlabel metal2 25530 13821 25530 13821 0 ct.ic.data_chain\[3\]
rlabel metal1 21942 13940 21942 13940 0 ct.ic.data_chain\[4\]
rlabel metal1 29532 9010 29532 9010 0 ct.ic.data_chain\[5\]
rlabel via2 18538 21403 18538 21403 0 ct.ic.data_chain\[6\]
rlabel via2 14582 18819 14582 18819 0 ct.ic.data_chain\[7\]
rlabel metal2 15962 21760 15962 21760 0 ct.ic.data_chain\[8\]
rlabel metal1 18998 21522 18998 21522 0 ct.ic.data_chain\[9\]
rlabel metal1 27830 21114 27830 21114 0 ct.ic.trig_chain\[0\]
rlabel metal1 17572 18802 17572 18802 0 ct.ic.trig_chain\[10\]
rlabel metal2 14030 19890 14030 19890 0 ct.ic.trig_chain\[11\]
rlabel metal1 15134 20434 15134 20434 0 ct.ic.trig_chain\[12\]
rlabel metal1 21942 13838 21942 13838 0 ct.ic.trig_chain\[1\]
rlabel metal2 19274 14144 19274 14144 0 ct.ic.trig_chain\[2\]
rlabel metal2 16882 21828 16882 21828 0 ct.ic.trig_chain\[3\]
rlabel metal1 19366 21454 19366 21454 0 ct.ic.trig_chain\[4\]
rlabel metal1 27554 17102 27554 17102 0 ct.ic.trig_chain\[5\]
rlabel metal1 23782 18904 23782 18904 0 ct.ic.trig_chain\[6\]
rlabel metal1 21160 19890 21160 19890 0 ct.ic.trig_chain\[7\]
rlabel metal1 20516 18802 20516 18802 0 ct.ic.trig_chain\[8\]
rlabel metal1 18814 18258 18814 18258 0 ct.ic.trig_chain\[9\]
rlabel metal2 12834 18836 12834 18836 0 ct.oc.capture_buffer\[0\]
rlabel metal1 29900 12954 29900 12954 0 ct.oc.capture_buffer\[100\]
rlabel metal1 29854 12886 29854 12886 0 ct.oc.capture_buffer\[101\]
rlabel metal1 28934 19244 28934 19244 0 ct.oc.capture_buffer\[102\]
rlabel metal2 25898 17408 25898 17408 0 ct.oc.capture_buffer\[103\]
rlabel metal1 24978 13294 24978 13294 0 ct.oc.capture_buffer\[104\]
rlabel metal1 24472 14450 24472 14450 0 ct.oc.capture_buffer\[105\]
rlabel metal1 24748 13906 24748 13906 0 ct.oc.capture_buffer\[106\]
rlabel metal1 27278 13294 27278 13294 0 ct.oc.capture_buffer\[107\]
rlabel metal1 30406 15640 30406 15640 0 ct.oc.capture_buffer\[108\]
rlabel metal1 29256 12954 29256 12954 0 ct.oc.capture_buffer\[109\]
rlabel metal1 13800 16218 13800 16218 0 ct.oc.capture_buffer\[10\]
rlabel metal1 29302 13872 29302 13872 0 ct.oc.capture_buffer\[110\]
rlabel metal2 29670 16388 29670 16388 0 ct.oc.capture_buffer\[111\]
rlabel metal1 22908 12954 22908 12954 0 ct.oc.capture_buffer\[112\]
rlabel metal1 24297 12750 24297 12750 0 ct.oc.capture_buffer\[113\]
rlabel via1 24150 13141 24150 13141 0 ct.oc.capture_buffer\[114\]
rlabel metal1 24656 11662 24656 11662 0 ct.oc.capture_buffer\[115\]
rlabel metal1 28750 11866 28750 11866 0 ct.oc.capture_buffer\[116\]
rlabel metal1 27968 12750 27968 12750 0 ct.oc.capture_buffer\[117\]
rlabel metal2 27830 11764 27830 11764 0 ct.oc.capture_buffer\[118\]
rlabel metal1 29256 11186 29256 11186 0 ct.oc.capture_buffer\[119\]
rlabel metal2 9430 18666 9430 18666 0 ct.oc.capture_buffer\[11\]
rlabel metal1 21735 12274 21735 12274 0 ct.oc.capture_buffer\[120\]
rlabel metal1 21574 11730 21574 11730 0 ct.oc.capture_buffer\[121\]
rlabel metal1 21298 12410 21298 12410 0 ct.oc.capture_buffer\[122\]
rlabel metal2 23046 11016 23046 11016 0 ct.oc.capture_buffer\[123\]
rlabel metal1 28106 7310 28106 7310 0 ct.oc.capture_buffer\[124\]
rlabel metal1 29164 6834 29164 6834 0 ct.oc.capture_buffer\[125\]
rlabel metal1 27370 11322 27370 11322 0 ct.oc.capture_buffer\[126\]
rlabel metal2 28474 9316 28474 9316 0 ct.oc.capture_buffer\[127\]
rlabel metal1 19274 11662 19274 11662 0 ct.oc.capture_buffer\[128\]
rlabel metal2 19458 12410 19458 12410 0 ct.oc.capture_buffer\[129\]
rlabel metal2 8970 13583 8970 13583 0 ct.oc.capture_buffer\[12\]
rlabel metal1 19412 13294 19412 13294 0 ct.oc.capture_buffer\[130\]
rlabel metal2 22402 10268 22402 10268 0 ct.oc.capture_buffer\[131\]
rlabel metal1 27600 8398 27600 8398 0 ct.oc.capture_buffer\[132\]
rlabel metal2 28014 10132 28014 10132 0 ct.oc.capture_buffer\[133\]
rlabel metal1 24518 10642 24518 10642 0 ct.oc.capture_buffer\[134\]
rlabel metal1 27692 9622 27692 9622 0 ct.oc.capture_buffer\[135\]
rlabel metal1 16885 11662 16885 11662 0 ct.oc.capture_buffer\[136\]
rlabel metal1 17158 11186 17158 11186 0 ct.oc.capture_buffer\[137\]
rlabel metal1 17848 12274 17848 12274 0 ct.oc.capture_buffer\[138\]
rlabel metal1 20930 9962 20930 9962 0 ct.oc.capture_buffer\[139\]
rlabel metal1 1909 17850 1909 17850 0 ct.oc.capture_buffer\[13\]
rlabel metal1 26864 9010 26864 9010 0 ct.oc.capture_buffer\[140\]
rlabel metal1 26864 9622 26864 9622 0 ct.oc.capture_buffer\[141\]
rlabel metal2 20378 10778 20378 10778 0 ct.oc.capture_buffer\[142\]
rlabel metal2 25714 9316 25714 9316 0 ct.oc.capture_buffer\[143\]
rlabel metal2 18170 8772 18170 8772 0 ct.oc.capture_buffer\[144\]
rlabel metal1 19596 9486 19596 9486 0 ct.oc.capture_buffer\[145\]
rlabel metal1 16284 9622 16284 9622 0 ct.oc.capture_buffer\[146\]
rlabel metal1 20930 9146 20930 9146 0 ct.oc.capture_buffer\[147\]
rlabel metal1 24288 8398 24288 8398 0 ct.oc.capture_buffer\[148\]
rlabel metal1 24518 7378 24518 7378 0 ct.oc.capture_buffer\[149\]
rlabel metal1 10534 13974 10534 13974 0 ct.oc.capture_buffer\[14\]
rlabel metal1 21482 9010 21482 9010 0 ct.oc.capture_buffer\[150\]
rlabel metal1 23920 9010 23920 9010 0 ct.oc.capture_buffer\[151\]
rlabel metal1 18722 7514 18722 7514 0 ct.oc.capture_buffer\[152\]
rlabel metal1 19136 7310 19136 7310 0 ct.oc.capture_buffer\[153\]
rlabel metal1 17802 7412 17802 7412 0 ct.oc.capture_buffer\[154\]
rlabel metal1 19780 6086 19780 6086 0 ct.oc.capture_buffer\[155\]
rlabel via2 22310 8381 22310 8381 0 ct.oc.capture_buffer\[156\]
rlabel metal1 22448 6426 22448 6426 0 ct.oc.capture_buffer\[157\]
rlabel metal1 21620 7922 21620 7922 0 ct.oc.capture_buffer\[158\]
rlabel metal1 23552 7922 23552 7922 0 ct.oc.capture_buffer\[159\]
rlabel metal1 4784 20366 4784 20366 0 ct.oc.capture_buffer\[15\]
rlabel metal1 28750 3502 28750 3502 0 ct.oc.capture_buffer\[160\]
rlabel metal1 28244 5202 28244 5202 0 ct.oc.capture_buffer\[161\]
rlabel metal1 28428 5746 28428 5746 0 ct.oc.capture_buffer\[162\]
rlabel metal1 25300 6834 25300 6834 0 ct.oc.capture_buffer\[163\]
rlabel metal2 28290 6154 28290 6154 0 ct.oc.capture_buffer\[164\]
rlabel metal1 25622 6290 25622 6290 0 ct.oc.capture_buffer\[165\]
rlabel metal1 29118 7446 29118 7446 0 ct.oc.capture_buffer\[166\]
rlabel metal1 27140 6222 27140 6222 0 ct.oc.capture_buffer\[167\]
rlabel metal4 17940 7208 17940 7208 0 ct.oc.capture_buffer\[168\]
rlabel metal2 17802 7327 17802 7327 0 ct.oc.capture_buffer\[169\]
rlabel metal1 9476 13498 9476 13498 0 ct.oc.capture_buffer\[16\]
rlabel metal2 4830 425 4830 425 0 ct.oc.capture_buffer\[170\]
rlabel metal2 20654 6477 20654 6477 0 ct.oc.capture_buffer\[171\]
rlabel metal1 28244 1326 28244 1326 0 ct.oc.capture_buffer\[172\]
rlabel metal1 28290 782 28290 782 0 ct.oc.capture_buffer\[173\]
rlabel metal2 17894 2720 17894 2720 0 ct.oc.capture_buffer\[174\]
rlabel metal2 21574 4794 21574 4794 0 ct.oc.capture_buffer\[175\]
rlabel via2 1702 867 1702 867 0 ct.oc.capture_buffer\[176\]
rlabel via2 1702 1955 1702 1955 0 ct.oc.capture_buffer\[177\]
rlabel metal1 20194 782 20194 782 0 ct.oc.capture_buffer\[178\]
rlabel metal1 27048 1938 27048 1938 0 ct.oc.capture_buffer\[179\]
rlabel metal2 9246 14603 9246 14603 0 ct.oc.capture_buffer\[17\]
rlabel metal1 26910 4114 26910 4114 0 ct.oc.capture_buffer\[180\]
rlabel metal1 26818 2958 26818 2958 0 ct.oc.capture_buffer\[181\]
rlabel via2 2070 1309 2070 1309 0 ct.oc.capture_buffer\[182\]
rlabel metal1 19734 4624 19734 4624 0 ct.oc.capture_buffer\[183\]
rlabel metal1 13662 1258 13662 1258 0 ct.oc.capture_buffer\[184\]
rlabel metal2 17158 612 17158 612 0 ct.oc.capture_buffer\[185\]
rlabel metal1 24702 782 24702 782 0 ct.oc.capture_buffer\[186\]
rlabel metal2 24794 4726 24794 4726 0 ct.oc.capture_buffer\[187\]
rlabel metal1 24702 4658 24702 4658 0 ct.oc.capture_buffer\[188\]
rlabel metal1 24840 5746 24840 5746 0 ct.oc.capture_buffer\[189\]
rlabel metal1 9292 19278 9292 19278 0 ct.oc.capture_buffer\[18\]
rlabel metal1 14766 2482 14766 2482 0 ct.oc.capture_buffer\[190\]
rlabel metal1 25668 2414 25668 2414 0 ct.oc.capture_buffer\[191\]
rlabel metal1 24196 1394 24196 1394 0 ct.oc.capture_buffer\[192\]
rlabel metal1 26266 986 26266 986 0 ct.oc.capture_buffer\[193\]
rlabel metal1 24518 3026 24518 3026 0 ct.oc.capture_buffer\[194\]
rlabel metal1 24288 5134 24288 5134 0 ct.oc.capture_buffer\[195\]
rlabel metal2 22586 5100 22586 5100 0 ct.oc.capture_buffer\[196\]
rlabel metal1 22632 5746 22632 5746 0 ct.oc.capture_buffer\[197\]
rlabel metal1 22632 850 22632 850 0 ct.oc.capture_buffer\[198\]
rlabel metal1 23920 3570 23920 3570 0 ct.oc.capture_buffer\[199\]
rlabel metal1 9706 13498 9706 13498 0 ct.oc.capture_buffer\[19\]
rlabel metal1 12834 18802 12834 18802 0 ct.oc.capture_buffer\[1\]
rlabel metal1 23782 918 23782 918 0 ct.oc.capture_buffer\[200\]
rlabel metal2 22862 1530 22862 1530 0 ct.oc.capture_buffer\[201\]
rlabel metal1 21942 3570 21942 3570 0 ct.oc.capture_buffer\[202\]
rlabel metal1 21022 5882 21022 5882 0 ct.oc.capture_buffer\[203\]
rlabel metal1 21574 5202 21574 5202 0 ct.oc.capture_buffer\[204\]
rlabel metal1 20746 4114 20746 4114 0 ct.oc.capture_buffer\[205\]
rlabel metal1 22908 2074 22908 2074 0 ct.oc.capture_buffer\[206\]
rlabel metal1 21482 2958 21482 2958 0 ct.oc.capture_buffer\[207\]
rlabel metal1 21298 680 21298 680 0 ct.oc.capture_buffer\[208\]
rlabel metal1 19826 1326 19826 1326 0 ct.oc.capture_buffer\[209\]
rlabel metal1 6716 20774 6716 20774 0 ct.oc.capture_buffer\[20\]
rlabel metal1 19228 3570 19228 3570 0 ct.oc.capture_buffer\[210\]
rlabel metal1 18538 5746 18538 5746 0 ct.oc.capture_buffer\[211\]
rlabel metal1 19596 5134 19596 5134 0 ct.oc.capture_buffer\[212\]
rlabel metal1 18998 4658 18998 4658 0 ct.oc.capture_buffer\[213\]
rlabel metal1 20838 1326 20838 1326 0 ct.oc.capture_buffer\[214\]
rlabel metal1 19596 2958 19596 2958 0 ct.oc.capture_buffer\[215\]
rlabel metal1 17434 1326 17434 1326 0 ct.oc.capture_buffer\[216\]
rlabel metal1 16192 986 16192 986 0 ct.oc.capture_buffer\[217\]
rlabel metal1 16790 3570 16790 3570 0 ct.oc.capture_buffer\[218\]
rlabel metal1 17296 4658 17296 4658 0 ct.oc.capture_buffer\[219\]
rlabel metal1 4738 19822 4738 19822 0 ct.oc.capture_buffer\[21\]
rlabel metal1 16928 5746 16928 5746 0 ct.oc.capture_buffer\[220\]
rlabel metal1 17020 5202 17020 5202 0 ct.oc.capture_buffer\[221\]
rlabel metal1 17342 1938 17342 1938 0 ct.oc.capture_buffer\[222\]
rlabel metal1 16514 3026 16514 3026 0 ct.oc.capture_buffer\[223\]
rlabel metal2 14490 2465 14490 2465 0 ct.oc.capture_buffer\[224\]
rlabel metal2 14490 1445 14490 1445 0 ct.oc.capture_buffer\[225\]
rlabel metal1 14030 3570 14030 3570 0 ct.oc.capture_buffer\[226\]
rlabel metal1 14490 5746 14490 5746 0 ct.oc.capture_buffer\[227\]
rlabel metal1 14490 5134 14490 5134 0 ct.oc.capture_buffer\[228\]
rlabel metal1 14536 4658 14536 4658 0 ct.oc.capture_buffer\[229\]
rlabel metal2 3036 12852 3036 12852 0 ct.oc.capture_buffer\[22\]
rlabel metal1 14306 1938 14306 1938 0 ct.oc.capture_buffer\[230\]
rlabel metal1 13202 3094 13202 3094 0 ct.oc.capture_buffer\[231\]
rlabel metal1 8556 2006 8556 2006 0 ct.oc.capture_buffer\[232\]
rlabel metal1 9108 1394 9108 1394 0 ct.oc.capture_buffer\[233\]
rlabel metal1 11684 2958 11684 2958 0 ct.oc.capture_buffer\[234\]
rlabel metal2 12650 5916 12650 5916 0 ct.oc.capture_buffer\[235\]
rlabel metal1 12098 5202 12098 5202 0 ct.oc.capture_buffer\[236\]
rlabel metal2 12374 5372 12374 5372 0 ct.oc.capture_buffer\[237\]
rlabel metal2 5842 544 5842 544 0 ct.oc.capture_buffer\[238\]
rlabel metal1 10350 2584 10350 2584 0 ct.oc.capture_buffer\[239\]
rlabel metal2 7866 14841 7866 14841 0 ct.oc.capture_buffer\[23\]
rlabel metal1 9108 782 9108 782 0 ct.oc.capture_buffer\[240\]
rlabel metal1 6532 782 6532 782 0 ct.oc.capture_buffer\[241\]
rlabel metal1 9752 3026 9752 3026 0 ct.oc.capture_buffer\[242\]
rlabel metal2 9430 5134 9430 5134 0 ct.oc.capture_buffer\[243\]
rlabel metal2 9798 5372 9798 5372 0 ct.oc.capture_buffer\[244\]
rlabel metal1 10580 4114 10580 4114 0 ct.oc.capture_buffer\[245\]
rlabel metal1 4876 918 4876 918 0 ct.oc.capture_buffer\[246\]
rlabel metal1 9384 3570 9384 3570 0 ct.oc.capture_buffer\[247\]
rlabel metal2 14306 612 14306 612 0 ct.oc.capture_buffer\[248\]
rlabel metal4 16652 5848 16652 5848 0 ct.oc.capture_buffer\[249\]
rlabel metal1 13202 16762 13202 16762 0 ct.oc.capture_buffer\[24\]
rlabel metal1 10580 918 10580 918 0 ct.oc.capture_buffer\[250\]
rlabel metal1 7360 2618 7360 2618 0 ct.oc.capture_buffer\[251\]
rlabel metal1 7682 5134 7682 5134 0 ct.oc.capture_buffer\[252\]
rlabel metal1 8510 3910 8510 3910 0 ct.oc.capture_buffer\[253\]
rlabel metal2 7314 2108 7314 2108 0 ct.oc.capture_buffer\[254\]
rlabel metal1 8188 2482 8188 2482 0 ct.oc.capture_buffer\[255\]
rlabel metal1 16560 12954 16560 12954 0 ct.oc.capture_buffer\[256\]
rlabel metal1 9338 6426 9338 6426 0 ct.oc.capture_buffer\[257\]
rlabel metal1 8004 918 8004 918 0 ct.oc.capture_buffer\[258\]
rlabel metal2 6670 4556 6670 4556 0 ct.oc.capture_buffer\[259\]
rlabel via2 13294 17221 13294 17221 0 ct.oc.capture_buffer\[25\]
rlabel metal1 4600 4590 4600 4590 0 ct.oc.capture_buffer\[260\]
rlabel metal1 6348 4046 6348 4046 0 ct.oc.capture_buffer\[261\]
rlabel metal1 8648 6426 8648 6426 0 ct.oc.capture_buffer\[262\]
rlabel metal2 7452 1972 7452 1972 0 ct.oc.capture_buffer\[263\]
rlabel metal2 1702 10829 1702 10829 0 ct.oc.capture_buffer\[264\]
rlabel metal1 2162 13838 2162 13838 0 ct.oc.capture_buffer\[265\]
rlabel via2 1702 20995 1702 20995 0 ct.oc.capture_buffer\[266\]
rlabel metal1 3956 4046 3956 4046 0 ct.oc.capture_buffer\[267\]
rlabel metal1 4830 2958 4830 2958 0 ct.oc.capture_buffer\[268\]
rlabel metal1 2070 3672 2070 3672 0 ct.oc.capture_buffer\[269\]
rlabel via3 6739 18020 6739 18020 0 ct.oc.capture_buffer\[26\]
rlabel via2 1794 9027 1794 9027 0 ct.oc.capture_buffer\[270\]
rlabel metal4 16836 5848 16836 5848 0 ct.oc.capture_buffer\[271\]
rlabel metal1 10028 13838 10028 13838 0 ct.oc.capture_buffer\[272\]
rlabel metal1 2208 4114 2208 4114 0 ct.oc.capture_buffer\[273\]
rlabel metal1 3082 4658 3082 4658 0 ct.oc.capture_buffer\[274\]
rlabel metal2 18722 1955 18722 1955 0 ct.oc.capture_buffer\[275\]
rlabel metal1 15548 986 15548 986 0 ct.oc.capture_buffer\[276\]
rlabel metal1 2024 5134 2024 5134 0 ct.oc.capture_buffer\[277\]
rlabel metal1 9338 8568 9338 8568 0 ct.oc.capture_buffer\[278\]
rlabel metal2 1702 3009 1702 3009 0 ct.oc.capture_buffer\[279\]
rlabel metal1 966 16728 966 16728 0 ct.oc.capture_buffer\[27\]
rlabel metal1 2231 7310 2231 7310 0 ct.oc.capture_buffer\[280\]
rlabel metal1 1058 1530 1058 1530 0 ct.oc.capture_buffer\[281\]
rlabel metal2 2162 2094 2162 2094 0 ct.oc.capture_buffer\[282\]
rlabel metal1 4462 6222 4462 6222 0 ct.oc.capture_buffer\[283\]
rlabel metal1 4646 6834 4646 6834 0 ct.oc.capture_buffer\[284\]
rlabel metal2 6394 6868 6394 6868 0 ct.oc.capture_buffer\[285\]
rlabel metal1 2323 6766 2323 6766 0 ct.oc.capture_buffer\[286\]
rlabel metal1 3496 7310 3496 7310 0 ct.oc.capture_buffer\[287\]
rlabel metal2 9430 8058 9430 8058 0 ct.oc.capture_buffer\[288\]
rlabel metal1 7176 7922 7176 7922 0 ct.oc.capture_buffer\[289\]
rlabel via2 1702 20451 1702 20451 0 ct.oc.capture_buffer\[28\]
rlabel metal1 7314 7378 7314 7378 0 ct.oc.capture_buffer\[290\]
rlabel metal1 8004 6834 8004 6834 0 ct.oc.capture_buffer\[291\]
rlabel metal1 6808 6290 6808 6290 0 ct.oc.capture_buffer\[292\]
rlabel metal1 9936 6222 9936 6222 0 ct.oc.capture_buffer\[293\]
rlabel metal1 9522 7310 9522 7310 0 ct.oc.capture_buffer\[294\]
rlabel metal1 10350 6732 10350 6732 0 ct.oc.capture_buffer\[295\]
rlabel metal1 15778 7514 15778 7514 0 ct.oc.capture_buffer\[296\]
rlabel metal1 15594 6970 15594 6970 0 ct.oc.capture_buffer\[297\]
rlabel metal1 15640 6698 15640 6698 0 ct.oc.capture_buffer\[298\]
rlabel metal2 15410 6732 15410 6732 0 ct.oc.capture_buffer\[299\]
rlabel metal1 11362 13260 11362 13260 0 ct.oc.capture_buffer\[29\]
rlabel metal1 9614 21930 9614 21930 0 ct.oc.capture_buffer\[2\]
rlabel metal1 14858 6936 14858 6936 0 ct.oc.capture_buffer\[300\]
rlabel metal1 13156 6086 13156 6086 0 ct.oc.capture_buffer\[301\]
rlabel metal2 12834 8092 12834 8092 0 ct.oc.capture_buffer\[302\]
rlabel metal2 12926 7684 12926 7684 0 ct.oc.capture_buffer\[303\]
rlabel metal1 14720 10642 14720 10642 0 ct.oc.capture_buffer\[304\]
rlabel metal1 14309 9486 14309 9486 0 ct.oc.capture_buffer\[305\]
rlabel metal1 14398 8466 14398 8466 0 ct.oc.capture_buffer\[306\]
rlabel metal1 14674 9010 14674 9010 0 ct.oc.capture_buffer\[307\]
rlabel metal2 14582 9962 14582 9962 0 ct.oc.capture_buffer\[308\]
rlabel metal1 10994 8806 10994 8806 0 ct.oc.capture_buffer\[309\]
rlabel metal1 17112 15674 17112 15674 0 ct.oc.capture_buffer\[30\]
rlabel metal1 11592 9010 11592 9010 0 ct.oc.capture_buffer\[310\]
rlabel metal1 12052 8602 12052 8602 0 ct.oc.capture_buffer\[311\]
rlabel metal1 13248 12274 13248 12274 0 ct.oc.capture_buffer\[312\]
rlabel metal2 13294 12682 13294 12682 0 ct.oc.capture_buffer\[313\]
rlabel metal1 13984 12750 13984 12750 0 ct.oc.capture_buffer\[314\]
rlabel metal1 14214 11662 14214 11662 0 ct.oc.capture_buffer\[315\]
rlabel metal1 13018 12614 13018 12614 0 ct.oc.capture_buffer\[316\]
rlabel metal1 9890 9146 9890 9146 0 ct.oc.capture_buffer\[317\]
rlabel metal1 10856 8466 10856 8466 0 ct.oc.capture_buffer\[318\]
rlabel metal1 10028 10098 10028 10098 0 ct.oc.capture_buffer\[319\]
rlabel metal2 1702 19601 1702 19601 0 ct.oc.capture_buffer\[31\]
rlabel viali 10350 12817 10350 12817 0 ct.oc.capture_buffer\[320\]
rlabel metal1 10672 10642 10672 10642 0 ct.oc.capture_buffer\[321\]
rlabel metal1 10028 11186 10028 11186 0 ct.oc.capture_buffer\[322\]
rlabel metal1 9384 12274 9384 12274 0 ct.oc.capture_buffer\[323\]
rlabel metal1 10166 13158 10166 13158 0 ct.oc.capture_buffer\[324\]
rlabel metal1 8096 9010 8096 9010 0 ct.oc.capture_buffer\[325\]
rlabel metal2 6854 9537 6854 9537 0 ct.oc.capture_buffer\[326\]
rlabel metal2 8418 9316 8418 9316 0 ct.oc.capture_buffer\[327\]
rlabel metal1 6903 12274 6903 12274 0 ct.oc.capture_buffer\[328\]
rlabel metal1 6808 13498 6808 13498 0 ct.oc.capture_buffer\[329\]
rlabel metal1 4876 17102 4876 17102 0 ct.oc.capture_buffer\[32\]
rlabel metal1 8464 12886 8464 12886 0 ct.oc.capture_buffer\[330\]
rlabel metal1 8142 12954 8142 12954 0 ct.oc.capture_buffer\[331\]
rlabel metal1 6808 12818 6808 12818 0 ct.oc.capture_buffer\[332\]
rlabel metal1 6256 10574 6256 10574 0 ct.oc.capture_buffer\[333\]
rlabel metal1 6256 8466 6256 8466 0 ct.oc.capture_buffer\[334\]
rlabel metal1 6302 6970 6302 6970 0 ct.oc.capture_buffer\[335\]
rlabel metal1 5060 13294 5060 13294 0 ct.oc.capture_buffer\[336\]
rlabel metal1 5658 13158 5658 13158 0 ct.oc.capture_buffer\[337\]
rlabel metal1 4646 13838 4646 13838 0 ct.oc.capture_buffer\[338\]
rlabel metal2 4646 13362 4646 13362 0 ct.oc.capture_buffer\[339\]
rlabel metal2 4738 8347 4738 8347 0 ct.oc.capture_buffer\[33\]
rlabel metal1 4278 14246 4278 14246 0 ct.oc.capture_buffer\[340\]
rlabel metal1 3864 9486 3864 9486 0 ct.oc.capture_buffer\[341\]
rlabel metal1 3910 10098 3910 10098 0 ct.oc.capture_buffer\[342\]
rlabel metal1 3910 9010 3910 9010 0 ct.oc.capture_buffer\[343\]
rlabel metal1 1472 6630 1472 6630 0 ct.oc.capture_buffer\[344\]
rlabel metal1 2208 11186 2208 11186 0 ct.oc.capture_buffer\[345\]
rlabel metal1 3358 12954 3358 12954 0 ct.oc.capture_buffer\[346\]
rlabel metal2 3266 13226 3266 13226 0 ct.oc.capture_buffer\[347\]
rlabel metal1 2116 12206 2116 12206 0 ct.oc.capture_buffer\[348\]
rlabel metal1 1380 5882 1380 5882 0 ct.oc.capture_buffer\[349\]
rlabel metal4 5428 15980 5428 15980 0 ct.oc.capture_buffer\[34\]
rlabel metal1 828 2618 828 2618 0 ct.oc.capture_buffer\[350\]
rlabel metal1 1656 3434 1656 3434 0 ct.oc.capture_buffer\[351\]
rlabel metal1 1909 13158 1909 13158 0 ct.oc.capture_buffer\[35\]
rlabel via2 7958 13141 7958 13141 0 ct.oc.capture_buffer\[36\]
rlabel metal2 2070 17034 2070 17034 0 ct.oc.capture_buffer\[37\]
rlabel metal2 2162 17629 2162 17629 0 ct.oc.capture_buffer\[38\]
rlabel metal1 16376 15334 16376 15334 0 ct.oc.capture_buffer\[39\]
rlabel metal1 10810 15062 10810 15062 0 ct.oc.capture_buffer\[3\]
rlabel metal2 4462 14807 4462 14807 0 ct.oc.capture_buffer\[40\]
rlabel metal1 4646 14586 4646 14586 0 ct.oc.capture_buffer\[41\]
rlabel metal1 966 14348 966 14348 0 ct.oc.capture_buffer\[42\]
rlabel metal2 5014 15300 5014 15300 0 ct.oc.capture_buffer\[43\]
rlabel metal1 1288 13498 1288 13498 0 ct.oc.capture_buffer\[44\]
rlabel via2 2070 15453 2070 15453 0 ct.oc.capture_buffer\[45\]
rlabel metal1 1932 16558 1932 16558 0 ct.oc.capture_buffer\[46\]
rlabel metal1 1104 16082 1104 16082 0 ct.oc.capture_buffer\[47\]
rlabel metal1 6624 13838 6624 13838 0 ct.oc.capture_buffer\[48\]
rlabel metal1 6211 14586 6211 14586 0 ct.oc.capture_buffer\[49\]
rlabel metal3 10373 19380 10373 19380 0 ct.oc.capture_buffer\[4\]
rlabel metal2 6394 14756 6394 14756 0 ct.oc.capture_buffer\[50\]
rlabel metal2 5474 15266 5474 15266 0 ct.oc.capture_buffer\[51\]
rlabel metal1 9384 14586 9384 14586 0 ct.oc.capture_buffer\[52\]
rlabel metal1 9292 16082 9292 16082 0 ct.oc.capture_buffer\[53\]
rlabel metal2 9706 14756 9706 14756 0 ct.oc.capture_buffer\[54\]
rlabel metal2 9982 15606 9982 15606 0 ct.oc.capture_buffer\[55\]
rlabel metal1 11178 14586 11178 14586 0 ct.oc.capture_buffer\[56\]
rlabel metal1 12236 13498 12236 13498 0 ct.oc.capture_buffer\[57\]
rlabel metal1 11684 13838 11684 13838 0 ct.oc.capture_buffer\[58\]
rlabel metal1 12144 13158 12144 13158 0 ct.oc.capture_buffer\[59\]
rlabel metal3 10143 21012 10143 21012 0 ct.oc.capture_buffer\[5\]
rlabel metal1 11960 17646 11960 17646 0 ct.oc.capture_buffer\[60\]
rlabel metal1 11684 16014 11684 16014 0 ct.oc.capture_buffer\[61\]
rlabel metal2 12006 16864 12006 16864 0 ct.oc.capture_buffer\[62\]
rlabel metal1 8602 16966 8602 16966 0 ct.oc.capture_buffer\[63\]
rlabel metal2 13662 14416 13662 14416 0 ct.oc.capture_buffer\[64\]
rlabel metal2 16146 12818 16146 12818 0 ct.oc.capture_buffer\[65\]
rlabel metal1 14720 13838 14720 13838 0 ct.oc.capture_buffer\[66\]
rlabel metal1 14674 13498 14674 13498 0 ct.oc.capture_buffer\[67\]
rlabel metal1 14904 16626 14904 16626 0 ct.oc.capture_buffer\[68\]
rlabel metal1 14904 16218 14904 16218 0 ct.oc.capture_buffer\[69\]
rlabel metal3 6095 16660 6095 16660 0 ct.oc.capture_buffer\[6\]
rlabel metal1 14996 15470 14996 15470 0 ct.oc.capture_buffer\[70\]
rlabel metal2 16698 17204 16698 17204 0 ct.oc.capture_buffer\[71\]
rlabel metal1 17940 13906 17940 13906 0 ct.oc.capture_buffer\[72\]
rlabel metal1 18952 13974 18952 13974 0 ct.oc.capture_buffer\[73\]
rlabel metal1 18124 12954 18124 12954 0 ct.oc.capture_buffer\[74\]
rlabel metal1 18630 14382 18630 14382 0 ct.oc.capture_buffer\[75\]
rlabel metal1 17342 16218 17342 16218 0 ct.oc.capture_buffer\[76\]
rlabel metal1 19136 16014 19136 16014 0 ct.oc.capture_buffer\[77\]
rlabel metal1 17848 16218 17848 16218 0 ct.oc.capture_buffer\[78\]
rlabel metal1 18676 15130 18676 15130 0 ct.oc.capture_buffer\[79\]
rlabel metal2 15870 13158 15870 13158 0 ct.oc.capture_buffer\[7\]
rlabel metal1 21666 14450 21666 14450 0 ct.oc.capture_buffer\[80\]
rlabel metal1 20746 15130 20746 15130 0 ct.oc.capture_buffer\[81\]
rlabel metal1 20332 13838 20332 13838 0 ct.oc.capture_buffer\[82\]
rlabel metal1 20470 14586 20470 14586 0 ct.oc.capture_buffer\[83\]
rlabel metal1 21735 18258 21735 18258 0 ct.oc.capture_buffer\[84\]
rlabel metal1 23506 17612 23506 17612 0 ct.oc.capture_buffer\[85\]
rlabel metal1 23230 16694 23230 16694 0 ct.oc.capture_buffer\[86\]
rlabel metal1 21735 17170 21735 17170 0 ct.oc.capture_buffer\[87\]
rlabel metal2 22494 15249 22494 15249 0 ct.oc.capture_buffer\[88\]
rlabel metal1 22586 15130 22586 15130 0 ct.oc.capture_buffer\[89\]
rlabel metal1 3910 19142 3910 19142 0 ct.oc.capture_buffer\[8\]
rlabel metal1 24472 14926 24472 14926 0 ct.oc.capture_buffer\[90\]
rlabel metal1 23644 15130 23644 15130 0 ct.oc.capture_buffer\[91\]
rlabel metal2 24886 17833 24886 17833 0 ct.oc.capture_buffer\[92\]
rlabel metal1 27094 16558 27094 16558 0 ct.oc.capture_buffer\[93\]
rlabel metal1 25576 17170 25576 17170 0 ct.oc.capture_buffer\[94\]
rlabel metal1 28382 18088 28382 18088 0 ct.oc.capture_buffer\[95\]
rlabel metal1 27094 15538 27094 15538 0 ct.oc.capture_buffer\[96\]
rlabel metal1 29210 15130 29210 15130 0 ct.oc.capture_buffer\[97\]
rlabel metal1 29376 16081 29376 16081 0 ct.oc.capture_buffer\[98\]
rlabel metal2 30406 11713 30406 11713 0 ct.oc.capture_buffer\[99\]
rlabel metal1 9016 16762 9016 16762 0 ct.oc.capture_buffer\[9\]
rlabel metal1 13984 18190 13984 18190 0 ct.oc.data_chain\[0\]
rlabel viali 24611 17648 24611 17648 0 ct.oc.data_chain\[100\]
rlabel metal1 26913 16593 26913 16593 0 ct.oc.data_chain\[101\]
rlabel via1 25347 17170 25347 17170 0 ct.oc.data_chain\[102\]
rlabel metal1 25691 18258 25691 18258 0 ct.oc.data_chain\[103\]
rlabel metal1 26542 13498 26542 13498 0 ct.oc.data_chain\[104\]
rlabel metal1 26359 14994 26359 14994 0 ct.oc.data_chain\[105\]
rlabel metal1 26451 16082 26451 16082 0 ct.oc.data_chain\[106\]
rlabel metal2 22034 15487 22034 15487 0 ct.oc.data_chain\[107\]
rlabel metal1 28957 20910 28957 20910 0 ct.oc.data_chain\[108\]
rlabel metal1 28267 20434 28267 20434 0 ct.oc.data_chain\[109\]
rlabel metal1 11363 21522 11363 21522 0 ct.oc.data_chain\[10\]
rlabel metal1 27301 19346 27301 19346 0 ct.oc.data_chain\[110\]
rlabel metal1 24725 18734 24725 18734 0 ct.oc.data_chain\[111\]
rlabel metal1 24496 13312 24496 13312 0 ct.oc.data_chain\[112\]
rlabel via1 24519 14382 24519 14382 0 ct.oc.data_chain\[113\]
rlabel via1 24610 13905 24610 13905 0 ct.oc.data_chain\[114\]
rlabel metal1 26542 11866 26542 11866 0 ct.oc.data_chain\[115\]
rlabel metal1 28957 17646 28957 17646 0 ct.oc.data_chain\[116\]
rlabel metal1 28842 12954 28842 12954 0 ct.oc.data_chain\[117\]
rlabel metal1 27301 13906 27301 13906 0 ct.oc.data_chain\[118\]
rlabel metal2 27968 15300 27968 15300 0 ct.oc.data_chain\[119\]
rlabel metal1 11317 20434 11317 20434 0 ct.oc.data_chain\[11\]
rlabel via1 22471 13294 22471 13294 0 ct.oc.data_chain\[120\]
rlabel metal1 23645 12818 23645 12818 0 ct.oc.data_chain\[121\]
rlabel metal1 23875 12206 23875 12206 0 ct.oc.data_chain\[122\]
rlabel metal1 25047 11730 25047 11730 0 ct.oc.data_chain\[123\]
rlabel metal1 28681 14382 28681 14382 0 ct.oc.data_chain\[124\]
rlabel metal1 29210 12818 29210 12818 0 ct.oc.data_chain\[125\]
rlabel via1 26911 12206 26911 12206 0 ct.oc.data_chain\[126\]
rlabel metal1 29095 11118 29095 11118 0 ct.oc.data_chain\[127\]
rlabel metal1 21252 11866 21252 11866 0 ct.oc.data_chain\[128\]
rlabel metal1 21115 11730 21115 11730 0 ct.oc.data_chain\[129\]
rlabel via1 8971 19822 8971 19822 0 ct.oc.data_chain\[12\]
rlabel metal1 20885 12818 20885 12818 0 ct.oc.data_chain\[130\]
rlabel metal1 23644 10234 23644 10234 0 ct.oc.data_chain\[131\]
rlabel metal1 27531 7378 27531 7378 0 ct.oc.data_chain\[132\]
rlabel metal1 28313 6766 28313 6766 0 ct.oc.data_chain\[133\]
rlabel metal1 26451 11730 26451 11730 0 ct.oc.data_chain\[134\]
rlabel metal1 28244 9894 28244 9894 0 ct.oc.data_chain\[135\]
rlabel metal1 18861 11730 18861 11730 0 ct.oc.data_chain\[136\]
rlabel metal1 18953 12818 18953 12818 0 ct.oc.data_chain\[137\]
rlabel via1 18815 13294 18815 13294 0 ct.oc.data_chain\[138\]
rlabel metal1 21873 10030 21873 10030 0 ct.oc.data_chain\[139\]
rlabel metal1 8142 19754 8142 19754 0 ct.oc.data_chain\[13\]
rlabel metal1 27577 8466 27577 8466 0 ct.oc.data_chain\[140\]
rlabel metal1 26729 10605 26729 10605 0 ct.oc.data_chain\[141\]
rlabel metal1 24059 10642 24059 10642 0 ct.oc.data_chain\[142\]
rlabel metal1 26772 9690 26772 9690 0 ct.oc.data_chain\[143\]
rlabel metal1 17503 11730 17503 11730 0 ct.oc.data_chain\[144\]
rlabel metal1 18193 11118 18193 11118 0 ct.oc.data_chain\[145\]
rlabel viali 17435 12208 17435 12208 0 ct.oc.data_chain\[146\]
rlabel metal1 21045 10642 21045 10642 0 ct.oc.data_chain\[147\]
rlabel metal1 26404 8602 26404 8602 0 ct.oc.data_chain\[148\]
rlabel metal1 24725 10030 24725 10030 0 ct.oc.data_chain\[149\]
rlabel metal2 6716 19142 6716 19142 0 ct.oc.data_chain\[14\]
rlabel metal1 21942 11152 21942 11152 0 ct.oc.data_chain\[150\]
rlabel metal1 25185 9554 25185 9554 0 ct.oc.data_chain\[151\]
rlabel metal1 18009 8942 18009 8942 0 ct.oc.data_chain\[152\]
rlabel metal1 19987 9554 19987 9554 0 ct.oc.data_chain\[153\]
rlabel metal1 18607 10030 18607 10030 0 ct.oc.data_chain\[154\]
rlabel metal2 22770 8534 22770 8534 0 ct.oc.data_chain\[155\]
rlabel metal1 24013 8466 24013 8466 0 ct.oc.data_chain\[156\]
rlabel metal1 24197 7378 24197 7378 0 ct.oc.data_chain\[157\]
rlabel metal2 22678 8500 22678 8500 0 ct.oc.data_chain\[158\]
rlabel metal1 24679 8942 24679 8942 0 ct.oc.data_chain\[159\]
rlabel viali 8889 21504 8889 21504 0 ct.oc.data_chain\[15\]
rlabel metal2 18998 7565 18998 7565 0 ct.oc.data_chain\[160\]
rlabel metal1 20654 7446 20654 7446 0 ct.oc.data_chain\[161\]
rlabel metal2 21574 6273 21574 6273 0 ct.oc.data_chain\[162\]
rlabel metal1 23966 7344 23966 7344 0 ct.oc.data_chain\[163\]
rlabel metal1 29394 4488 29394 4488 0 ct.oc.data_chain\[164\]
rlabel metal1 22425 6766 22425 6766 0 ct.oc.data_chain\[165\]
rlabel metal2 30038 2890 30038 2890 0 ct.oc.data_chain\[166\]
rlabel metal1 25047 7854 25047 7854 0 ct.oc.data_chain\[167\]
rlabel metal2 18538 9707 18538 9707 0 ct.oc.data_chain\[168\]
rlabel metal2 19734 8381 19734 8381 0 ct.oc.data_chain\[169\]
rlabel metal2 10810 19278 10810 19278 0 ct.oc.data_chain\[16\]
rlabel metal2 13294 3111 13294 3111 0 ct.oc.data_chain\[170\]
rlabel metal1 24568 6766 24568 6766 0 ct.oc.data_chain\[171\]
rlabel metal1 29210 1530 29210 1530 0 ct.oc.data_chain\[172\]
rlabel metal1 25714 1326 25714 1326 0 ct.oc.data_chain\[173\]
rlabel metal1 28291 2414 28291 2414 0 ct.oc.data_chain\[174\]
rlabel metal2 18814 6477 18814 6477 0 ct.oc.data_chain\[175\]
rlabel via2 16606 10659 16606 10659 0 ct.oc.data_chain\[176\]
rlabel via2 16606 9571 16606 9571 0 ct.oc.data_chain\[177\]
rlabel metal2 18354 374 18354 374 0 ct.oc.data_chain\[178\]
rlabel metal2 21666 4488 21666 4488 0 ct.oc.data_chain\[179\]
rlabel metal1 11179 19346 11179 19346 0 ct.oc.data_chain\[17\]
rlabel metal1 28060 1326 28060 1326 0 ct.oc.data_chain\[180\]
rlabel metal1 27439 850 27439 850 0 ct.oc.data_chain\[181\]
rlabel metal1 3634 1530 3634 1530 0 ct.oc.data_chain\[182\]
rlabel via1 17251 6766 17251 6766 0 ct.oc.data_chain\[183\]
rlabel metal1 1610 340 1610 340 0 ct.oc.data_chain\[184\]
rlabel metal2 1518 1343 1518 1343 0 ct.oc.data_chain\[185\]
rlabel metal1 20746 918 20746 918 0 ct.oc.data_chain\[186\]
rlabel metal1 26589 1938 26589 1938 0 ct.oc.data_chain\[187\]
rlabel metal1 26405 4114 26405 4114 0 ct.oc.data_chain\[188\]
rlabel metal1 26451 3026 26451 3026 0 ct.oc.data_chain\[189\]
rlabel metal1 9637 20434 9637 20434 0 ct.oc.data_chain\[18\]
rlabel metal1 2162 1360 2162 1360 0 ct.oc.data_chain\[190\]
rlabel metal2 16974 3638 16974 3638 0 ct.oc.data_chain\[191\]
rlabel metal2 12190 833 12190 833 0 ct.oc.data_chain\[192\]
rlabel metal1 16882 408 16882 408 0 ct.oc.data_chain\[193\]
rlabel via1 24679 850 24679 850 0 ct.oc.data_chain\[194\]
rlabel metal1 24633 4114 24633 4114 0 ct.oc.data_chain\[195\]
rlabel viali 24519 4592 24519 4592 0 ct.oc.data_chain\[196\]
rlabel metal1 24335 5678 24335 5678 0 ct.oc.data_chain\[197\]
rlabel via2 15134 3043 15134 3043 0 ct.oc.data_chain\[198\]
rlabel metal1 25070 2482 25070 2482 0 ct.oc.data_chain\[199\]
rlabel metal1 9269 18734 9269 18734 0 ct.oc.data_chain\[19\]
rlabel metal1 13754 21386 13754 21386 0 ct.oc.data_chain\[1\]
rlabel metal1 23783 1326 23783 1326 0 ct.oc.data_chain\[200\]
rlabel metal1 24289 1938 24289 1938 0 ct.oc.data_chain\[201\]
rlabel metal1 23829 3026 23829 3026 0 ct.oc.data_chain\[202\]
rlabel metal1 24197 5202 24197 5202 0 ct.oc.data_chain\[203\]
rlabel metal1 22425 4590 22425 4590 0 ct.oc.data_chain\[204\]
rlabel metal2 22402 4896 22402 4896 0 ct.oc.data_chain\[205\]
rlabel metal1 22149 850 22149 850 0 ct.oc.data_chain\[206\]
rlabel metal1 23414 3094 23414 3094 0 ct.oc.data_chain\[207\]
rlabel metal1 21207 1938 21207 1938 0 ct.oc.data_chain\[208\]
rlabel viali 21761 1335 21761 1335 0 ct.oc.data_chain\[209\]
rlabel metal1 6211 20910 6211 20910 0 ct.oc.data_chain\[20\]
rlabel metal1 21575 3502 21575 3502 0 ct.oc.data_chain\[210\]
rlabel metal1 20425 6290 20425 6290 0 ct.oc.data_chain\[211\]
rlabel metal1 21115 5202 21115 5202 0 ct.oc.data_chain\[212\]
rlabel via1 20379 4114 20379 4114 0 ct.oc.data_chain\[213\]
rlabel viali 21785 2432 21785 2432 0 ct.oc.data_chain\[214\]
rlabel metal1 21115 3026 21115 3026 0 ct.oc.data_chain\[215\]
rlabel metal1 18999 1938 18999 1938 0 ct.oc.data_chain\[216\]
rlabel via1 18815 1326 18815 1326 0 ct.oc.data_chain\[217\]
rlabel viali 18815 3502 18815 3502 0 ct.oc.data_chain\[218\]
rlabel metal1 18446 4794 18446 4794 0 ct.oc.data_chain\[219\]
rlabel metal1 6257 19824 6257 19824 0 ct.oc.data_chain\[21\]
rlabel metal1 18677 5202 18677 5202 0 ct.oc.data_chain\[220\]
rlabel metal1 18769 4590 18769 4590 0 ct.oc.data_chain\[221\]
rlabel metal1 17940 2074 17940 2074 0 ct.oc.data_chain\[222\]
rlabel metal1 18585 3026 18585 3026 0 ct.oc.data_chain\[223\]
rlabel metal1 16285 1326 16285 1326 0 ct.oc.data_chain\[224\]
rlabel metal1 15916 1530 15916 1530 0 ct.oc.data_chain\[225\]
rlabel metal1 16609 3537 16609 3537 0 ct.oc.data_chain\[226\]
rlabel metal1 16515 4590 16515 4590 0 ct.oc.data_chain\[227\]
rlabel metal1 16192 5338 16192 5338 0 ct.oc.data_chain\[228\]
rlabel metal1 16239 5202 16239 5202 0 ct.oc.data_chain\[229\]
rlabel metal1 5613 19346 5613 19346 0 ct.oc.data_chain\[22\]
rlabel metal1 16055 1938 16055 1938 0 ct.oc.data_chain\[230\]
rlabel metal1 16193 3026 16193 3026 0 ct.oc.data_chain\[231\]
rlabel viali 14260 2415 14260 2415 0 ct.oc.data_chain\[232\]
rlabel metal1 14031 1326 14031 1326 0 ct.oc.data_chain\[233\]
rlabel metal1 13800 3162 13800 3162 0 ct.oc.data_chain\[234\]
rlabel viali 14307 5678 14307 5678 0 ct.oc.data_chain\[235\]
rlabel metal1 13755 5202 13755 5202 0 ct.oc.data_chain\[236\]
rlabel viali 14307 4590 14307 4590 0 ct.oc.data_chain\[237\]
rlabel metal1 13755 1938 13755 1938 0 ct.oc.data_chain\[238\]
rlabel metal1 14309 4079 14309 4079 0 ct.oc.data_chain\[239\]
rlabel metal1 5359 20434 5359 20434 0 ct.oc.data_chain\[23\]
rlabel metal1 10902 986 10902 986 0 ct.oc.data_chain\[240\]
rlabel metal1 8648 986 8648 986 0 ct.oc.data_chain\[241\]
rlabel metal1 11455 3026 11455 3026 0 ct.oc.data_chain\[242\]
rlabel metal1 11086 4794 11086 4794 0 ct.oc.data_chain\[243\]
rlabel metal1 11455 5202 11455 5202 0 ct.oc.data_chain\[244\]
rlabel metal1 12052 4250 12052 4250 0 ct.oc.data_chain\[245\]
rlabel metal1 11455 1938 11455 1938 0 ct.oc.data_chain\[246\]
rlabel metal1 12101 3537 12101 3537 0 ct.oc.data_chain\[247\]
rlabel metal1 11086 748 11086 748 0 ct.oc.data_chain\[248\]
rlabel metal1 5751 850 5751 850 0 ct.oc.data_chain\[249\]
rlabel metal1 9157 17681 9157 17681 0 ct.oc.data_chain\[24\]
rlabel metal1 9477 3026 9477 3026 0 ct.oc.data_chain\[250\]
rlabel viali 9155 4590 9155 4590 0 ct.oc.data_chain\[251\]
rlabel viali 9525 5201 9525 5201 0 ct.oc.data_chain\[252\]
rlabel metal1 10213 4114 10213 4114 0 ct.oc.data_chain\[253\]
rlabel viali 9526 1936 9526 1936 0 ct.oc.data_chain\[254\]
rlabel metal1 9499 3502 9499 3502 0 ct.oc.data_chain\[255\]
rlabel via1 14099 850 14099 850 0 ct.oc.data_chain\[256\]
rlabel metal2 1886 2465 1886 2465 0 ct.oc.data_chain\[257\]
rlabel viali 6581 3017 6581 3017 0 ct.oc.data_chain\[258\]
rlabel metal1 7061 4590 7061 4590 0 ct.oc.data_chain\[259\]
rlabel via1 9063 18258 9063 18258 0 ct.oc.data_chain\[25\]
rlabel metal1 6441 5202 6441 5202 0 ct.oc.data_chain\[260\]
rlabel metal1 8234 4114 8234 4114 0 ct.oc.data_chain\[261\]
rlabel metal1 6992 1326 6992 1326 0 ct.oc.data_chain\[262\]
rlabel metal1 8050 2074 8050 2074 0 ct.oc.data_chain\[263\]
rlabel via2 16606 13277 16606 13277 0 ct.oc.data_chain\[264\]
rlabel metal2 15226 13311 15226 13311 0 ct.oc.data_chain\[265\]
rlabel via3 3979 2380 3979 2380 0 ct.oc.data_chain\[266\]
rlabel metal1 6509 3502 6509 3502 0 ct.oc.data_chain\[267\]
rlabel metal1 4117 4590 4117 4590 0 ct.oc.data_chain\[268\]
rlabel metal1 5981 4114 5981 4114 0 ct.oc.data_chain\[269\]
rlabel metal1 8741 19346 8741 19346 0 ct.oc.data_chain\[26\]
rlabel metal1 3451 10642 3451 10642 0 ct.oc.data_chain\[270\]
rlabel viali 6305 1937 6305 1937 0 ct.oc.data_chain\[271\]
rlabel metal1 10350 13906 10350 13906 0 ct.oc.data_chain\[272\]
rlabel metal2 2346 13175 2346 13175 0 ct.oc.data_chain\[273\]
rlabel metal2 1932 16388 1932 16388 0 ct.oc.data_chain\[274\]
rlabel metal1 3681 4114 3681 4114 0 ct.oc.data_chain\[275\]
rlabel metal1 4439 3026 4439 3026 0 ct.oc.data_chain\[276\]
rlabel metal1 3937 5202 3937 5202 0 ct.oc.data_chain\[277\]
rlabel metal1 2162 8942 2162 8942 0 ct.oc.data_chain\[278\]
rlabel metal2 4048 1292 4048 1292 0 ct.oc.data_chain\[279\]
rlabel viali 9200 17169 9200 17169 0 ct.oc.data_chain\[27\]
rlabel metal1 8833 13906 8833 13906 0 ct.oc.data_chain\[280\]
rlabel metal2 1518 5916 1518 5916 0 ct.oc.data_chain\[281\]
rlabel metal1 1978 4624 1978 4624 0 ct.oc.data_chain\[282\]
rlabel metal1 1978 5712 1978 5712 0 ct.oc.data_chain\[283\]
rlabel metal1 3358 6358 3358 6358 0 ct.oc.data_chain\[284\]
rlabel metal1 2047 5202 2047 5202 0 ct.oc.data_chain\[285\]
rlabel viali 3729 8457 3729 8457 0 ct.oc.data_chain\[286\]
rlabel viali 1472 3017 1472 3017 0 ct.oc.data_chain\[287\]
rlabel metal2 2162 7174 2162 7174 0 ct.oc.data_chain\[288\]
rlabel metal1 1817 7854 1817 7854 0 ct.oc.data_chain\[289\]
rlabel metal1 3312 20570 3312 20570 0 ct.oc.data_chain\[28\]
rlabel metal1 2001 8466 2001 8466 0 ct.oc.data_chain\[290\]
rlabel metal1 4991 6290 4991 6290 0 ct.oc.data_chain\[291\]
rlabel metal1 5083 6766 5083 6766 0 ct.oc.data_chain\[292\]
rlabel metal1 4117 7854 4117 7854 0 ct.oc.data_chain\[293\]
rlabel metal2 1794 7021 1794 7021 0 ct.oc.data_chain\[294\]
rlabel metal1 4991 7378 4991 7378 0 ct.oc.data_chain\[295\]
rlabel via2 15686 7803 15686 7803 0 ct.oc.data_chain\[296\]
rlabel metal3 15916 7888 15916 7888 0 ct.oc.data_chain\[297\]
rlabel metal2 16330 8109 16330 8109 0 ct.oc.data_chain\[298\]
rlabel metal3 16468 6664 16468 6664 0 ct.oc.data_chain\[299\]
rlabel metal1 3542 18394 3542 18394 0 ct.oc.data_chain\[29\]
rlabel metal2 13018 20944 13018 20944 0 ct.oc.data_chain\[2\]
rlabel metal2 17986 7497 17986 7497 0 ct.oc.data_chain\[300\]
rlabel metal2 12650 6732 12650 6732 0 ct.oc.data_chain\[301\]
rlabel metal2 13478 7616 13478 7616 0 ct.oc.data_chain\[302\]
rlabel metal1 9338 6800 9338 6800 0 ct.oc.data_chain\[303\]
rlabel metal1 14421 7854 14421 7854 0 ct.oc.data_chain\[304\]
rlabel metal1 15341 7378 15341 7378 0 ct.oc.data_chain\[305\]
rlabel metal1 16147 8466 16147 8466 0 ct.oc.data_chain\[306\]
rlabel via1 15135 6290 15135 6290 0 ct.oc.data_chain\[307\]
rlabel metal1 16330 10030 16330 10030 0 ct.oc.data_chain\[308\]
rlabel metal2 12374 8636 12374 8636 0 ct.oc.data_chain\[309\]
rlabel metal1 3405 21522 3405 21522 0 ct.oc.data_chain\[30\]
rlabel metal2 12742 8330 12742 8330 0 ct.oc.data_chain\[310\]
rlabel metal1 12857 6766 12857 6766 0 ct.oc.data_chain\[311\]
rlabel metal1 14513 10642 14513 10642 0 ct.oc.data_chain\[312\]
rlabel metal2 14398 12789 14398 12789 0 ct.oc.data_chain\[313\]
rlabel via1 14215 8466 14215 8466 0 ct.oc.data_chain\[314\]
rlabel metal1 14605 8942 14605 8942 0 ct.oc.data_chain\[315\]
rlabel metal1 14031 10030 14031 10030 0 ct.oc.data_chain\[316\]
rlabel metal1 11040 9622 11040 9622 0 ct.oc.data_chain\[317\]
rlabel viali 11639 8944 11639 8944 0 ct.oc.data_chain\[318\]
rlabel metal1 11363 9554 11363 9554 0 ct.oc.data_chain\[319\]
rlabel metal1 5199 21522 5199 21522 0 ct.oc.data_chain\[31\]
rlabel metal1 12973 12224 12973 12224 0 ct.oc.data_chain\[320\]
rlabel metal1 11684 10710 11684 10710 0 ct.oc.data_chain\[321\]
rlabel metal1 13985 12818 13985 12818 0 ct.oc.data_chain\[322\]
rlabel viali 14033 11721 14033 11721 0 ct.oc.data_chain\[323\]
rlabel metal1 12927 11118 12927 11118 0 ct.oc.data_chain\[324\]
rlabel metal1 9495 9554 9495 9554 0 ct.oc.data_chain\[325\]
rlabel metal1 9200 8262 9200 8262 0 ct.oc.data_chain\[326\]
rlabel metal1 9157 10065 9157 10065 0 ct.oc.data_chain\[327\]
rlabel metal1 9937 12818 9937 12818 0 ct.oc.data_chain\[328\]
rlabel metal2 10074 12444 10074 12444 0 ct.oc.data_chain\[329\]
rlabel metal1 6440 17306 6440 17306 0 ct.oc.data_chain\[32\]
rlabel metal1 9157 11153 9157 11153 0 ct.oc.data_chain\[330\]
rlabel metal1 9157 12241 9157 12241 0 ct.oc.data_chain\[331\]
rlabel via2 8878 12597 8878 12597 0 ct.oc.data_chain\[332\]
rlabel via1 8143 8942 8143 8942 0 ct.oc.data_chain\[333\]
rlabel metal1 6785 9554 6785 9554 0 ct.oc.data_chain\[334\]
rlabel metal1 7061 10030 7061 10030 0 ct.oc.data_chain\[335\]
rlabel metal1 6901 12206 6901 12206 0 ct.oc.data_chain\[336\]
rlabel metal1 7245 14382 7245 14382 0 ct.oc.data_chain\[337\]
rlabel metal1 6257 11730 6257 11730 0 ct.oc.data_chain\[338\]
rlabel metal1 6578 12954 6578 12954 0 ct.oc.data_chain\[339\]
rlabel via1 6579 17170 6579 17170 0 ct.oc.data_chain\[33\]
rlabel metal2 6716 12614 6716 12614 0 ct.oc.data_chain\[340\]
rlabel metal1 5658 9554 5658 9554 0 ct.oc.data_chain\[341\]
rlabel metal1 5981 8466 5981 8466 0 ct.oc.data_chain\[342\]
rlabel metal1 5796 9146 5796 9146 0 ct.oc.data_chain\[343\]
rlabel metal1 4005 13329 4005 13329 0 ct.oc.data_chain\[344\]
rlabel via1 4279 11730 4279 11730 0 ct.oc.data_chain\[345\]
rlabel metal1 4049 13906 4049 13906 0 ct.oc.data_chain\[346\]
rlabel metal1 3727 12818 3727 12818 0 ct.oc.data_chain\[347\]
rlabel metal1 4005 12241 4005 12241 0 ct.oc.data_chain\[348\]
rlabel metal1 3451 9554 3451 9554 0 ct.oc.data_chain\[349\]
rlabel metal1 6210 18394 6210 18394 0 ct.oc.data_chain\[34\]
rlabel metal1 3543 10030 3543 10030 0 ct.oc.data_chain\[350\]
rlabel viali 3727 8944 3727 8944 0 ct.oc.data_chain\[351\]
rlabel metal1 6303 18258 6303 18258 0 ct.oc.data_chain\[35\]
rlabel metal2 1610 18870 1610 18870 0 ct.oc.data_chain\[36\]
rlabel viali 1462 18249 1462 18249 0 ct.oc.data_chain\[37\]
rlabel metal1 1610 21488 1610 21488 0 ct.oc.data_chain\[38\]
rlabel metal1 1610 19856 1610 19856 0 ct.oc.data_chain\[39\]
rlabel metal2 13110 20128 13110 20128 0 ct.oc.data_chain\[3\]
rlabel metal1 4991 17170 4991 17170 0 ct.oc.data_chain\[40\]
rlabel metal1 6118 15130 6118 15130 0 ct.oc.data_chain\[41\]
rlabel metal1 5037 18258 5037 18258 0 ct.oc.data_chain\[42\]
rlabel metal1 4117 17646 4117 17646 0 ct.oc.data_chain\[43\]
rlabel metal2 2806 16150 2806 16150 0 ct.oc.data_chain\[44\]
rlabel metal1 1978 17680 1978 17680 0 ct.oc.data_chain\[45\]
rlabel metal2 3082 18054 3082 18054 0 ct.oc.data_chain\[46\]
rlabel metal1 1840 18769 1840 18769 0 ct.oc.data_chain\[47\]
rlabel viali 4005 15471 4005 15471 0 ct.oc.data_chain\[48\]
rlabel metal1 5313 14994 5313 14994 0 ct.oc.data_chain\[49\]
rlabel metal1 17894 21454 17894 21454 0 ct.oc.data_chain\[4\]
rlabel via1 4003 16558 4003 16558 0 ct.oc.data_chain\[50\]
rlabel metal1 5221 16082 5221 16082 0 ct.oc.data_chain\[51\]
rlabel via2 2162 15011 2162 15011 0 ct.oc.data_chain\[52\]
rlabel metal1 1978 15504 1978 15504 0 ct.oc.data_chain\[53\]
rlabel metal2 1794 16677 1794 16677 0 ct.oc.data_chain\[54\]
rlabel metal2 10442 16337 10442 16337 0 ct.oc.data_chain\[55\]
rlabel metal1 11086 14824 11086 14824 0 ct.oc.data_chain\[56\]
rlabel metal2 13478 15623 13478 15623 0 ct.oc.data_chain\[57\]
rlabel metal2 10534 14586 10534 14586 0 ct.oc.data_chain\[58\]
rlabel metal2 13478 14739 13478 14739 0 ct.oc.data_chain\[59\]
rlabel metal1 8280 21114 8280 21114 0 ct.oc.data_chain\[5\]
rlabel metal2 13110 16694 13110 16694 0 ct.oc.data_chain\[60\]
rlabel metal1 9098 16047 9098 16047 0 ct.oc.data_chain\[61\]
rlabel metal2 12742 15606 12742 15606 0 ct.oc.data_chain\[62\]
rlabel metal1 11178 18360 11178 18360 0 ct.oc.data_chain\[63\]
rlabel metal1 11845 14994 11845 14994 0 ct.oc.data_chain\[64\]
rlabel metal1 12213 15470 12213 15470 0 ct.oc.data_chain\[65\]
rlabel metal1 13846 13974 13846 13974 0 ct.oc.data_chain\[66\]
rlabel metal1 12134 14417 12134 14417 0 ct.oc.data_chain\[67\]
rlabel metal1 11776 17681 11776 17681 0 ct.oc.data_chain\[68\]
rlabel metal2 13570 17204 13570 17204 0 ct.oc.data_chain\[69\]
rlabel metal2 4738 19720 4738 19720 0 ct.oc.data_chain\[6\]
rlabel metal2 15962 16133 15962 16133 0 ct.oc.data_chain\[70\]
rlabel metal1 14582 18224 14582 18224 0 ct.oc.data_chain\[71\]
rlabel metal1 15157 14994 15157 14994 0 ct.oc.data_chain\[72\]
rlabel metal1 15893 16082 15893 16082 0 ct.oc.data_chain\[73\]
rlabel metal1 14927 13906 14927 13906 0 ct.oc.data_chain\[74\]
rlabel metal1 14421 14382 14421 14382 0 ct.oc.data_chain\[75\]
rlabel metal1 14697 16558 14697 16558 0 ct.oc.data_chain\[76\]
rlabel viali 14951 18256 14951 18256 0 ct.oc.data_chain\[77\]
rlabel metal1 14421 15470 14421 15470 0 ct.oc.data_chain\[78\]
rlabel metal1 14421 17646 14421 17646 0 ct.oc.data_chain\[79\]
rlabel metal1 5290 18904 5290 18904 0 ct.oc.data_chain\[7\]
rlabel metal1 18814 13940 18814 13940 0 ct.oc.data_chain\[80\]
rlabel metal2 19826 15164 19826 15164 0 ct.oc.data_chain\[81\]
rlabel metal1 17825 15470 17825 15470 0 ct.oc.data_chain\[82\]
rlabel metal1 17733 14382 17733 14382 0 ct.oc.data_chain\[83\]
rlabel metal2 21850 17578 21850 17578 0 ct.oc.data_chain\[84\]
rlabel metal1 20654 16150 20654 16150 0 ct.oc.data_chain\[85\]
rlabel metal2 21666 17255 21666 17255 0 ct.oc.data_chain\[86\]
rlabel metal1 19550 16694 19550 16694 0 ct.oc.data_chain\[87\]
rlabel metal2 22954 14705 22954 14705 0 ct.oc.data_chain\[88\]
rlabel metal1 21804 15504 21804 15504 0 ct.oc.data_chain\[89\]
rlabel metal1 12673 19822 12673 19822 0 ct.oc.data_chain\[8\]
rlabel metal2 20654 14127 20654 14127 0 ct.oc.data_chain\[90\]
rlabel metal2 20562 15079 20562 15079 0 ct.oc.data_chain\[91\]
rlabel metal1 21229 18258 21229 18258 0 ct.oc.data_chain\[92\]
rlabel metal2 21942 17493 21942 17493 0 ct.oc.data_chain\[93\]
rlabel via1 22034 16949 22034 16949 0 ct.oc.data_chain\[94\]
rlabel metal2 21298 17391 21298 17391 0 ct.oc.data_chain\[95\]
rlabel metal1 24337 16047 24337 16047 0 ct.oc.data_chain\[96\]
rlabel viali 23985 16559 23985 16559 0 ct.oc.data_chain\[97\]
rlabel metal1 25134 14994 25134 14994 0 ct.oc.data_chain\[98\]
rlabel metal1 23969 15505 23969 15505 0 ct.oc.data_chain\[99\]
rlabel metal1 12420 18769 12420 18769 0 ct.oc.data_chain\[9\]
rlabel metal1 12926 21386 12926 21386 0 ct.oc.mode_buffer\[0\]
rlabel metal1 20335 14790 20335 14790 0 ct.oc.mode_buffer\[10\]
rlabel metal1 25303 18054 25303 18054 0 ct.oc.mode_buffer\[11\]
rlabel metal1 26981 20434 26981 20434 0 ct.oc.mode_buffer\[12\]
rlabel via1 28821 19822 28821 19822 0 ct.oc.mode_buffer\[13\]
rlabel metal1 27511 12614 27511 12614 0 ct.oc.mode_buffer\[14\]
rlabel metal1 21577 12614 21577 12614 0 ct.oc.mode_buffer\[15\]
rlabel metal1 19001 13498 19001 13498 0 ct.oc.mode_buffer\[16\]
rlabel metal1 21117 10438 21117 10438 0 ct.oc.mode_buffer\[17\]
rlabel metal1 21715 9350 21715 9350 0 ct.oc.mode_buffer\[18\]
rlabel via1 19069 7378 19069 7378 0 ct.oc.mode_buffer\[19\]
rlabel metal1 6075 20026 6075 20026 0 ct.oc.mode_buffer\[1\]
rlabel via1 28269 3502 28269 3502 0 ct.oc.mode_buffer\[20\]
rlabel metal1 17045 6766 17045 6766 0 ct.oc.mode_buffer\[21\]
rlabel metal1 2073 646 2073 646 0 ct.oc.mode_buffer\[22\]
rlabel metal1 17437 646 17437 646 0 ct.oc.mode_buffer\[23\]
rlabel viali 23833 1396 23833 1396 0 ct.oc.mode_buffer\[24\]
rlabel metal1 21669 2618 21669 2618 0 ct.oc.mode_buffer\[25\]
rlabel metal1 19093 1734 19093 1734 0 ct.oc.mode_buffer\[26\]
rlabel metal1 16885 5882 16885 5882 0 ct.oc.mode_buffer\[27\]
rlabel metal1 14125 2618 14125 2618 0 ct.oc.mode_buffer\[28\]
rlabel metal1 11319 1734 11319 1734 0 ct.oc.mode_buffer\[29\]
rlabel metal1 6213 21318 6213 21318 0 ct.oc.mode_buffer\[2\]
rlabel metal1 7872 646 7872 646 0 ct.oc.mode_buffer\[30\]
rlabel metal1 13941 646 13941 646 0 ct.oc.mode_buffer\[31\]
rlabel metal1 16263 12750 16263 12750 0 ct.oc.mode_buffer\[32\]
rlabel via1 1313 13906 1313 13906 0 ct.oc.mode_buffer\[33\]
rlabel metal2 7176 12852 7176 12852 0 ct.oc.mode_buffer\[34\]
rlabel metal1 1521 8262 1521 8262 0 ct.oc.mode_buffer\[35\]
rlabel metal1 9341 6970 9341 6970 0 ct.oc.mode_buffer\[36\]
rlabel metal1 16517 8058 16517 8058 0 ct.oc.mode_buffer\[37\]
rlabel via1 14309 9350 14309 9350 0 ct.oc.mode_buffer\[38\]
rlabel via1 9317 9554 9317 9554 0 ct.oc.mode_buffer\[39\]
rlabel via1 1313 20434 1313 20434 0 ct.oc.mode_buffer\[3\]
rlabel metal1 7961 9146 7961 9146 0 ct.oc.mode_buffer\[40\]
rlabel via1 6029 8262 6029 8262 0 ct.oc.mode_buffer\[41\]
rlabel metal1 3959 9350 3959 9350 0 ct.oc.mode_buffer\[42\]
rlabel metal1 1613 9350 1613 9350 0 ct.oc.mode_buffer\[43\]
rlabel via1 1681 17714 1681 17714 0 ct.oc.mode_buffer\[4\]
rlabel via1 1681 15470 1681 15470 0 ct.oc.mode_buffer\[5\]
rlabel metal1 6535 14790 6535 14790 0 ct.oc.mode_buffer\[6\]
rlabel via1 11617 17714 11617 17714 0 ct.oc.mode_buffer\[7\]
rlabel metal1 14769 13702 14769 13702 0 ct.oc.mode_buffer\[8\]
rlabel metal1 16839 14790 16839 14790 0 ct.oc.mode_buffer\[9\]
rlabel metal1 16560 14246 16560 14246 0 ct.oc.trig_chain\[10\]
rlabel metal2 19918 14416 19918 14416 0 ct.oc.trig_chain\[11\]
rlabel metal1 23690 15470 23690 15470 0 ct.oc.trig_chain\[12\]
rlabel metal1 26726 20502 26726 20502 0 ct.oc.trig_chain\[13\]
rlabel metal1 28474 17646 28474 17646 0 ct.oc.trig_chain\[14\]
rlabel metal1 23782 12750 23782 12750 0 ct.oc.trig_chain\[15\]
rlabel metal1 26588 7310 26588 7310 0 ct.oc.trig_chain\[16\]
rlabel metal2 18676 12444 18676 12444 0 ct.oc.trig_chain\[17\]
rlabel metal1 20930 9078 20930 9078 0 ct.oc.trig_chain\[18\]
rlabel metal2 17434 9520 17434 9520 0 ct.oc.trig_chain\[19\]
rlabel metal1 5336 19142 5336 19142 0 ct.oc.trig_chain\[1\]
rlabel metal1 18906 8398 18906 8398 0 ct.oc.trig_chain\[20\]
rlabel metal1 28106 2482 28106 2482 0 ct.oc.trig_chain\[21\]
rlabel metal1 16790 6698 16790 6698 0 ct.oc.trig_chain\[22\]
rlabel metal2 1334 1156 1334 1156 0 ct.oc.trig_chain\[23\]
rlabel metal2 24150 476 24150 476 0 ct.oc.trig_chain\[24\]
rlabel metal1 23230 1326 23230 1326 0 ct.oc.trig_chain\[25\]
rlabel metal1 20838 5134 20838 5134 0 ct.oc.trig_chain\[26\]
rlabel metal1 18630 5134 18630 5134 0 ct.oc.trig_chain\[27\]
rlabel metal1 16008 1870 16008 1870 0 ct.oc.trig_chain\[28\]
rlabel metal2 12558 4420 12558 4420 0 ct.oc.trig_chain\[29\]
rlabel metal1 5658 19822 5658 19822 0 ct.oc.trig_chain\[2\]
rlabel metal1 8694 1258 8694 1258 0 ct.oc.trig_chain\[30\]
rlabel metal1 8694 748 8694 748 0 ct.oc.trig_chain\[31\]
rlabel metal1 6351 2482 6351 2482 0 ct.oc.trig_chain\[32\]
rlabel metal1 15226 12750 15226 12750 0 ct.oc.trig_chain\[33\]
rlabel metal2 966 17408 966 17408 0 ct.oc.trig_chain\[34\]
rlabel metal1 6394 5746 6394 5746 0 ct.oc.trig_chain\[35\]
rlabel metal2 3542 7956 3542 7956 0 ct.oc.trig_chain\[36\]
rlabel metal2 9062 7616 9062 7616 0 ct.oc.trig_chain\[37\]
rlabel metal1 16054 7922 16054 7922 0 ct.oc.trig_chain\[38\]
rlabel metal1 13892 10098 13892 10098 0 ct.oc.trig_chain\[39\]
rlabel metal1 5152 19482 5152 19482 0 ct.oc.trig_chain\[3\]
rlabel metal1 8970 9520 8970 9520 0 ct.oc.trig_chain\[40\]
rlabel metal1 6256 9554 6256 9554 0 ct.oc.trig_chain\[41\]
rlabel metal2 5520 9044 5520 9044 0 ct.oc.trig_chain\[42\]
rlabel metal1 3312 9486 3312 9486 0 ct.oc.trig_chain\[43\]
rlabel metal1 1426 13294 1426 13294 0 ct.oc.trig_chain\[44\]
rlabel metal1 920 19822 920 19822 0 ct.oc.trig_chain\[4\]
rlabel metal1 1334 17748 1334 17748 0 ct.oc.trig_chain\[5\]
rlabel metal1 1334 15402 1334 15402 0 ct.oc.trig_chain\[6\]
rlabel metal1 9982 15368 9982 15368 0 ct.oc.trig_chain\[7\]
rlabel metal1 11592 14926 11592 14926 0 ct.oc.trig_chain\[8\]
rlabel metal1 13846 14314 13846 14314 0 ct.oc.trig_chain\[9\]
rlabel metal1 21252 19822 21252 19822 0 ct.ro.counter\[0\]
rlabel metal1 21390 21386 21390 21386 0 ct.ro.counter\[1\]
rlabel metal1 21206 20264 21206 20264 0 ct.ro.counter\[2\]
rlabel metal2 22310 21284 22310 21284 0 ct.ro.counter\[3\]
rlabel metal1 24058 21386 24058 21386 0 ct.ro.counter\[4\]
rlabel metal1 23920 21522 23920 21522 0 ct.ro.counter\[5\]
rlabel via1 23403 20366 23403 20366 0 ct.ro.counter\[6\]
rlabel metal2 25714 20876 25714 20876 0 ct.ro.counter\[7\]
rlabel metal2 21758 19584 21758 19584 0 ct.ro.counter_n\[0\]
rlabel metal1 20148 20910 20148 20910 0 ct.ro.counter_n\[1\]
rlabel metal1 21160 20366 21160 20366 0 ct.ro.counter_n\[2\]
rlabel metal1 23322 20944 23322 20944 0 ct.ro.counter_n\[3\]
rlabel metal1 23690 20910 23690 20910 0 ct.ro.counter_n\[4\]
rlabel metal1 21574 19822 21574 19822 0 ct.ro.counter_n\[5\]
rlabel metal1 23598 20400 23598 20400 0 ct.ro.counter_n\[6\]
rlabel metal1 25898 20400 25898 20400 0 ct.ro.counter_n\[7\]
rlabel metal1 20470 19958 20470 19958 0 ct.ro.gate
rlabel metal2 20654 20876 20654 20876 0 ct.ro.ring\[0\]
rlabel metal1 20470 18734 20470 18734 0 ct.ro.ring\[1\]
rlabel metal1 23506 18938 23506 18938 0 ct.ro.ring\[2\]
rlabel metal1 20976 14246 20976 14246 0 net1
rlabel metal2 4508 14450 4508 14450 0 net10
rlabel metal1 12466 8296 12466 8296 0 net11
rlabel metal2 1426 18751 1426 18751 0 net12
rlabel metal1 18262 1428 18262 1428 0 net13
rlabel metal2 18630 15776 18630 15776 0 net14
rlabel metal1 1058 5712 1058 5712 0 net15
rlabel metal1 8786 7310 8786 7310 0 net16
rlabel metal1 1242 17612 1242 17612 0 net17
rlabel metal1 29578 10710 29578 10710 0 net18
rlabel metal1 18906 6256 18906 6256 0 net19
rlabel metal3 28497 12444 28497 12444 0 net2
rlabel metal2 20746 15895 20746 15895 0 net20
rlabel metal1 15272 782 15272 782 0 net21
rlabel metal1 13938 6222 13938 6222 0 net22
rlabel metal1 9614 14484 9614 14484 0 net23
rlabel metal1 29578 10472 29578 10472 0 net24
rlabel metal1 29118 12614 29118 12614 0 net25
rlabel metal1 20930 16456 20930 16456 0 net26
rlabel metal1 6808 5746 6808 5746 0 net27
rlabel metal1 1196 13362 1196 13362 0 net28
rlabel metal3 7452 19788 7452 19788 0 net29
rlabel metal2 25070 21862 25070 21862 0 net3
rlabel metal1 20516 9010 20516 9010 0 net30
rlabel metal1 30820 14790 30820 14790 0 net31
rlabel metal1 29164 13974 29164 13974 0 net32
rlabel metal1 1426 14518 1426 14518 0 net33
rlabel metal2 9062 8670 9062 8670 0 net34
rlabel metal1 5428 20978 5428 20978 0 net35
rlabel metal1 16330 9418 16330 9418 0 net36
rlabel metal3 19228 14280 19228 14280 0 net37
rlabel metal2 21022 13158 21022 13158 0 net38
rlabel metal2 13662 17289 13662 17289 0 net39
rlabel metal2 23598 19516 23598 19516 0 net4
rlabel metal2 18262 7072 18262 7072 0 net40
rlabel metal1 12604 19278 12604 19278 0 net41
rlabel metal1 18216 7310 18216 7310 0 net42
rlabel metal1 17250 12274 17250 12274 0 net43
rlabel metal1 19182 13906 19182 13906 0 net44
rlabel via2 2346 6851 2346 6851 0 net45
rlabel metal2 13386 11968 13386 11968 0 net46
rlabel metal1 13432 18122 13432 18122 0 net47
rlabel metal1 18538 1938 18538 1938 0 net48
rlabel metal1 16100 11662 16100 11662 0 net49
rlabel metal2 1150 5780 1150 5780 0 net5
rlabel metal2 12650 19788 12650 19788 0 net50
rlabel metal1 13248 4046 13248 4046 0 net51
rlabel metal2 16146 21760 16146 21760 0 net52
rlabel metal1 20562 3536 20562 3536 0 net53
rlabel metal2 18906 20196 18906 20196 0 net54
rlabel metal1 19458 14280 19458 14280 0 net55
rlabel metal4 8188 22137 8188 22137 0 net56
rlabel metal1 10028 19890 10028 19890 0 net57
rlabel metal1 10258 13770 10258 13770 0 net58
rlabel metal4 6532 20165 6532 20165 0 net59
rlabel metal2 9246 3876 9246 3876 0 net6
rlabel metal3 7636 17340 7636 17340 0 net60
rlabel metal1 15226 15368 15226 15368 0 net61
rlabel metal4 4876 22137 4876 22137 0 net62
rlabel metal1 12098 12852 12098 12852 0 net63
rlabel metal1 1150 4726 1150 4726 0 net7
rlabel metal1 16790 4080 16790 4080 0 net8
rlabel metal2 20010 16167 20010 16167 0 net9
rlabel metal2 19918 19061 19918 19061 0 rst_n
rlabel metal1 17802 19278 17802 19278 0 ui_in[0]
rlabel metal1 17158 20978 17158 20978 0 ui_in[1]
rlabel metal1 18170 19414 18170 19414 0 ui_in[2]
rlabel metal1 21114 14348 21114 14348 0 ui_in[3]
rlabel metal2 18722 21250 18722 21250 0 ui_in[4]
rlabel metal4 23092 22137 23092 22137 0 ui_in[5]
rlabel metal4 22540 20097 22540 20097 0 ui_in[6]
rlabel metal4 21988 21049 21988 21049 0 ui_in[7]
rlabel metal4 12604 20709 12604 20709 0 uio_out[0]
rlabel metal2 12558 21743 12558 21743 0 uio_out[1]
rlabel metal1 10994 20502 10994 20502 0 uio_out[2]
rlabel metal2 8326 19584 8326 19584 0 uio_out[3]
rlabel metal2 18906 21964 18906 21964 0 uio_out[4]
rlabel metal1 8050 17510 8050 17510 0 uio_out[5]
rlabel via2 5106 18853 5106 18853 0 uio_out[6]
rlabel metal1 6486 18598 6486 18598 0 uio_out[7]
rlabel metal2 17158 21335 17158 21335 0 uo_out[0]
rlabel metal1 16836 17850 16836 17850 0 uo_out[1]
rlabel metal1 17342 19142 17342 19142 0 uo_out[2]
rlabel metal4 15364 21457 15364 21457 0 uo_out[3]
rlabel metal1 15410 17306 15410 17306 0 uo_out[4]
rlabel via2 13386 16405 13386 16405 0 uo_out[5]
rlabel metal1 15042 20570 15042 20570 0 uo_out[6]
rlabel metal4 13156 22137 13156 22137 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 31464 22304
<< end >>
