magic
tech sky130A
magscale 1 2
timestamp 1698890999
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1931 203
rect 29 -17 63 21
<< locali >>
rect 1809 59 1903 93
rect 1869 93 1903 451
rect 1809 451 1903 485
rect 29 215 117 249
rect 29 249 63 323
rect 1593 153 1627 215
rect 1593 215 1749 249
rect 1685 249 1719 255
rect 305 215 373 249
rect 305 249 339 255
<< obsli1 >>
rect 121 435 155 527
rect 63 527 121 561
rect 155 527 213 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 1093 51 1127 127
rect 1029 127 1127 161
rect 1029 161 1063 199
rect 767 199 801 215
rect 1029 199 1063 215
rect 767 215 803 265
rect 1029 215 1063 265
rect 769 265 803 299
rect 1029 265 1063 299
rect 769 299 1063 333
rect 1029 333 1063 357
rect 1029 357 1111 391
rect 1077 391 1111 427
rect 1077 427 1223 477
rect 1105 477 1223 493
rect 37 51 71 143
rect 37 143 195 177
rect 161 177 195 199
rect 161 199 197 265
rect 161 265 195 289
rect 121 289 195 323
rect 161 323 195 359
rect 37 359 71 367
rect 161 359 195 367
rect 37 367 195 401
rect 37 401 71 493
rect 393 427 523 493
rect 1557 59 1707 93
rect 1673 93 1707 143
rect 1673 143 1819 177
rect 1785 177 1819 199
rect 1785 199 1829 265
rect 1785 265 1819 289
rect 1777 289 1819 323
rect 1785 323 1819 357
rect 1657 357 1819 391
rect 1657 391 1691 493
rect 737 375 939 409
rect 737 409 771 493
rect 905 409 939 493
rect 1173 127 1535 161
rect 1501 161 1535 199
rect 1501 199 1553 265
rect 1501 265 1535 357
rect 1393 357 1535 391
rect 1393 391 1427 451
rect 1269 451 1427 485
rect 473 127 991 161
rect 697 161 731 199
rect 957 161 991 199
rect 697 199 731 249
rect 957 199 993 249
rect 697 249 731 265
rect 959 249 993 265
rect 697 265 731 299
rect 669 299 731 333
rect 669 333 703 451
rect 557 451 703 485
rect 189 67 267 101
rect 233 101 267 199
rect 233 199 267 215
rect 627 199 661 215
rect 233 215 267 249
rect 419 215 485 249
rect 601 215 661 249
rect 233 249 267 265
rect 421 249 455 265
rect 601 249 661 265
rect 233 265 267 299
rect 421 265 455 299
rect 601 265 635 299
rect 233 299 455 333
rect 601 299 635 333
rect 233 333 267 357
rect 421 333 455 357
rect 601 333 635 357
rect 233 357 267 391
rect 421 357 635 391
rect 233 391 267 443
rect 189 443 267 477
rect 1135 199 1169 215
rect 1327 199 1361 215
rect 1135 215 1179 265
rect 1317 215 1361 265
rect 1145 265 1179 357
rect 1317 265 1351 357
rect 1145 357 1351 391
rect 1231 199 1265 215
rect 1225 215 1265 265
rect 1225 265 1259 323
rect 1423 199 1457 215
rect 1409 215 1457 265
rect 1409 265 1443 323
rect 531 199 565 215
rect 529 215 565 265
rect 529 265 563 289
rect 489 289 563 323
rect 863 199 897 221
rect 857 221 897 255
rect 863 255 897 265
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 1269 59 1419 93
rect 557 59 707 93
rect 0 527 29 561
rect 805 451 871 527
rect 799 527 857 561
rect 707 527 765 561
rect 615 527 673 561
rect 523 527 581 561
rect 431 527 489 561
rect 1009 427 1043 527
rect 983 527 1041 561
rect 891 527 949 561
rect 1573 367 1607 435
rect 1469 435 1607 527
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1351 527 1409 561
rect 1259 527 1317 561
rect 1167 527 1225 561
rect 1075 527 1133 561
rect 1741 435 1775 527
rect 1719 527 1777 561
rect 1627 527 1685 561
rect 309 367 343 527
rect 339 527 397 561
rect 247 527 305 561
rect 1719 -17 1777 17
rect 1741 17 1775 109
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1453 17 1519 93
rect 1351 -17 1409 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 889 17 1059 93
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 309 17 343 177
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 121 17 155 109
rect 0 -17 29 17
<< obsli1c >>
rect 1593 527 1627 561
rect 1041 527 1075 561
rect 1685 527 1719 561
rect 1133 527 1167 561
rect 489 527 523 561
rect 1317 527 1351 561
rect 213 527 247 561
rect 765 527 799 561
rect 29 527 63 561
rect 397 527 431 561
rect 949 527 983 561
rect 121 527 155 561
rect 305 527 339 561
rect 1869 527 1903 561
rect 581 527 615 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 857 527 891 561
rect 1225 527 1259 561
rect 673 527 707 561
rect 1777 527 1811 561
rect 213 -17 247 17
rect 1869 -17 1903 17
rect 1777 -17 1811 17
rect 1593 -17 1627 17
rect 581 -17 615 17
rect 1501 -17 1535 17
rect 1409 -17 1443 17
rect 673 -17 707 17
rect 1041 -17 1075 17
rect 1225 -17 1259 17
rect 397 -17 431 17
rect 1317 -17 1351 17
rect 121 -17 155 17
rect 765 -17 799 17
rect 29 -17 63 17
rect 949 -17 983 17
rect 1133 -17 1167 17
rect 305 -17 339 17
rect 489 -17 523 17
rect 857 -17 891 17
rect 1685 -17 1719 17
<< metal1 >>
rect 0 496 1932 527
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 561 1932 592
rect 0 -48 1932 -17
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 17 1932 48
<< obsm1 >>
rect 569 351 627 360
rect 1305 351 1363 360
rect 569 360 1363 388
rect 569 388 627 397
rect 1305 388 1363 397
rect 109 283 167 292
rect 477 283 535 292
rect 1213 283 1271 292
rect 109 292 1271 320
rect 109 320 167 329
rect 477 320 535 329
rect 1213 320 1271 329
rect 1397 283 1455 292
rect 1765 283 1823 292
rect 1397 292 1823 320
rect 1397 320 1455 329
rect 1765 320 1823 329
rect 845 215 903 224
rect 1673 215 1731 224
rect 845 224 1731 252
rect 845 252 903 261
rect 1673 252 1731 261
<< labels >>
rlabel locali s 29 215 117 249 6 CLK
port 5 nsew signal input
rlabel locali s 29 249 63 323 6 CLK
port 5 nsew signal input
rlabel locali s 305 215 373 249 6 D
port 6 nsew signal input
rlabel locali s 305 249 339 255 6 D
port 6 nsew signal input
rlabel locali s 1593 153 1627 215 6 RESET_B
port 7 nsew signal input
rlabel locali s 1593 215 1749 249 6 RESET_B
port 7 nsew signal input
rlabel locali s 1685 249 1719 255 6 RESET_B
port 7 nsew signal input
rlabel locali s 1809 59 1903 93 6 Q
port 8 nsew signal output
rlabel locali s 1869 93 1903 451 6 Q
port 8 nsew signal output
rlabel locali s 1809 451 1903 485 6 Q
port 8 nsew signal output
rlabel pwell s 30 -17 64 21 6 VNB
port 1 nsew ground bidirectional
rlabel pwell s 1 21 1931 203 6 VNB
port 1 nsew ground bidirectional
rlabel nwell s -38 261 1970 582 6 VPB
port 2 nsew power bidirectional
rlabel metal1 s 0 -48 1932 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ht_sc_tt05.gds
string GDS_START 24132
string GDS_END 38260
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
