magic
tech sky130A
magscale 1 2
timestamp 1698890999
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 1 21 1379 203
rect 29 -17 63 21
<< scnmos >>
rect 1057 47 1087 177
rect 1153 47 1183 177
rect 1249 47 1279 177
rect 81 47 111 177
rect 165 47 195 177
rect 353 47 383 177
rect 449 47 479 177
rect 557 47 587 177
rect 665 47 695 177
rect 773 47 803 177
rect 869 47 899 177
<< scpmoshvt >>
rect 1057 297 1087 497
rect 1153 297 1183 497
rect 1249 297 1279 497
rect 81 297 111 497
rect 165 297 195 497
rect 353 297 383 497
rect 449 297 479 497
rect 557 297 587 497
rect 665 297 695 497
rect 773 297 803 497
rect 869 297 899 497
<< ndiff >>
rect 803 47 869 59
rect 803 59 825 93
rect 859 59 869 93
rect 803 93 869 177
rect 899 47 951 59
rect 899 59 909 93
rect 943 59 951 93
rect 899 93 951 177
rect 695 47 773 59
rect 695 59 729 93
rect 763 59 773 93
rect 695 93 773 177
rect 587 47 665 127
rect 587 127 621 161
rect 655 127 665 161
rect 587 161 665 177
rect 479 47 557 177
rect 383 47 449 59
rect 383 59 405 93
rect 439 59 449 93
rect 383 93 449 177
rect 195 47 247 67
rect 195 67 205 101
rect 239 67 247 101
rect 195 101 247 177
rect 111 47 165 59
rect 111 59 121 93
rect 155 59 165 93
rect 111 93 165 177
rect 1279 47 1331 59
rect 1279 59 1289 93
rect 1323 59 1331 93
rect 1279 93 1331 177
rect 1183 47 1249 59
rect 1183 59 1205 93
rect 1239 59 1249 93
rect 1183 93 1249 177
rect 1087 47 1153 177
rect 1005 47 1057 59
rect 1005 59 1013 93
rect 1047 59 1057 93
rect 1005 93 1057 177
rect 29 47 81 127
rect 29 127 37 161
rect 71 127 81 161
rect 29 161 81 177
rect 301 47 353 67
rect 301 67 309 101
rect 343 67 353 101
rect 301 101 353 177
<< pdiff >>
rect 803 297 869 497
rect 899 297 951 451
rect 899 451 909 485
rect 943 451 951 485
rect 899 485 951 497
rect 301 297 353 375
rect 301 375 309 409
rect 343 375 353 409
rect 301 409 353 443
rect 301 443 309 477
rect 343 443 353 477
rect 301 477 353 497
rect 29 297 81 375
rect 29 375 37 409
rect 71 375 81 409
rect 29 409 81 443
rect 29 443 37 477
rect 71 443 81 477
rect 29 477 81 497
rect 1005 297 1057 451
rect 1005 451 1013 485
rect 1047 451 1057 485
rect 1005 485 1057 497
rect 1087 297 1153 357
rect 1087 357 1109 391
rect 1143 357 1153 391
rect 1087 391 1153 451
rect 1087 451 1109 485
rect 1143 451 1153 485
rect 1087 485 1153 497
rect 1183 297 1249 451
rect 1183 451 1205 485
rect 1239 451 1249 485
rect 1183 485 1249 497
rect 1279 297 1331 383
rect 1279 383 1289 417
rect 1323 383 1331 417
rect 1279 417 1331 451
rect 1279 451 1289 485
rect 1323 451 1331 485
rect 1279 485 1331 497
rect 111 297 165 451
rect 111 451 121 485
rect 155 451 165 485
rect 111 485 165 497
rect 195 297 247 375
rect 195 375 205 409
rect 239 375 247 409
rect 195 409 247 443
rect 195 443 205 477
rect 239 443 247 477
rect 195 477 247 497
rect 383 297 449 383
rect 383 383 405 417
rect 439 383 449 417
rect 383 417 449 451
rect 383 451 405 485
rect 439 451 449 485
rect 383 485 449 497
rect 479 297 557 451
rect 479 451 513 485
rect 547 451 557 485
rect 479 485 557 497
rect 587 297 665 451
rect 587 451 621 485
rect 655 451 665 485
rect 587 485 665 497
rect 695 297 773 451
rect 695 451 729 485
rect 763 451 773 485
rect 695 485 773 497
<< ndiffc >>
rect 621 127 655 161
rect 37 127 71 161
rect 309 67 343 101
rect 205 67 239 101
rect 729 59 763 93
rect 1013 59 1047 93
rect 1289 59 1323 93
rect 909 59 943 93
rect 1205 59 1239 93
rect 121 59 155 93
rect 825 59 859 93
rect 405 59 439 93
<< pdiffc >>
rect 1013 451 1047 485
rect 513 451 547 485
rect 1205 451 1239 485
rect 405 451 439 485
rect 621 451 655 485
rect 121 451 155 485
rect 909 451 943 485
rect 1109 451 1143 485
rect 729 451 763 485
rect 1289 451 1323 485
rect 37 443 71 477
rect 205 443 239 477
rect 309 443 343 477
rect 1289 383 1323 417
rect 405 383 439 417
rect 37 375 71 409
rect 309 375 343 409
rect 205 375 239 409
rect 1109 357 1143 391
<< poly >>
rect 81 497 111 523
rect 1249 497 1279 523
rect 1153 497 1183 523
rect 1057 497 1087 523
rect 773 497 803 523
rect 665 497 695 523
rect 557 497 587 523
rect 449 497 479 523
rect 353 497 383 523
rect 165 497 195 523
rect 869 497 899 523
rect 1057 177 1087 199
rect 1033 199 1087 215
rect 1033 215 1043 249
rect 1077 215 1087 249
rect 1033 249 1087 265
rect 1057 265 1087 297
rect 81 177 111 199
rect 21 199 111 215
rect 21 215 31 249
rect 65 215 111 249
rect 21 249 111 265
rect 81 265 111 297
rect 869 177 899 199
rect 869 199 983 215
rect 869 215 939 249
rect 973 215 983 249
rect 869 249 983 265
rect 869 265 899 297
rect 773 177 803 199
rect 761 199 815 215
rect 761 215 771 249
rect 805 215 815 249
rect 761 249 815 265
rect 773 265 803 297
rect 665 177 695 199
rect 653 199 707 215
rect 653 215 663 249
rect 697 215 707 249
rect 653 249 707 265
rect 665 265 695 297
rect 557 177 587 199
rect 545 199 599 215
rect 545 215 555 249
rect 589 215 599 249
rect 545 249 599 265
rect 557 265 587 297
rect 353 177 383 199
rect 309 199 383 215
rect 309 215 319 249
rect 353 215 383 249
rect 309 249 383 265
rect 353 265 383 297
rect 165 177 195 199
rect 153 199 207 215
rect 153 215 163 249
rect 197 215 207 249
rect 153 249 207 265
rect 165 265 195 297
rect 1153 177 1183 199
rect 1141 199 1195 215
rect 1141 215 1151 249
rect 1185 215 1195 249
rect 1141 249 1195 265
rect 1153 265 1183 297
rect 449 177 479 199
rect 437 199 491 215
rect 437 215 447 249
rect 481 215 491 249
rect 437 249 491 265
rect 449 265 479 297
rect 1249 177 1279 199
rect 1249 199 1303 215
rect 1249 215 1259 249
rect 1293 215 1303 249
rect 1249 249 1303 265
rect 1249 265 1279 297
rect 81 21 111 47
rect 869 21 899 47
rect 773 21 803 47
rect 665 21 695 47
rect 557 21 587 47
rect 449 21 479 47
rect 353 21 383 47
rect 1249 21 1279 47
rect 1153 21 1183 47
rect 1057 21 1087 47
rect 165 21 195 47
<< polycont >>
rect 555 215 589 249
rect 663 215 697 249
rect 771 215 805 249
rect 319 215 353 249
rect 1259 215 1293 249
rect 939 215 973 249
rect 1151 215 1185 249
rect 447 215 481 249
rect 31 215 65 249
rect 163 215 197 249
rect 1043 215 1077 249
<< locali >>
rect 105 451 121 485
rect 155 451 171 485
rect 105 485 171 527
rect 63 527 121 561
rect 155 527 213 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 205 351 251 357
rect 205 357 213 375
rect 247 357 251 375
rect 247 375 251 391
rect 239 391 251 409
rect 205 409 251 443
rect 239 443 251 477
rect 205 477 251 493
rect 309 477 343 493
rect 37 477 71 493
rect 891 289 895 323
rect 857 323 891 357
rect 841 357 891 391
rect 841 391 875 451
rect 763 451 875 485
rect 1143 451 1159 485
rect 1273 59 1289 93
rect 1323 59 1363 93
rect 1273 93 1363 119
rect 1329 119 1363 357
rect 1273 357 1363 383
rect 1273 383 1289 417
rect 1323 383 1363 417
rect 1273 417 1363 451
rect 1273 451 1289 485
rect 1323 451 1363 485
rect 655 451 671 485
rect 713 451 729 485
rect 1093 451 1109 485
rect 547 451 621 485
rect 497 451 513 485
rect 1205 435 1239 451
rect 405 417 439 451
rect 309 409 343 443
rect 1259 199 1293 215
rect 1257 215 1259 249
rect 1257 249 1293 265
rect 1257 265 1291 289
rect 1133 289 1291 323
rect 1133 323 1167 357
rect 1143 357 1167 391
rect 977 59 1013 93
rect 977 93 1011 143
rect 941 143 1011 177
rect 941 177 975 199
rect 939 199 975 215
rect 973 215 975 249
rect 939 249 975 265
rect 941 265 975 357
rect 941 357 1109 391
rect 405 367 439 383
rect 309 101 343 143
rect 309 143 439 177
rect 405 177 439 199
rect 405 199 481 215
rect 405 215 447 249
rect 405 249 481 265
rect 405 265 439 289
rect 309 289 439 323
rect 309 323 343 375
rect 1027 215 1043 249
rect 1041 249 1075 289
rect 647 215 663 249
rect 697 215 713 249
rect 647 249 713 255
rect 673 255 711 289
rect 707 289 711 323
rect 29 221 31 249
rect 29 249 65 265
rect 29 265 63 323
rect 71 127 155 161
rect 121 161 155 199
rect 121 199 197 215
rect 121 215 163 249
rect 121 249 197 265
rect 121 265 159 289
rect 155 289 159 323
rect 121 323 155 375
rect 21 375 37 409
rect 71 375 155 409
rect 37 409 71 443
rect 1075 289 1079 323
rect 303 215 319 249
rect 353 215 369 249
rect 303 249 369 255
rect 1133 85 1167 215
rect 1133 215 1151 249
rect 1133 249 1167 255
rect 755 215 771 249
rect 589 215 605 249
rect 1185 215 1201 249
rect 1077 215 1093 249
rect 31 199 65 215
rect 21 127 37 161
rect 205 51 251 67
rect 239 67 251 85
rect 247 85 251 101
rect 205 101 213 119
rect 247 101 251 119
rect 205 119 251 125
rect 523 85 551 119
rect 517 119 551 215
rect 517 215 555 249
rect 805 215 821 249
rect 517 249 551 357
rect 773 249 807 357
rect 523 357 807 391
rect 1205 93 1239 109
rect 909 93 943 109
rect 1351 -17 1380 17
rect 859 59 875 93
rect 763 59 825 93
rect 1047 59 1063 93
rect 713 59 729 93
rect 309 51 343 67
rect 0 527 29 561
rect 1205 485 1239 527
rect 1167 527 1225 561
rect 1075 527 1133 561
rect 405 485 439 527
rect 431 527 489 561
rect 339 527 397 561
rect 247 527 305 561
rect 909 435 1047 451
rect 943 451 1013 485
rect 909 485 1047 527
rect 891 527 949 561
rect 983 527 1041 561
rect 799 527 857 561
rect 707 527 765 561
rect 615 527 673 561
rect 523 527 581 561
rect 605 127 621 143
rect 655 127 671 143
rect 605 143 621 161
rect 655 143 891 161
rect 605 161 891 177
rect 857 177 891 289
rect 1259 -17 1317 17
rect 1167 -17 1225 17
rect 1205 17 1239 59
rect 1075 -17 1133 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 909 17 943 59
rect 799 -17 857 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 389 17 455 59
rect 389 59 405 93
rect 439 59 455 93
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 105 17 171 59
rect 105 59 121 93
rect 155 59 171 93
rect 0 -17 29 17
<< viali >>
rect 1317 527 1351 561
rect 1225 527 1259 561
rect 1133 527 1167 561
rect 1041 527 1075 561
rect 949 527 983 561
rect 857 527 891 561
rect 765 527 799 561
rect 673 527 707 561
rect 581 527 615 561
rect 489 527 523 561
rect 397 527 431 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 527 63 561
rect 213 357 247 391
rect 489 357 523 391
rect 673 289 707 323
rect 857 289 891 323
rect 1041 289 1075 323
rect 121 289 155 323
rect 489 85 523 119
rect 213 85 247 119
rect 857 -17 891 17
rect 1133 -17 1167 17
rect 673 -17 707 17
rect 949 -17 983 17
rect 581 -17 615 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 121 -17 155 17
rect 29 -17 63 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 1041 -17 1075 17
rect 765 -17 799 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 496 1380 527
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 561 1380 592
rect 201 351 259 357
rect 477 351 535 357
rect 201 357 213 360
rect 247 357 259 360
rect 477 357 489 360
rect 523 357 535 360
rect 201 360 213 388
rect 247 360 489 388
rect 523 360 535 388
rect 201 388 213 391
rect 247 388 259 391
rect 477 388 489 391
rect 523 388 535 391
rect 201 391 259 397
rect 477 391 535 397
rect 845 283 903 289
rect 1029 283 1087 289
rect 845 289 857 292
rect 891 289 903 292
rect 1029 289 1041 292
rect 1075 289 1087 292
rect 845 292 857 320
rect 891 292 1041 320
rect 1075 292 1087 320
rect 845 320 857 323
rect 891 320 903 323
rect 1029 320 1041 323
rect 1075 320 1087 323
rect 845 323 903 329
rect 1029 323 1087 329
rect 109 283 167 289
rect 661 283 719 289
rect 109 289 121 292
rect 155 289 167 292
rect 661 289 673 292
rect 707 289 719 292
rect 109 292 121 320
rect 155 292 673 320
rect 707 292 719 320
rect 109 320 121 323
rect 155 320 167 323
rect 661 320 673 323
rect 707 320 719 323
rect 109 323 167 329
rect 661 323 719 329
rect 201 79 259 85
rect 477 79 535 85
rect 201 85 213 88
rect 247 85 259 88
rect 477 85 489 88
rect 523 85 535 88
rect 201 88 213 116
rect 247 88 489 116
rect 523 88 535 116
rect 201 116 213 119
rect 247 116 259 119
rect 477 116 489 119
rect 523 116 535 119
rect 201 119 259 125
rect 477 119 535 125
rect 0 -48 1380 -17
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 17 1380 48
<< labels >>
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 GATE
port 5 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 GATE
port 5 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 D
port 6 nsew signal input
flabel locali s 1133 85 1167 119 0 FreeSans 200 0 0 0 RESET_B
port 7 nsew signal input
flabel locali s 1133 153 1167 187 0 FreeSans 200 0 0 0 RESET_B
port 7 nsew signal input
flabel locali s 1133 221 1167 255 0 FreeSans 200 0 0 0 RESET_B
port 7 nsew signal input
flabel locali s 1317 85 1351 119 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1317 357 1351 391 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1317 425 1351 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 -48 1380 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1380 592 1 VPWR
port 4 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 dlrtp_1
<< properties >>
string FIXED_BBOX 0 0 1380 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ht_sc_tt05.gds
string GDS_START 13210
string GDS_END 24074
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
