magic
tech sky130A
magscale 1 2
timestamp 1699030165
<< viali >>
rect 3249 21641 3283 21675
rect 13185 21641 13219 21675
rect 25881 21641 25915 21675
rect 29653 21641 29687 21675
rect 30389 21641 30423 21675
rect 8401 21573 8435 21607
rect 15945 21573 15979 21607
rect 20729 21573 20763 21607
rect 23213 21573 23247 21607
rect 1455 21505 1489 21539
rect 3988 21503 4022 21537
rect 4261 21505 4295 21539
rect 5825 21505 5859 21539
rect 6288 21505 6322 21539
rect 9004 21505 9038 21539
rect 9140 21505 9174 21539
rect 11440 21505 11474 21539
rect 14016 21505 14050 21539
rect 21465 21505 21499 21539
rect 21925 21505 21959 21539
rect 22477 21505 22511 21539
rect 24501 21505 24535 21539
rect 949 21437 983 21471
rect 1685 21437 1719 21471
rect 3433 21437 3467 21471
rect 3525 21437 3559 21471
rect 6152 21437 6186 21471
rect 6561 21437 6595 21471
rect 8217 21437 8251 21471
rect 8585 21437 8619 21471
rect 8677 21437 8711 21471
rect 9413 21437 9447 21471
rect 10977 21437 11011 21471
rect 11713 21437 11747 21471
rect 13369 21437 13403 21471
rect 13553 21437 13587 21471
rect 14289 21437 14323 21471
rect 15669 21437 15703 21471
rect 15761 21437 15795 21471
rect 16129 21437 16163 21471
rect 16405 21437 16439 21471
rect 18705 21437 18739 21471
rect 18981 21437 19015 21471
rect 21281 21437 21315 21471
rect 22201 21437 22235 21471
rect 22318 21437 22352 21471
rect 23397 21437 23431 21471
rect 23673 21437 23707 21471
rect 23857 21437 23891 21471
rect 24041 21437 24075 21471
rect 24777 21437 24811 21471
rect 24915 21437 24949 21471
rect 25053 21437 25087 21471
rect 25789 21437 25823 21471
rect 26433 21437 26467 21471
rect 26709 21437 26743 21471
rect 28273 21437 28307 21471
rect 29101 21437 29135 21471
rect 29285 21437 29319 21471
rect 29377 21437 29411 21471
rect 30573 21437 30607 21471
rect 3065 21369 3099 21403
rect 17969 21369 18003 21403
rect 20545 21369 20579 21403
rect 29929 21369 29963 21403
rect 1415 21301 1449 21335
rect 3991 21301 4025 21335
rect 5549 21301 5583 21335
rect 7849 21301 7883 21335
rect 8033 21301 8067 21335
rect 10517 21301 10551 21335
rect 11443 21301 11477 21335
rect 12817 21301 12851 21335
rect 14019 21301 14053 21335
rect 17509 21301 17543 21335
rect 18061 21301 18095 21335
rect 20085 21301 20119 21335
rect 23121 21301 23155 21335
rect 23581 21301 23615 21335
rect 25697 21301 25731 21335
rect 27813 21301 27847 21335
rect 28365 21301 28399 21335
rect 30021 21301 30055 21335
rect 1783 21097 1817 21131
rect 6291 21097 6325 21131
rect 8499 21097 8533 21131
rect 10977 21097 11011 21131
rect 11719 21097 11753 21131
rect 15301 21097 15335 21131
rect 17969 21097 18003 21131
rect 20821 21097 20855 21131
rect 23121 21097 23155 21131
rect 25329 21097 25363 21131
rect 27813 21097 27847 21131
rect 30389 21097 30423 21131
rect 10425 21029 10459 21063
rect 10793 21029 10827 21063
rect 13369 21029 13403 21063
rect 3852 20961 3886 20995
rect 5641 20961 5675 20995
rect 5825 20961 5859 20995
rect 8769 20961 8803 20995
rect 11161 20985 11195 21019
rect 11989 20961 12023 20995
rect 13461 20961 13495 20995
rect 13788 20961 13822 20995
rect 15761 20961 15795 20995
rect 16406 20961 16440 20995
rect 18245 20961 18279 20995
rect 18521 20961 18555 20995
rect 18981 20961 19015 20995
rect 21005 20961 21039 20995
rect 23305 20961 23339 20995
rect 25513 20961 25547 20995
rect 25789 20961 25823 20995
rect 26709 20961 26743 20995
rect 28508 20961 28542 20995
rect 30573 20961 30607 20995
rect 1317 20893 1351 20927
rect 1823 20893 1857 20927
rect 2053 20893 2087 20927
rect 3525 20893 3559 20927
rect 3988 20893 4022 20927
rect 4261 20893 4295 20927
rect 6288 20911 6322 20945
rect 6561 20893 6595 20927
rect 8033 20893 8067 20927
rect 8496 20893 8530 20927
rect 11253 20893 11287 20927
rect 11716 20893 11750 20927
rect 13924 20893 13958 20927
rect 14197 20893 14231 20927
rect 16129 20893 16163 20927
rect 19257 20893 19291 20927
rect 21281 20893 21315 20927
rect 21557 20893 21591 20927
rect 23489 20893 23523 20927
rect 23765 20893 23799 20927
rect 26433 20893 26467 20927
rect 28181 20893 28215 20927
rect 28644 20893 28678 20927
rect 28917 20893 28951 20927
rect 17693 20825 17727 20859
rect 25973 20825 26007 20859
rect 1133 20757 1167 20791
rect 3157 20757 3191 20791
rect 7665 20757 7699 20791
rect 9873 20757 9907 20791
rect 15853 20757 15887 20791
rect 18061 20757 18095 20791
rect 18797 20757 18831 20791
rect 30021 20757 30055 20791
rect 2973 20553 3007 20587
rect 7113 20553 7147 20587
rect 7481 20553 7515 20587
rect 10517 20553 10551 20587
rect 28549 20553 28583 20587
rect 3525 20485 3559 20519
rect 8125 20485 8159 20519
rect 18061 20485 18095 20519
rect 18337 20485 18371 20519
rect 26341 20485 26375 20519
rect 1455 20417 1489 20451
rect 5736 20417 5770 20451
rect 8999 20417 9033 20451
rect 9229 20417 9263 20451
rect 11759 20417 11793 20451
rect 13369 20417 13403 20451
rect 14049 20399 14083 20433
rect 16224 20417 16258 20451
rect 19257 20417 19291 20451
rect 19533 20417 19567 20451
rect 21278 20417 21312 20451
rect 21833 20417 21867 20451
rect 24133 20417 24167 20451
rect 27215 20417 27249 20451
rect 949 20349 983 20383
rect 1685 20349 1719 20383
rect 4169 20349 4203 20383
rect 5273 20349 5307 20383
rect 6009 20349 6043 20383
rect 7665 20349 7699 20383
rect 8493 20349 8527 20383
rect 10701 20349 10735 20383
rect 10977 20349 11011 20383
rect 11253 20349 11287 20383
rect 11989 20349 12023 20383
rect 13553 20349 13587 20383
rect 14289 20349 14323 20383
rect 15761 20349 15795 20383
rect 16497 20349 16531 20383
rect 18245 20349 18279 20383
rect 18521 20349 18555 20383
rect 21557 20349 21591 20383
rect 23581 20349 23615 20383
rect 23857 20349 23891 20383
rect 25881 20349 25915 20383
rect 26157 20349 26191 20383
rect 26709 20349 26743 20383
rect 27445 20349 27479 20383
rect 29469 20349 29503 20383
rect 29837 20349 29871 20383
rect 4721 20281 4755 20315
rect 7849 20281 7883 20315
rect 18797 20281 18831 20315
rect 29101 20281 29135 20315
rect 30113 20281 30147 20315
rect 1415 20213 1449 20247
rect 3893 20213 3927 20247
rect 4445 20213 4479 20247
rect 4997 20213 5031 20247
rect 5739 20213 5773 20247
rect 8959 20213 8993 20247
rect 11719 20213 11753 20247
rect 14019 20213 14053 20247
rect 15393 20213 15427 20247
rect 16227 20213 16261 20247
rect 17601 20213 17635 20247
rect 18889 20213 18923 20247
rect 21097 20213 21131 20247
rect 23397 20213 23431 20247
rect 25697 20213 25731 20247
rect 27175 20213 27209 20247
rect 29929 20213 29963 20247
rect 30205 20213 30239 20247
rect 1783 20009 1817 20043
rect 3341 20009 3375 20043
rect 10333 20009 10367 20043
rect 20913 20009 20947 20043
rect 23949 20009 23983 20043
rect 28181 20009 28215 20043
rect 3617 19941 3651 19975
rect 4169 19941 4203 19975
rect 4537 19941 4571 19975
rect 4721 19941 4755 19975
rect 5089 19941 5123 19975
rect 5273 19941 5307 19975
rect 8401 19941 8435 19975
rect 11713 19941 11747 19975
rect 15945 19941 15979 19975
rect 19809 19941 19843 19975
rect 1225 19873 1259 19907
rect 1317 19873 1351 19907
rect 5825 19873 5859 19907
rect 6469 19873 6503 19907
rect 6745 19873 6779 19907
rect 7021 19873 7055 19907
rect 8493 19873 8527 19907
rect 8820 19873 8854 19907
rect 9229 19873 9263 19907
rect 11161 19873 11195 19907
rect 11345 19873 11379 19907
rect 12541 19873 12575 19907
rect 14197 19873 14231 19907
rect 14565 19873 14599 19907
rect 20177 19873 20211 19907
rect 21097 19873 21131 19907
rect 21281 19873 21315 19907
rect 22017 19873 22051 19907
rect 22109 19873 22143 19907
rect 24133 19873 24167 19907
rect 24593 19873 24627 19907
rect 26249 19873 26283 19907
rect 26709 19873 26743 19907
rect 28365 19873 28399 19907
rect 1813 19823 1847 19857
rect 2053 19805 2087 19839
rect 8956 19805 8990 19839
rect 11805 19805 11839 19839
rect 12132 19805 12166 19839
rect 12311 19805 12345 19839
rect 14289 19805 14323 19839
rect 16129 19805 16163 19839
rect 16405 19805 16439 19839
rect 17969 19805 18003 19839
rect 18245 19805 18279 19839
rect 20545 19805 20579 19839
rect 21649 19805 21683 19839
rect 22385 19805 22419 19839
rect 24317 19805 24351 19839
rect 26433 19805 26467 19839
rect 28457 19805 28491 19839
rect 28784 19805 28818 19839
rect 28920 19807 28954 19841
rect 29193 19805 29227 19839
rect 1041 19669 1075 19703
rect 3893 19669 3927 19703
rect 5549 19669 5583 19703
rect 6009 19669 6043 19703
rect 10977 19669 11011 19703
rect 13645 19669 13679 19703
rect 14013 19669 14047 19703
rect 17877 19669 17911 19703
rect 19349 19669 19383 19703
rect 20637 19669 20671 19703
rect 25697 19669 25731 19703
rect 26065 19669 26099 19703
rect 27997 19669 28031 19703
rect 30481 19669 30515 19703
rect 2973 19465 3007 19499
rect 3893 19465 3927 19499
rect 10241 19465 10275 19499
rect 13093 19465 13127 19499
rect 17877 19465 17911 19499
rect 23581 19465 23615 19499
rect 5549 19397 5583 19431
rect 11069 19397 11103 19431
rect 24133 19397 24167 19431
rect 30297 19397 30331 19431
rect 6288 19329 6322 19363
rect 8401 19329 8435 19363
rect 8864 19329 8898 19363
rect 11580 19329 11614 19363
rect 11759 19329 11793 19363
rect 14841 19329 14875 19363
rect 18153 19329 18187 19363
rect 21833 19329 21867 19363
rect 25007 19329 25041 19363
rect 27215 19327 27249 19361
rect 27399 19329 27433 19363
rect 857 19261 891 19295
rect 1133 19261 1167 19295
rect 2513 19261 2547 19295
rect 3433 19261 3467 19295
rect 4077 19261 4111 19295
rect 4353 19261 4387 19295
rect 5365 19261 5399 19295
rect 5825 19261 5859 19295
rect 6561 19261 6595 19295
rect 8217 19261 8251 19295
rect 9137 19261 9171 19295
rect 11253 19261 11287 19295
rect 11989 19261 12023 19295
rect 13829 19261 13863 19295
rect 15117 19261 15151 19295
rect 16129 19261 16163 19295
rect 16405 19261 16439 19295
rect 18061 19261 18095 19295
rect 18337 19261 18371 19295
rect 18521 19261 18555 19295
rect 18705 19261 18739 19295
rect 18981 19261 19015 19295
rect 20361 19261 20395 19295
rect 20453 19261 20487 19295
rect 20729 19261 20763 19295
rect 24501 19261 24535 19295
rect 25237 19261 25271 19295
rect 26709 19261 26743 19295
rect 27036 19261 27070 19295
rect 29009 19261 29043 19295
rect 29285 19261 29319 19295
rect 30205 19261 30239 19295
rect 2697 19193 2731 19227
rect 3617 19193 3651 19227
rect 7941 19193 7975 19227
rect 10793 19193 10827 19227
rect 15485 19193 15519 19227
rect 15853 19193 15887 19227
rect 17785 19193 17819 19227
rect 22477 19193 22511 19227
rect 23949 19193 23983 19227
rect 3249 19125 3283 19159
rect 4997 19125 5031 19159
rect 5181 19125 5215 19159
rect 6291 19125 6325 19159
rect 8033 19125 8067 19159
rect 8867 19125 8901 19159
rect 14473 19125 14507 19159
rect 14933 19125 14967 19159
rect 15945 19125 15979 19159
rect 24967 19125 25001 19159
rect 26341 19125 26375 19159
rect 28549 19125 28583 19159
rect 29929 19125 29963 19159
rect 30113 19125 30147 19159
rect 1783 18921 1817 18955
rect 7941 18921 7975 18955
rect 9143 18921 9177 18955
rect 14019 18921 14053 18955
rect 15393 18921 15427 18955
rect 23397 18921 23431 18955
rect 23489 18921 23523 18955
rect 28831 18921 28865 18955
rect 30205 18921 30239 18955
rect 3433 18853 3467 18887
rect 5641 18853 5675 18887
rect 8401 18853 8435 18887
rect 1225 18785 1259 18819
rect 6244 18785 6278 18819
rect 8125 18785 8159 18819
rect 10793 18785 10827 18819
rect 13461 18785 13495 18819
rect 14289 18785 14323 18819
rect 15945 18785 15979 18819
rect 16129 18785 16163 18819
rect 18613 18785 18647 18819
rect 20177 18785 20211 18819
rect 20545 18785 20579 18819
rect 21557 18785 21591 18819
rect 24041 18785 24075 18819
rect 24460 18785 24494 18819
rect 26709 18785 26743 18819
rect 28365 18785 28399 18819
rect 1317 18717 1351 18751
rect 1813 18735 1847 18769
rect 2053 18717 2087 18751
rect 3525 18717 3559 18751
rect 3852 18717 3886 18751
rect 3988 18719 4022 18753
rect 4261 18717 4295 18751
rect 5917 18717 5951 18751
rect 6380 18717 6414 18751
rect 6653 18717 6687 18751
rect 8677 18717 8711 18751
rect 9140 18717 9174 18751
rect 9413 18717 9447 18751
rect 10977 18717 11011 18751
rect 11304 18717 11338 18751
rect 11483 18719 11517 18753
rect 11713 18717 11747 18751
rect 13553 18717 13587 18751
rect 14016 18735 14050 18769
rect 16456 18717 16490 18751
rect 16592 18717 16626 18751
rect 16865 18717 16899 18751
rect 18337 18717 18371 18751
rect 19993 18717 20027 18751
rect 20913 18717 20947 18751
rect 21288 18717 21322 18751
rect 23581 18717 23615 18751
rect 24133 18717 24167 18751
rect 24639 18717 24673 18751
rect 24869 18717 24903 18751
rect 26433 18717 26467 18751
rect 28828 18717 28862 18751
rect 29101 18717 29135 18751
rect 12817 18649 12851 18683
rect 23029 18649 23063 18683
rect 27997 18649 28031 18683
rect 1041 18581 1075 18615
rect 13277 18581 13311 18615
rect 15761 18581 15795 18615
rect 18153 18581 18187 18615
rect 21005 18581 21039 18615
rect 22845 18581 22879 18615
rect 23857 18581 23891 18615
rect 25973 18581 26007 18615
rect 28273 18581 28307 18615
rect 5917 18377 5951 18411
rect 22753 18377 22787 18411
rect 28457 18377 28491 18411
rect 30297 18377 30331 18411
rect 2973 18309 3007 18343
rect 20085 18309 20119 18343
rect 24409 18309 24443 18343
rect 1455 18241 1489 18275
rect 4399 18241 4433 18275
rect 6564 18241 6598 18275
rect 8585 18241 8619 18275
rect 9091 18239 9125 18273
rect 9321 18241 9355 18275
rect 10701 18241 10735 18275
rect 11256 18241 11290 18275
rect 11529 18241 11563 18275
rect 14156 18241 14190 18275
rect 14335 18241 14369 18275
rect 17141 18241 17175 18275
rect 18705 18241 18739 18275
rect 20361 18241 20395 18275
rect 20867 18241 20901 18275
rect 24685 18241 24719 18275
rect 25191 18241 25225 18275
rect 27169 18241 27203 18275
rect 29009 18241 29043 18275
rect 949 18173 983 18207
rect 1685 18173 1719 18207
rect 3249 18173 3283 18207
rect 3893 18173 3927 18207
rect 4629 18173 4663 18207
rect 6101 18173 6135 18207
rect 6837 18173 6871 18207
rect 10793 18173 10827 18207
rect 13369 18173 13403 18207
rect 13829 18173 13863 18207
rect 14565 18173 14599 18207
rect 16313 18173 16347 18207
rect 16773 18173 16807 18207
rect 16865 18173 16899 18207
rect 18981 18173 19015 18207
rect 20269 18173 20303 18207
rect 21097 18173 21131 18207
rect 24593 18173 24627 18207
rect 25421 18173 25455 18207
rect 26893 18173 26927 18207
rect 28825 18173 28859 18207
rect 29285 18173 29319 18207
rect 30113 18173 30147 18207
rect 30573 18173 30607 18207
rect 3525 18105 3559 18139
rect 18521 18105 18555 18139
rect 19809 18105 19843 18139
rect 22661 18105 22695 18139
rect 23213 18105 23247 18139
rect 23581 18105 23615 18139
rect 23949 18105 23983 18139
rect 1415 18037 1449 18071
rect 4359 18037 4393 18071
rect 6567 18037 6601 18071
rect 8125 18037 8159 18071
rect 9051 18037 9085 18071
rect 11259 18037 11293 18071
rect 12633 18037 12667 18071
rect 13185 18037 13219 18071
rect 15669 18037 15703 18071
rect 16589 18037 16623 18071
rect 19993 18037 20027 18071
rect 20827 18037 20861 18071
rect 22201 18037 22235 18071
rect 24041 18037 24075 18071
rect 25151 18037 25185 18071
rect 26525 18037 26559 18071
rect 28641 18037 28675 18071
rect 30389 18037 30423 18071
rect 949 17833 983 17867
rect 1783 17833 1817 17867
rect 3157 17833 3191 17867
rect 9143 17833 9177 17867
rect 11995 17833 12029 17867
rect 15669 17833 15703 17867
rect 16773 17833 16807 17867
rect 23121 17833 23155 17867
rect 25973 17833 26007 17867
rect 26899 17833 26933 17867
rect 5641 17765 5675 17799
rect 6101 17765 6135 17799
rect 8585 17765 8619 17799
rect 10793 17765 10827 17799
rect 1133 17697 1167 17731
rect 3525 17697 3559 17731
rect 5825 17697 5859 17731
rect 6796 17697 6830 17731
rect 7205 17697 7239 17731
rect 9413 17697 9447 17731
rect 11069 17697 11103 17731
rect 11529 17697 11563 17731
rect 14565 17697 14599 17731
rect 16313 17697 16347 17731
rect 16497 17697 16531 17731
rect 17284 17697 17318 17731
rect 19165 17697 19199 17731
rect 19441 17697 19475 17731
rect 21097 17697 21131 17731
rect 22017 17697 22051 17731
rect 23673 17697 23707 17731
rect 24133 17697 24167 17731
rect 24460 17697 24494 17731
rect 28641 17697 28675 17731
rect 1317 17629 1351 17663
rect 1823 17631 1857 17665
rect 2053 17629 2087 17663
rect 3852 17629 3886 17663
rect 4021 17647 4055 17681
rect 4261 17629 4295 17663
rect 6469 17629 6503 17663
rect 6932 17631 6966 17665
rect 8677 17629 8711 17663
rect 9140 17629 9174 17663
rect 12035 17629 12069 17663
rect 12265 17629 12299 17663
rect 13829 17629 13863 17663
rect 14156 17629 14190 17663
rect 14335 17629 14369 17663
rect 16221 17629 16255 17663
rect 16957 17629 16991 17663
rect 17453 17647 17487 17681
rect 17693 17629 17727 17663
rect 21281 17629 21315 17663
rect 21608 17629 21642 17663
rect 21787 17629 21821 17663
rect 24639 17629 24673 17663
rect 24869 17629 24903 17663
rect 26433 17629 26467 17663
rect 26896 17629 26930 17663
rect 27169 17629 27203 17663
rect 28917 17629 28951 17663
rect 20913 17561 20947 17595
rect 23949 17561 23983 17595
rect 28457 17561 28491 17595
rect 30389 17561 30423 17595
rect 11161 17493 11195 17527
rect 13369 17493 13403 17527
rect 18797 17493 18831 17527
rect 20729 17493 20763 17527
rect 2973 17289 3007 17323
rect 5825 17289 5859 17323
rect 10517 17289 10551 17323
rect 14197 17289 14231 17323
rect 16129 17289 16163 17323
rect 25789 17289 25823 17323
rect 27997 17289 28031 17323
rect 28733 17289 28767 17323
rect 29929 17289 29963 17323
rect 8401 17221 8435 17255
rect 11069 17221 11103 17255
rect 30297 17221 30331 17255
rect 30389 17221 30423 17255
rect 949 17153 983 17187
rect 1445 17135 1479 17169
rect 1685 17153 1719 17187
rect 3341 17153 3375 17187
rect 3847 17153 3881 17187
rect 5457 17153 5491 17187
rect 6564 17153 6598 17187
rect 6837 17153 6871 17187
rect 8677 17153 8711 17187
rect 9140 17153 9174 17187
rect 9413 17153 9447 17187
rect 11580 17153 11614 17187
rect 11759 17153 11793 17187
rect 16911 17153 16945 17187
rect 17141 17153 17175 17187
rect 20959 17153 20993 17187
rect 21189 17153 21223 17187
rect 22845 17153 22879 17187
rect 23949 17153 23983 17187
rect 24455 17153 24489 17187
rect 26620 17153 26654 17187
rect 26893 17153 26927 17187
rect 3668 17085 3702 17119
rect 4077 17085 4111 17119
rect 6009 17085 6043 17119
rect 6101 17085 6135 17119
rect 6428 17085 6462 17119
rect 8585 17085 8619 17119
rect 10885 17085 10919 17119
rect 11253 17085 11287 17119
rect 11989 17085 12023 17119
rect 13737 17085 13771 17119
rect 13921 17085 13955 17119
rect 14013 17085 14047 17119
rect 14565 17085 14599 17119
rect 14841 17085 14875 17119
rect 16405 17085 16439 17119
rect 18705 17085 18739 17119
rect 18981 17085 19015 17119
rect 20453 17085 20487 17119
rect 20780 17085 20814 17119
rect 22661 17085 22695 17119
rect 23213 17085 23247 17119
rect 24685 17085 24719 17119
rect 26157 17085 26191 17119
rect 28457 17085 28491 17119
rect 29101 17085 29135 17119
rect 29653 17085 29687 17119
rect 29837 17085 29871 17119
rect 30573 17085 30607 17119
rect 8217 17017 8251 17051
rect 23489 17017 23523 17051
rect 30113 17017 30147 17051
rect 1415 16949 1449 16983
rect 9143 16949 9177 16983
rect 13093 16949 13127 16983
rect 16871 16949 16905 16983
rect 18245 16949 18279 16983
rect 20085 16949 20119 16983
rect 22293 16949 22327 16983
rect 24415 16949 24449 16983
rect 26623 16949 26657 16983
rect 3065 16745 3099 16779
rect 5549 16745 5583 16779
rect 6291 16745 6325 16779
rect 7665 16745 7699 16779
rect 8493 16745 8527 16779
rect 9143 16745 9177 16779
rect 10517 16745 10551 16779
rect 15669 16745 15703 16779
rect 16129 16745 16163 16779
rect 18797 16745 18831 16779
rect 23857 16745 23891 16779
rect 24599 16745 24633 16779
rect 30389 16745 30423 16779
rect 8217 16677 8251 16711
rect 23581 16677 23615 16711
rect 1133 16609 1167 16643
rect 4261 16609 4295 16643
rect 5825 16609 5859 16643
rect 6561 16609 6595 16643
rect 9413 16609 9447 16643
rect 11069 16609 11103 16643
rect 12357 16609 12391 16643
rect 14156 16609 14190 16643
rect 16313 16609 16347 16643
rect 16865 16609 16899 16643
rect 17284 16609 17318 16643
rect 17693 16609 17727 16643
rect 19349 16609 19383 16643
rect 19441 16609 19475 16643
rect 19717 16609 19751 16643
rect 21097 16609 21131 16643
rect 22017 16609 22051 16643
rect 24133 16609 24167 16643
rect 24869 16609 24903 16643
rect 27169 16609 27203 16643
rect 28641 16609 28675 16643
rect 28917 16609 28951 16643
rect 30573 16609 30607 16643
rect 1225 16541 1259 16575
rect 1552 16541 1586 16575
rect 1731 16543 1765 16577
rect 1961 16541 1995 16575
rect 3525 16541 3559 16575
rect 3852 16541 3886 16575
rect 4031 16543 4065 16577
rect 6288 16541 6322 16575
rect 8677 16541 8711 16575
rect 9173 16559 9207 16593
rect 11621 16541 11655 16575
rect 11948 16541 11982 16575
rect 12127 16541 12161 16575
rect 13829 16541 13863 16575
rect 14335 16543 14369 16577
rect 14565 16541 14599 16575
rect 16957 16541 16991 16575
rect 17453 16559 17487 16593
rect 21281 16541 21315 16575
rect 21608 16541 21642 16575
rect 21787 16541 21821 16575
rect 24596 16559 24630 16593
rect 26433 16541 26467 16575
rect 26760 16541 26794 16575
rect 26896 16543 26930 16577
rect 30021 16541 30055 16575
rect 11345 16473 11379 16507
rect 23121 16473 23155 16507
rect 25973 16473 26007 16507
rect 949 16405 983 16439
rect 13461 16405 13495 16439
rect 16681 16405 16715 16439
rect 19165 16405 19199 16439
rect 28273 16405 28307 16439
rect 2973 16201 3007 16235
rect 5641 16201 5675 16235
rect 7941 16201 7975 16235
rect 8401 16201 8435 16235
rect 13829 16201 13863 16235
rect 16405 16201 16439 16235
rect 25697 16201 25731 16235
rect 28457 16201 28491 16235
rect 30297 16201 30331 16235
rect 10517 16133 10551 16167
rect 10977 16133 11011 16167
rect 14473 16133 14507 16167
rect 20729 16133 20763 16167
rect 23213 16133 23247 16167
rect 29653 16133 29687 16167
rect 1455 16065 1489 16099
rect 4307 16065 4341 16099
rect 6597 16047 6631 16081
rect 9183 16065 9217 16099
rect 11253 16065 11287 16099
rect 11759 16065 11793 16099
rect 15028 16065 15062 16099
rect 18245 16065 18279 16099
rect 19211 16065 19245 16099
rect 21240 16065 21274 16099
rect 21419 16065 21453 16099
rect 23857 16065 23891 16099
rect 24184 16065 24218 16099
rect 24363 16065 24397 16099
rect 26392 16065 26426 16099
rect 26528 16063 26562 16097
rect 26801 16065 26835 16099
rect 29469 16065 29503 16099
rect 949 15997 983 16031
rect 1685 15997 1719 16031
rect 3801 15997 3835 16031
rect 4537 15997 4571 16031
rect 6101 15997 6135 16031
rect 6837 15997 6871 16031
rect 8585 15997 8619 16031
rect 8677 15997 8711 16031
rect 9413 15997 9447 16031
rect 11161 15997 11195 16031
rect 11989 15997 12023 16031
rect 14565 15997 14599 16031
rect 15301 15997 15335 16031
rect 16865 15997 16899 16031
rect 17141 15997 17175 16031
rect 18705 15997 18739 16031
rect 19441 15997 19475 16031
rect 20913 15997 20947 16031
rect 21649 15997 21683 16031
rect 23121 15997 23155 16031
rect 24593 15997 24627 16031
rect 26065 15997 26099 16031
rect 28273 15997 28307 16031
rect 28825 15997 28859 16031
rect 29193 15997 29227 16031
rect 29359 15975 29393 16009
rect 30021 15997 30055 16031
rect 30205 15997 30239 16031
rect 3341 15929 3375 15963
rect 13737 15929 13771 15963
rect 14289 15929 14323 15963
rect 1415 15861 1449 15895
rect 3617 15861 3651 15895
rect 4267 15861 4301 15895
rect 6567 15861 6601 15895
rect 9143 15861 9177 15895
rect 11719 15861 11753 15895
rect 13093 15861 13127 15895
rect 15031 15861 15065 15895
rect 19171 15861 19205 15895
rect 22753 15861 22787 15895
rect 27905 15861 27939 15895
rect 28641 15861 28675 15895
rect 29837 15861 29871 15895
rect 3157 15657 3191 15691
rect 10517 15657 10551 15691
rect 11437 15657 11471 15691
rect 14295 15657 14329 15691
rect 23955 15657 23989 15691
rect 28463 15657 28497 15691
rect 29837 15657 29871 15691
rect 27169 15589 27203 15623
rect 1041 15521 1075 15555
rect 5917 15521 5951 15555
rect 6796 15521 6830 15555
rect 11161 15521 11195 15555
rect 11621 15521 11655 15555
rect 11948 15521 11982 15555
rect 13829 15521 13863 15555
rect 14565 15521 14599 15555
rect 16221 15521 16255 15555
rect 17049 15521 17083 15555
rect 17468 15521 17502 15555
rect 17877 15521 17911 15555
rect 19717 15521 19751 15555
rect 21608 15521 21642 15555
rect 24225 15521 24259 15555
rect 25789 15521 25823 15555
rect 26525 15521 26559 15555
rect 26893 15521 26927 15555
rect 27629 15521 27663 15555
rect 30205 15521 30239 15555
rect 1317 15453 1351 15487
rect 1644 15453 1678 15487
rect 1813 15471 1847 15505
rect 2053 15453 2087 15487
rect 3525 15453 3559 15487
rect 3852 15453 3886 15487
rect 3988 15453 4022 15487
rect 4261 15453 4295 15487
rect 5641 15453 5675 15487
rect 6469 15453 6503 15487
rect 6965 15471 6999 15505
rect 7205 15453 7239 15487
rect 8677 15453 8711 15487
rect 9004 15453 9038 15487
rect 9140 15453 9174 15487
rect 9413 15453 9447 15487
rect 12127 15453 12161 15487
rect 12357 15453 12391 15487
rect 14335 15453 14369 15487
rect 17141 15453 17175 15487
rect 17637 15471 17671 15505
rect 19441 15453 19475 15487
rect 21281 15453 21315 15487
rect 21787 15455 21821 15489
rect 22017 15453 22051 15487
rect 23489 15453 23523 15487
rect 23985 15471 24019 15505
rect 26065 15453 26099 15487
rect 27997 15453 28031 15487
rect 28503 15453 28537 15487
rect 28733 15453 28767 15487
rect 25329 15385 25363 15419
rect 27813 15385 27847 15419
rect 30389 15385 30423 15419
rect 857 15317 891 15351
rect 6193 15317 6227 15351
rect 8309 15317 8343 15351
rect 13461 15317 13495 15351
rect 15669 15317 15703 15351
rect 16497 15317 16531 15351
rect 16865 15317 16899 15351
rect 18981 15317 19015 15351
rect 21005 15317 21039 15351
rect 23121 15317 23155 15351
rect 26709 15317 26743 15351
rect 2789 15113 2823 15147
rect 5825 15113 5859 15147
rect 13093 15113 13127 15147
rect 14289 15113 14323 15147
rect 23397 15113 23431 15147
rect 25697 15113 25731 15147
rect 26065 15113 26099 15147
rect 28549 15113 28583 15147
rect 10977 15045 11011 15079
rect 18429 15045 18463 15079
rect 26525 15045 26559 15079
rect 29837 15045 29871 15079
rect 949 14977 983 15011
rect 1455 14977 1489 15011
rect 3801 14977 3835 15011
rect 4307 14977 4341 15011
rect 6607 14977 6641 15011
rect 9004 14977 9038 15011
rect 9183 14977 9217 15011
rect 11253 14977 11287 15011
rect 11759 14977 11793 15011
rect 13553 14977 13587 15011
rect 14984 14977 15018 15011
rect 15163 14977 15197 15011
rect 17141 14977 17175 15011
rect 18889 14977 18923 15011
rect 19717 14977 19751 15011
rect 20223 14977 20257 15011
rect 22293 14977 22327 15011
rect 23857 14977 23891 15011
rect 24184 14977 24218 15011
rect 24363 14977 24397 15011
rect 27036 14977 27070 15011
rect 27215 14975 27249 15009
rect 27445 14977 27479 15011
rect 1685 14909 1719 14943
rect 3249 14909 3283 14943
rect 4128 14909 4162 14943
rect 4537 14909 4571 14943
rect 6101 14909 6135 14943
rect 6428 14909 6462 14943
rect 6837 14909 6871 14943
rect 8585 14909 8619 14943
rect 8677 14909 8711 14943
rect 9413 14909 9447 14943
rect 11161 14909 11195 14943
rect 11989 14909 12023 14943
rect 14013 14909 14047 14943
rect 14657 14909 14691 14943
rect 15393 14909 15427 14943
rect 16865 14909 16899 14943
rect 18705 14909 18739 14943
rect 19441 14909 19475 14943
rect 20453 14909 20487 14943
rect 22017 14909 22051 14943
rect 24593 14909 24627 14943
rect 26249 14909 26283 14943
rect 26341 14909 26375 14943
rect 26709 14909 26743 14943
rect 29101 14909 29135 14943
rect 29653 14909 29687 14943
rect 30205 14909 30239 14943
rect 30389 14909 30423 14943
rect 3525 14841 3559 14875
rect 14197 14841 14231 14875
rect 1415 14773 1449 14807
rect 7941 14773 7975 14807
rect 8401 14773 8435 14807
rect 10517 14773 10551 14807
rect 11719 14773 11753 14807
rect 13829 14773 13863 14807
rect 16497 14773 16531 14807
rect 19257 14773 19291 14807
rect 20183 14773 20217 14807
rect 21557 14773 21591 14807
rect 29193 14773 29227 14807
rect 4077 14569 4111 14603
rect 4629 14569 4663 14603
rect 5181 14569 5215 14603
rect 5457 14569 5491 14603
rect 6285 14569 6319 14603
rect 6561 14569 6595 14603
rect 9137 14569 9171 14603
rect 9413 14569 9447 14603
rect 10517 14569 10551 14603
rect 11069 14569 11103 14603
rect 11345 14569 11379 14603
rect 12087 14569 12121 14603
rect 13461 14569 13495 14603
rect 18521 14569 18555 14603
rect 22115 14569 22149 14603
rect 25697 14569 25731 14603
rect 28463 14569 28497 14603
rect 29837 14569 29871 14603
rect 1225 14501 1259 14535
rect 10057 14501 10091 14535
rect 15945 14501 15979 14535
rect 19073 14501 19107 14535
rect 21097 14501 21131 14535
rect 23765 14501 23799 14535
rect 26985 14501 27019 14535
rect 27353 14501 27387 14535
rect 27721 14501 27755 14535
rect 949 14433 983 14467
rect 2237 14433 2271 14467
rect 3985 14433 4019 14467
rect 4261 14433 4295 14467
rect 4537 14433 4571 14467
rect 4813 14433 4847 14467
rect 5089 14433 5123 14467
rect 5365 14433 5399 14467
rect 5641 14433 5675 14467
rect 6193 14433 6227 14467
rect 6469 14433 6503 14467
rect 6745 14433 6779 14467
rect 9321 14433 9355 14467
rect 9597 14433 9631 14467
rect 9873 14433 9907 14467
rect 10701 14433 10735 14467
rect 11253 14433 11287 14467
rect 11529 14433 11563 14467
rect 13829 14433 13863 14467
rect 16129 14433 16163 14467
rect 17008 14433 17042 14467
rect 17417 14433 17451 14467
rect 23857 14433 23891 14467
rect 24184 14433 24218 14467
rect 26241 14433 26275 14467
rect 26617 14433 26651 14467
rect 26719 14433 26753 14467
rect 27997 14433 28031 14467
rect 30389 14433 30423 14467
rect 1501 14365 1535 14399
rect 1828 14365 1862 14399
rect 2007 14367 2041 14401
rect 6837 14365 6871 14399
rect 7164 14365 7198 14399
rect 7300 14365 7334 14399
rect 7573 14365 7607 14399
rect 10333 14365 10367 14399
rect 11621 14365 11655 14399
rect 12127 14365 12161 14399
rect 12357 14365 12391 14399
rect 14156 14365 14190 14399
rect 14335 14365 14369 14399
rect 14565 14365 14599 14399
rect 16681 14365 16715 14399
rect 17187 14365 17221 14399
rect 19441 14365 19475 14399
rect 19717 14365 19751 14399
rect 21649 14365 21683 14399
rect 22128 14365 22162 14399
rect 22385 14365 22419 14399
rect 24353 14383 24387 14417
rect 24593 14365 24627 14399
rect 28460 14365 28494 14399
rect 28733 14365 28767 14399
rect 3801 14297 3835 14331
rect 4905 14297 4939 14331
rect 6009 14297 6043 14331
rect 9689 14297 9723 14331
rect 30205 14297 30239 14331
rect 3525 14229 3559 14263
rect 4353 14229 4387 14263
rect 8861 14229 8895 14263
rect 16313 14229 16347 14263
rect 21465 14229 21499 14263
rect 26065 14229 26099 14263
rect 26433 14229 26467 14263
rect 5917 14025 5951 14059
rect 12449 14025 12483 14059
rect 13001 14025 13035 14059
rect 13921 14025 13955 14059
rect 18245 14025 18279 14059
rect 19073 14025 19107 14059
rect 22477 14025 22511 14059
rect 26525 14025 26559 14059
rect 29009 14025 29043 14059
rect 29285 14025 29319 14059
rect 29561 14025 29595 14059
rect 29837 14025 29871 14059
rect 30297 14025 30331 14059
rect 8953 13957 8987 13991
rect 12725 13957 12759 13991
rect 13645 13957 13679 13991
rect 16037 13957 16071 13991
rect 19533 13957 19567 13991
rect 22201 13957 22235 13991
rect 22753 13957 22787 13991
rect 28549 13957 28583 13991
rect 30573 13957 30607 13991
rect 949 13889 983 13923
rect 1455 13889 1489 13923
rect 3893 13889 3927 13923
rect 4356 13889 4390 13923
rect 6428 13889 6462 13923
rect 6607 13889 6641 13923
rect 8585 13889 8619 13923
rect 10152 13889 10186 13923
rect 12081 13889 12115 13923
rect 14660 13887 14694 13921
rect 14933 13889 14967 13923
rect 16732 13889 16766 13923
rect 16911 13889 16945 13923
rect 20499 13887 20533 13921
rect 22109 13889 22143 13923
rect 25007 13889 25041 13923
rect 25237 13889 25271 13923
rect 26709 13889 26743 13923
rect 27172 13889 27206 13923
rect 1685 13821 1719 13855
rect 3065 13821 3099 13855
rect 3525 13821 3559 13855
rect 3801 13797 3835 13831
rect 4629 13821 4663 13855
rect 6101 13821 6135 13855
rect 6837 13821 6871 13855
rect 8401 13821 8435 13855
rect 9137 13821 9171 13855
rect 9689 13821 9723 13855
rect 10016 13821 10050 13855
rect 10425 13821 10459 13855
rect 11897 13821 11931 13855
rect 12633 13821 12667 13855
rect 12909 13821 12943 13855
rect 13185 13821 13219 13855
rect 13829 13821 13863 13855
rect 14105 13821 14139 13855
rect 14197 13821 14231 13855
rect 16405 13821 16439 13855
rect 17141 13821 17175 13855
rect 19441 13821 19475 13855
rect 19717 13821 19751 13855
rect 19993 13821 20027 13855
rect 20729 13821 20763 13855
rect 22385 13821 22419 13855
rect 22661 13821 22695 13855
rect 22937 13821 22971 13855
rect 23213 13821 23247 13855
rect 23397 13821 23431 13855
rect 24041 13821 24075 13855
rect 24317 13821 24351 13855
rect 24501 13821 24535 13855
rect 27445 13821 27479 13855
rect 29193 13821 29227 13855
rect 29469 13821 29503 13855
rect 29745 13821 29779 13855
rect 30021 13821 30055 13855
rect 30113 13821 30147 13855
rect 30389 13821 30423 13855
rect 9229 13753 9263 13787
rect 11805 13753 11839 13787
rect 18797 13753 18831 13787
rect 1415 13685 1449 13719
rect 3341 13685 3375 13719
rect 3617 13685 3651 13719
rect 4359 13685 4393 13719
rect 7941 13685 7975 13719
rect 14663 13685 14697 13719
rect 19257 13685 19291 13719
rect 20459 13685 20493 13719
rect 23029 13685 23063 13719
rect 23581 13685 23615 13719
rect 23857 13685 23891 13719
rect 24133 13685 24167 13719
rect 24967 13685 25001 13719
rect 27175 13685 27209 13719
rect 1783 13481 1817 13515
rect 3991 13481 4025 13515
rect 5825 13481 5859 13515
rect 6101 13481 6135 13515
rect 7303 13481 7337 13515
rect 9045 13481 9079 13515
rect 9505 13481 9539 13515
rect 11161 13481 11195 13515
rect 16129 13481 16163 13515
rect 18981 13481 19015 13515
rect 21557 13481 21591 13515
rect 23949 13481 23983 13515
rect 28273 13481 28307 13515
rect 9597 13413 9631 13447
rect 15025 13413 15059 13447
rect 1225 13345 1259 13379
rect 1317 13345 1351 13379
rect 2053 13345 2087 13379
rect 3525 13345 3559 13379
rect 6009 13345 6043 13379
rect 6285 13345 6319 13379
rect 6745 13345 6779 13379
rect 6837 13345 6871 13379
rect 9321 13345 9355 13379
rect 9873 13345 9907 13379
rect 10149 13345 10183 13379
rect 10425 13329 10459 13363
rect 10977 13345 11011 13379
rect 11805 13345 11839 13379
rect 12081 13345 12115 13379
rect 14749 13345 14783 13379
rect 15393 13345 15427 13379
rect 16313 13345 16347 13379
rect 16497 13345 16531 13379
rect 17468 13345 17502 13379
rect 17877 13345 17911 13379
rect 21465 13345 21499 13379
rect 21741 13345 21775 13379
rect 21925 13345 21959 13379
rect 22252 13345 22286 13379
rect 24133 13345 24167 13379
rect 24869 13345 24903 13379
rect 26249 13345 26283 13379
rect 27169 13345 27203 13379
rect 30573 13345 30607 13379
rect 1823 13277 1857 13311
rect 3433 13277 3467 13311
rect 3988 13277 4022 13311
rect 4261 13277 4295 13311
rect 5641 13277 5675 13311
rect 7300 13277 7334 13311
rect 7573 13277 7607 13311
rect 11253 13277 11287 13311
rect 11529 13277 11563 13311
rect 12449 13277 12483 13311
rect 12776 13277 12810 13311
rect 12912 13279 12946 13313
rect 13185 13277 13219 13311
rect 17141 13277 17175 13311
rect 17647 13277 17681 13311
rect 19441 13277 19475 13311
rect 19717 13277 19751 13311
rect 21097 13277 21131 13311
rect 22388 13277 22422 13311
rect 22661 13277 22695 13311
rect 24460 13277 24494 13311
rect 24596 13279 24630 13313
rect 26433 13277 26467 13311
rect 26760 13277 26794 13311
rect 26896 13279 26930 13313
rect 28641 13277 28675 13311
rect 28917 13277 28951 13311
rect 8861 13209 8895 13243
rect 10057 13209 10091 13243
rect 10333 13209 10367 13243
rect 11989 13209 12023 13243
rect 30389 13209 30423 13243
rect 1041 13141 1075 13175
rect 6561 13141 6595 13175
rect 10609 13141 10643 13175
rect 12265 13141 12299 13175
rect 14289 13141 14323 13175
rect 15485 13141 15519 13175
rect 16681 13141 16715 13175
rect 21281 13141 21315 13175
rect 30021 13141 30055 13175
rect 2973 12937 3007 12971
rect 5917 12937 5951 12971
rect 8769 12937 8803 12971
rect 12081 12937 12115 12971
rect 12173 12937 12207 12971
rect 22201 12937 22235 12971
rect 22753 12937 22787 12971
rect 25697 12937 25731 12971
rect 29929 12937 29963 12971
rect 30389 12937 30423 12971
rect 3249 12869 3283 12903
rect 3617 12869 3651 12903
rect 8585 12869 8619 12903
rect 9045 12869 9079 12903
rect 12633 12869 12667 12903
rect 13185 12869 13219 12903
rect 18429 12869 18463 12903
rect 19717 12869 19751 12903
rect 22017 12869 22051 12903
rect 949 12801 983 12835
rect 1455 12799 1489 12833
rect 1685 12801 1719 12835
rect 4356 12801 4390 12835
rect 6564 12801 6598 12835
rect 6837 12801 6871 12835
rect 9689 12801 9723 12835
rect 10152 12801 10186 12835
rect 14059 12799 14093 12833
rect 16868 12801 16902 12835
rect 19993 12801 20027 12835
rect 20456 12801 20490 12835
rect 24320 12801 24354 12835
rect 26528 12801 26562 12835
rect 26801 12801 26835 12835
rect 3433 12733 3467 12767
rect 3801 12733 3835 12767
rect 3893 12733 3927 12767
rect 4629 12733 4663 12767
rect 6101 12733 6135 12767
rect 8401 12733 8435 12767
rect 8953 12733 8987 12767
rect 9229 12733 9263 12767
rect 10425 12733 10459 12767
rect 11897 12733 11931 12767
rect 12357 12733 12391 12767
rect 12817 12733 12851 12767
rect 13093 12733 13127 12767
rect 13369 12733 13403 12767
rect 13553 12733 13587 12767
rect 14289 12733 14323 12767
rect 16405 12733 16439 12767
rect 17141 12733 17175 12767
rect 19073 12733 19107 12767
rect 19349 12733 19383 12767
rect 19625 12733 19659 12767
rect 19901 12733 19935 12767
rect 20729 12733 20763 12767
rect 22385 12733 22419 12767
rect 22937 12733 22971 12767
rect 23397 12733 23431 12767
rect 23673 12733 23707 12767
rect 23857 12733 23891 12767
rect 24593 12733 24627 12767
rect 26065 12733 26099 12767
rect 28365 12733 28399 12767
rect 29469 12733 29503 12767
rect 30113 12733 30147 12767
rect 30573 12733 30607 12767
rect 8217 12665 8251 12699
rect 15669 12665 15703 12699
rect 16313 12665 16347 12699
rect 29101 12665 29135 12699
rect 29653 12665 29687 12699
rect 1415 12597 1449 12631
rect 4359 12597 4393 12631
rect 6567 12597 6601 12631
rect 9321 12597 9355 12631
rect 10155 12597 10189 12631
rect 11713 12597 11747 12631
rect 12909 12597 12943 12631
rect 14019 12597 14053 12631
rect 16871 12597 16905 12631
rect 18889 12597 18923 12631
rect 19165 12597 19199 12631
rect 19441 12597 19475 12631
rect 20459 12597 20493 12631
rect 23213 12597 23247 12631
rect 23489 12597 23523 12631
rect 24323 12597 24357 12631
rect 26531 12597 26565 12631
rect 27905 12597 27939 12631
rect 28457 12597 28491 12631
rect 29745 12597 29779 12631
rect 3991 12393 4025 12427
rect 5549 12393 5583 12427
rect 11253 12393 11287 12427
rect 15393 12393 15427 12427
rect 16313 12393 16347 12427
rect 16681 12393 16715 12427
rect 19993 12393 20027 12427
rect 20269 12393 20303 12427
rect 20729 12393 20763 12427
rect 21747 12393 21781 12427
rect 23121 12393 23155 12427
rect 25513 12393 25547 12427
rect 28273 12393 28307 12427
rect 30389 12393 30423 12427
rect 14933 12325 14967 12359
rect 1225 12257 1259 12291
rect 1317 12257 1351 12291
rect 1644 12257 1678 12291
rect 3433 12257 3467 12291
rect 6009 12257 6043 12291
rect 6285 12257 6319 12291
rect 6469 12257 6503 12291
rect 7205 12257 7239 12291
rect 9004 12257 9038 12291
rect 11161 12257 11195 12291
rect 11437 12257 11471 12291
rect 11713 12257 11747 12291
rect 11989 12257 12023 12291
rect 12357 12257 12391 12291
rect 12449 12257 12483 12291
rect 12776 12257 12810 12291
rect 13185 12257 13219 12291
rect 14657 12257 14691 12291
rect 17233 12257 17267 12291
rect 17417 12257 17451 12291
rect 17693 12257 17727 12291
rect 18296 12257 18330 12291
rect 18705 12257 18739 12291
rect 20453 12257 20487 12291
rect 20913 12257 20947 12291
rect 22017 12257 22051 12291
rect 23489 12257 23523 12291
rect 23816 12257 23850 12291
rect 24225 12257 24259 12291
rect 25789 12257 25823 12291
rect 26433 12257 26467 12291
rect 27169 12257 27203 12291
rect 28917 12257 28951 12291
rect 30573 12257 30607 12291
rect 1813 12207 1847 12241
rect 2053 12189 2087 12223
rect 3525 12189 3559 12223
rect 3988 12189 4022 12223
rect 4261 12189 4295 12223
rect 6796 12189 6830 12223
rect 6932 12189 6966 12223
rect 8677 12189 8711 12223
rect 9140 12189 9174 12223
rect 9413 12189 9447 12223
rect 12912 12189 12946 12223
rect 15853 12189 15887 12223
rect 17969 12189 18003 12223
rect 18432 12189 18466 12223
rect 21281 12189 21315 12223
rect 21787 12189 21821 12223
rect 23952 12189 23986 12223
rect 26760 12189 26794 12223
rect 26896 12189 26930 12223
rect 28641 12189 28675 12223
rect 5825 12121 5859 12155
rect 10701 12121 10735 12155
rect 11529 12121 11563 12155
rect 1041 12053 1075 12087
rect 6101 12053 6135 12087
rect 8493 12053 8527 12087
rect 10977 12053 11011 12087
rect 11805 12053 11839 12087
rect 12173 12053 12207 12087
rect 14289 12053 14323 12087
rect 17049 12053 17083 12087
rect 26065 12053 26099 12087
rect 30021 12053 30055 12087
rect 8033 11849 8067 11883
rect 8861 11849 8895 11883
rect 9137 11849 9171 11883
rect 9413 11849 9447 11883
rect 11529 11849 11563 11883
rect 12357 11849 12391 11883
rect 12817 11849 12851 11883
rect 18429 11849 18463 11883
rect 20545 11849 20579 11883
rect 23581 11849 23615 11883
rect 26525 11849 26559 11883
rect 28733 11849 28767 11883
rect 13369 11781 13403 11815
rect 30113 11781 30147 11815
rect 1455 11713 1489 11747
rect 3065 11713 3099 11747
rect 3804 11713 3838 11747
rect 4077 11713 4111 11747
rect 5457 11713 5491 11747
rect 6012 11711 6046 11745
rect 10152 11713 10186 11747
rect 10425 11713 10459 11747
rect 13880 11713 13914 11747
rect 14059 11713 14093 11747
rect 14289 11713 14323 11747
rect 16911 11711 16945 11745
rect 17141 11713 17175 11747
rect 18705 11713 18739 11747
rect 19168 11713 19202 11747
rect 19441 11713 19475 11747
rect 21557 11713 21591 11747
rect 22063 11713 22097 11747
rect 24225 11713 24259 11747
rect 24501 11713 24535 11747
rect 25007 11713 25041 11747
rect 26709 11713 26743 11747
rect 27215 11713 27249 11747
rect 27445 11713 27479 11747
rect 949 11645 983 11679
rect 1685 11645 1719 11679
rect 3341 11645 3375 11679
rect 5549 11645 5583 11679
rect 6285 11645 6319 11679
rect 7941 11645 7975 11679
rect 8217 11645 8251 11679
rect 8677 11645 8711 11679
rect 8953 11645 8987 11679
rect 9229 11645 9263 11679
rect 9689 11645 9723 11679
rect 12081 11645 12115 11679
rect 13001 11645 13035 11679
rect 13185 11645 13219 11679
rect 13553 11645 13587 11679
rect 16313 11645 16347 11679
rect 16405 11645 16439 11679
rect 22293 11645 22327 11679
rect 23949 11645 23983 11679
rect 25237 11645 25271 11679
rect 29469 11645 29503 11679
rect 29561 11645 29595 11679
rect 30297 11645 30331 11679
rect 30573 11645 30607 11679
rect 8401 11577 8435 11611
rect 29101 11577 29135 11611
rect 29837 11577 29871 11611
rect 1415 11509 1449 11543
rect 3807 11509 3841 11543
rect 6015 11509 6049 11543
rect 7389 11509 7423 11543
rect 7757 11509 7791 11543
rect 10155 11509 10189 11543
rect 11897 11509 11931 11543
rect 15393 11509 15427 11543
rect 15945 11509 15979 11543
rect 16129 11509 16163 11543
rect 16871 11509 16905 11543
rect 19171 11509 19205 11543
rect 21097 11509 21131 11543
rect 22023 11509 22057 11543
rect 24967 11509 25001 11543
rect 27175 11509 27209 11543
rect 30389 11509 30423 11543
rect 1409 11305 1443 11339
rect 1967 11305 2001 11339
rect 3525 11305 3559 11339
rect 4813 11305 4847 11339
rect 5457 11305 5491 11339
rect 5825 11305 5859 11339
rect 8861 11305 8895 11339
rect 9689 11305 9723 11339
rect 10241 11305 10275 11339
rect 15761 11305 15795 11339
rect 16681 11305 16715 11339
rect 18797 11305 18831 11339
rect 21005 11305 21039 11339
rect 22207 11305 22241 11339
rect 24415 11305 24449 11339
rect 25789 11305 25823 11339
rect 3985 11237 4019 11271
rect 12265 11237 12299 11271
rect 1501 11169 1535 11203
rect 2237 11169 2271 11203
rect 3709 11169 3743 11203
rect 4445 11169 4479 11203
rect 4721 11169 4755 11203
rect 5365 11169 5399 11203
rect 5641 11169 5675 11203
rect 6009 11169 6043 11203
rect 6377 11169 6411 11203
rect 7164 11169 7198 11203
rect 7573 11169 7607 11203
rect 9045 11169 9079 11203
rect 9597 11169 9631 11203
rect 10425 11169 10459 11203
rect 10701 11169 10735 11203
rect 11161 11169 11195 11203
rect 11437 11169 11471 11203
rect 11713 11169 11747 11203
rect 11989 11169 12023 11203
rect 13185 11169 13219 11203
rect 14841 11169 14875 11203
rect 15117 11169 15151 11203
rect 17509 11169 17543 11203
rect 19308 11169 19342 11203
rect 19717 11169 19751 11203
rect 21465 11169 21499 11203
rect 23857 11169 23891 11203
rect 26760 11169 26794 11203
rect 28641 11169 28675 11203
rect 28917 11169 28951 11203
rect 30573 11169 30607 11203
rect 2007 11101 2041 11135
rect 6837 11101 6871 11135
rect 7300 11103 7334 11137
rect 12449 11101 12483 11135
rect 12776 11101 12810 11135
rect 12912 11103 12946 11137
rect 16773 11101 16807 11135
rect 17100 11101 17134 11135
rect 17279 11101 17313 11135
rect 18981 11101 19015 11135
rect 19444 11101 19478 11135
rect 21741 11101 21775 11135
rect 22247 11101 22281 11135
rect 22477 11101 22511 11135
rect 23949 11101 23983 11135
rect 24412 11101 24446 11135
rect 24685 11101 24719 11135
rect 26433 11101 26467 11135
rect 26896 11101 26930 11135
rect 27169 11101 27203 11135
rect 5181 11033 5215 11067
rect 9229 11033 9263 11067
rect 10517 11033 10551 11067
rect 10977 11033 11011 11067
rect 11253 11033 11287 11067
rect 11805 11033 11839 11067
rect 14657 11033 14691 11067
rect 14933 11033 14967 11067
rect 15485 11033 15519 11067
rect 28273 11033 28307 11067
rect 30021 11033 30055 11067
rect 30389 11033 30423 11067
rect 4261 10965 4295 10999
rect 6469 10965 6503 10999
rect 11529 10965 11563 10999
rect 14289 10965 14323 10999
rect 21281 10965 21315 10999
rect 5273 10761 5307 10795
rect 8125 10761 8159 10795
rect 16037 10761 16071 10795
rect 19257 10761 19291 10795
rect 21741 10761 21775 10795
rect 26617 10761 26651 10795
rect 28641 10761 28675 10795
rect 19073 10693 19107 10727
rect 949 10625 983 10659
rect 1455 10623 1489 10657
rect 3065 10625 3099 10659
rect 3712 10625 3746 10659
rect 6012 10625 6046 10659
rect 9689 10625 9723 10659
rect 10016 10625 10050 10659
rect 10152 10625 10186 10659
rect 10425 10625 10459 10659
rect 11805 10625 11839 10659
rect 14059 10625 14093 10659
rect 16901 10607 16935 10641
rect 19533 10625 19567 10659
rect 20039 10623 20073 10657
rect 21649 10625 21683 10659
rect 22017 10625 22051 10659
rect 23489 10625 23523 10659
rect 24920 10625 24954 10659
rect 25099 10625 25133 10659
rect 26801 10625 26835 10659
rect 1685 10557 1719 10591
rect 3249 10557 3283 10591
rect 3985 10557 4019 10591
rect 5549 10557 5583 10591
rect 6285 10557 6319 10591
rect 7941 10557 7975 10591
rect 8401 10557 8435 10591
rect 8861 10557 8895 10591
rect 9597 10533 9631 10567
rect 12449 10557 12483 10591
rect 13369 10557 13403 10591
rect 13553 10557 13587 10591
rect 14289 10557 14323 10591
rect 16405 10557 16439 10591
rect 17141 10557 17175 10591
rect 19441 10557 19475 10591
rect 20269 10557 20303 10591
rect 21925 10557 21959 10591
rect 22293 10557 22327 10591
rect 23949 10557 23983 10591
rect 24593 10557 24627 10591
rect 25329 10557 25363 10591
rect 27077 10557 27111 10591
rect 28825 10557 28859 10591
rect 30113 10557 30147 10591
rect 7665 10489 7699 10523
rect 9137 10489 9171 10523
rect 11989 10489 12023 10523
rect 18521 10489 18555 10523
rect 18797 10489 18831 10523
rect 29101 10489 29135 10523
rect 29653 10489 29687 10523
rect 1415 10421 1449 10455
rect 3715 10421 3749 10455
rect 6015 10421 6049 10455
rect 8585 10421 8619 10455
rect 9413 10421 9447 10455
rect 12081 10421 12115 10455
rect 12633 10421 12667 10455
rect 12909 10421 12943 10455
rect 13185 10421 13219 10455
rect 14019 10421 14053 10455
rect 15393 10421 15427 10455
rect 16871 10421 16905 10455
rect 19999 10421 20033 10455
rect 24041 10421 24075 10455
rect 28181 10421 28215 10455
rect 29193 10421 29227 10455
rect 29745 10421 29779 10455
rect 30297 10421 30331 10455
rect 1599 10217 1633 10251
rect 3807 10217 3841 10251
rect 6935 10217 6969 10251
rect 13369 10217 13403 10251
rect 16865 10217 16899 10251
rect 17607 10217 17641 10251
rect 19165 10217 19199 10251
rect 19993 10217 20027 10251
rect 21005 10217 21039 10251
rect 23121 10217 23155 10251
rect 23489 10217 23523 10251
rect 23857 10217 23891 10251
rect 30021 10217 30055 10251
rect 5457 10149 5491 10183
rect 6193 10149 6227 10183
rect 19625 10149 19659 10183
rect 1041 10081 1075 10115
rect 3249 10081 3283 10115
rect 4077 10081 4111 10115
rect 5917 10081 5951 10115
rect 6469 10081 6503 10115
rect 8585 10081 8619 10115
rect 9413 10081 9447 10115
rect 11713 10081 11747 10115
rect 13277 10081 13311 10115
rect 13553 10081 13587 10115
rect 15953 10081 15987 10115
rect 16313 10081 16347 10115
rect 16773 10081 16807 10115
rect 17049 10081 17083 10115
rect 17877 10081 17911 10115
rect 19349 10081 19383 10115
rect 20177 10081 20211 10115
rect 20453 10081 20487 10115
rect 21608 10081 21642 10115
rect 22017 10081 22051 10115
rect 23673 10081 23707 10115
rect 24041 10081 24075 10115
rect 24460 10081 24494 10115
rect 26249 10081 26283 10115
rect 28641 10081 28675 10115
rect 28917 10081 28951 10115
rect 30573 10081 30607 10115
rect 1133 10013 1167 10047
rect 1639 10013 1673 10047
rect 1869 10013 1903 10047
rect 3341 10013 3375 10047
rect 3804 10013 3838 10047
rect 6975 10013 7009 10047
rect 7205 10013 7239 10047
rect 8677 10013 8711 10047
rect 9004 10013 9038 10047
rect 9140 10013 9174 10047
rect 10977 10013 11011 10047
rect 11304 10013 11338 10047
rect 11440 10013 11474 10047
rect 13880 10013 13914 10047
rect 14032 10015 14066 10049
rect 14289 10013 14323 10047
rect 17141 10013 17175 10047
rect 17647 10013 17681 10047
rect 21281 10013 21315 10047
rect 21744 10013 21778 10047
rect 24133 10013 24167 10047
rect 24612 10013 24646 10047
rect 24869 10013 24903 10047
rect 26433 10013 26467 10047
rect 26760 10013 26794 10047
rect 26896 10013 26930 10047
rect 27169 10013 27203 10047
rect 15761 9945 15795 9979
rect 857 9877 891 9911
rect 10701 9877 10735 9911
rect 12817 9877 12851 9911
rect 15393 9877 15427 9911
rect 16129 9877 16163 9911
rect 16589 9877 16623 9911
rect 28273 9877 28307 9911
rect 30389 9877 30423 9911
rect 5825 9673 5859 9707
rect 25697 9673 25731 9707
rect 28273 9673 28307 9707
rect 18245 9605 18279 9639
rect 20545 9605 20579 9639
rect 22753 9605 22787 9639
rect 23213 9605 23247 9639
rect 23489 9605 23523 9639
rect 28549 9605 28583 9639
rect 30021 9605 30055 9639
rect 949 9537 983 9571
rect 1455 9537 1489 9571
rect 3065 9537 3099 9571
rect 4080 9537 4114 9571
rect 6607 9537 6641 9571
rect 8585 9537 8619 9571
rect 9091 9537 9125 9571
rect 10701 9537 10735 9571
rect 11120 9537 11154 9571
rect 11256 9537 11290 9571
rect 13553 9537 13587 9571
rect 14016 9535 14050 9569
rect 14289 9537 14323 9571
rect 16868 9537 16902 9571
rect 19211 9537 19245 9571
rect 21376 9535 21410 9569
rect 21649 9537 21683 9571
rect 23857 9537 23891 9571
rect 24363 9537 24397 9571
rect 26528 9537 26562 9571
rect 1685 9469 1719 9503
rect 3617 9469 3651 9503
rect 3944 9469 3978 9503
rect 4353 9469 4387 9503
rect 6009 9469 6043 9503
rect 6101 9469 6135 9503
rect 6837 9469 6871 9503
rect 9321 9469 9355 9503
rect 10793 9469 10827 9503
rect 11529 9469 11563 9503
rect 13093 9469 13127 9503
rect 15761 9469 15795 9503
rect 16405 9469 16439 9503
rect 17141 9469 17175 9503
rect 18705 9469 18739 9503
rect 19441 9469 19475 9503
rect 20913 9469 20947 9503
rect 23397 9469 23431 9503
rect 23673 9469 23707 9503
rect 24593 9469 24627 9503
rect 26065 9469 26099 9503
rect 26801 9469 26835 9503
rect 28457 9469 28491 9503
rect 28733 9469 28767 9503
rect 29193 9469 29227 9503
rect 30205 9469 30239 9503
rect 30481 9469 30515 9503
rect 5733 9401 5767 9435
rect 8217 9401 8251 9435
rect 13277 9401 13311 9435
rect 15669 9401 15703 9435
rect 16037 9401 16071 9435
rect 1415 9333 1449 9367
rect 3525 9333 3559 9367
rect 6567 9333 6601 9367
rect 9051 9333 9085 9367
rect 12633 9333 12667 9367
rect 14019 9333 14053 9367
rect 16871 9333 16905 9367
rect 19171 9333 19205 9367
rect 21379 9333 21413 9367
rect 24323 9333 24357 9367
rect 26531 9333 26565 9367
rect 27905 9333 27939 9367
rect 29009 9333 29043 9367
rect 30297 9333 30331 9367
rect 1317 9129 1351 9163
rect 2887 9129 2921 9163
rect 4629 9129 4663 9163
rect 7297 9129 7331 9163
rect 8039 9129 8073 9163
rect 9413 9129 9447 9163
rect 10333 9129 10367 9163
rect 13369 9129 13403 9163
rect 14019 9129 14053 9163
rect 16589 9129 16623 9163
rect 17331 9129 17365 9163
rect 18705 9129 18739 9163
rect 19073 9129 19107 9163
rect 20269 9129 20303 9163
rect 21281 9129 21315 9163
rect 24961 9129 24995 9163
rect 25697 9129 25731 9163
rect 25973 9129 26007 9163
rect 30021 9129 30055 9163
rect 30389 9129 30423 9163
rect 1041 9061 1075 9095
rect 4537 9061 4571 9095
rect 20637 9061 20671 9095
rect 1685 8993 1719 9027
rect 2421 8993 2455 9027
rect 4813 8993 4847 9027
rect 5089 8993 5123 9027
rect 5373 8993 5407 9027
rect 5641 8993 5675 9027
rect 6009 8993 6043 9027
rect 6377 8993 6411 9027
rect 6653 8993 6687 9027
rect 6929 8993 6963 9027
rect 7205 8993 7239 9027
rect 7481 8993 7515 9027
rect 9873 8993 9907 9027
rect 10517 8993 10551 9027
rect 10793 8993 10827 9027
rect 11304 8993 11338 9027
rect 11713 8993 11747 9027
rect 13185 8993 13219 9027
rect 13553 8993 13587 9027
rect 14289 8993 14323 9027
rect 15945 8993 15979 9027
rect 16773 8993 16807 9027
rect 17601 8993 17635 9027
rect 19257 8993 19291 9027
rect 19533 8993 19567 9027
rect 20361 8993 20395 9027
rect 21465 8993 21499 9027
rect 22201 8993 22235 9027
rect 22477 8993 22511 9027
rect 22937 8993 22971 9027
rect 23264 8993 23298 9027
rect 25329 8993 25363 9027
rect 25605 8993 25639 9027
rect 25881 8993 25915 9027
rect 26157 8993 26191 9027
rect 26433 8993 26467 9027
rect 28641 8993 28675 9027
rect 28917 8993 28951 9027
rect 30573 8993 30607 9027
rect 1869 8925 1903 8959
rect 2927 8927 2961 8961
rect 3157 8925 3191 8959
rect 7573 8925 7607 8959
rect 8036 8943 8070 8977
rect 8309 8925 8343 8959
rect 10977 8925 11011 8959
rect 11440 8927 11474 8961
rect 14059 8925 14093 8959
rect 16865 8925 16899 8959
rect 17371 8925 17405 8959
rect 23443 8925 23477 8959
rect 23673 8925 23707 8959
rect 26760 8925 26794 8959
rect 26939 8925 26973 8959
rect 27169 8925 27203 8959
rect 5457 8857 5491 8891
rect 6193 8857 6227 8891
rect 6745 8857 6779 8891
rect 10609 8857 10643 8891
rect 15761 8857 15795 8891
rect 19901 8857 19935 8891
rect 22661 8857 22695 8891
rect 25145 8857 25179 8891
rect 4905 8789 4939 8823
rect 5181 8789 5215 8823
rect 5825 8789 5859 8823
rect 6469 8789 6503 8823
rect 7021 8789 7055 8823
rect 10149 8789 10183 8823
rect 12817 8789 12851 8823
rect 15577 8789 15611 8823
rect 16405 8789 16439 8823
rect 19349 8789 19383 8823
rect 22017 8789 22051 8823
rect 25421 8789 25455 8823
rect 28273 8789 28307 8823
rect 2789 8585 2823 8619
rect 7389 8585 7423 8619
rect 8033 8585 8067 8619
rect 8401 8585 8435 8619
rect 11529 8585 11563 8619
rect 12081 8585 12115 8619
rect 13369 8585 13403 8619
rect 17601 8585 17635 8619
rect 20729 8585 20763 8619
rect 25881 8585 25915 8619
rect 26065 8585 26099 8619
rect 28549 8585 28583 8619
rect 30297 8585 30331 8619
rect 5089 8517 5123 8551
rect 7757 8517 7791 8551
rect 12817 8517 12851 8551
rect 13093 8517 13127 8551
rect 15393 8517 15427 8551
rect 29837 8517 29871 8551
rect 1455 8449 1489 8483
rect 3712 8449 3746 8483
rect 5549 8449 5583 8483
rect 6012 8449 6046 8483
rect 9968 8449 10002 8483
rect 10241 8449 10275 8483
rect 13553 8449 13587 8483
rect 13880 8449 13914 8483
rect 14059 8449 14093 8483
rect 16224 8449 16258 8483
rect 18705 8449 18739 8483
rect 19032 8449 19066 8483
rect 19168 8449 19202 8483
rect 19441 8449 19475 8483
rect 22063 8449 22097 8483
rect 22293 8449 22327 8483
rect 23673 8449 23707 8483
rect 24320 8449 24354 8483
rect 24593 8449 24627 8483
rect 27036 8449 27070 8483
rect 27215 8449 27249 8483
rect 949 8381 983 8415
rect 1276 8381 1310 8415
rect 1685 8381 1719 8415
rect 3249 8381 3283 8415
rect 3576 8381 3610 8415
rect 3985 8381 4019 8415
rect 6285 8381 6319 8415
rect 7941 8381 7975 8415
rect 8217 8381 8251 8415
rect 8585 8381 8619 8415
rect 9045 8381 9079 8415
rect 9321 8381 9355 8415
rect 9505 8381 9539 8415
rect 9832 8381 9866 8415
rect 12357 8381 12391 8415
rect 12633 8381 12667 8415
rect 12909 8381 12943 8415
rect 13185 8381 13219 8415
rect 14289 8381 14323 8415
rect 15761 8381 15795 8415
rect 16497 8381 16531 8415
rect 18061 8381 18095 8415
rect 18429 8381 18463 8415
rect 21557 8381 21591 8415
rect 23857 8381 23891 8415
rect 24184 8381 24218 8415
rect 26249 8381 26283 8415
rect 26709 8381 26743 8415
rect 27445 8381 27479 8415
rect 29101 8381 29135 8415
rect 29653 8381 29687 8415
rect 30113 8381 30147 8415
rect 11805 8313 11839 8347
rect 6015 8245 6049 8279
rect 8861 8245 8895 8279
rect 9137 8245 9171 8279
rect 12449 8245 12483 8279
rect 16227 8245 16261 8279
rect 22023 8245 22057 8279
rect 29193 8245 29227 8279
rect 1409 8041 1443 8075
rect 2887 8041 2921 8075
rect 5181 8041 5215 8075
rect 7665 8041 7699 8075
rect 13553 8041 13587 8075
rect 14295 8041 14329 8075
rect 17049 8041 17083 8075
rect 17601 8041 17635 8075
rect 18527 8041 18561 8075
rect 19901 8041 19935 8075
rect 23121 8041 23155 8075
rect 25329 8041 25363 8075
rect 28187 8041 28221 8075
rect 29561 8041 29595 8075
rect 16221 7973 16255 8007
rect 1041 7905 1075 7939
rect 1685 7905 1719 7939
rect 3157 7905 3191 7939
rect 4721 7905 4755 7939
rect 5365 7905 5399 7939
rect 5641 7905 5675 7939
rect 6561 7905 6595 7939
rect 8217 7905 8251 7939
rect 8309 7905 8343 7939
rect 9045 7905 9079 7939
rect 10517 7905 10551 7939
rect 10977 7905 11011 7939
rect 12081 7905 12115 7939
rect 13737 7905 13771 7939
rect 14565 7905 14599 7939
rect 16773 7905 16807 7939
rect 17233 7905 17267 7939
rect 17785 7905 17819 7939
rect 20545 7905 20579 7939
rect 21097 7905 21131 7939
rect 22017 7905 22051 7939
rect 23816 7905 23850 7939
rect 25697 7905 25731 7939
rect 27629 7905 27663 7939
rect 28457 7905 28491 7939
rect 30297 7905 30331 7939
rect 30573 7905 30607 7939
rect 1869 7837 1903 7871
rect 2421 7837 2455 7871
rect 2927 7837 2961 7871
rect 5825 7837 5859 7871
rect 6152 7837 6186 7871
rect 6331 7837 6365 7871
rect 8636 7837 8670 7871
rect 8815 7837 8849 7871
rect 11345 7837 11379 7871
rect 11672 7837 11706 7871
rect 11841 7837 11875 7871
rect 13829 7837 13863 7871
rect 14335 7837 14369 7871
rect 18061 7837 18095 7871
rect 18557 7855 18591 7889
rect 18797 7837 18831 7871
rect 21281 7837 21315 7871
rect 21608 7837 21642 7871
rect 21787 7837 21821 7871
rect 23489 7837 23523 7871
rect 23995 7837 24029 7871
rect 24225 7837 24259 7871
rect 25881 7837 25915 7871
rect 27721 7837 27755 7871
rect 28184 7837 28218 7871
rect 4997 7769 5031 7803
rect 5457 7769 5491 7803
rect 17417 7769 17451 7803
rect 20361 7769 20395 7803
rect 30113 7769 30147 7803
rect 857 7701 891 7735
rect 4261 7701 4295 7735
rect 8033 7701 8067 7735
rect 10333 7701 10367 7735
rect 10701 7701 10735 7735
rect 11161 7701 11195 7735
rect 13185 7701 13219 7735
rect 15669 7701 15703 7735
rect 16313 7701 16347 7735
rect 20913 7701 20947 7735
rect 27445 7701 27479 7735
rect 30389 7701 30423 7735
rect 10241 7497 10275 7531
rect 16221 7497 16255 7531
rect 17785 7497 17819 7531
rect 20729 7497 20763 7531
rect 21281 7497 21315 7531
rect 23581 7497 23615 7531
rect 29009 7497 29043 7531
rect 7389 7429 7423 7463
rect 10977 7429 11011 7463
rect 14105 7429 14139 7463
rect 25973 7429 26007 7463
rect 1455 7361 1489 7395
rect 3576 7361 3610 7395
rect 3755 7361 3789 7395
rect 5549 7361 5583 7395
rect 5876 7361 5910 7395
rect 6055 7361 6089 7395
rect 7941 7361 7975 7395
rect 8728 7361 8762 7395
rect 8907 7359 8941 7393
rect 9137 7361 9171 7395
rect 11759 7361 11793 7395
rect 14887 7361 14921 7395
rect 18337 7361 18371 7395
rect 19032 7361 19066 7395
rect 19201 7361 19235 7395
rect 21884 7361 21918 7395
rect 22020 7343 22054 7377
rect 22293 7361 22327 7395
rect 24133 7361 24167 7395
rect 24596 7361 24630 7395
rect 26804 7361 26838 7395
rect 949 7293 983 7327
rect 1276 7293 1310 7327
rect 1685 7293 1719 7327
rect 3249 7293 3283 7327
rect 3985 7293 4019 7327
rect 6285 7293 6319 7327
rect 7757 7293 7791 7327
rect 8401 7293 8435 7327
rect 10885 7293 10919 7327
rect 11161 7293 11195 7327
rect 11253 7293 11287 7327
rect 11989 7293 12023 7327
rect 13553 7293 13587 7327
rect 14289 7293 14323 7327
rect 14381 7293 14415 7327
rect 15117 7293 15151 7327
rect 16681 7293 16715 7327
rect 17141 7293 17175 7327
rect 17417 7293 17451 7327
rect 17969 7293 18003 7327
rect 18061 7293 18095 7327
rect 18705 7293 18739 7327
rect 19441 7293 19475 7327
rect 21465 7293 21499 7327
rect 21557 7293 21591 7327
rect 24869 7293 24903 7327
rect 26341 7293 26375 7327
rect 27077 7293 27111 7327
rect 28733 7293 28767 7327
rect 29193 7293 29227 7327
rect 29469 7293 29503 7327
rect 3065 7225 3099 7259
rect 13829 7225 13863 7259
rect 5089 7157 5123 7191
rect 10701 7157 10735 7191
rect 11719 7157 11753 7191
rect 13093 7157 13127 7191
rect 14847 7157 14881 7191
rect 16773 7157 16807 7191
rect 17325 7157 17359 7191
rect 17601 7157 17635 7191
rect 24599 7157 24633 7191
rect 26807 7157 26841 7191
rect 28181 7157 28215 7191
rect 28549 7157 28583 7191
rect 29285 7157 29319 7191
rect 5181 6953 5215 6987
rect 8683 6953 8717 6987
rect 11161 6953 11195 6987
rect 11903 6953 11937 6987
rect 17785 6953 17819 6987
rect 18527 6953 18561 6987
rect 1777 6885 1811 6919
rect 4537 6885 4571 6919
rect 27261 6885 27295 6919
rect 27629 6885 27663 6919
rect 1133 6817 1167 6851
rect 1409 6817 1443 6851
rect 1501 6817 1535 6851
rect 2380 6817 2414 6851
rect 4261 6817 4295 6851
rect 5089 6817 5123 6851
rect 5365 6817 5399 6851
rect 5641 6817 5675 6851
rect 5825 6817 5859 6851
rect 6152 6817 6186 6851
rect 8217 6817 8251 6851
rect 10609 6817 10643 6851
rect 11345 6817 11379 6851
rect 12173 6817 12207 6851
rect 13829 6817 13863 6851
rect 14156 6817 14190 6851
rect 16313 6817 16347 6851
rect 16405 6817 16439 6851
rect 16673 6817 16707 6851
rect 16957 6817 16991 6851
rect 17233 6817 17267 6851
rect 17693 6817 17727 6851
rect 17969 6817 18003 6851
rect 18797 6817 18831 6851
rect 20453 6817 20487 6851
rect 20729 6817 20763 6851
rect 21005 6817 21039 6851
rect 24501 6817 24535 6851
rect 24593 6817 24627 6851
rect 26525 6817 26559 6851
rect 27721 6817 27755 6851
rect 28048 6817 28082 6851
rect 28457 6817 28491 6851
rect 2053 6749 2087 6783
rect 2549 6767 2583 6801
rect 2789 6749 2823 6783
rect 6288 6767 6322 6801
rect 6561 6749 6595 6783
rect 8723 6749 8757 6783
rect 8953 6749 8987 6783
rect 11437 6749 11471 6783
rect 11943 6751 11977 6785
rect 14335 6749 14369 6783
rect 14565 6749 14599 6783
rect 18061 6749 18095 6783
rect 18567 6751 18601 6785
rect 22109 6749 22143 6783
rect 22436 6749 22470 6783
rect 22615 6749 22649 6783
rect 22845 6749 22879 6783
rect 24869 6749 24903 6783
rect 26157 6749 26191 6783
rect 28217 6767 28251 6801
rect 15669 6681 15703 6715
rect 16129 6681 16163 6715
rect 17141 6681 17175 6715
rect 17509 6681 17543 6715
rect 26801 6681 26835 6715
rect 29561 6681 29595 6715
rect 949 6613 983 6647
rect 1225 6613 1259 6647
rect 3893 6613 3927 6647
rect 4905 6613 4939 6647
rect 5457 6613 5491 6647
rect 7665 6613 7699 6647
rect 10057 6613 10091 6647
rect 10425 6613 10459 6647
rect 13277 6613 13311 6647
rect 16589 6613 16623 6647
rect 16865 6613 16899 6647
rect 17417 6613 17451 6647
rect 19901 6613 19935 6647
rect 20269 6613 20303 6647
rect 20545 6613 20579 6647
rect 20821 6613 20855 6647
rect 24133 6613 24167 6647
rect 24317 6613 24351 6647
rect 2789 6409 2823 6443
rect 13829 6409 13863 6443
rect 16221 6409 16255 6443
rect 20729 6409 20763 6443
rect 22753 6409 22787 6443
rect 17693 6341 17727 6375
rect 28549 6341 28583 6375
rect 1455 6273 1489 6307
rect 3755 6273 3789 6307
rect 5876 6273 5910 6307
rect 6055 6273 6089 6307
rect 6285 6273 6319 6307
rect 8728 6273 8762 6307
rect 8907 6273 8941 6307
rect 11072 6273 11106 6307
rect 14381 6273 14415 6307
rect 14887 6273 14921 6307
rect 19211 6273 19245 6307
rect 21376 6273 21410 6307
rect 24504 6273 24538 6307
rect 26709 6273 26743 6307
rect 27172 6273 27206 6307
rect 27445 6273 27479 6307
rect 949 6205 983 6239
rect 1276 6205 1310 6239
rect 1685 6205 1719 6239
rect 3249 6205 3283 6239
rect 3985 6205 4019 6239
rect 5549 6205 5583 6239
rect 8401 6205 8435 6239
rect 9137 6205 9171 6239
rect 10609 6205 10643 6239
rect 11345 6205 11379 6239
rect 13001 6205 13035 6239
rect 13277 6205 13311 6239
rect 13737 6205 13771 6239
rect 14013 6205 14047 6239
rect 14289 6205 14323 6239
rect 15117 6205 15151 6239
rect 16865 6205 16899 6239
rect 17141 6205 17175 6239
rect 17393 6201 17427 6235
rect 17509 6205 17543 6239
rect 17969 6205 18003 6239
rect 18061 6205 18095 6239
rect 18521 6205 18555 6239
rect 18705 6205 18739 6239
rect 19441 6205 19475 6239
rect 20913 6205 20947 6239
rect 21649 6205 21683 6239
rect 23305 6205 23339 6239
rect 24041 6205 24075 6239
rect 24777 6205 24811 6239
rect 26617 6205 26651 6239
rect 7849 6137 7883 6171
rect 3715 6069 3749 6103
rect 5089 6069 5123 6103
rect 7389 6069 7423 6103
rect 7941 6069 7975 6103
rect 10241 6069 10275 6103
rect 11075 6069 11109 6103
rect 12449 6069 12483 6103
rect 12817 6069 12851 6103
rect 13093 6069 13127 6103
rect 13553 6069 13587 6103
rect 14105 6069 14139 6103
rect 14847 6069 14881 6103
rect 16681 6069 16715 6103
rect 16957 6069 16991 6103
rect 17233 6069 17267 6103
rect 17785 6069 17819 6103
rect 18245 6069 18279 6103
rect 18337 6069 18371 6103
rect 19171 6069 19205 6103
rect 21379 6069 21413 6103
rect 23121 6069 23155 6103
rect 24507 6069 24541 6103
rect 25881 6069 25915 6103
rect 26433 6069 26467 6103
rect 27175 6069 27209 6103
rect 949 5865 983 5899
rect 1783 5865 1817 5899
rect 3991 5865 4025 5899
rect 6291 5865 6325 5899
rect 8499 5865 8533 5899
rect 10977 5865 11011 5899
rect 21747 5865 21781 5899
rect 23955 5865 23989 5899
rect 25697 5865 25731 5899
rect 26899 5865 26933 5899
rect 1133 5729 1167 5763
rect 6561 5729 6595 5763
rect 10425 5729 10459 5763
rect 10793 5729 10827 5763
rect 11161 5729 11195 5763
rect 11437 5729 11471 5763
rect 11948 5729 11982 5763
rect 14565 5729 14599 5763
rect 15945 5729 15979 5763
rect 16957 5729 16991 5763
rect 18337 5729 18371 5763
rect 19165 5729 19199 5763
rect 20821 5729 20855 5763
rect 21089 5729 21123 5763
rect 21281 5729 21315 5763
rect 22017 5729 22051 5763
rect 23397 5729 23431 5763
rect 25881 5729 25915 5763
rect 26157 5729 26191 5763
rect 26433 5729 26467 5763
rect 28641 5729 28675 5763
rect 29193 5729 29227 5763
rect 29469 5729 29503 5763
rect 1317 5661 1351 5695
rect 1813 5679 1847 5713
rect 2053 5661 2087 5695
rect 3525 5661 3559 5695
rect 4031 5661 4065 5695
rect 4261 5661 4295 5695
rect 5825 5661 5859 5695
rect 6288 5661 6322 5695
rect 8033 5661 8067 5695
rect 8496 5661 8530 5695
rect 8769 5661 8803 5695
rect 11621 5661 11655 5695
rect 12127 5661 12161 5695
rect 12357 5661 12391 5695
rect 13829 5661 13863 5695
rect 14156 5661 14190 5695
rect 14308 5679 14342 5713
rect 16221 5661 16255 5695
rect 16548 5661 16582 5695
rect 16684 5661 16718 5695
rect 18429 5661 18463 5695
rect 18756 5661 18790 5695
rect 18892 5661 18926 5695
rect 20545 5661 20579 5695
rect 21744 5661 21778 5695
rect 23489 5661 23523 5695
rect 23952 5661 23986 5695
rect 24225 5661 24259 5695
rect 26896 5661 26930 5695
rect 27169 5661 27203 5695
rect 10609 5593 10643 5627
rect 20637 5593 20671 5627
rect 3341 5525 3375 5559
rect 5549 5525 5583 5559
rect 7665 5525 7699 5559
rect 9873 5525 9907 5559
rect 10241 5525 10275 5559
rect 11253 5525 11287 5559
rect 13645 5525 13679 5559
rect 20913 5525 20947 5559
rect 25329 5525 25363 5559
rect 25973 5525 26007 5559
rect 28273 5525 28307 5559
rect 28825 5525 28859 5559
rect 29009 5525 29043 5559
rect 29285 5525 29319 5559
rect 2973 5321 3007 5355
rect 5917 5321 5951 5355
rect 13277 5321 13311 5355
rect 23397 5321 23431 5355
rect 29193 5321 29227 5355
rect 3525 5253 3559 5287
rect 23121 5253 23155 5287
rect 26249 5253 26283 5287
rect 949 5185 983 5219
rect 1445 5167 1479 5201
rect 4399 5185 4433 5219
rect 6607 5185 6641 5219
rect 8585 5185 8619 5219
rect 9372 5185 9406 5219
rect 9508 5183 9542 5217
rect 11253 5185 11287 5219
rect 11716 5185 11750 5219
rect 11989 5185 12023 5219
rect 14013 5185 14047 5219
rect 14476 5185 14510 5219
rect 14749 5185 14783 5219
rect 16129 5185 16163 5219
rect 16684 5185 16718 5219
rect 16957 5185 16991 5219
rect 18337 5185 18371 5219
rect 19168 5185 19202 5219
rect 19441 5185 19475 5219
rect 20821 5185 20855 5219
rect 21376 5185 21410 5219
rect 21649 5185 21683 5219
rect 24547 5185 24581 5219
rect 27036 5185 27070 5219
rect 27205 5167 27239 5201
rect 27445 5185 27479 5219
rect 1685 5117 1719 5151
rect 3893 5117 3927 5151
rect 4629 5117 4663 5151
rect 6101 5117 6135 5151
rect 6837 5117 6871 5151
rect 8401 5117 8435 5151
rect 9045 5117 9079 5151
rect 9781 5117 9815 5151
rect 13921 5117 13955 5151
rect 16221 5117 16255 5151
rect 18705 5117 18739 5151
rect 20913 5117 20947 5151
rect 23305 5117 23339 5151
rect 23581 5117 23615 5151
rect 24041 5117 24075 5151
rect 24777 5117 24811 5151
rect 26433 5117 26467 5151
rect 26709 5117 26743 5151
rect 29001 5117 29035 5151
rect 29285 5117 29319 5151
rect 3341 5049 3375 5083
rect 11161 5049 11195 5083
rect 26157 5049 26191 5083
rect 1415 4981 1449 5015
rect 4359 4981 4393 5015
rect 6567 4981 6601 5015
rect 8125 4981 8159 5015
rect 11719 4981 11753 5015
rect 13737 4981 13771 5015
rect 14479 4981 14513 5015
rect 16687 4981 16721 5015
rect 19171 4981 19205 5015
rect 21379 4981 21413 5015
rect 22753 4981 22787 5015
rect 24507 4981 24541 5015
rect 28549 4981 28583 5015
rect 29469 4981 29503 5015
rect 1041 4777 1075 4811
rect 3991 4777 4025 4811
rect 6291 4777 6325 4811
rect 8499 4777 8533 4811
rect 10609 4777 10643 4811
rect 12087 4777 12121 4811
rect 13645 4777 13679 4811
rect 16687 4777 16721 4811
rect 21741 4777 21775 4811
rect 22017 4777 22051 4811
rect 22575 4777 22609 4811
rect 24501 4777 24535 4811
rect 29745 4777 29779 4811
rect 20545 4709 20579 4743
rect 24225 4709 24259 4743
rect 1225 4641 1259 4675
rect 5641 4641 5675 4675
rect 7941 4641 7975 4675
rect 10425 4641 10459 4675
rect 10793 4641 10827 4675
rect 11253 4641 11287 4675
rect 11529 4641 11563 4675
rect 12357 4641 12391 4675
rect 14565 4641 14599 4675
rect 15945 4641 15979 4675
rect 16957 4641 16991 4675
rect 18337 4641 18371 4675
rect 19165 4641 19199 4675
rect 20821 4641 20855 4675
rect 21097 4641 21131 4675
rect 21465 4641 21499 4675
rect 21557 4641 21591 4675
rect 21833 4641 21867 4675
rect 22109 4641 22143 4675
rect 22845 4641 22879 4675
rect 24685 4641 24719 4675
rect 26617 4641 26651 4675
rect 26893 4641 26927 4675
rect 27077 4641 27111 4675
rect 27905 4641 27939 4675
rect 28641 4641 28675 4675
rect 1317 4573 1351 4607
rect 1644 4573 1678 4607
rect 1813 4591 1847 4625
rect 2053 4573 2087 4607
rect 3525 4573 3559 4607
rect 3988 4573 4022 4607
rect 4261 4573 4295 4607
rect 5825 4573 5859 4607
rect 6288 4575 6322 4609
rect 6561 4573 6595 4607
rect 8033 4573 8067 4607
rect 8496 4573 8530 4607
rect 8769 4573 8803 4607
rect 11621 4573 11655 4607
rect 12084 4575 12118 4609
rect 13829 4573 13863 4607
rect 14156 4573 14190 4607
rect 14292 4573 14326 4607
rect 16221 4573 16255 4607
rect 16684 4573 16718 4607
rect 18429 4573 18463 4607
rect 18756 4573 18790 4607
rect 18892 4573 18926 4607
rect 22615 4573 22649 4607
rect 28232 4573 28266 4607
rect 28384 4575 28418 4609
rect 10241 4505 10275 4539
rect 11069 4505 11103 4539
rect 20637 4505 20671 4539
rect 3157 4437 3191 4471
rect 10057 4437 10091 4471
rect 11345 4437 11379 4471
rect 20913 4437 20947 4471
rect 21281 4437 21315 4471
rect 26433 4437 26467 4471
rect 26709 4437 26743 4471
rect 27261 4437 27295 4471
rect 11989 4233 12023 4267
rect 857 4097 891 4131
rect 1353 4079 1387 4113
rect 1593 4097 1627 4131
rect 4264 4095 4298 4129
rect 4537 4097 4571 4131
rect 5917 4097 5951 4131
rect 6336 4097 6370 4131
rect 6472 4095 6506 4129
rect 10612 4097 10646 4131
rect 10885 4097 10919 4131
rect 13277 4097 13311 4131
rect 13921 4097 13955 4131
rect 14703 4097 14737 4131
rect 16901 4079 16935 4113
rect 18521 4097 18555 4131
rect 19993 4097 20027 4131
rect 20361 4097 20395 4131
rect 20824 4097 20858 4131
rect 21097 4097 21131 4131
rect 22845 4097 22879 4131
rect 25007 4097 25041 4131
rect 27036 4097 27070 4131
rect 27205 4095 27239 4129
rect 27445 4097 27479 4131
rect 2973 4029 3007 4063
rect 3801 4029 3835 4063
rect 6009 4029 6043 4063
rect 6745 4029 6779 4063
rect 8401 4029 8435 4063
rect 9597 4029 9631 4063
rect 10149 4029 10183 4063
rect 14197 4029 14231 4063
rect 14524 4029 14558 4063
rect 14933 4029 14967 4063
rect 16405 4029 16439 4063
rect 17141 4029 17175 4063
rect 18705 4029 18739 4063
rect 19809 4029 19843 4063
rect 22661 4029 22695 4063
rect 23397 4029 23431 4063
rect 23673 4029 23707 4063
rect 24501 4029 24535 4063
rect 25237 4029 25271 4063
rect 26709 4029 26743 4063
rect 29009 4029 29043 4063
rect 8677 3961 8711 3995
rect 9045 3961 9079 3995
rect 9873 3961 9907 3995
rect 12449 3961 12483 3995
rect 13001 3961 13035 3995
rect 16313 3961 16347 3995
rect 18981 3961 19015 3995
rect 19349 3961 19383 3995
rect 1323 3893 1357 3927
rect 3433 3893 3467 3927
rect 4267 3893 4301 3927
rect 7849 3893 7883 3927
rect 9137 3893 9171 3927
rect 10615 3893 10649 3927
rect 12541 3893 12575 3927
rect 16871 3893 16905 3927
rect 19625 3893 19659 3927
rect 20827 3893 20861 3927
rect 22385 3893 22419 3927
rect 23213 3893 23247 3927
rect 23489 3893 23523 3927
rect 24041 3893 24075 3927
rect 24967 3893 25001 3927
rect 26525 3893 26559 3927
rect 28549 3893 28583 3927
rect 29193 3893 29227 3927
rect 30205 3893 30239 3927
rect 1041 3689 1075 3723
rect 3991 3689 4025 3723
rect 8401 3689 8435 3723
rect 9143 3689 9177 3723
rect 12087 3689 12121 3723
rect 16595 3689 16629 3723
rect 20361 3689 20395 3723
rect 22759 3689 22793 3723
rect 26065 3689 26099 3723
rect 29837 3689 29871 3723
rect 8125 3621 8159 3655
rect 10793 3621 10827 3655
rect 21557 3621 21591 3655
rect 25053 3621 25087 3655
rect 26985 3621 27019 3655
rect 1225 3553 1259 3587
rect 1644 3553 1678 3587
rect 8585 3553 8619 3587
rect 9413 3553 9447 3587
rect 11069 3553 11103 3587
rect 11621 3553 11655 3587
rect 12357 3553 12391 3587
rect 13737 3553 13771 3587
rect 15945 3553 15979 3587
rect 18245 3553 18279 3587
rect 19073 3553 19107 3587
rect 20637 3553 20671 3587
rect 21281 3553 21315 3587
rect 22017 3553 22051 3587
rect 22293 3553 22327 3587
rect 23029 3553 23063 3587
rect 24777 3553 24811 3587
rect 25513 3553 25547 3587
rect 25789 3553 25823 3587
rect 26617 3553 26651 3587
rect 26709 3553 26743 3587
rect 27353 3553 27387 3587
rect 27997 3553 28031 3587
rect 28733 3553 28767 3587
rect 1317 3485 1351 3519
rect 1823 3485 1857 3519
rect 2053 3485 2087 3519
rect 3525 3485 3559 3519
rect 3988 3485 4022 3519
rect 4261 3485 4295 3519
rect 6009 3485 6043 3519
rect 6336 3485 6370 3519
rect 6472 3485 6506 3519
rect 6745 3485 6779 3519
rect 8677 3485 8711 3519
rect 9183 3485 9217 3519
rect 11345 3485 11379 3519
rect 12084 3485 12118 3519
rect 13829 3485 13863 3519
rect 14156 3485 14190 3519
rect 14292 3487 14326 3521
rect 14565 3485 14599 3519
rect 16129 3485 16163 3519
rect 16592 3487 16626 3521
rect 16865 3485 16899 3519
rect 18337 3485 18371 3519
rect 18664 3485 18698 3519
rect 18800 3487 18834 3521
rect 22756 3487 22790 3521
rect 27629 3485 27663 3519
rect 28324 3485 28358 3519
rect 28460 3485 28494 3519
rect 30389 3485 30423 3519
rect 26433 3417 26467 3451
rect 3341 3349 3375 3383
rect 5549 3349 5583 3383
rect 20729 3349 20763 3383
rect 21833 3349 21867 3383
rect 24317 3349 24351 3383
rect 25329 3349 25363 3383
rect 25605 3349 25639 3383
rect 3249 3145 3283 3179
rect 5733 3145 5767 3179
rect 8125 3145 8159 3179
rect 23397 3145 23431 3179
rect 30205 3145 30239 3179
rect 3617 3077 3651 3111
rect 1455 3009 1489 3043
rect 4389 2991 4423 3025
rect 6607 3007 6641 3041
rect 9372 3009 9406 3043
rect 9551 3007 9585 3041
rect 11161 3009 11195 3043
rect 11716 3009 11750 3043
rect 13369 3009 13403 3043
rect 14476 3009 14510 3043
rect 16129 3009 16163 3043
rect 16684 3009 16718 3043
rect 18337 3009 18371 3043
rect 19168 3009 19202 3043
rect 19441 3009 19475 3043
rect 20821 3009 20855 3043
rect 21376 3009 21410 3043
rect 21649 3009 21683 3043
rect 23857 3009 23891 3043
rect 24320 3009 24354 3043
rect 26528 3009 26562 3043
rect 26801 3009 26835 3043
rect 29285 3009 29319 3043
rect 949 2941 983 2975
rect 1685 2941 1719 2975
rect 3433 2941 3467 2975
rect 3801 2941 3835 2975
rect 3893 2941 3927 2975
rect 4629 2941 4663 2975
rect 6101 2941 6135 2975
rect 6837 2941 6871 2975
rect 9045 2941 9079 2975
rect 9781 2941 9815 2975
rect 11253 2941 11287 2975
rect 11989 2941 12023 2975
rect 13737 2941 13771 2975
rect 14013 2941 14047 2975
rect 14749 2941 14783 2975
rect 16221 2941 16255 2975
rect 16957 2941 16991 2975
rect 18705 2941 18739 2975
rect 20913 2941 20947 2975
rect 21240 2941 21274 2975
rect 24593 2941 24627 2975
rect 26065 2941 26099 2975
rect 29009 2941 29043 2975
rect 3065 2873 3099 2907
rect 8585 2873 8619 2907
rect 23029 2873 23063 2907
rect 23305 2873 23339 2907
rect 1415 2805 1449 2839
rect 4359 2805 4393 2839
rect 6567 2805 6601 2839
rect 8677 2805 8711 2839
rect 11719 2805 11753 2839
rect 13553 2805 13587 2839
rect 14479 2805 14513 2839
rect 16687 2805 16721 2839
rect 19171 2805 19205 2839
rect 24323 2805 24357 2839
rect 25697 2805 25731 2839
rect 26531 2805 26565 2839
rect 28089 2805 28123 2839
rect 949 2601 983 2635
rect 1783 2601 1817 2635
rect 3341 2601 3375 2635
rect 3991 2601 4025 2635
rect 5549 2601 5583 2635
rect 6383 2601 6417 2635
rect 9965 2601 9999 2635
rect 14295 2601 14329 2635
rect 16595 2601 16629 2635
rect 18803 2601 18837 2635
rect 20821 2601 20855 2635
rect 21747 2601 21781 2635
rect 23489 2601 23523 2635
rect 26617 2601 26651 2635
rect 30021 2601 30055 2635
rect 11345 2533 11379 2567
rect 1133 2465 1167 2499
rect 4261 2465 4295 2499
rect 6653 2465 6687 2499
rect 8033 2465 8067 2499
rect 8452 2465 8486 2499
rect 8861 2465 8895 2499
rect 10425 2465 10459 2499
rect 11069 2465 11103 2499
rect 11948 2465 11982 2499
rect 13737 2465 13771 2499
rect 14565 2465 14599 2499
rect 15945 2465 15979 2499
rect 18245 2465 18279 2499
rect 20729 2465 20763 2499
rect 23673 2465 23707 2499
rect 23949 2465 23983 2499
rect 24869 2465 24903 2499
rect 26525 2465 26559 2499
rect 27353 2465 27387 2499
rect 27997 2465 28031 2499
rect 28324 2465 28358 2499
rect 28733 2465 28767 2499
rect 1317 2397 1351 2431
rect 1823 2397 1857 2431
rect 2053 2397 2087 2431
rect 3525 2397 3559 2431
rect 4031 2399 4065 2433
rect 5917 2397 5951 2431
rect 6423 2399 6457 2433
rect 8125 2397 8159 2431
rect 8588 2397 8622 2431
rect 10701 2397 10735 2431
rect 11621 2397 11655 2431
rect 12084 2397 12118 2431
rect 12357 2397 12391 2431
rect 13829 2397 13863 2431
rect 14292 2397 14326 2431
rect 16129 2397 16163 2431
rect 16592 2397 16626 2431
rect 16865 2397 16899 2431
rect 18337 2397 18371 2431
rect 18800 2397 18834 2431
rect 19073 2397 19107 2431
rect 21281 2397 21315 2431
rect 21744 2397 21778 2431
rect 22017 2397 22051 2431
rect 24133 2397 24167 2431
rect 24460 2397 24494 2431
rect 24596 2397 24630 2431
rect 28460 2399 28494 2433
rect 20361 2329 20395 2363
rect 30389 2329 30423 2363
rect 23121 2261 23155 2295
rect 23765 2261 23799 2295
rect 25973 2261 26007 2295
rect 27445 2261 27479 2295
rect 3249 2057 3283 2091
rect 5457 2057 5491 2091
rect 7665 2057 7699 2091
rect 8033 2057 8067 2091
rect 8769 2057 8803 2091
rect 13645 2057 13679 2091
rect 18337 2057 18371 2091
rect 28089 2057 28123 2091
rect 29193 2057 29227 2091
rect 29653 2057 29687 2091
rect 23121 1989 23155 2023
rect 30113 1989 30147 2023
rect 1455 1921 1489 1955
rect 3617 1921 3651 1955
rect 3944 1921 3978 1955
rect 4123 1919 4157 1953
rect 4353 1921 4387 1955
rect 6288 1921 6322 1955
rect 9508 1921 9542 1955
rect 11161 1921 11195 1955
rect 11716 1921 11750 1955
rect 13369 1921 13403 1955
rect 14384 1921 14418 1955
rect 16129 1921 16163 1955
rect 16592 1921 16626 1955
rect 18245 1921 18279 1955
rect 19168 1921 19202 1955
rect 21240 1921 21274 1955
rect 21392 1919 21426 1953
rect 21649 1921 21683 1955
rect 23857 1921 23891 1955
rect 24184 1921 24218 1955
rect 24320 1919 24354 1953
rect 24593 1921 24627 1955
rect 26249 1921 26283 1955
rect 26745 1903 26779 1937
rect 26985 1921 27019 1955
rect 949 1853 983 1887
rect 1685 1853 1719 1887
rect 3433 1853 3467 1887
rect 5825 1853 5859 1887
rect 6561 1853 6595 1887
rect 8217 1853 8251 1887
rect 9045 1853 9079 1887
rect 9781 1853 9815 1887
rect 11253 1853 11287 1887
rect 11580 1853 11614 1887
rect 11989 1853 12023 1887
rect 13829 1853 13863 1887
rect 13921 1853 13955 1887
rect 14248 1853 14282 1887
rect 14657 1853 14691 1887
rect 16865 1853 16899 1887
rect 18521 1853 18555 1887
rect 18705 1853 18739 1887
rect 19032 1853 19066 1887
rect 19441 1853 19475 1887
rect 20913 1853 20947 1887
rect 23305 1853 23339 1887
rect 23581 1853 23615 1887
rect 26576 1853 26610 1887
rect 28641 1853 28675 1887
rect 29001 1853 29035 1887
rect 3065 1785 3099 1819
rect 8493 1785 8527 1819
rect 16037 1785 16071 1819
rect 20821 1785 20855 1819
rect 23029 1785 23063 1819
rect 30389 1785 30423 1819
rect 1415 1717 1449 1751
rect 6291 1717 6325 1751
rect 9511 1717 9545 1751
rect 16595 1717 16629 1751
rect 23397 1717 23431 1751
rect 25697 1717 25731 1751
rect 28825 1717 28859 1751
rect 1041 1513 1075 1547
rect 1783 1513 1817 1547
rect 5549 1513 5583 1547
rect 5917 1513 5951 1547
rect 6935 1513 6969 1547
rect 8493 1513 8527 1547
rect 12087 1513 12121 1547
rect 14295 1513 14329 1547
rect 16595 1513 16629 1547
rect 18803 1513 18837 1547
rect 20821 1513 20855 1547
rect 21747 1513 21781 1547
rect 23489 1513 23523 1547
rect 23765 1513 23799 1547
rect 26893 1513 26927 1547
rect 27261 1513 27295 1547
rect 27537 1513 27571 1547
rect 29469 1513 29503 1547
rect 11069 1445 11103 1479
rect 20453 1445 20487 1479
rect 1225 1377 1259 1411
rect 1317 1377 1351 1411
rect 3433 1377 3467 1411
rect 6101 1377 6135 1411
rect 6377 1377 6411 1411
rect 8677 1377 8711 1411
rect 11437 1377 11471 1411
rect 13737 1377 13771 1411
rect 15945 1377 15979 1411
rect 18245 1377 18279 1411
rect 20729 1377 20763 1411
rect 21005 1377 21039 1411
rect 21281 1377 21315 1411
rect 23673 1377 23707 1411
rect 23949 1377 23983 1411
rect 24133 1377 24167 1411
rect 24460 1377 24494 1411
rect 26617 1377 26651 1411
rect 26709 1377 26743 1411
rect 27077 1377 27111 1411
rect 27353 1377 27387 1411
rect 27629 1377 27663 1411
rect 27956 1377 27990 1411
rect 30021 1377 30055 1411
rect 1813 1327 1847 1361
rect 2053 1309 2087 1343
rect 3525 1309 3559 1343
rect 3852 1309 3886 1343
rect 4031 1309 4065 1343
rect 4261 1309 4295 1343
rect 6469 1309 6503 1343
rect 6965 1327 6999 1361
rect 7205 1309 7239 1343
rect 9004 1309 9038 1343
rect 9140 1309 9174 1343
rect 9413 1309 9447 1343
rect 10793 1309 10827 1343
rect 11621 1309 11655 1343
rect 12084 1327 12118 1361
rect 12357 1309 12391 1343
rect 13829 1309 13863 1343
rect 14292 1309 14326 1343
rect 14565 1309 14599 1343
rect 16129 1309 16163 1343
rect 16592 1309 16626 1343
rect 16865 1309 16899 1343
rect 18337 1309 18371 1343
rect 18800 1309 18834 1343
rect 19073 1309 19107 1343
rect 21744 1309 21778 1343
rect 22017 1309 22051 1343
rect 24629 1327 24663 1361
rect 24869 1309 24903 1343
rect 28092 1309 28126 1343
rect 28365 1309 28399 1343
rect 30389 1309 30423 1343
rect 6193 1241 6227 1275
rect 20545 1241 20579 1275
rect 23305 1241 23339 1275
rect 25973 1241 26007 1275
rect 26433 1173 26467 1207
rect 2789 969 2823 1003
rect 3249 969 3283 1003
rect 3617 969 3651 1003
rect 4721 969 4755 1003
rect 5089 969 5123 1003
rect 5181 969 5215 1003
rect 8401 969 8435 1003
rect 10517 969 10551 1003
rect 11529 969 11563 1003
rect 11989 969 12023 1003
rect 13185 969 13219 1003
rect 13553 969 13587 1003
rect 16129 969 16163 1003
rect 18705 969 18739 1003
rect 20821 969 20855 1003
rect 21281 969 21315 1003
rect 23581 969 23615 1003
rect 26617 969 26651 1003
rect 28549 969 28583 1003
rect 29469 969 29503 1003
rect 29837 969 29871 1003
rect 30205 969 30239 1003
rect 3893 901 3927 935
rect 4169 901 4203 935
rect 5825 901 5859 935
rect 11253 901 11287 935
rect 12909 901 12943 935
rect 18429 901 18463 935
rect 949 833 983 867
rect 1455 833 1489 867
rect 1685 833 1719 867
rect 6428 833 6462 867
rect 6607 831 6641 865
rect 6837 833 6871 867
rect 8217 833 8251 867
rect 9183 831 9217 865
rect 13829 833 13863 867
rect 14335 831 14369 865
rect 16868 833 16902 867
rect 17141 833 17175 867
rect 19308 833 19342 867
rect 19487 833 19521 867
rect 19717 833 19751 867
rect 21557 833 21591 867
rect 22063 833 22097 867
rect 22293 833 22327 867
rect 23857 833 23891 867
rect 24320 833 24354 867
rect 24593 833 24627 867
rect 27172 833 27206 867
rect 27445 833 27479 867
rect 3433 765 3467 799
rect 3801 765 3835 799
rect 4077 765 4111 799
rect 4353 765 4387 799
rect 5365 765 5399 799
rect 5641 765 5675 799
rect 6009 765 6043 799
rect 6101 765 6135 799
rect 8585 765 8619 799
rect 8677 765 8711 799
rect 9004 765 9038 799
rect 9413 765 9447 799
rect 12265 765 12299 799
rect 13093 765 13127 799
rect 13369 765 13403 799
rect 13737 765 13771 799
rect 14565 765 14599 799
rect 16313 765 16347 799
rect 16405 765 16439 799
rect 18889 765 18923 799
rect 18981 765 19015 799
rect 21465 765 21499 799
rect 21884 765 21918 799
rect 26249 765 26283 799
rect 26433 765 26467 799
rect 26709 765 26743 799
rect 29009 765 29043 799
rect 1415 629 1449 663
rect 5457 629 5491 663
rect 12817 629 12851 663
rect 14295 629 14329 663
rect 15669 629 15703 663
rect 16871 629 16905 663
rect 24323 629 24357 663
rect 25697 629 25731 663
rect 26065 629 26099 663
rect 27175 629 27209 663
rect 29193 629 29227 663
<< metal1 >>
rect 7650 22284 7656 22296
rect 5368 22256 7656 22284
rect 5368 22228 5396 22256
rect 7650 22244 7656 22256
rect 7708 22244 7714 22296
rect 7742 22244 7748 22296
rect 7800 22284 7806 22296
rect 14918 22284 14924 22296
rect 7800 22256 14924 22284
rect 7800 22244 7806 22256
rect 14918 22244 14924 22256
rect 14976 22244 14982 22296
rect 22278 22284 22284 22296
rect 18984 22256 22284 22284
rect 18984 22228 19012 22256
rect 22278 22244 22284 22256
rect 22336 22244 22342 22296
rect 22370 22244 22376 22296
rect 22428 22284 22434 22296
rect 23658 22284 23664 22296
rect 22428 22256 23664 22284
rect 22428 22244 22434 22256
rect 23658 22244 23664 22256
rect 23716 22244 23722 22296
rect 23750 22244 23756 22296
rect 23808 22284 23814 22296
rect 28534 22284 28540 22296
rect 23808 22256 28540 22284
rect 23808 22244 23814 22256
rect 28534 22244 28540 22256
rect 28592 22244 28598 22296
rect 5350 22176 5356 22228
rect 5408 22176 5414 22228
rect 5442 22176 5448 22228
rect 5500 22216 5506 22228
rect 14366 22216 14372 22228
rect 5500 22188 14372 22216
rect 5500 22176 5506 22188
rect 14366 22176 14372 22188
rect 14424 22176 14430 22228
rect 18966 22176 18972 22228
rect 19024 22176 19030 22228
rect 21726 22176 21732 22228
rect 21784 22216 21790 22228
rect 30374 22216 30380 22228
rect 21784 22188 30380 22216
rect 21784 22176 21790 22188
rect 30374 22176 30380 22188
rect 30432 22176 30438 22228
rect 1762 22108 1768 22160
rect 1820 22148 1826 22160
rect 7282 22148 7288 22160
rect 1820 22120 7288 22148
rect 1820 22108 1826 22120
rect 7282 22108 7288 22120
rect 7340 22108 7346 22160
rect 7650 22108 7656 22160
rect 7708 22148 7714 22160
rect 9950 22148 9956 22160
rect 7708 22120 9956 22148
rect 7708 22108 7714 22120
rect 9950 22108 9956 22120
rect 10008 22108 10014 22160
rect 13170 22108 13176 22160
rect 13228 22148 13234 22160
rect 22462 22148 22468 22160
rect 13228 22120 22468 22148
rect 13228 22108 13234 22120
rect 22462 22108 22468 22120
rect 22520 22108 22526 22160
rect 22738 22108 22744 22160
rect 22796 22148 22802 22160
rect 25590 22148 25596 22160
rect 22796 22120 25596 22148
rect 22796 22108 22802 22120
rect 25590 22108 25596 22120
rect 25648 22108 25654 22160
rect 3602 22040 3608 22092
rect 3660 22080 3666 22092
rect 18506 22080 18512 22092
rect 3660 22052 12940 22080
rect 3660 22040 3666 22052
rect 12912 22024 12940 22052
rect 13924 22052 18512 22080
rect 1946 21972 1952 22024
rect 2004 22012 2010 22024
rect 7742 22012 7748 22024
rect 2004 21984 7748 22012
rect 2004 21972 2010 21984
rect 7742 21972 7748 21984
rect 7800 21972 7806 22024
rect 12710 22012 12716 22024
rect 7852 21984 12716 22012
rect 3970 21904 3976 21956
rect 4028 21944 4034 21956
rect 7852 21944 7880 21984
rect 12710 21972 12716 21984
rect 12768 21972 12774 22024
rect 12894 21972 12900 22024
rect 12952 21972 12958 22024
rect 13078 21972 13084 22024
rect 13136 22012 13142 22024
rect 13924 22012 13952 22052
rect 18506 22040 18512 22052
rect 18564 22040 18570 22092
rect 18598 22040 18604 22092
rect 18656 22080 18662 22092
rect 23750 22080 23756 22092
rect 18656 22052 23756 22080
rect 18656 22040 18662 22052
rect 23750 22040 23756 22052
rect 23808 22040 23814 22092
rect 25038 22040 25044 22092
rect 25096 22080 25102 22092
rect 25096 22052 31248 22080
rect 25096 22040 25102 22052
rect 31220 22024 31248 22052
rect 13136 21984 13952 22012
rect 13136 21972 13142 21984
rect 13998 21972 14004 22024
rect 14056 22012 14062 22024
rect 16666 22012 16672 22024
rect 14056 21984 16672 22012
rect 14056 21972 14062 21984
rect 16666 21972 16672 21984
rect 16724 21972 16730 22024
rect 21818 22012 21824 22024
rect 17236 21984 21824 22012
rect 17236 21944 17264 21984
rect 21818 21972 21824 21984
rect 21876 21972 21882 22024
rect 27890 22012 27896 22024
rect 22756 21984 27896 22012
rect 4028 21916 7880 21944
rect 8312 21916 17264 21944
rect 4028 21904 4034 21916
rect 1670 21836 1676 21888
rect 1728 21876 1734 21888
rect 4982 21876 4988 21888
rect 1728 21848 4988 21876
rect 1728 21836 1734 21848
rect 4982 21836 4988 21848
rect 5040 21836 5046 21888
rect 6822 21836 6828 21888
rect 6880 21876 6886 21888
rect 8312 21876 8340 21916
rect 17310 21904 17316 21956
rect 17368 21944 17374 21956
rect 20806 21944 20812 21956
rect 17368 21916 20812 21944
rect 17368 21904 17374 21916
rect 20806 21904 20812 21916
rect 20864 21904 20870 21956
rect 21358 21904 21364 21956
rect 21416 21944 21422 21956
rect 22756 21944 22784 21984
rect 27890 21972 27896 21984
rect 27948 21972 27954 22024
rect 31202 21972 31208 22024
rect 31260 21972 31266 22024
rect 21416 21916 22784 21944
rect 21416 21904 21422 21916
rect 22830 21904 22836 21956
rect 22888 21944 22894 21956
rect 25774 21944 25780 21956
rect 22888 21916 25780 21944
rect 22888 21904 22894 21916
rect 25774 21904 25780 21916
rect 25832 21904 25838 21956
rect 6880 21848 8340 21876
rect 6880 21836 6886 21848
rect 8386 21836 8392 21888
rect 8444 21876 8450 21888
rect 10686 21876 10692 21888
rect 8444 21848 10692 21876
rect 8444 21836 8450 21848
rect 10686 21836 10692 21848
rect 10744 21836 10750 21888
rect 10962 21836 10968 21888
rect 11020 21876 11026 21888
rect 20714 21876 20720 21888
rect 11020 21848 20720 21876
rect 11020 21836 11026 21848
rect 20714 21836 20720 21848
rect 20772 21836 20778 21888
rect 21450 21836 21456 21888
rect 21508 21876 21514 21888
rect 22370 21876 22376 21888
rect 21508 21848 22376 21876
rect 21508 21836 21514 21848
rect 22370 21836 22376 21848
rect 22428 21836 22434 21888
rect 22554 21836 22560 21888
rect 22612 21876 22618 21888
rect 25866 21876 25872 21888
rect 22612 21848 25872 21876
rect 22612 21836 22618 21848
rect 25866 21836 25872 21848
rect 25924 21836 25930 21888
rect 552 21786 30912 21808
rect 552 21734 4193 21786
rect 4245 21734 4257 21786
rect 4309 21734 4321 21786
rect 4373 21734 4385 21786
rect 4437 21734 4449 21786
rect 4501 21734 11783 21786
rect 11835 21734 11847 21786
rect 11899 21734 11911 21786
rect 11963 21734 11975 21786
rect 12027 21734 12039 21786
rect 12091 21734 19373 21786
rect 19425 21734 19437 21786
rect 19489 21734 19501 21786
rect 19553 21734 19565 21786
rect 19617 21734 19629 21786
rect 19681 21734 26963 21786
rect 27015 21734 27027 21786
rect 27079 21734 27091 21786
rect 27143 21734 27155 21786
rect 27207 21734 27219 21786
rect 27271 21734 30912 21786
rect 552 21712 30912 21734
rect 3237 21675 3295 21681
rect 3237 21641 3249 21675
rect 3283 21672 3295 21675
rect 8570 21672 8576 21684
rect 3283 21644 8576 21672
rect 3283 21641 3295 21644
rect 3237 21635 3295 21641
rect 8570 21632 8576 21644
rect 8628 21632 8634 21684
rect 10134 21672 10140 21684
rect 8680 21644 10140 21672
rect 7282 21564 7288 21616
rect 7340 21564 7346 21616
rect 8389 21607 8447 21613
rect 8389 21573 8401 21607
rect 8435 21604 8447 21607
rect 8680 21604 8708 21644
rect 10134 21632 10140 21644
rect 10192 21632 10198 21684
rect 10226 21632 10232 21684
rect 10284 21672 10290 21684
rect 10284 21644 12388 21672
rect 10284 21632 10290 21644
rect 8435 21576 8708 21604
rect 12360 21604 12388 21644
rect 13170 21632 13176 21684
rect 13228 21632 13234 21684
rect 13280 21644 14964 21672
rect 13280 21604 13308 21644
rect 12360 21576 13308 21604
rect 8435 21573 8447 21576
rect 8389 21567 8447 21573
rect 1443 21539 1501 21545
rect 1443 21505 1455 21539
rect 1489 21536 1501 21539
rect 3142 21536 3148 21548
rect 1489 21508 3148 21536
rect 1489 21505 1501 21508
rect 1443 21499 1501 21505
rect 3142 21496 3148 21508
rect 3200 21496 3206 21548
rect 3976 21537 4034 21543
rect 3976 21503 3988 21537
rect 4022 21536 4034 21537
rect 4062 21536 4068 21548
rect 4022 21508 4068 21536
rect 4022 21503 4034 21508
rect 3976 21497 4034 21503
rect 4062 21496 4068 21508
rect 4120 21496 4126 21548
rect 4249 21539 4307 21545
rect 4249 21505 4261 21539
rect 4295 21536 4307 21539
rect 5350 21536 5356 21548
rect 4295 21508 5356 21536
rect 4295 21505 4307 21508
rect 4249 21499 4307 21505
rect 5350 21496 5356 21508
rect 5408 21496 5414 21548
rect 5813 21539 5871 21545
rect 5813 21536 5825 21539
rect 5460 21508 5825 21536
rect 937 21471 995 21477
rect 937 21437 949 21471
rect 983 21468 995 21471
rect 1210 21468 1216 21480
rect 983 21440 1216 21468
rect 983 21437 995 21440
rect 937 21431 995 21437
rect 1210 21428 1216 21440
rect 1268 21428 1274 21480
rect 1670 21428 1676 21480
rect 1728 21428 1734 21480
rect 2774 21428 2780 21480
rect 2832 21468 2838 21480
rect 3421 21471 3479 21477
rect 3421 21468 3433 21471
rect 2832 21440 3433 21468
rect 2832 21428 2838 21440
rect 3421 21437 3433 21440
rect 3467 21437 3479 21471
rect 3421 21431 3479 21437
rect 3513 21471 3571 21477
rect 3513 21437 3525 21471
rect 3559 21468 3571 21471
rect 5258 21468 5264 21480
rect 3559 21440 5264 21468
rect 3559 21437 3571 21440
rect 3513 21431 3571 21437
rect 5258 21428 5264 21440
rect 5316 21428 5322 21480
rect 5460 21468 5488 21508
rect 5813 21505 5825 21508
rect 5859 21505 5871 21539
rect 5813 21499 5871 21505
rect 5994 21496 6000 21548
rect 6052 21536 6058 21548
rect 6276 21539 6334 21545
rect 6276 21536 6288 21539
rect 6052 21508 6288 21536
rect 6052 21496 6058 21508
rect 6276 21505 6288 21508
rect 6322 21505 6334 21539
rect 7300 21536 7328 21564
rect 8992 21539 9050 21545
rect 8992 21536 9004 21539
rect 7300 21508 9004 21536
rect 6276 21499 6334 21505
rect 8992 21505 9004 21508
rect 9038 21505 9050 21539
rect 8992 21499 9050 21505
rect 9122 21496 9128 21548
rect 9180 21536 9186 21548
rect 9180 21508 9225 21536
rect 9180 21496 9186 21508
rect 10778 21496 10784 21548
rect 10836 21536 10842 21548
rect 11428 21539 11486 21545
rect 11428 21536 11440 21539
rect 10836 21508 11440 21536
rect 10836 21496 10842 21508
rect 11428 21505 11440 21508
rect 11474 21505 11486 21539
rect 12986 21536 12992 21548
rect 11428 21499 11486 21505
rect 11532 21508 12992 21536
rect 5368 21440 5488 21468
rect 5368 21412 5396 21440
rect 5534 21428 5540 21480
rect 5592 21468 5598 21480
rect 6140 21471 6198 21477
rect 6140 21468 6152 21471
rect 5592 21440 6152 21468
rect 5592 21428 5598 21440
rect 6140 21437 6152 21440
rect 6186 21437 6198 21471
rect 6140 21431 6198 21437
rect 6546 21428 6552 21480
rect 6604 21428 6610 21480
rect 7190 21428 7196 21480
rect 7248 21468 7254 21480
rect 8205 21471 8263 21477
rect 8205 21468 8217 21471
rect 7248 21440 8217 21468
rect 7248 21428 7254 21440
rect 8205 21437 8217 21440
rect 8251 21468 8263 21471
rect 8294 21468 8300 21480
rect 8251 21440 8300 21468
rect 8251 21437 8263 21440
rect 8205 21431 8263 21437
rect 8294 21428 8300 21440
rect 8352 21428 8358 21480
rect 8573 21471 8631 21477
rect 8573 21437 8585 21471
rect 8619 21437 8631 21471
rect 8573 21431 8631 21437
rect 3050 21360 3056 21412
rect 3108 21360 3114 21412
rect 5350 21360 5356 21412
rect 5408 21360 5414 21412
rect 5902 21400 5908 21412
rect 5460 21372 5908 21400
rect 1403 21335 1461 21341
rect 1403 21301 1415 21335
rect 1449 21332 1461 21335
rect 2314 21332 2320 21344
rect 1449 21304 2320 21332
rect 1449 21301 1461 21304
rect 1403 21295 1461 21301
rect 2314 21292 2320 21304
rect 2372 21292 2378 21344
rect 3979 21335 4037 21341
rect 3979 21301 3991 21335
rect 4025 21332 4037 21335
rect 5460 21332 5488 21372
rect 5902 21360 5908 21372
rect 5960 21360 5966 21412
rect 8386 21400 8392 21412
rect 8036 21372 8392 21400
rect 4025 21304 5488 21332
rect 5537 21335 5595 21341
rect 4025 21301 4037 21304
rect 3979 21295 4037 21301
rect 5537 21301 5549 21335
rect 5583 21332 5595 21335
rect 7282 21332 7288 21344
rect 5583 21304 7288 21332
rect 5583 21301 5595 21304
rect 5537 21295 5595 21301
rect 7282 21292 7288 21304
rect 7340 21292 7346 21344
rect 7834 21292 7840 21344
rect 7892 21292 7898 21344
rect 8036 21341 8064 21372
rect 8386 21360 8392 21372
rect 8444 21360 8450 21412
rect 8588 21400 8616 21431
rect 8662 21428 8668 21480
rect 8720 21468 8726 21480
rect 9214 21468 9220 21480
rect 8720 21440 9220 21468
rect 8720 21428 8726 21440
rect 9214 21428 9220 21440
rect 9272 21428 9278 21480
rect 9401 21471 9459 21477
rect 9401 21437 9413 21471
rect 9447 21468 9459 21471
rect 10042 21468 10048 21480
rect 9447 21440 10048 21468
rect 9447 21437 9459 21440
rect 9401 21431 9459 21437
rect 10042 21428 10048 21440
rect 10100 21428 10106 21480
rect 10962 21428 10968 21480
rect 11020 21428 11026 21480
rect 11532 21468 11560 21508
rect 12986 21496 12992 21508
rect 13044 21496 13050 21548
rect 14004 21539 14062 21545
rect 14004 21505 14016 21539
rect 14050 21536 14062 21539
rect 14182 21536 14188 21548
rect 14050 21508 14188 21536
rect 14050 21505 14062 21508
rect 14004 21499 14062 21505
rect 14182 21496 14188 21508
rect 14240 21496 14246 21548
rect 11072 21440 11560 21468
rect 8754 21400 8760 21412
rect 8588 21372 8760 21400
rect 8754 21360 8760 21372
rect 8812 21360 8818 21412
rect 10594 21360 10600 21412
rect 10652 21400 10658 21412
rect 11072 21400 11100 21440
rect 11698 21428 11704 21480
rect 11756 21428 11762 21480
rect 13078 21428 13084 21480
rect 13136 21468 13142 21480
rect 13357 21471 13415 21477
rect 13357 21468 13369 21471
rect 13136 21440 13369 21468
rect 13136 21428 13142 21440
rect 13357 21437 13369 21440
rect 13403 21437 13415 21471
rect 13357 21431 13415 21437
rect 13538 21428 13544 21480
rect 13596 21428 13602 21480
rect 14277 21471 14335 21477
rect 14277 21468 14289 21471
rect 13648 21440 14289 21468
rect 10652 21372 11100 21400
rect 10652 21360 10658 21372
rect 13262 21360 13268 21412
rect 13320 21400 13326 21412
rect 13648 21400 13676 21440
rect 14277 21437 14289 21440
rect 14323 21437 14335 21471
rect 14277 21431 14335 21437
rect 13320 21372 13676 21400
rect 14936 21400 14964 21644
rect 15746 21632 15752 21684
rect 15804 21672 15810 21684
rect 21910 21672 21916 21684
rect 15804 21644 21916 21672
rect 15804 21632 15810 21644
rect 21910 21632 21916 21644
rect 21968 21632 21974 21684
rect 22020 21644 25544 21672
rect 15933 21607 15991 21613
rect 15933 21573 15945 21607
rect 15979 21573 15991 21607
rect 15933 21567 15991 21573
rect 15378 21496 15384 21548
rect 15436 21536 15442 21548
rect 15948 21536 15976 21567
rect 17954 21564 17960 21616
rect 18012 21604 18018 21616
rect 18598 21604 18604 21616
rect 18012 21576 18604 21604
rect 18012 21564 18018 21576
rect 18598 21564 18604 21576
rect 18656 21564 18662 21616
rect 20714 21564 20720 21616
rect 20772 21564 20778 21616
rect 20806 21564 20812 21616
rect 20864 21604 20870 21616
rect 22020 21604 22048 21644
rect 25516 21616 25544 21644
rect 25590 21632 25596 21684
rect 25648 21672 25654 21684
rect 25869 21675 25927 21681
rect 25869 21672 25881 21675
rect 25648 21644 25881 21672
rect 25648 21632 25654 21644
rect 25869 21641 25881 21644
rect 25915 21641 25927 21675
rect 25869 21635 25927 21641
rect 25958 21632 25964 21684
rect 26016 21672 26022 21684
rect 26016 21644 28994 21672
rect 26016 21632 26022 21644
rect 20864 21576 22048 21604
rect 23201 21607 23259 21613
rect 20864 21564 20870 21576
rect 23201 21573 23213 21607
rect 23247 21604 23259 21607
rect 23247 21576 24624 21604
rect 23247 21573 23259 21576
rect 23201 21567 23259 21573
rect 15436 21508 15884 21536
rect 15948 21508 21404 21536
rect 15436 21496 15442 21508
rect 15010 21428 15016 21480
rect 15068 21468 15074 21480
rect 15657 21471 15715 21477
rect 15657 21468 15669 21471
rect 15068 21440 15669 21468
rect 15068 21428 15074 21440
rect 15657 21437 15669 21440
rect 15703 21437 15715 21471
rect 15657 21431 15715 21437
rect 15746 21428 15752 21480
rect 15804 21428 15810 21480
rect 15856 21468 15884 21508
rect 16114 21468 16120 21480
rect 15856 21440 16120 21468
rect 16114 21428 16120 21440
rect 16172 21428 16178 21480
rect 16393 21471 16451 21477
rect 16393 21437 16405 21471
rect 16439 21468 16451 21471
rect 17678 21468 17684 21480
rect 16439 21440 17684 21468
rect 16439 21437 16451 21440
rect 16393 21431 16451 21437
rect 17678 21428 17684 21440
rect 17736 21428 17742 21480
rect 18322 21428 18328 21480
rect 18380 21468 18386 21480
rect 18693 21471 18751 21477
rect 18693 21468 18705 21471
rect 18380 21440 18705 21468
rect 18380 21428 18386 21440
rect 18693 21437 18705 21440
rect 18739 21437 18751 21471
rect 18693 21431 18751 21437
rect 18969 21471 19027 21477
rect 18969 21437 18981 21471
rect 19015 21464 19027 21471
rect 19058 21464 19064 21480
rect 19015 21437 19064 21464
rect 18969 21436 19064 21437
rect 18969 21431 19027 21436
rect 19058 21428 19064 21436
rect 19116 21428 19122 21480
rect 19334 21428 19340 21480
rect 19392 21468 19398 21480
rect 20438 21468 20444 21480
rect 19392 21440 20444 21468
rect 19392 21428 19398 21440
rect 20438 21428 20444 21440
rect 20496 21428 20502 21480
rect 21269 21471 21327 21477
rect 21269 21468 21281 21471
rect 20824 21440 21281 21468
rect 16206 21400 16212 21412
rect 14936 21372 16212 21400
rect 13320 21360 13326 21372
rect 16206 21360 16212 21372
rect 16264 21360 16270 21412
rect 17954 21360 17960 21412
rect 18012 21360 18018 21412
rect 20533 21403 20591 21409
rect 20533 21400 20545 21403
rect 19628 21372 20545 21400
rect 8021 21335 8079 21341
rect 8021 21301 8033 21335
rect 8067 21301 8079 21335
rect 8021 21295 8079 21301
rect 8938 21292 8944 21344
rect 8996 21332 9002 21344
rect 10318 21332 10324 21344
rect 8996 21304 10324 21332
rect 8996 21292 9002 21304
rect 10318 21292 10324 21304
rect 10376 21292 10382 21344
rect 10502 21292 10508 21344
rect 10560 21292 10566 21344
rect 10962 21292 10968 21344
rect 11020 21332 11026 21344
rect 11431 21335 11489 21341
rect 11431 21332 11443 21335
rect 11020 21304 11443 21332
rect 11020 21292 11026 21304
rect 11431 21301 11443 21304
rect 11477 21301 11489 21335
rect 11431 21295 11489 21301
rect 12802 21292 12808 21344
rect 12860 21292 12866 21344
rect 13998 21292 14004 21344
rect 14056 21341 14062 21344
rect 14056 21295 14065 21341
rect 14056 21292 14062 21295
rect 15470 21292 15476 21344
rect 15528 21332 15534 21344
rect 17497 21335 17555 21341
rect 17497 21332 17509 21335
rect 15528 21304 17509 21332
rect 15528 21292 15534 21304
rect 17497 21301 17509 21304
rect 17543 21301 17555 21335
rect 17497 21295 17555 21301
rect 17586 21292 17592 21344
rect 17644 21332 17650 21344
rect 18049 21335 18107 21341
rect 18049 21332 18061 21335
rect 17644 21304 18061 21332
rect 17644 21292 17650 21304
rect 18049 21301 18061 21304
rect 18095 21301 18107 21335
rect 18049 21295 18107 21301
rect 18230 21292 18236 21344
rect 18288 21332 18294 21344
rect 19628 21332 19656 21372
rect 20533 21369 20545 21372
rect 20579 21369 20591 21403
rect 20533 21363 20591 21369
rect 20824 21344 20852 21440
rect 21269 21437 21281 21440
rect 21315 21437 21327 21471
rect 21269 21431 21327 21437
rect 18288 21304 19656 21332
rect 18288 21292 18294 21304
rect 20070 21292 20076 21344
rect 20128 21292 20134 21344
rect 20806 21292 20812 21344
rect 20864 21292 20870 21344
rect 21376 21332 21404 21508
rect 21450 21496 21456 21548
rect 21508 21496 21514 21548
rect 21913 21539 21971 21545
rect 21913 21505 21925 21539
rect 21959 21536 21971 21539
rect 22002 21536 22008 21548
rect 21959 21508 22008 21536
rect 21959 21505 21971 21508
rect 21913 21499 21971 21505
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 22465 21539 22523 21545
rect 22465 21505 22477 21539
rect 22511 21536 22523 21539
rect 23290 21536 23296 21548
rect 22511 21508 23296 21536
rect 22511 21505 22523 21508
rect 22465 21499 22523 21505
rect 23290 21496 23296 21508
rect 23348 21496 23354 21548
rect 24486 21496 24492 21548
rect 24544 21496 24550 21548
rect 24596 21536 24624 21576
rect 25498 21564 25504 21616
rect 25556 21564 25562 21616
rect 28966 21604 28994 21644
rect 29454 21632 29460 21684
rect 29512 21672 29518 21684
rect 29641 21675 29699 21681
rect 29641 21672 29653 21675
rect 29512 21644 29653 21672
rect 29512 21632 29518 21644
rect 29641 21641 29653 21644
rect 29687 21641 29699 21675
rect 29641 21635 29699 21641
rect 30374 21632 30380 21684
rect 30432 21632 30438 21684
rect 28966 21576 31156 21604
rect 31128 21548 31156 21576
rect 29822 21536 29828 21548
rect 24596 21508 28304 21536
rect 22186 21428 22192 21480
rect 22244 21428 22250 21480
rect 22303 21428 22309 21480
rect 22361 21428 22367 21480
rect 23106 21428 23112 21480
rect 23164 21468 23170 21480
rect 23385 21471 23443 21477
rect 23385 21468 23397 21471
rect 23164 21440 23397 21468
rect 23164 21428 23170 21440
rect 23385 21437 23397 21440
rect 23431 21437 23443 21471
rect 23385 21431 23443 21437
rect 23566 21428 23572 21480
rect 23624 21468 23630 21480
rect 23661 21471 23719 21477
rect 23661 21468 23673 21471
rect 23624 21440 23673 21468
rect 23624 21428 23630 21440
rect 23661 21437 23673 21440
rect 23707 21437 23719 21471
rect 23661 21431 23719 21437
rect 23842 21428 23848 21480
rect 23900 21428 23906 21480
rect 23934 21428 23940 21480
rect 23992 21468 23998 21480
rect 24029 21471 24087 21477
rect 24029 21468 24041 21471
rect 23992 21440 24041 21468
rect 23992 21428 23998 21440
rect 24029 21437 24041 21440
rect 24075 21437 24087 21471
rect 24029 21431 24087 21437
rect 24762 21428 24768 21480
rect 24820 21428 24826 21480
rect 24946 21477 24952 21480
rect 24903 21471 24952 21477
rect 24903 21437 24915 21471
rect 24949 21437 24952 21471
rect 24903 21431 24952 21437
rect 24946 21428 24952 21431
rect 25004 21428 25010 21480
rect 25038 21428 25044 21480
rect 25096 21428 25102 21480
rect 25774 21428 25780 21480
rect 25832 21428 25838 21480
rect 26050 21428 26056 21480
rect 26108 21468 26114 21480
rect 26421 21471 26479 21477
rect 26421 21468 26433 21471
rect 26108 21440 26433 21468
rect 26108 21428 26114 21440
rect 26421 21437 26433 21440
rect 26467 21437 26479 21471
rect 26421 21431 26479 21437
rect 26694 21428 26700 21480
rect 26752 21428 26758 21480
rect 28276 21477 28304 21508
rect 29380 21508 29828 21536
rect 28261 21471 28319 21477
rect 28261 21437 28273 21471
rect 28307 21437 28319 21471
rect 28261 21431 28319 21437
rect 29086 21428 29092 21480
rect 29144 21428 29150 21480
rect 29270 21428 29276 21480
rect 29328 21428 29334 21480
rect 29380 21477 29408 21508
rect 29822 21496 29828 21508
rect 29880 21496 29886 21548
rect 31110 21496 31116 21548
rect 31168 21496 31174 21548
rect 29365 21471 29423 21477
rect 29365 21437 29377 21471
rect 29411 21437 29423 21471
rect 30561 21471 30619 21477
rect 30561 21468 30573 21471
rect 29365 21431 29423 21437
rect 29472 21440 30573 21468
rect 28442 21360 28448 21412
rect 28500 21400 28506 21412
rect 29472 21400 29500 21440
rect 30561 21437 30573 21440
rect 30607 21437 30619 21471
rect 30561 21431 30619 21437
rect 28500 21372 29500 21400
rect 29917 21403 29975 21409
rect 28500 21360 28506 21372
rect 29917 21369 29929 21403
rect 29963 21369 29975 21403
rect 29917 21363 29975 21369
rect 22002 21332 22008 21344
rect 21376 21304 22008 21332
rect 22002 21292 22008 21304
rect 22060 21292 22066 21344
rect 23106 21292 23112 21344
rect 23164 21292 23170 21344
rect 23569 21335 23627 21341
rect 23569 21301 23581 21335
rect 23615 21332 23627 21335
rect 23750 21332 23756 21344
rect 23615 21304 23756 21332
rect 23615 21301 23627 21304
rect 23569 21295 23627 21301
rect 23750 21292 23756 21304
rect 23808 21292 23814 21344
rect 23934 21292 23940 21344
rect 23992 21332 23998 21344
rect 25314 21332 25320 21344
rect 23992 21304 25320 21332
rect 23992 21292 23998 21304
rect 25314 21292 25320 21304
rect 25372 21292 25378 21344
rect 25682 21292 25688 21344
rect 25740 21292 25746 21344
rect 27798 21292 27804 21344
rect 27856 21292 27862 21344
rect 28350 21292 28356 21344
rect 28408 21332 28414 21344
rect 29932 21332 29960 21363
rect 28408 21304 29960 21332
rect 30009 21335 30067 21341
rect 28408 21292 28414 21304
rect 30009 21301 30021 21335
rect 30055 21332 30067 21335
rect 30098 21332 30104 21344
rect 30055 21304 30104 21332
rect 30055 21301 30067 21304
rect 30009 21295 30067 21301
rect 30098 21292 30104 21304
rect 30156 21292 30162 21344
rect 552 21242 31072 21264
rect 552 21190 7988 21242
rect 8040 21190 8052 21242
rect 8104 21190 8116 21242
rect 8168 21190 8180 21242
rect 8232 21190 8244 21242
rect 8296 21190 15578 21242
rect 15630 21190 15642 21242
rect 15694 21190 15706 21242
rect 15758 21190 15770 21242
rect 15822 21190 15834 21242
rect 15886 21190 23168 21242
rect 23220 21190 23232 21242
rect 23284 21190 23296 21242
rect 23348 21190 23360 21242
rect 23412 21190 23424 21242
rect 23476 21190 30758 21242
rect 30810 21190 30822 21242
rect 30874 21190 30886 21242
rect 30938 21190 30950 21242
rect 31002 21190 31014 21242
rect 31066 21190 31072 21242
rect 552 21168 31072 21190
rect 1762 21128 1768 21140
rect 1820 21137 1826 21140
rect 1729 21100 1768 21128
rect 1762 21088 1768 21100
rect 1820 21091 1829 21137
rect 5810 21128 5816 21140
rect 3620 21100 5816 21128
rect 1820 21088 1826 21091
rect 3620 20992 3648 21100
rect 5810 21088 5816 21100
rect 5868 21088 5874 21140
rect 5902 21088 5908 21140
rect 5960 21128 5966 21140
rect 6279 21131 6337 21137
rect 6279 21128 6291 21131
rect 5960 21100 6291 21128
rect 5960 21088 5966 21100
rect 6279 21097 6291 21100
rect 6325 21128 6337 21131
rect 8487 21131 8545 21137
rect 8487 21128 8499 21131
rect 6325 21100 8499 21128
rect 6325 21097 6337 21100
rect 6279 21091 6337 21097
rect 5258 21020 5264 21072
rect 5316 21060 5322 21072
rect 5316 21032 5856 21060
rect 5316 21020 5322 21032
rect 5828 21004 5856 21032
rect 7484 21004 7512 21100
rect 8487 21097 8499 21100
rect 8533 21097 8545 21131
rect 8487 21091 8545 21097
rect 8662 21088 8668 21140
rect 8720 21128 8726 21140
rect 8720 21100 9444 21128
rect 8720 21088 8726 21100
rect 9416 21060 9444 21100
rect 9490 21088 9496 21140
rect 9548 21128 9554 21140
rect 9766 21128 9772 21140
rect 9548 21100 9772 21128
rect 9548 21088 9554 21100
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 10965 21131 11023 21137
rect 10965 21097 10977 21131
rect 11011 21128 11023 21131
rect 11514 21128 11520 21140
rect 11011 21100 11520 21128
rect 11011 21097 11023 21100
rect 10965 21091 11023 21097
rect 11514 21088 11520 21100
rect 11572 21088 11578 21140
rect 11606 21088 11612 21140
rect 11664 21128 11670 21140
rect 11707 21131 11765 21137
rect 11707 21128 11719 21131
rect 11664 21100 11719 21128
rect 11664 21088 11670 21100
rect 11707 21097 11719 21100
rect 11753 21097 11765 21131
rect 11707 21091 11765 21097
rect 14918 21088 14924 21140
rect 14976 21128 14982 21140
rect 15289 21131 15347 21137
rect 15289 21128 15301 21131
rect 14976 21100 15301 21128
rect 14976 21088 14982 21100
rect 15289 21097 15301 21100
rect 15335 21097 15347 21131
rect 15289 21091 15347 21097
rect 16666 21088 16672 21140
rect 16724 21128 16730 21140
rect 17957 21131 18015 21137
rect 17957 21128 17969 21131
rect 16724 21100 17969 21128
rect 16724 21088 16730 21100
rect 17957 21097 17969 21100
rect 18003 21097 18015 21131
rect 17957 21091 18015 21097
rect 19058 21088 19064 21140
rect 19116 21128 19122 21140
rect 20162 21128 20168 21140
rect 19116 21100 20168 21128
rect 19116 21088 19122 21100
rect 20162 21088 20168 21100
rect 20220 21088 20226 21140
rect 20806 21088 20812 21140
rect 20864 21088 20870 21140
rect 22186 21088 22192 21140
rect 22244 21128 22250 21140
rect 23109 21131 23167 21137
rect 23109 21128 23121 21131
rect 22244 21100 23121 21128
rect 22244 21088 22250 21100
rect 23109 21097 23121 21100
rect 23155 21097 23167 21131
rect 23109 21091 23167 21097
rect 23382 21088 23388 21140
rect 23440 21128 23446 21140
rect 25038 21128 25044 21140
rect 23440 21100 25044 21128
rect 23440 21088 23446 21100
rect 25038 21088 25044 21100
rect 25096 21088 25102 21140
rect 25314 21088 25320 21140
rect 25372 21088 25378 21140
rect 25498 21088 25504 21140
rect 25556 21128 25562 21140
rect 27801 21131 27859 21137
rect 27801 21128 27813 21131
rect 25556 21100 27813 21128
rect 25556 21088 25562 21100
rect 27801 21097 27813 21100
rect 27847 21097 27859 21131
rect 27801 21091 27859 21097
rect 27890 21088 27896 21140
rect 27948 21128 27954 21140
rect 30377 21131 30435 21137
rect 30377 21128 30389 21131
rect 27948 21100 30389 21128
rect 27948 21088 27954 21100
rect 30377 21097 30389 21100
rect 30423 21097 30435 21131
rect 30377 21091 30435 21097
rect 10226 21060 10232 21072
rect 9416 21032 10232 21060
rect 10226 21020 10232 21032
rect 10284 21020 10290 21072
rect 10410 21020 10416 21072
rect 10468 21020 10474 21072
rect 10781 21063 10839 21069
rect 10781 21029 10793 21063
rect 10827 21060 10839 21063
rect 10870 21060 10876 21072
rect 10827 21032 10876 21060
rect 10827 21029 10839 21032
rect 10781 21023 10839 21029
rect 10870 21020 10876 21032
rect 10928 21020 10934 21072
rect 11149 21019 11207 21025
rect 12894 21020 12900 21072
rect 12952 21060 12958 21072
rect 13357 21063 13415 21069
rect 13357 21060 13369 21063
rect 12952 21032 13369 21060
rect 12952 21020 12958 21032
rect 13357 21029 13369 21032
rect 13403 21029 13415 21063
rect 13357 21023 13415 21029
rect 16592 21032 18276 21060
rect 11149 21016 11161 21019
rect 1320 20964 3648 20992
rect 3840 20995 3898 21001
rect 750 20884 756 20936
rect 808 20924 814 20936
rect 1320 20933 1348 20964
rect 3840 20961 3852 20995
rect 3886 20992 3898 20995
rect 5534 20992 5540 21004
rect 3886 20964 5540 20992
rect 3886 20961 3898 20964
rect 3840 20955 3898 20961
rect 5534 20952 5540 20964
rect 5592 20952 5598 21004
rect 5629 20995 5687 21001
rect 5629 20961 5641 20995
rect 5675 20961 5687 20995
rect 5629 20955 5687 20961
rect 1305 20927 1363 20933
rect 1305 20924 1317 20927
rect 808 20896 1317 20924
rect 808 20884 814 20896
rect 1305 20893 1317 20896
rect 1351 20893 1363 20927
rect 1305 20887 1363 20893
rect 1486 20884 1492 20936
rect 1544 20924 1550 20936
rect 1811 20927 1869 20933
rect 1811 20924 1823 20927
rect 1544 20896 1823 20924
rect 1544 20884 1550 20896
rect 1811 20893 1823 20896
rect 1857 20893 1869 20927
rect 1811 20887 1869 20893
rect 2041 20927 2099 20933
rect 2041 20893 2053 20927
rect 2087 20924 2099 20927
rect 2406 20924 2412 20936
rect 2087 20896 2412 20924
rect 2087 20893 2099 20896
rect 2041 20887 2099 20893
rect 2406 20884 2412 20896
rect 2464 20884 2470 20936
rect 3513 20927 3571 20933
rect 3513 20893 3525 20927
rect 3559 20924 3571 20927
rect 3694 20924 3700 20936
rect 3559 20896 3700 20924
rect 3559 20893 3571 20896
rect 3513 20887 3571 20893
rect 3694 20884 3700 20896
rect 3752 20884 3758 20936
rect 3970 20884 3976 20936
rect 4028 20884 4034 20936
rect 4246 20884 4252 20936
rect 4304 20884 4310 20936
rect 5644 20924 5672 20955
rect 5810 20952 5816 21004
rect 5868 20952 5874 21004
rect 6472 20964 6914 20992
rect 6276 20945 6334 20951
rect 6276 20942 6288 20945
rect 6104 20924 6288 20942
rect 5644 20914 6288 20924
rect 5644 20896 6132 20914
rect 6276 20911 6288 20914
rect 6322 20911 6334 20945
rect 6472 20936 6500 20964
rect 6276 20905 6334 20911
rect 6454 20884 6460 20936
rect 6512 20884 6518 20936
rect 6549 20927 6607 20933
rect 6549 20893 6561 20927
rect 6595 20924 6607 20927
rect 6730 20924 6736 20936
rect 6595 20896 6736 20924
rect 6595 20893 6607 20896
rect 6549 20887 6607 20893
rect 6730 20884 6736 20896
rect 6788 20884 6794 20936
rect 6886 20924 6914 20964
rect 7466 20952 7472 21004
rect 7524 20952 7530 21004
rect 8570 20952 8576 21004
rect 8628 20992 8634 21004
rect 8757 20995 8815 21001
rect 8757 20992 8769 20995
rect 8628 20964 8769 20992
rect 8628 20952 8634 20964
rect 8757 20961 8769 20964
rect 8803 20961 8815 20995
rect 8757 20955 8815 20961
rect 9582 20952 9588 21004
rect 9640 20992 9646 21004
rect 9640 20952 9674 20992
rect 10686 20952 10692 21004
rect 10744 20992 10750 21004
rect 11072 20992 11161 21016
rect 10744 20988 11161 20992
rect 10744 20964 11100 20988
rect 11149 20985 11161 20988
rect 11195 20985 11207 21019
rect 11149 20979 11207 20985
rect 11977 20995 12035 21001
rect 10744 20952 10750 20964
rect 7834 20924 7840 20936
rect 6886 20896 7840 20924
rect 7834 20884 7840 20896
rect 7892 20924 7898 20936
rect 8021 20927 8079 20933
rect 8021 20924 8033 20927
rect 7892 20896 8033 20924
rect 7892 20884 7898 20896
rect 8021 20893 8033 20896
rect 8067 20893 8079 20927
rect 8021 20887 8079 20893
rect 8386 20884 8392 20936
rect 8444 20924 8450 20936
rect 8484 20927 8542 20933
rect 8484 20924 8496 20927
rect 8444 20896 8496 20924
rect 8444 20884 8450 20896
rect 8484 20893 8496 20896
rect 8530 20893 8542 20927
rect 8484 20887 8542 20893
rect 8846 20884 8852 20936
rect 8904 20924 8910 20936
rect 9490 20924 9496 20936
rect 8904 20896 9496 20924
rect 8904 20884 8910 20896
rect 9490 20884 9496 20896
rect 9548 20884 9554 20936
rect 9646 20856 9674 20952
rect 11072 20924 11100 20964
rect 11977 20961 11989 20995
rect 12023 20961 12035 20995
rect 13449 20995 13507 21001
rect 13449 20992 13461 20995
rect 11977 20955 12035 20961
rect 13372 20964 13461 20992
rect 11146 20924 11152 20936
rect 11072 20896 11152 20924
rect 11146 20884 11152 20896
rect 11204 20884 11210 20936
rect 11238 20884 11244 20936
rect 11296 20884 11302 20936
rect 11514 20884 11520 20936
rect 11572 20924 11578 20936
rect 11704 20927 11762 20933
rect 11704 20924 11716 20927
rect 11572 20896 11716 20924
rect 11572 20884 11578 20896
rect 11704 20893 11716 20896
rect 11750 20893 11762 20927
rect 11704 20887 11762 20893
rect 11790 20884 11796 20936
rect 11848 20924 11854 20936
rect 11992 20924 12020 20955
rect 13372 20936 13400 20964
rect 13449 20961 13461 20964
rect 13495 20961 13507 20995
rect 13449 20955 13507 20961
rect 13776 20995 13834 21001
rect 13776 20961 13788 20995
rect 13822 20992 13834 20995
rect 13998 20992 14004 21004
rect 13822 20964 14004 20992
rect 13822 20961 13834 20964
rect 13776 20955 13834 20961
rect 13998 20952 14004 20964
rect 14056 20992 14062 21004
rect 15102 20992 15108 21004
rect 14056 20964 15108 20992
rect 14056 20952 14062 20964
rect 15102 20952 15108 20964
rect 15160 20952 15166 21004
rect 15746 20952 15752 21004
rect 15804 20952 15810 21004
rect 16022 20952 16028 21004
rect 16080 20992 16086 21004
rect 16394 20995 16452 21001
rect 16394 20992 16406 20995
rect 16080 20964 16406 20992
rect 16080 20952 16086 20964
rect 16394 20961 16406 20964
rect 16440 20961 16452 20995
rect 16394 20955 16452 20961
rect 16482 20952 16488 21004
rect 16540 20992 16546 21004
rect 16592 20992 16620 21032
rect 18248 21001 18276 21032
rect 18322 21020 18328 21072
rect 18380 21060 18386 21072
rect 19334 21060 19340 21072
rect 18380 21032 19340 21060
rect 18380 21020 18386 21032
rect 19334 21020 19340 21032
rect 19392 21020 19398 21072
rect 20254 21020 20260 21072
rect 20312 21020 20318 21072
rect 25222 21060 25228 21072
rect 24978 21032 25228 21060
rect 25222 21020 25228 21032
rect 25280 21060 25286 21072
rect 26142 21060 26148 21072
rect 25280 21032 26148 21060
rect 25280 21020 25286 21032
rect 26142 21020 26148 21032
rect 26200 21020 26206 21072
rect 16540 20964 16620 20992
rect 18233 20995 18291 21001
rect 16540 20952 16546 20964
rect 18233 20961 18245 20995
rect 18279 20961 18291 20995
rect 18233 20955 18291 20961
rect 18509 20995 18567 21001
rect 18509 20961 18521 20995
rect 18555 20992 18567 20995
rect 18782 20992 18788 21004
rect 18555 20964 18788 20992
rect 18555 20961 18567 20964
rect 18509 20955 18567 20961
rect 18782 20952 18788 20964
rect 18840 20952 18846 21004
rect 18966 20952 18972 21004
rect 19024 20952 19030 21004
rect 20993 20995 21051 21001
rect 20993 20961 21005 20995
rect 21039 20961 21051 20995
rect 20993 20955 21051 20961
rect 11848 20896 12020 20924
rect 11848 20884 11854 20896
rect 13354 20884 13360 20936
rect 13412 20884 13418 20936
rect 13912 20927 13970 20933
rect 13912 20924 13924 20927
rect 13464 20896 13924 20924
rect 7208 20828 7788 20856
rect 9646 20828 11192 20856
rect 842 20748 848 20800
rect 900 20788 906 20800
rect 1121 20791 1179 20797
rect 1121 20788 1133 20791
rect 900 20760 1133 20788
rect 900 20748 906 20760
rect 1121 20757 1133 20760
rect 1167 20757 1179 20791
rect 1121 20751 1179 20757
rect 2682 20748 2688 20800
rect 2740 20788 2746 20800
rect 3145 20791 3203 20797
rect 3145 20788 3157 20791
rect 2740 20760 3157 20788
rect 2740 20748 2746 20760
rect 3145 20757 3157 20760
rect 3191 20757 3203 20791
rect 3145 20751 3203 20757
rect 4706 20748 4712 20800
rect 4764 20788 4770 20800
rect 7208 20788 7236 20828
rect 4764 20760 7236 20788
rect 4764 20748 4770 20760
rect 7650 20748 7656 20800
rect 7708 20748 7714 20800
rect 7760 20788 7788 20828
rect 9861 20791 9919 20797
rect 9861 20788 9873 20791
rect 7760 20760 9873 20788
rect 9861 20757 9873 20760
rect 9907 20757 9919 20791
rect 11164 20788 11192 20828
rect 12986 20816 12992 20868
rect 13044 20856 13050 20868
rect 13464 20856 13492 20896
rect 13912 20893 13924 20896
rect 13958 20893 13970 20927
rect 13912 20887 13970 20893
rect 14090 20884 14096 20936
rect 14148 20924 14154 20936
rect 14185 20927 14243 20933
rect 14185 20924 14197 20927
rect 14148 20896 14197 20924
rect 14148 20884 14154 20896
rect 14185 20893 14197 20896
rect 14231 20893 14243 20927
rect 14185 20887 14243 20893
rect 14274 20884 14280 20936
rect 14332 20924 14338 20936
rect 15010 20924 15016 20936
rect 14332 20896 15016 20924
rect 14332 20884 14338 20896
rect 15010 20884 15016 20896
rect 15068 20884 15074 20936
rect 16114 20884 16120 20936
rect 16172 20884 16178 20936
rect 19242 20884 19248 20936
rect 19300 20924 19306 20936
rect 21008 20924 21036 20955
rect 22554 20952 22560 21004
rect 22612 20992 22618 21004
rect 23293 20995 23351 21001
rect 22612 20964 22678 20992
rect 22612 20952 22618 20964
rect 23293 20961 23305 20995
rect 23339 20961 23351 20995
rect 23293 20955 23351 20961
rect 25501 20995 25559 21001
rect 25501 20961 25513 20995
rect 25547 20961 25559 20995
rect 25501 20955 25559 20961
rect 19300 20896 21036 20924
rect 19300 20884 19306 20896
rect 21174 20884 21180 20936
rect 21232 20924 21238 20936
rect 21269 20927 21327 20933
rect 21269 20924 21281 20927
rect 21232 20896 21281 20924
rect 21232 20884 21238 20896
rect 21269 20893 21281 20896
rect 21315 20893 21327 20927
rect 21269 20887 21327 20893
rect 21545 20927 21603 20933
rect 21545 20893 21557 20927
rect 21591 20924 21603 20927
rect 23308 20924 23336 20955
rect 23477 20927 23535 20933
rect 23477 20924 23489 20927
rect 21591 20896 23489 20924
rect 21591 20893 21603 20896
rect 21545 20887 21603 20893
rect 23477 20893 23489 20896
rect 23523 20893 23535 20927
rect 23753 20927 23811 20933
rect 23753 20924 23765 20927
rect 23477 20887 23535 20893
rect 23584 20896 23765 20924
rect 13044 20828 13492 20856
rect 13044 20816 13050 20828
rect 17678 20816 17684 20868
rect 17736 20816 17742 20868
rect 17880 20828 19012 20856
rect 11790 20788 11796 20800
rect 11164 20760 11796 20788
rect 9861 20751 9919 20757
rect 11790 20748 11796 20760
rect 11848 20748 11854 20800
rect 15841 20791 15899 20797
rect 15841 20757 15853 20791
rect 15887 20788 15899 20791
rect 17880 20788 17908 20828
rect 15887 20760 17908 20788
rect 15887 20757 15899 20760
rect 15841 20751 15899 20757
rect 18046 20748 18052 20800
rect 18104 20748 18110 20800
rect 18690 20748 18696 20800
rect 18748 20788 18754 20800
rect 18785 20791 18843 20797
rect 18785 20788 18797 20791
rect 18748 20760 18797 20788
rect 18748 20748 18754 20760
rect 18785 20757 18797 20760
rect 18831 20757 18843 20791
rect 18984 20788 19012 20828
rect 22646 20816 22652 20868
rect 22704 20856 22710 20868
rect 23584 20856 23612 20896
rect 23753 20893 23765 20896
rect 23799 20924 23811 20927
rect 25516 20924 25544 20955
rect 25774 20952 25780 21004
rect 25832 20952 25838 21004
rect 25866 20952 25872 21004
rect 25924 20992 25930 21004
rect 26697 20995 26755 21001
rect 26697 20992 26709 20995
rect 25924 20964 26709 20992
rect 25924 20952 25930 20964
rect 26697 20961 26709 20964
rect 26743 20961 26755 20995
rect 26697 20955 26755 20961
rect 27338 20952 27344 21004
rect 27396 20992 27402 21004
rect 28496 20995 28554 21001
rect 28496 20992 28508 20995
rect 27396 20964 28508 20992
rect 27396 20952 27402 20964
rect 28496 20961 28508 20964
rect 28542 20961 28554 20995
rect 28496 20955 28554 20961
rect 30561 20995 30619 21001
rect 30561 20961 30573 20995
rect 30607 20961 30619 20995
rect 30561 20955 30619 20961
rect 23799 20896 25544 20924
rect 23799 20893 23811 20896
rect 23753 20887 23811 20893
rect 26050 20884 26056 20936
rect 26108 20884 26114 20936
rect 26418 20884 26424 20936
rect 26476 20884 26482 20936
rect 26786 20884 26792 20936
rect 26844 20924 26850 20936
rect 28169 20927 28227 20933
rect 28169 20924 28181 20927
rect 26844 20896 28181 20924
rect 26844 20884 26850 20896
rect 28169 20893 28181 20896
rect 28215 20893 28227 20927
rect 28169 20887 28227 20893
rect 28626 20884 28632 20936
rect 28684 20924 28690 20936
rect 28905 20927 28963 20933
rect 28684 20896 28729 20924
rect 28684 20884 28690 20896
rect 28905 20893 28917 20927
rect 28951 20924 28963 20927
rect 30466 20924 30472 20936
rect 28951 20896 30472 20924
rect 28951 20893 28963 20896
rect 28905 20887 28963 20893
rect 30466 20884 30472 20896
rect 30524 20884 30530 20936
rect 22704 20828 23612 20856
rect 22704 20816 22710 20828
rect 25958 20816 25964 20868
rect 26016 20816 26022 20868
rect 23566 20788 23572 20800
rect 18984 20760 23572 20788
rect 18785 20751 18843 20757
rect 23566 20748 23572 20760
rect 23624 20748 23630 20800
rect 24118 20748 24124 20800
rect 24176 20788 24182 20800
rect 26068 20788 26096 20884
rect 29730 20816 29736 20868
rect 29788 20856 29794 20868
rect 30576 20856 30604 20955
rect 29788 20828 30604 20856
rect 29788 20816 29794 20828
rect 24176 20760 26096 20788
rect 24176 20748 24182 20760
rect 26602 20748 26608 20800
rect 26660 20788 26666 20800
rect 30009 20791 30067 20797
rect 30009 20788 30021 20791
rect 26660 20760 30021 20788
rect 26660 20748 26666 20760
rect 30009 20757 30021 20760
rect 30055 20757 30067 20791
rect 30009 20751 30067 20757
rect 552 20698 30912 20720
rect 552 20646 4193 20698
rect 4245 20646 4257 20698
rect 4309 20646 4321 20698
rect 4373 20646 4385 20698
rect 4437 20646 4449 20698
rect 4501 20646 11783 20698
rect 11835 20646 11847 20698
rect 11899 20646 11911 20698
rect 11963 20646 11975 20698
rect 12027 20646 12039 20698
rect 12091 20646 19373 20698
rect 19425 20646 19437 20698
rect 19489 20646 19501 20698
rect 19553 20646 19565 20698
rect 19617 20646 19629 20698
rect 19681 20646 26963 20698
rect 27015 20646 27027 20698
rect 27079 20646 27091 20698
rect 27143 20646 27155 20698
rect 27207 20646 27219 20698
rect 27271 20646 30912 20698
rect 552 20624 30912 20646
rect 2961 20587 3019 20593
rect 2961 20553 2973 20587
rect 3007 20584 3019 20587
rect 5994 20584 6000 20596
rect 3007 20556 6000 20584
rect 3007 20553 3019 20556
rect 2961 20547 3019 20553
rect 5994 20544 6000 20556
rect 6052 20544 6058 20596
rect 7098 20544 7104 20596
rect 7156 20544 7162 20596
rect 7469 20587 7527 20593
rect 7469 20553 7481 20587
rect 7515 20584 7527 20587
rect 9582 20584 9588 20596
rect 7515 20556 9588 20584
rect 7515 20553 7527 20556
rect 7469 20547 7527 20553
rect 9582 20544 9588 20556
rect 9640 20544 9646 20596
rect 10505 20587 10563 20593
rect 10505 20553 10517 20587
rect 10551 20584 10563 20587
rect 10870 20584 10876 20596
rect 10551 20556 10876 20584
rect 10551 20553 10563 20556
rect 10505 20547 10563 20553
rect 10870 20544 10876 20556
rect 10928 20544 10934 20596
rect 13354 20544 13360 20596
rect 13412 20584 13418 20596
rect 21910 20584 21916 20596
rect 13412 20556 14964 20584
rect 13412 20544 13418 20556
rect 3510 20516 3516 20528
rect 2746 20488 3516 20516
rect 1443 20451 1501 20457
rect 1443 20417 1455 20451
rect 1489 20448 1501 20451
rect 2746 20448 2774 20488
rect 3510 20476 3516 20488
rect 3568 20476 3574 20528
rect 3694 20476 3700 20528
rect 3752 20516 3758 20528
rect 5258 20516 5264 20528
rect 3752 20488 5264 20516
rect 3752 20476 3758 20488
rect 5258 20476 5264 20488
rect 5316 20476 5322 20528
rect 7742 20476 7748 20528
rect 7800 20516 7806 20528
rect 8113 20519 8171 20525
rect 8113 20516 8125 20519
rect 7800 20488 8125 20516
rect 7800 20476 7806 20488
rect 8113 20485 8125 20488
rect 8159 20516 8171 20519
rect 8478 20516 8484 20528
rect 8159 20488 8484 20516
rect 8159 20485 8171 20488
rect 8113 20479 8171 20485
rect 8478 20476 8484 20488
rect 8536 20476 8542 20528
rect 10686 20476 10692 20528
rect 10744 20516 10750 20528
rect 11054 20516 11060 20528
rect 10744 20488 11060 20516
rect 10744 20476 10750 20488
rect 11054 20476 11060 20488
rect 11112 20476 11118 20528
rect 5724 20451 5782 20457
rect 5724 20448 5736 20451
rect 1489 20420 2774 20448
rect 3344 20420 5736 20448
rect 1489 20417 1501 20420
rect 1443 20411 1501 20417
rect 937 20383 995 20389
rect 937 20349 949 20383
rect 983 20380 995 20383
rect 1302 20380 1308 20392
rect 983 20352 1308 20380
rect 983 20349 995 20352
rect 937 20343 995 20349
rect 1302 20340 1308 20352
rect 1360 20340 1366 20392
rect 1670 20340 1676 20392
rect 1728 20340 1734 20392
rect 3344 20256 3372 20420
rect 5724 20417 5736 20420
rect 5770 20417 5782 20451
rect 8846 20448 8852 20460
rect 5724 20411 5782 20417
rect 5920 20420 8852 20448
rect 3786 20340 3792 20392
rect 3844 20380 3850 20392
rect 4157 20383 4215 20389
rect 4157 20380 4169 20383
rect 3844 20352 4169 20380
rect 3844 20340 3850 20352
rect 4157 20349 4169 20352
rect 4203 20380 4215 20383
rect 4890 20380 4896 20392
rect 4203 20352 4896 20380
rect 4203 20349 4215 20352
rect 4157 20343 4215 20349
rect 4890 20340 4896 20352
rect 4948 20340 4954 20392
rect 5258 20340 5264 20392
rect 5316 20340 5322 20392
rect 5920 20380 5948 20420
rect 8846 20408 8852 20420
rect 8904 20408 8910 20460
rect 8938 20408 8944 20460
rect 8996 20457 9002 20460
rect 8996 20451 9045 20457
rect 8996 20417 8999 20451
rect 9033 20417 9045 20451
rect 8996 20411 9045 20417
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20448 9275 20451
rect 9398 20448 9404 20460
rect 9263 20420 9404 20448
rect 9263 20417 9275 20420
rect 9217 20411 9275 20417
rect 8996 20408 9002 20411
rect 9398 20408 9404 20420
rect 9456 20408 9462 20460
rect 9582 20408 9588 20460
rect 9640 20448 9646 20460
rect 10226 20448 10232 20460
rect 9640 20420 10232 20448
rect 9640 20408 9646 20420
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 10318 20408 10324 20460
rect 10376 20448 10382 20460
rect 10376 20420 11376 20448
rect 10376 20408 10382 20420
rect 5368 20352 5948 20380
rect 4709 20315 4767 20321
rect 4709 20281 4721 20315
rect 4755 20312 4767 20315
rect 5368 20312 5396 20352
rect 5994 20340 6000 20392
rect 6052 20340 6058 20392
rect 6454 20340 6460 20392
rect 6512 20380 6518 20392
rect 7653 20383 7711 20389
rect 7653 20380 7665 20383
rect 6512 20352 7665 20380
rect 6512 20340 6518 20352
rect 7653 20349 7665 20352
rect 7699 20380 7711 20383
rect 8294 20380 8300 20392
rect 7699 20352 8300 20380
rect 7699 20349 7711 20352
rect 7653 20343 7711 20349
rect 8294 20340 8300 20352
rect 8352 20340 8358 20392
rect 8386 20340 8392 20392
rect 8444 20380 8450 20392
rect 8481 20383 8539 20389
rect 8481 20380 8493 20383
rect 8444 20352 8493 20380
rect 8444 20340 8450 20352
rect 8481 20349 8493 20352
rect 8527 20349 8539 20383
rect 8481 20343 8539 20349
rect 8570 20340 8576 20392
rect 8628 20380 8634 20392
rect 10689 20383 10747 20389
rect 10689 20380 10701 20383
rect 8628 20352 10701 20380
rect 8628 20340 8634 20352
rect 10689 20349 10701 20352
rect 10735 20349 10747 20383
rect 10689 20343 10747 20349
rect 10962 20340 10968 20392
rect 11020 20340 11026 20392
rect 11238 20340 11244 20392
rect 11296 20340 11302 20392
rect 11348 20380 11376 20420
rect 11422 20408 11428 20460
rect 11480 20448 11486 20460
rect 11606 20448 11612 20460
rect 11480 20420 11612 20448
rect 11480 20408 11486 20420
rect 11606 20408 11612 20420
rect 11664 20408 11670 20460
rect 11747 20451 11805 20457
rect 11747 20417 11759 20451
rect 11793 20448 11805 20451
rect 12802 20448 12808 20460
rect 11793 20420 12808 20448
rect 11793 20417 11805 20420
rect 11747 20411 11805 20417
rect 12802 20408 12808 20420
rect 12860 20408 12866 20460
rect 13357 20451 13415 20457
rect 13357 20417 13369 20451
rect 13403 20448 13415 20451
rect 13814 20448 13820 20460
rect 13403 20420 13820 20448
rect 13403 20417 13415 20420
rect 13357 20411 13415 20417
rect 13814 20408 13820 20420
rect 13872 20408 13878 20460
rect 13998 20408 14004 20460
rect 14056 20439 14062 20460
rect 14056 20433 14095 20439
rect 14016 20402 14049 20408
rect 14037 20399 14049 20402
rect 14083 20399 14095 20433
rect 14037 20393 14095 20399
rect 11977 20383 12035 20389
rect 11977 20380 11989 20383
rect 11348 20352 11989 20380
rect 11977 20349 11989 20352
rect 12023 20349 12035 20383
rect 11977 20343 12035 20349
rect 12066 20340 12072 20392
rect 12124 20380 12130 20392
rect 12618 20380 12624 20392
rect 12124 20352 12624 20380
rect 12124 20340 12130 20352
rect 12618 20340 12624 20352
rect 12676 20340 12682 20392
rect 12894 20340 12900 20392
rect 12952 20380 12958 20392
rect 13541 20383 13599 20389
rect 13541 20380 13553 20383
rect 12952 20352 13553 20380
rect 12952 20340 12958 20352
rect 13541 20349 13553 20352
rect 13587 20349 13599 20383
rect 13541 20343 13599 20349
rect 14277 20383 14335 20389
rect 14277 20349 14289 20383
rect 14323 20380 14335 20383
rect 14642 20380 14648 20392
rect 14323 20352 14648 20380
rect 14323 20349 14335 20352
rect 14277 20343 14335 20349
rect 14642 20340 14648 20352
rect 14700 20340 14706 20392
rect 14936 20380 14964 20556
rect 18064 20556 21916 20584
rect 18064 20525 18092 20556
rect 21910 20544 21916 20556
rect 21968 20544 21974 20596
rect 22002 20544 22008 20596
rect 22060 20584 22066 20596
rect 24302 20584 24308 20596
rect 22060 20556 24308 20584
rect 22060 20544 22066 20556
rect 24302 20544 24308 20556
rect 24360 20544 24366 20596
rect 25130 20544 25136 20596
rect 25188 20584 25194 20596
rect 28537 20587 28595 20593
rect 28537 20584 28549 20587
rect 25188 20556 28549 20584
rect 25188 20544 25194 20556
rect 28537 20553 28549 20556
rect 28583 20553 28595 20587
rect 28537 20547 28595 20553
rect 18049 20519 18107 20525
rect 18049 20485 18061 20519
rect 18095 20485 18107 20519
rect 18049 20479 18107 20485
rect 18325 20519 18383 20525
rect 18325 20485 18337 20519
rect 18371 20516 18383 20519
rect 18371 20488 19196 20516
rect 18371 20485 18383 20488
rect 18325 20479 18383 20485
rect 15194 20408 15200 20460
rect 15252 20448 15258 20460
rect 16212 20451 16270 20457
rect 16212 20448 16224 20451
rect 15252 20420 16224 20448
rect 15252 20408 15258 20420
rect 16212 20417 16224 20420
rect 16258 20417 16270 20451
rect 19058 20448 19064 20460
rect 16212 20411 16270 20417
rect 18248 20420 19064 20448
rect 15749 20383 15807 20389
rect 15749 20380 15761 20383
rect 14936 20352 15761 20380
rect 15749 20349 15761 20352
rect 15795 20349 15807 20383
rect 15749 20343 15807 20349
rect 16114 20340 16120 20392
rect 16172 20380 16178 20392
rect 18248 20389 18276 20420
rect 19058 20408 19064 20420
rect 19116 20408 19122 20460
rect 16485 20383 16543 20389
rect 16485 20380 16497 20383
rect 16172 20352 16497 20380
rect 16172 20340 16178 20352
rect 16485 20349 16497 20352
rect 16531 20349 16543 20383
rect 16485 20343 16543 20349
rect 18233 20383 18291 20389
rect 18233 20349 18245 20383
rect 18279 20349 18291 20383
rect 18233 20343 18291 20349
rect 18509 20383 18567 20389
rect 18509 20349 18521 20383
rect 18555 20380 18567 20383
rect 18598 20380 18604 20392
rect 18555 20352 18604 20380
rect 18555 20349 18567 20352
rect 18509 20343 18567 20349
rect 18598 20340 18604 20352
rect 18656 20340 18662 20392
rect 19168 20380 19196 20488
rect 26234 20476 26240 20528
rect 26292 20516 26298 20528
rect 26329 20519 26387 20525
rect 26329 20516 26341 20519
rect 26292 20488 26341 20516
rect 26292 20476 26298 20488
rect 26329 20485 26341 20488
rect 26375 20485 26387 20519
rect 26329 20479 26387 20485
rect 19242 20408 19248 20460
rect 19300 20408 19306 20460
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20448 19579 20451
rect 21174 20448 21180 20460
rect 19567 20420 21180 20448
rect 19567 20417 19579 20420
rect 19521 20411 19579 20417
rect 21174 20408 21180 20420
rect 21232 20448 21238 20460
rect 21266 20451 21324 20457
rect 21266 20448 21278 20451
rect 21232 20420 21278 20448
rect 21232 20408 21238 20420
rect 21266 20417 21278 20420
rect 21312 20417 21324 20451
rect 21266 20411 21324 20417
rect 21821 20451 21879 20457
rect 21821 20417 21833 20451
rect 21867 20448 21879 20451
rect 24121 20451 24179 20457
rect 21867 20420 23612 20448
rect 21867 20417 21879 20420
rect 21821 20411 21879 20417
rect 19168 20352 19288 20380
rect 4755 20284 5396 20312
rect 4755 20281 4767 20284
rect 4709 20275 4767 20281
rect 7558 20272 7564 20324
rect 7616 20312 7622 20324
rect 7837 20315 7895 20321
rect 7837 20312 7849 20315
rect 7616 20284 7849 20312
rect 7616 20272 7622 20284
rect 7837 20281 7849 20284
rect 7883 20281 7895 20315
rect 7837 20275 7895 20281
rect 1403 20247 1461 20253
rect 1403 20213 1415 20247
rect 1449 20244 1461 20247
rect 1578 20244 1584 20256
rect 1449 20216 1584 20244
rect 1449 20213 1461 20216
rect 1403 20207 1461 20213
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 3326 20204 3332 20256
rect 3384 20204 3390 20256
rect 3878 20204 3884 20256
rect 3936 20204 3942 20256
rect 4430 20204 4436 20256
rect 4488 20204 4494 20256
rect 4985 20247 5043 20253
rect 4985 20213 4997 20247
rect 5031 20244 5043 20247
rect 5350 20244 5356 20256
rect 5031 20216 5356 20244
rect 5031 20213 5043 20216
rect 4985 20207 5043 20213
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 5534 20204 5540 20256
rect 5592 20244 5598 20256
rect 5727 20247 5785 20253
rect 5727 20244 5739 20247
rect 5592 20216 5739 20244
rect 5592 20204 5598 20216
rect 5727 20213 5739 20216
rect 5773 20213 5785 20247
rect 5727 20207 5785 20213
rect 5902 20204 5908 20256
rect 5960 20244 5966 20256
rect 8404 20244 8432 20340
rect 5960 20216 8432 20244
rect 8947 20247 9005 20253
rect 5960 20204 5966 20216
rect 8947 20213 8959 20247
rect 8993 20244 9005 20247
rect 10980 20244 11008 20340
rect 11146 20272 11152 20324
rect 11204 20312 11210 20324
rect 11330 20312 11336 20324
rect 11204 20284 11336 20312
rect 11204 20272 11210 20284
rect 11330 20272 11336 20284
rect 11388 20272 11394 20324
rect 15102 20272 15108 20324
rect 15160 20312 15166 20324
rect 15160 20284 15516 20312
rect 15160 20272 15166 20284
rect 8993 20216 11008 20244
rect 8993 20213 9005 20216
rect 8947 20207 9005 20213
rect 11514 20204 11520 20256
rect 11572 20244 11578 20256
rect 11707 20247 11765 20253
rect 11707 20244 11719 20247
rect 11572 20216 11719 20244
rect 11572 20204 11578 20216
rect 11707 20213 11719 20216
rect 11753 20213 11765 20247
rect 11707 20207 11765 20213
rect 14007 20247 14065 20253
rect 14007 20213 14019 20247
rect 14053 20244 14065 20247
rect 14366 20244 14372 20256
rect 14053 20216 14372 20244
rect 14053 20213 14065 20216
rect 14007 20207 14065 20213
rect 14366 20204 14372 20216
rect 14424 20204 14430 20256
rect 15378 20204 15384 20256
rect 15436 20204 15442 20256
rect 15488 20244 15516 20284
rect 18690 20272 18696 20324
rect 18748 20312 18754 20324
rect 18785 20315 18843 20321
rect 18785 20312 18797 20315
rect 18748 20284 18797 20312
rect 18748 20272 18754 20284
rect 18785 20281 18797 20284
rect 18831 20312 18843 20315
rect 19150 20312 19156 20324
rect 18831 20284 19156 20312
rect 18831 20281 18843 20284
rect 18785 20275 18843 20281
rect 19150 20272 19156 20284
rect 19208 20272 19214 20324
rect 19260 20312 19288 20352
rect 21542 20340 21548 20392
rect 21600 20340 21606 20392
rect 23382 20340 23388 20392
rect 23440 20340 23446 20392
rect 23584 20389 23612 20420
rect 24121 20417 24133 20451
rect 24167 20448 24179 20451
rect 27203 20451 27261 20457
rect 24167 20420 25912 20448
rect 24167 20417 24179 20420
rect 24121 20411 24179 20417
rect 23569 20383 23627 20389
rect 23569 20349 23581 20383
rect 23615 20380 23627 20383
rect 23845 20383 23903 20389
rect 23845 20380 23857 20383
rect 23615 20352 23857 20380
rect 23615 20349 23627 20352
rect 23569 20343 23627 20349
rect 23845 20349 23857 20352
rect 23891 20349 23903 20383
rect 23845 20343 23903 20349
rect 25222 20340 25228 20392
rect 25280 20340 25286 20392
rect 25884 20389 25912 20420
rect 27203 20417 27215 20451
rect 27249 20448 27261 20451
rect 27249 20420 30236 20448
rect 27249 20417 27261 20420
rect 27203 20411 27261 20417
rect 30208 20392 30236 20420
rect 25869 20383 25927 20389
rect 25869 20349 25881 20383
rect 25915 20349 25927 20383
rect 25869 20343 25927 20349
rect 26145 20383 26203 20389
rect 26145 20349 26157 20383
rect 26191 20349 26203 20383
rect 26145 20343 26203 20349
rect 19260 20284 19932 20312
rect 16215 20247 16273 20253
rect 16215 20244 16227 20247
rect 15488 20216 16227 20244
rect 16215 20213 16227 20216
rect 16261 20213 16273 20247
rect 16215 20207 16273 20213
rect 16758 20204 16764 20256
rect 16816 20244 16822 20256
rect 17218 20244 17224 20256
rect 16816 20216 17224 20244
rect 16816 20204 16822 20216
rect 17218 20204 17224 20216
rect 17276 20244 17282 20256
rect 17589 20247 17647 20253
rect 17589 20244 17601 20247
rect 17276 20216 17601 20244
rect 17276 20204 17282 20216
rect 17589 20213 17601 20216
rect 17635 20213 17647 20247
rect 17589 20207 17647 20213
rect 17954 20204 17960 20256
rect 18012 20244 18018 20256
rect 18877 20247 18935 20253
rect 18877 20244 18889 20247
rect 18012 20216 18889 20244
rect 18012 20204 18018 20216
rect 18877 20213 18889 20216
rect 18923 20213 18935 20247
rect 19904 20244 19932 20284
rect 20254 20272 20260 20324
rect 20312 20272 20318 20324
rect 21818 20312 21824 20324
rect 20824 20284 21824 20312
rect 20824 20244 20852 20284
rect 21818 20272 21824 20284
rect 21876 20272 21882 20324
rect 22554 20272 22560 20324
rect 22612 20272 22618 20324
rect 19904 20216 20852 20244
rect 21085 20247 21143 20253
rect 18877 20207 18935 20213
rect 21085 20213 21097 20247
rect 21131 20244 21143 20247
rect 22186 20244 22192 20256
rect 21131 20216 22192 20244
rect 21131 20213 21143 20216
rect 21085 20207 21143 20213
rect 22186 20204 22192 20216
rect 22244 20204 22250 20256
rect 23400 20253 23428 20340
rect 26160 20256 26188 20343
rect 26418 20340 26424 20392
rect 26476 20380 26482 20392
rect 26697 20383 26755 20389
rect 26697 20380 26709 20383
rect 26476 20352 26709 20380
rect 26476 20340 26482 20352
rect 26697 20349 26709 20352
rect 26743 20380 26755 20383
rect 26786 20380 26792 20392
rect 26743 20352 26792 20380
rect 26743 20349 26755 20352
rect 26697 20343 26755 20349
rect 26786 20340 26792 20352
rect 26844 20340 26850 20392
rect 27433 20383 27491 20389
rect 27433 20349 27445 20383
rect 27479 20380 27491 20383
rect 29270 20380 29276 20392
rect 27479 20352 29276 20380
rect 27479 20349 27491 20352
rect 27433 20343 27491 20349
rect 29270 20340 29276 20352
rect 29328 20340 29334 20392
rect 29362 20340 29368 20392
rect 29420 20380 29426 20392
rect 29457 20383 29515 20389
rect 29457 20380 29469 20383
rect 29420 20352 29469 20380
rect 29420 20340 29426 20352
rect 29457 20349 29469 20352
rect 29503 20349 29515 20383
rect 29457 20343 29515 20349
rect 29822 20340 29828 20392
rect 29880 20340 29886 20392
rect 30190 20340 30196 20392
rect 30248 20340 30254 20392
rect 29086 20272 29092 20324
rect 29144 20272 29150 20324
rect 29840 20284 30052 20312
rect 23385 20247 23443 20253
rect 23385 20213 23397 20247
rect 23431 20213 23443 20247
rect 23385 20207 23443 20213
rect 24762 20204 24768 20256
rect 24820 20244 24826 20256
rect 25685 20247 25743 20253
rect 25685 20244 25697 20247
rect 24820 20216 25697 20244
rect 24820 20204 24826 20216
rect 25685 20213 25697 20216
rect 25731 20213 25743 20247
rect 25685 20207 25743 20213
rect 26142 20204 26148 20256
rect 26200 20204 26206 20256
rect 26786 20204 26792 20256
rect 26844 20244 26850 20256
rect 27163 20247 27221 20253
rect 27163 20244 27175 20247
rect 26844 20216 27175 20244
rect 26844 20204 26850 20216
rect 27163 20213 27175 20216
rect 27209 20244 27221 20247
rect 27338 20244 27344 20256
rect 27209 20216 27344 20244
rect 27209 20213 27221 20216
rect 27163 20207 27221 20213
rect 27338 20204 27344 20216
rect 27396 20204 27402 20256
rect 27798 20204 27804 20256
rect 27856 20244 27862 20256
rect 29840 20244 29868 20284
rect 27856 20216 29868 20244
rect 27856 20204 27862 20216
rect 29914 20204 29920 20256
rect 29972 20204 29978 20256
rect 30024 20244 30052 20284
rect 30098 20272 30104 20324
rect 30156 20312 30162 20324
rect 30650 20312 30656 20324
rect 30156 20284 30656 20312
rect 30156 20272 30162 20284
rect 30650 20272 30656 20284
rect 30708 20272 30714 20324
rect 30193 20247 30251 20253
rect 30193 20244 30205 20247
rect 30024 20216 30205 20244
rect 30193 20213 30205 20216
rect 30239 20213 30251 20247
rect 30193 20207 30251 20213
rect 552 20154 31072 20176
rect 552 20102 7988 20154
rect 8040 20102 8052 20154
rect 8104 20102 8116 20154
rect 8168 20102 8180 20154
rect 8232 20102 8244 20154
rect 8296 20102 15578 20154
rect 15630 20102 15642 20154
rect 15694 20102 15706 20154
rect 15758 20102 15770 20154
rect 15822 20102 15834 20154
rect 15886 20102 23168 20154
rect 23220 20102 23232 20154
rect 23284 20102 23296 20154
rect 23348 20102 23360 20154
rect 23412 20102 23424 20154
rect 23476 20102 30758 20154
rect 30810 20102 30822 20154
rect 30874 20102 30886 20154
rect 30938 20102 30950 20154
rect 31002 20102 31014 20154
rect 31066 20102 31072 20154
rect 552 20080 31072 20102
rect 1578 20000 1584 20052
rect 1636 20040 1642 20052
rect 1771 20043 1829 20049
rect 1771 20040 1783 20043
rect 1636 20012 1783 20040
rect 1636 20000 1642 20012
rect 1771 20009 1783 20012
rect 1817 20040 1829 20043
rect 1817 20012 2774 20040
rect 1817 20009 1829 20012
rect 1771 20003 1829 20009
rect 1213 19907 1271 19913
rect 1213 19873 1225 19907
rect 1259 19873 1271 19907
rect 1213 19867 1271 19873
rect 1228 19836 1256 19867
rect 1302 19864 1308 19916
rect 1360 19864 1366 19916
rect 2746 19904 2774 20012
rect 3326 20000 3332 20052
rect 3384 20000 3390 20052
rect 10321 20043 10379 20049
rect 10321 20040 10333 20043
rect 4172 20012 10333 20040
rect 3602 19932 3608 19984
rect 3660 19932 3666 19984
rect 4172 19981 4200 20012
rect 10321 20009 10333 20012
rect 10367 20009 10379 20043
rect 18874 20040 18880 20052
rect 10321 20003 10379 20009
rect 11072 20012 15792 20040
rect 4157 19975 4215 19981
rect 4157 19941 4169 19975
rect 4203 19941 4215 19975
rect 4157 19935 4215 19941
rect 4522 19932 4528 19984
rect 4580 19932 4586 19984
rect 4706 19932 4712 19984
rect 4764 19932 4770 19984
rect 5074 19932 5080 19984
rect 5132 19932 5138 19984
rect 5258 19932 5264 19984
rect 5316 19972 5322 19984
rect 5902 19972 5908 19984
rect 5316 19944 5908 19972
rect 5316 19932 5322 19944
rect 5902 19932 5908 19944
rect 5960 19932 5966 19984
rect 8389 19975 8447 19981
rect 8389 19941 8401 19975
rect 8435 19972 8447 19975
rect 8570 19972 8576 19984
rect 8435 19944 8576 19972
rect 8435 19941 8447 19944
rect 8389 19935 8447 19941
rect 8570 19932 8576 19944
rect 8628 19932 8634 19984
rect 3694 19904 3700 19916
rect 2746 19876 3700 19904
rect 3694 19864 3700 19876
rect 3752 19864 3758 19916
rect 3878 19864 3884 19916
rect 3936 19904 3942 19916
rect 5626 19904 5632 19916
rect 3936 19876 5632 19904
rect 3936 19864 3942 19876
rect 5626 19864 5632 19876
rect 5684 19864 5690 19916
rect 5810 19864 5816 19916
rect 5868 19864 5874 19916
rect 6457 19907 6515 19913
rect 6457 19873 6469 19907
rect 6503 19904 6515 19907
rect 6733 19907 6791 19913
rect 6733 19904 6745 19907
rect 6503 19876 6745 19904
rect 6503 19873 6515 19876
rect 6457 19867 6515 19873
rect 6733 19873 6745 19876
rect 6779 19904 6791 19907
rect 6822 19904 6828 19916
rect 6779 19876 6828 19904
rect 6779 19873 6791 19876
rect 6733 19867 6791 19873
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 7006 19864 7012 19916
rect 7064 19864 7070 19916
rect 7834 19864 7840 19916
rect 7892 19904 7898 19916
rect 8481 19907 8539 19913
rect 8481 19904 8493 19907
rect 7892 19876 8493 19904
rect 7892 19864 7898 19876
rect 1801 19857 1859 19863
rect 1578 19836 1584 19848
rect 1228 19808 1584 19836
rect 1578 19796 1584 19808
rect 1636 19796 1642 19848
rect 1801 19823 1813 19857
rect 1847 19836 1859 19857
rect 1946 19836 1952 19848
rect 1847 19823 1952 19836
rect 1801 19817 1952 19823
rect 1826 19808 1952 19817
rect 1946 19796 1952 19808
rect 2004 19796 2010 19848
rect 2038 19796 2044 19848
rect 2096 19796 2102 19848
rect 3326 19796 3332 19848
rect 3384 19836 3390 19848
rect 3896 19836 3924 19864
rect 3384 19808 3924 19836
rect 8312 19836 8340 19876
rect 8481 19873 8493 19876
rect 8527 19873 8539 19907
rect 8481 19867 8539 19873
rect 8808 19907 8866 19913
rect 8808 19873 8820 19907
rect 8854 19904 8866 19907
rect 9217 19907 9275 19913
rect 8854 19876 9174 19904
rect 8854 19873 8866 19876
rect 8808 19867 8866 19873
rect 8386 19836 8392 19848
rect 8312 19808 8392 19836
rect 3384 19796 3390 19808
rect 8386 19796 8392 19808
rect 8444 19796 8450 19848
rect 8938 19796 8944 19848
rect 8996 19796 9002 19848
rect 9146 19836 9174 19876
rect 9217 19873 9229 19907
rect 9263 19904 9275 19907
rect 11072 19904 11100 20012
rect 15764 19984 15792 20012
rect 15948 20012 18880 20040
rect 11606 19932 11612 19984
rect 11664 19972 11670 19984
rect 11701 19975 11759 19981
rect 11701 19972 11713 19975
rect 11664 19944 11713 19972
rect 11664 19932 11670 19944
rect 11701 19941 11713 19944
rect 11747 19941 11759 19975
rect 11701 19935 11759 19941
rect 14108 19944 14412 19972
rect 9263 19876 11100 19904
rect 11149 19907 11207 19913
rect 9263 19873 9275 19876
rect 9217 19867 9275 19873
rect 11149 19873 11161 19907
rect 11195 19873 11207 19907
rect 11149 19867 11207 19873
rect 11333 19907 11391 19913
rect 11333 19873 11345 19907
rect 11379 19904 11391 19907
rect 11882 19904 11888 19916
rect 11379 19876 11888 19904
rect 11379 19873 11391 19876
rect 11333 19867 11391 19873
rect 9306 19836 9312 19848
rect 9146 19808 9312 19836
rect 9306 19796 9312 19808
rect 9364 19796 9370 19848
rect 9398 19796 9404 19848
rect 9456 19836 9462 19848
rect 9582 19836 9588 19848
rect 9456 19808 9588 19836
rect 9456 19796 9462 19808
rect 9582 19796 9588 19808
rect 9640 19796 9646 19848
rect 5258 19768 5264 19780
rect 2746 19740 5264 19768
rect 1029 19703 1087 19709
rect 1029 19669 1041 19703
rect 1075 19700 1087 19703
rect 2746 19700 2774 19740
rect 5258 19728 5264 19740
rect 5316 19728 5322 19780
rect 5718 19728 5724 19780
rect 5776 19768 5782 19780
rect 11164 19768 11192 19867
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 12434 19864 12440 19916
rect 12492 19904 12498 19916
rect 12529 19907 12587 19913
rect 12529 19904 12541 19907
rect 12492 19876 12541 19904
rect 12492 19864 12498 19876
rect 12529 19873 12541 19876
rect 12575 19873 12587 19907
rect 12529 19867 12587 19873
rect 11606 19796 11612 19848
rect 11664 19836 11670 19848
rect 12158 19845 12164 19848
rect 11793 19839 11851 19845
rect 11793 19836 11805 19839
rect 11664 19808 11805 19836
rect 11664 19796 11670 19808
rect 11793 19805 11805 19808
rect 11839 19805 11851 19839
rect 11793 19799 11851 19805
rect 12120 19839 12164 19845
rect 12120 19805 12132 19839
rect 12120 19799 12164 19805
rect 12158 19796 12164 19799
rect 12216 19796 12222 19848
rect 12299 19839 12357 19845
rect 12299 19805 12311 19839
rect 12345 19836 12357 19839
rect 14108 19836 14136 19944
rect 14182 19864 14188 19916
rect 14240 19864 14246 19916
rect 12345 19808 14136 19836
rect 14277 19839 14335 19845
rect 12345 19805 12357 19808
rect 12299 19799 12357 19805
rect 14277 19805 14289 19839
rect 14323 19805 14335 19839
rect 14384 19836 14412 19944
rect 15746 19932 15752 19984
rect 15804 19932 15810 19984
rect 15948 19981 15976 20012
rect 18874 20000 18880 20012
rect 18932 20000 18938 20052
rect 19058 20000 19064 20052
rect 19116 20040 19122 20052
rect 20714 20040 20720 20052
rect 19116 20012 20720 20040
rect 19116 20000 19122 20012
rect 20714 20000 20720 20012
rect 20772 20000 20778 20052
rect 20901 20043 20959 20049
rect 20901 20009 20913 20043
rect 20947 20009 20959 20043
rect 22554 20040 22560 20052
rect 20901 20003 20959 20009
rect 21284 20012 22560 20040
rect 15933 19975 15991 19981
rect 15933 19941 15945 19975
rect 15979 19941 15991 19975
rect 16298 19972 16304 19984
rect 15933 19935 15991 19941
rect 16132 19944 16304 19972
rect 14553 19907 14611 19913
rect 14553 19873 14565 19907
rect 14599 19904 14611 19907
rect 15470 19904 15476 19916
rect 14599 19876 15476 19904
rect 14599 19873 14611 19876
rect 14553 19867 14611 19873
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 15286 19836 15292 19848
rect 14384 19808 15292 19836
rect 14277 19799 14335 19805
rect 11330 19768 11336 19780
rect 5776 19740 6776 19768
rect 11164 19740 11336 19768
rect 5776 19728 5782 19740
rect 1075 19672 2774 19700
rect 3881 19703 3939 19709
rect 1075 19669 1087 19672
rect 1029 19663 1087 19669
rect 3881 19669 3893 19703
rect 3927 19700 3939 19703
rect 4062 19700 4068 19712
rect 3927 19672 4068 19700
rect 3927 19669 3939 19672
rect 3881 19663 3939 19669
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 5534 19660 5540 19712
rect 5592 19660 5598 19712
rect 5997 19703 6055 19709
rect 5997 19669 6009 19703
rect 6043 19700 6055 19703
rect 6454 19700 6460 19712
rect 6043 19672 6460 19700
rect 6043 19669 6055 19672
rect 5997 19663 6055 19669
rect 6454 19660 6460 19672
rect 6512 19660 6518 19712
rect 6748 19700 6776 19740
rect 11330 19728 11336 19740
rect 11388 19728 11394 19780
rect 11422 19728 11428 19780
rect 11480 19768 11486 19780
rect 11698 19768 11704 19780
rect 11480 19740 11704 19768
rect 11480 19728 11486 19740
rect 11698 19728 11704 19740
rect 11756 19728 11762 19780
rect 13906 19728 13912 19780
rect 13964 19768 13970 19780
rect 14090 19768 14096 19780
rect 13964 19740 14096 19768
rect 13964 19728 13970 19740
rect 14090 19728 14096 19740
rect 14148 19768 14154 19780
rect 14292 19768 14320 19799
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 16132 19845 16160 19944
rect 16298 19932 16304 19944
rect 16356 19932 16362 19984
rect 17678 19972 17684 19984
rect 17618 19944 17684 19972
rect 17678 19932 17684 19944
rect 17736 19932 17742 19984
rect 19794 19932 19800 19984
rect 19852 19932 19858 19984
rect 20622 19932 20628 19984
rect 20680 19972 20686 19984
rect 20916 19972 20944 20003
rect 20680 19944 20944 19972
rect 20680 19932 20686 19944
rect 17696 19904 17724 19932
rect 19812 19904 19840 19932
rect 17696 19876 19840 19904
rect 20070 19864 20076 19916
rect 20128 19864 20134 19916
rect 20162 19864 20168 19916
rect 20220 19864 20226 19916
rect 20254 19864 20260 19916
rect 20312 19904 20318 19916
rect 20312 19876 21036 19904
rect 20312 19864 20318 19876
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19805 16175 19839
rect 16393 19839 16451 19845
rect 16393 19836 16405 19839
rect 16117 19799 16175 19805
rect 16230 19808 16405 19836
rect 14148 19740 14320 19768
rect 14148 19728 14154 19740
rect 9030 19700 9036 19712
rect 6748 19672 9036 19700
rect 9030 19660 9036 19672
rect 9088 19660 9094 19712
rect 9122 19660 9128 19712
rect 9180 19700 9186 19712
rect 9398 19700 9404 19712
rect 9180 19672 9404 19700
rect 9180 19660 9186 19672
rect 9398 19660 9404 19672
rect 9456 19660 9462 19712
rect 10965 19703 11023 19709
rect 10965 19669 10977 19703
rect 11011 19700 11023 19703
rect 12250 19700 12256 19712
rect 11011 19672 12256 19700
rect 11011 19669 11023 19672
rect 10965 19663 11023 19669
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 12434 19660 12440 19712
rect 12492 19700 12498 19712
rect 13262 19700 13268 19712
rect 12492 19672 13268 19700
rect 12492 19660 12498 19672
rect 13262 19660 13268 19672
rect 13320 19660 13326 19712
rect 13630 19660 13636 19712
rect 13688 19660 13694 19712
rect 14001 19703 14059 19709
rect 14001 19669 14013 19703
rect 14047 19700 14059 19703
rect 14458 19700 14464 19712
rect 14047 19672 14464 19700
rect 14047 19669 14059 19672
rect 14001 19663 14059 19669
rect 14458 19660 14464 19672
rect 14516 19660 14522 19712
rect 16022 19660 16028 19712
rect 16080 19700 16086 19712
rect 16230 19700 16258 19808
rect 16393 19805 16405 19808
rect 16439 19805 16451 19839
rect 16393 19799 16451 19805
rect 16482 19796 16488 19848
rect 16540 19836 16546 19848
rect 17954 19836 17960 19848
rect 16540 19808 17960 19836
rect 16540 19796 16546 19808
rect 17954 19796 17960 19808
rect 18012 19796 18018 19848
rect 18233 19839 18291 19845
rect 18233 19805 18245 19839
rect 18279 19836 18291 19839
rect 20088 19836 20116 19864
rect 20533 19839 20591 19845
rect 20533 19836 20545 19839
rect 18279 19808 20116 19836
rect 20180 19808 20545 19836
rect 18279 19805 18291 19808
rect 18233 19799 18291 19805
rect 20180 19712 20208 19808
rect 20533 19805 20545 19808
rect 20579 19805 20591 19839
rect 21008 19836 21036 19876
rect 21082 19864 21088 19916
rect 21140 19864 21146 19916
rect 21284 19913 21312 20012
rect 22554 20000 22560 20012
rect 22612 20040 22618 20052
rect 22612 20012 23704 20040
rect 22612 20000 22618 20012
rect 21542 19932 21548 19984
rect 21600 19932 21606 19984
rect 22646 19972 22652 19984
rect 22112 19944 22652 19972
rect 21269 19907 21327 19913
rect 21269 19873 21281 19907
rect 21315 19873 21327 19907
rect 21560 19904 21588 19932
rect 21560 19876 21864 19904
rect 21269 19867 21327 19873
rect 21284 19836 21312 19867
rect 21008 19808 21312 19836
rect 21637 19839 21695 19845
rect 20533 19799 20591 19805
rect 21637 19805 21649 19839
rect 21683 19805 21695 19839
rect 21637 19799 21695 19805
rect 16080 19672 16258 19700
rect 16080 19660 16086 19672
rect 16758 19660 16764 19712
rect 16816 19700 16822 19712
rect 17865 19703 17923 19709
rect 17865 19700 17877 19703
rect 16816 19672 17877 19700
rect 16816 19660 16822 19672
rect 17865 19669 17877 19672
rect 17911 19669 17923 19703
rect 17865 19663 17923 19669
rect 18966 19660 18972 19712
rect 19024 19700 19030 19712
rect 19337 19703 19395 19709
rect 19337 19700 19349 19703
rect 19024 19672 19349 19700
rect 19024 19660 19030 19672
rect 19337 19669 19349 19672
rect 19383 19669 19395 19703
rect 19337 19663 19395 19669
rect 20162 19660 20168 19712
rect 20220 19660 20226 19712
rect 20622 19660 20628 19712
rect 20680 19660 20686 19712
rect 21652 19700 21680 19799
rect 21836 19768 21864 19876
rect 22002 19864 22008 19916
rect 22060 19864 22066 19916
rect 22112 19913 22140 19944
rect 22646 19932 22652 19944
rect 22704 19932 22710 19984
rect 23676 19972 23704 20012
rect 23842 20000 23848 20052
rect 23900 20040 23906 20052
rect 23937 20043 23995 20049
rect 23937 20040 23949 20043
rect 23900 20012 23949 20040
rect 23900 20000 23906 20012
rect 23937 20009 23949 20012
rect 23983 20009 23995 20043
rect 25222 20040 25228 20052
rect 23937 20003 23995 20009
rect 24044 20012 25228 20040
rect 24044 19972 24072 20012
rect 25222 20000 25228 20012
rect 25280 20000 25286 20052
rect 26234 20000 26240 20052
rect 26292 20040 26298 20052
rect 28169 20043 28227 20049
rect 28169 20040 28181 20043
rect 26292 20012 28181 20040
rect 26292 20000 26298 20012
rect 28169 20009 28181 20012
rect 28215 20009 28227 20043
rect 28169 20003 28227 20009
rect 29270 20000 29276 20052
rect 29328 20040 29334 20052
rect 30558 20040 30564 20052
rect 29328 20012 30564 20040
rect 29328 20000 29334 20012
rect 30558 20000 30564 20012
rect 30616 20000 30622 20052
rect 23598 19944 24072 19972
rect 22097 19907 22155 19913
rect 22097 19873 22109 19907
rect 22143 19873 22155 19907
rect 22097 19867 22155 19873
rect 24121 19907 24179 19913
rect 24121 19873 24133 19907
rect 24167 19873 24179 19907
rect 24581 19907 24639 19913
rect 24581 19904 24593 19907
rect 24121 19867 24179 19873
rect 24228 19876 24593 19904
rect 22373 19839 22431 19845
rect 22373 19836 22385 19839
rect 22204 19808 22385 19836
rect 22204 19768 22232 19808
rect 22373 19805 22385 19808
rect 22419 19836 22431 19839
rect 24136 19836 24164 19867
rect 22419 19808 24164 19836
rect 22419 19805 22431 19808
rect 22373 19799 22431 19805
rect 21836 19740 22232 19768
rect 23382 19728 23388 19780
rect 23440 19768 23446 19780
rect 24228 19768 24256 19876
rect 24581 19873 24593 19876
rect 24627 19873 24639 19907
rect 24581 19867 24639 19873
rect 26237 19907 26295 19913
rect 26237 19873 26249 19907
rect 26283 19873 26295 19907
rect 26237 19867 26295 19873
rect 24302 19796 24308 19848
rect 24360 19796 24366 19848
rect 23440 19740 24256 19768
rect 26252 19768 26280 19867
rect 26326 19864 26332 19916
rect 26384 19904 26390 19916
rect 26697 19907 26755 19913
rect 26697 19904 26709 19907
rect 26384 19876 26709 19904
rect 26384 19864 26390 19876
rect 26697 19873 26709 19876
rect 26743 19873 26755 19907
rect 26697 19867 26755 19873
rect 27614 19864 27620 19916
rect 27672 19904 27678 19916
rect 27982 19904 27988 19916
rect 27672 19876 27988 19904
rect 27672 19864 27678 19876
rect 27982 19864 27988 19876
rect 28040 19904 28046 19916
rect 28353 19907 28411 19913
rect 28353 19904 28365 19907
rect 28040 19876 28365 19904
rect 28040 19864 28046 19876
rect 28353 19873 28365 19876
rect 28399 19873 28411 19907
rect 28353 19867 28411 19873
rect 28534 19864 28540 19916
rect 28592 19904 28598 19916
rect 28592 19876 30328 19904
rect 28592 19864 28598 19876
rect 26421 19839 26479 19845
rect 26421 19805 26433 19839
rect 26467 19836 26479 19839
rect 27798 19836 27804 19848
rect 26467 19808 27804 19836
rect 26467 19805 26479 19808
rect 26421 19799 26479 19805
rect 26326 19768 26332 19780
rect 26252 19740 26332 19768
rect 23440 19728 23446 19740
rect 26326 19728 26332 19740
rect 26384 19728 26390 19780
rect 22094 19700 22100 19712
rect 21652 19672 22100 19700
rect 22094 19660 22100 19672
rect 22152 19660 22158 19712
rect 22186 19660 22192 19712
rect 22244 19700 22250 19712
rect 25685 19703 25743 19709
rect 25685 19700 25697 19703
rect 22244 19672 25697 19700
rect 22244 19660 22250 19672
rect 25685 19669 25697 19672
rect 25731 19669 25743 19703
rect 25685 19663 25743 19669
rect 26050 19660 26056 19712
rect 26108 19660 26114 19712
rect 26142 19660 26148 19712
rect 26200 19700 26206 19712
rect 26436 19700 26464 19799
rect 27798 19796 27804 19808
rect 27856 19796 27862 19848
rect 28258 19796 28264 19848
rect 28316 19836 28322 19848
rect 28810 19845 28816 19848
rect 28445 19839 28503 19845
rect 28445 19836 28457 19839
rect 28316 19808 28457 19836
rect 28316 19796 28322 19808
rect 28445 19805 28457 19808
rect 28491 19805 28503 19839
rect 28445 19799 28503 19805
rect 28772 19839 28816 19845
rect 28772 19805 28784 19839
rect 28772 19799 28816 19805
rect 28810 19796 28816 19799
rect 28868 19796 28874 19848
rect 28908 19841 28966 19847
rect 28908 19807 28920 19841
rect 28954 19836 28966 19841
rect 28994 19836 29000 19848
rect 28954 19808 29000 19836
rect 28954 19807 28966 19808
rect 28908 19801 28966 19807
rect 28994 19796 29000 19808
rect 29052 19796 29058 19848
rect 29181 19839 29239 19845
rect 29181 19805 29193 19839
rect 29227 19836 29239 19839
rect 29546 19836 29552 19848
rect 29227 19808 29552 19836
rect 29227 19805 29239 19808
rect 29181 19799 29239 19805
rect 29546 19796 29552 19808
rect 29604 19796 29610 19848
rect 30300 19712 30328 19876
rect 26200 19672 26464 19700
rect 27985 19703 28043 19709
rect 26200 19660 26206 19672
rect 27985 19669 27997 19703
rect 28031 19700 28043 19703
rect 30006 19700 30012 19712
rect 28031 19672 30012 19700
rect 28031 19669 28043 19672
rect 27985 19663 28043 19669
rect 30006 19660 30012 19672
rect 30064 19660 30070 19712
rect 30282 19660 30288 19712
rect 30340 19660 30346 19712
rect 30469 19703 30527 19709
rect 30469 19669 30481 19703
rect 30515 19700 30527 19703
rect 30515 19672 30972 19700
rect 30515 19669 30527 19672
rect 30469 19663 30527 19669
rect 552 19610 30912 19632
rect 552 19558 4193 19610
rect 4245 19558 4257 19610
rect 4309 19558 4321 19610
rect 4373 19558 4385 19610
rect 4437 19558 4449 19610
rect 4501 19558 11783 19610
rect 11835 19558 11847 19610
rect 11899 19558 11911 19610
rect 11963 19558 11975 19610
rect 12027 19558 12039 19610
rect 12091 19558 19373 19610
rect 19425 19558 19437 19610
rect 19489 19558 19501 19610
rect 19553 19558 19565 19610
rect 19617 19558 19629 19610
rect 19681 19558 26963 19610
rect 27015 19558 27027 19610
rect 27079 19558 27091 19610
rect 27143 19558 27155 19610
rect 27207 19558 27219 19610
rect 27271 19558 30912 19610
rect 552 19536 30912 19558
rect 1210 19456 1216 19508
rect 1268 19496 1274 19508
rect 2961 19499 3019 19505
rect 2961 19496 2973 19499
rect 1268 19468 2973 19496
rect 1268 19456 1274 19468
rect 2961 19465 2973 19468
rect 3007 19496 3019 19499
rect 3786 19496 3792 19508
rect 3007 19468 3792 19496
rect 3007 19465 3019 19468
rect 2961 19459 3019 19465
rect 3786 19456 3792 19468
rect 3844 19456 3850 19508
rect 3881 19499 3939 19505
rect 3881 19465 3893 19499
rect 3927 19496 3939 19499
rect 8202 19496 8208 19508
rect 3927 19468 8208 19496
rect 3927 19465 3939 19468
rect 3881 19459 3939 19465
rect 8202 19456 8208 19468
rect 8260 19456 8266 19508
rect 8294 19456 8300 19508
rect 8352 19496 8358 19508
rect 8352 19468 9812 19496
rect 8352 19456 8358 19468
rect 5166 19388 5172 19440
rect 5224 19428 5230 19440
rect 5537 19431 5595 19437
rect 5224 19400 5396 19428
rect 5224 19388 5230 19400
rect 1302 19320 1308 19372
rect 1360 19320 1366 19372
rect 1578 19320 1584 19372
rect 1636 19360 1642 19372
rect 2222 19360 2228 19372
rect 1636 19332 2228 19360
rect 1636 19320 1642 19332
rect 2222 19320 2228 19332
rect 2280 19320 2286 19372
rect 3786 19320 3792 19372
rect 3844 19360 3850 19372
rect 3844 19332 4108 19360
rect 3844 19320 3850 19332
rect 842 19252 848 19304
rect 900 19252 906 19304
rect 1121 19295 1179 19301
rect 1121 19292 1133 19295
rect 952 19264 1133 19292
rect 658 19184 664 19236
rect 716 19224 722 19236
rect 952 19224 980 19264
rect 1121 19261 1133 19264
rect 1167 19261 1179 19295
rect 1320 19292 1348 19320
rect 1320 19264 2452 19292
rect 1121 19255 1179 19261
rect 716 19196 980 19224
rect 2424 19224 2452 19264
rect 2498 19252 2504 19304
rect 2556 19252 2562 19304
rect 3421 19295 3479 19301
rect 3421 19261 3433 19295
rect 3467 19292 3479 19295
rect 3970 19292 3976 19304
rect 3467 19264 3976 19292
rect 3467 19261 3479 19264
rect 3421 19255 3479 19261
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 4080 19301 4108 19332
rect 4065 19295 4123 19301
rect 4065 19261 4077 19295
rect 4111 19261 4123 19295
rect 4065 19255 4123 19261
rect 4341 19295 4399 19301
rect 4341 19261 4353 19295
rect 4387 19292 4399 19295
rect 5166 19292 5172 19304
rect 4387 19264 5172 19292
rect 4387 19261 4399 19264
rect 4341 19255 4399 19261
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 5368 19301 5396 19400
rect 5537 19397 5549 19431
rect 5583 19428 5595 19431
rect 5810 19428 5816 19440
rect 5583 19400 5816 19428
rect 5583 19397 5595 19400
rect 5537 19391 5595 19397
rect 5353 19295 5411 19301
rect 5353 19261 5365 19295
rect 5399 19261 5411 19295
rect 5552 19292 5580 19391
rect 5810 19388 5816 19400
rect 5868 19388 5874 19440
rect 7650 19388 7656 19440
rect 7708 19388 7714 19440
rect 9784 19428 9812 19468
rect 10226 19456 10232 19508
rect 10284 19456 10290 19508
rect 11238 19496 11244 19508
rect 10336 19468 11244 19496
rect 10336 19428 10364 19468
rect 11238 19456 11244 19468
rect 11296 19496 11302 19508
rect 11790 19496 11796 19508
rect 11296 19468 11796 19496
rect 11296 19456 11302 19468
rect 11790 19456 11796 19468
rect 11848 19456 11854 19508
rect 12618 19456 12624 19508
rect 12676 19496 12682 19508
rect 13081 19499 13139 19505
rect 13081 19496 13093 19499
rect 12676 19468 13093 19496
rect 12676 19456 12682 19468
rect 13081 19465 13093 19468
rect 13127 19465 13139 19499
rect 13081 19459 13139 19465
rect 14090 19456 14096 19508
rect 14148 19496 14154 19508
rect 16482 19496 16488 19508
rect 14148 19468 16488 19496
rect 14148 19456 14154 19468
rect 9784 19400 10364 19428
rect 11057 19431 11115 19437
rect 11057 19397 11069 19431
rect 11103 19428 11115 19431
rect 11146 19428 11152 19440
rect 11103 19400 11152 19428
rect 11103 19397 11115 19400
rect 11057 19391 11115 19397
rect 11146 19388 11152 19400
rect 11204 19388 11210 19440
rect 15930 19428 15936 19440
rect 13648 19400 15936 19428
rect 5626 19320 5632 19372
rect 5684 19360 5690 19372
rect 6276 19363 6334 19369
rect 6276 19360 6288 19363
rect 5684 19332 6288 19360
rect 5684 19320 5690 19332
rect 6276 19329 6288 19332
rect 6322 19329 6334 19363
rect 7668 19360 7696 19388
rect 6276 19323 6334 19329
rect 6380 19332 7696 19360
rect 5813 19295 5871 19301
rect 5813 19292 5825 19295
rect 5552 19264 5825 19292
rect 5353 19255 5411 19261
rect 5813 19261 5825 19264
rect 5859 19261 5871 19295
rect 6380 19292 6408 19332
rect 8386 19320 8392 19372
rect 8444 19320 8450 19372
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 8852 19363 8910 19369
rect 8852 19360 8864 19363
rect 8628 19332 8864 19360
rect 8628 19320 8634 19332
rect 8852 19329 8864 19332
rect 8898 19329 8910 19363
rect 8852 19323 8910 19329
rect 9030 19320 9036 19372
rect 9088 19360 9094 19372
rect 9306 19360 9312 19372
rect 9088 19332 9312 19360
rect 9088 19320 9094 19332
rect 9306 19320 9312 19332
rect 9364 19360 9370 19372
rect 11422 19360 11428 19372
rect 9364 19332 11428 19360
rect 9364 19320 9370 19332
rect 11422 19320 11428 19332
rect 11480 19360 11486 19372
rect 11568 19363 11626 19369
rect 11568 19360 11580 19363
rect 11480 19332 11580 19360
rect 11480 19320 11486 19332
rect 11568 19329 11580 19332
rect 11614 19329 11626 19363
rect 11568 19323 11626 19329
rect 11747 19363 11805 19369
rect 11747 19329 11759 19363
rect 11793 19360 11805 19363
rect 11793 19332 12434 19360
rect 11793 19329 11805 19332
rect 11747 19323 11805 19329
rect 5813 19255 5871 19261
rect 5920 19264 6408 19292
rect 2685 19227 2743 19233
rect 2685 19224 2697 19227
rect 2424 19196 2697 19224
rect 716 19184 722 19196
rect 2685 19193 2697 19196
rect 2731 19224 2743 19227
rect 2958 19224 2964 19236
rect 2731 19196 2964 19224
rect 2731 19193 2743 19196
rect 2685 19187 2743 19193
rect 2958 19184 2964 19196
rect 3016 19184 3022 19236
rect 3605 19227 3663 19233
rect 3605 19193 3617 19227
rect 3651 19224 3663 19227
rect 5920 19224 5948 19264
rect 6546 19252 6552 19304
rect 6604 19252 6610 19304
rect 7190 19252 7196 19304
rect 7248 19292 7254 19304
rect 8205 19295 8263 19301
rect 8205 19292 8217 19295
rect 7248 19264 8217 19292
rect 7248 19252 7254 19264
rect 8205 19261 8217 19264
rect 8251 19261 8263 19295
rect 8662 19292 8668 19304
rect 8205 19255 8263 19261
rect 8502 19264 8668 19292
rect 3651 19196 5948 19224
rect 7929 19227 7987 19233
rect 3651 19193 3663 19196
rect 3605 19187 3663 19193
rect 7929 19193 7941 19227
rect 7975 19224 7987 19227
rect 8502 19224 8530 19264
rect 8662 19252 8668 19264
rect 8720 19252 8726 19304
rect 9125 19295 9183 19301
rect 9125 19261 9137 19295
rect 9171 19292 9183 19295
rect 9858 19292 9864 19304
rect 9171 19264 9864 19292
rect 9171 19261 9183 19264
rect 9125 19255 9183 19261
rect 9858 19252 9864 19264
rect 9916 19252 9922 19304
rect 10134 19252 10140 19304
rect 10192 19292 10198 19304
rect 10192 19264 11192 19292
rect 10192 19252 10198 19264
rect 7975 19196 8530 19224
rect 7975 19193 7987 19196
rect 7929 19187 7987 19193
rect 10226 19184 10232 19236
rect 10284 19224 10290 19236
rect 10781 19227 10839 19233
rect 10781 19224 10793 19227
rect 10284 19196 10793 19224
rect 10284 19184 10290 19196
rect 10781 19193 10793 19196
rect 10827 19193 10839 19227
rect 11164 19224 11192 19264
rect 11238 19252 11244 19304
rect 11296 19252 11302 19304
rect 11977 19295 12035 19301
rect 11977 19292 11989 19295
rect 11348 19264 11989 19292
rect 11348 19224 11376 19264
rect 11977 19261 11989 19264
rect 12023 19261 12035 19295
rect 12406 19292 12434 19332
rect 12894 19320 12900 19372
rect 12952 19360 12958 19372
rect 13648 19360 13676 19400
rect 15930 19388 15936 19400
rect 15988 19388 15994 19440
rect 12952 19332 13676 19360
rect 14829 19363 14887 19369
rect 12952 19320 12958 19332
rect 14829 19329 14841 19363
rect 14875 19360 14887 19363
rect 14875 19332 15240 19360
rect 14875 19329 14887 19332
rect 14829 19323 14887 19329
rect 13817 19295 13875 19301
rect 12406 19264 13032 19292
rect 11977 19255 12035 19261
rect 13004 19236 13032 19264
rect 13817 19261 13829 19295
rect 13863 19292 13875 19295
rect 14918 19292 14924 19304
rect 13863 19264 14924 19292
rect 13863 19261 13875 19264
rect 13817 19255 13875 19261
rect 14918 19252 14924 19264
rect 14976 19252 14982 19304
rect 15102 19252 15108 19304
rect 15160 19252 15166 19304
rect 11164 19196 11376 19224
rect 10781 19187 10839 19193
rect 12986 19184 12992 19236
rect 13044 19184 13050 19236
rect 14550 19184 14556 19236
rect 14608 19224 14614 19236
rect 15212 19224 15240 19332
rect 16132 19301 16160 19468
rect 16482 19456 16488 19468
rect 16540 19456 16546 19508
rect 16850 19456 16856 19508
rect 16908 19496 16914 19508
rect 17678 19496 17684 19508
rect 16908 19468 17684 19496
rect 16908 19456 16914 19468
rect 17678 19456 17684 19468
rect 17736 19456 17742 19508
rect 17865 19499 17923 19505
rect 17865 19465 17877 19499
rect 17911 19496 17923 19499
rect 17954 19496 17960 19508
rect 17911 19468 17960 19496
rect 17911 19465 17923 19468
rect 17865 19459 17923 19465
rect 17954 19456 17960 19468
rect 18012 19456 18018 19508
rect 19150 19456 19156 19508
rect 19208 19496 19214 19508
rect 21910 19496 21916 19508
rect 19208 19468 21916 19496
rect 19208 19456 19214 19468
rect 21910 19456 21916 19468
rect 21968 19456 21974 19508
rect 22094 19456 22100 19508
rect 22152 19496 22158 19508
rect 22830 19496 22836 19508
rect 22152 19468 22836 19496
rect 22152 19456 22158 19468
rect 22830 19456 22836 19468
rect 22888 19456 22894 19508
rect 23566 19456 23572 19508
rect 23624 19456 23630 19508
rect 26510 19496 26516 19508
rect 24136 19468 26516 19496
rect 24136 19437 24164 19468
rect 26510 19456 26516 19468
rect 26568 19456 26574 19508
rect 30944 19496 30972 19672
rect 26712 19468 30972 19496
rect 24121 19431 24179 19437
rect 24121 19428 24133 19431
rect 22848 19400 24133 19428
rect 22848 19372 22876 19400
rect 24121 19397 24133 19400
rect 24167 19397 24179 19431
rect 24121 19391 24179 19397
rect 18138 19320 18144 19372
rect 18196 19320 18202 19372
rect 18230 19320 18236 19372
rect 18288 19360 18294 19372
rect 18288 19332 19288 19360
rect 18288 19320 18294 19332
rect 16117 19295 16175 19301
rect 16117 19261 16129 19295
rect 16163 19261 16175 19295
rect 16117 19255 16175 19261
rect 16393 19295 16451 19301
rect 16393 19261 16405 19295
rect 16439 19292 16451 19295
rect 17310 19292 17316 19304
rect 16439 19264 17316 19292
rect 16439 19261 16451 19264
rect 16393 19255 16451 19261
rect 17310 19252 17316 19264
rect 17368 19252 17374 19304
rect 17402 19252 17408 19304
rect 17460 19292 17466 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17460 19264 18061 19292
rect 17460 19252 17466 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 18325 19295 18383 19301
rect 18325 19261 18337 19295
rect 18371 19292 18383 19295
rect 18414 19292 18420 19304
rect 18371 19264 18420 19292
rect 18371 19261 18383 19264
rect 18325 19255 18383 19261
rect 18414 19252 18420 19264
rect 18472 19252 18478 19304
rect 18506 19252 18512 19304
rect 18564 19252 18570 19304
rect 18690 19252 18696 19304
rect 18748 19252 18754 19304
rect 18969 19295 19027 19301
rect 18969 19292 18981 19295
rect 18800 19264 18981 19292
rect 15378 19224 15384 19236
rect 14608 19196 15384 19224
rect 14608 19184 14614 19196
rect 15378 19184 15384 19196
rect 15436 19184 15442 19236
rect 15473 19227 15531 19233
rect 15473 19193 15485 19227
rect 15519 19224 15531 19227
rect 15841 19227 15899 19233
rect 15841 19224 15853 19227
rect 15519 19196 15853 19224
rect 15519 19193 15531 19196
rect 15473 19187 15531 19193
rect 15841 19193 15853 19196
rect 15887 19224 15899 19227
rect 16206 19224 16212 19236
rect 15887 19196 16212 19224
rect 15887 19193 15899 19196
rect 15841 19187 15899 19193
rect 16206 19184 16212 19196
rect 16264 19184 16270 19236
rect 17773 19227 17831 19233
rect 17773 19193 17785 19227
rect 17819 19224 17831 19227
rect 18800 19224 18828 19264
rect 18969 19261 18981 19264
rect 19015 19261 19027 19295
rect 19260 19292 19288 19332
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 21821 19363 21879 19369
rect 21821 19360 21833 19363
rect 19392 19332 21833 19360
rect 19392 19320 19398 19332
rect 21821 19329 21833 19332
rect 21867 19329 21879 19363
rect 21821 19323 21879 19329
rect 22830 19320 22836 19372
rect 22888 19320 22894 19372
rect 24995 19363 25053 19369
rect 24995 19329 25007 19363
rect 25041 19360 25053 19363
rect 26712 19360 26740 19468
rect 30282 19388 30288 19440
rect 30340 19388 30346 19440
rect 27246 19367 27252 19372
rect 25041 19332 26740 19360
rect 27203 19361 27252 19367
rect 25041 19329 25053 19332
rect 24995 19323 25053 19329
rect 27203 19327 27215 19361
rect 27249 19327 27252 19361
rect 27203 19321 27252 19327
rect 27246 19320 27252 19321
rect 27304 19320 27310 19372
rect 27338 19320 27344 19372
rect 27396 19369 27402 19372
rect 27396 19363 27445 19369
rect 27396 19329 27399 19363
rect 27433 19329 27445 19363
rect 29822 19360 29828 19372
rect 27396 19323 27445 19329
rect 29564 19332 29828 19360
rect 27396 19320 27402 19323
rect 19886 19292 19892 19304
rect 19260 19264 19892 19292
rect 18969 19255 19027 19261
rect 19886 19252 19892 19264
rect 19944 19252 19950 19304
rect 20070 19252 20076 19304
rect 20128 19294 20134 19304
rect 20349 19295 20407 19301
rect 20128 19292 20300 19294
rect 20349 19292 20361 19295
rect 20128 19266 20361 19292
rect 20128 19252 20134 19266
rect 20272 19264 20361 19266
rect 20349 19261 20361 19264
rect 20395 19261 20407 19295
rect 20349 19255 20407 19261
rect 20438 19252 20444 19304
rect 20496 19252 20502 19304
rect 20717 19295 20775 19301
rect 20717 19292 20729 19295
rect 20548 19264 20729 19292
rect 17819 19196 18828 19224
rect 17819 19193 17831 19196
rect 17773 19187 17831 19193
rect 20162 19184 20168 19236
rect 20220 19224 20226 19236
rect 20548 19224 20576 19264
rect 20717 19261 20729 19264
rect 20763 19292 20775 19295
rect 20806 19292 20812 19304
rect 20763 19264 20812 19292
rect 20763 19261 20775 19264
rect 20717 19255 20775 19261
rect 20806 19252 20812 19264
rect 20864 19292 20870 19304
rect 20864 19264 22094 19292
rect 20864 19252 20870 19264
rect 20220 19196 20576 19224
rect 20220 19184 20226 19196
rect 3234 19116 3240 19168
rect 3292 19116 3298 19168
rect 4982 19116 4988 19168
rect 5040 19116 5046 19168
rect 5169 19159 5227 19165
rect 5169 19125 5181 19159
rect 5215 19156 5227 19159
rect 5442 19156 5448 19168
rect 5215 19128 5448 19156
rect 5215 19125 5227 19128
rect 5169 19119 5227 19125
rect 5442 19116 5448 19128
rect 5500 19116 5506 19168
rect 5718 19116 5724 19168
rect 5776 19156 5782 19168
rect 6279 19159 6337 19165
rect 6279 19156 6291 19159
rect 5776 19128 6291 19156
rect 5776 19116 5782 19128
rect 6279 19125 6291 19128
rect 6325 19125 6337 19159
rect 6279 19119 6337 19125
rect 8021 19159 8079 19165
rect 8021 19125 8033 19159
rect 8067 19156 8079 19159
rect 8662 19156 8668 19168
rect 8067 19128 8668 19156
rect 8067 19125 8079 19128
rect 8021 19119 8079 19125
rect 8662 19116 8668 19128
rect 8720 19116 8726 19168
rect 8855 19159 8913 19165
rect 8855 19125 8867 19159
rect 8901 19156 8913 19159
rect 9214 19156 9220 19168
rect 8901 19128 9220 19156
rect 8901 19125 8913 19128
rect 8855 19119 8913 19125
rect 9214 19116 9220 19128
rect 9272 19156 9278 19168
rect 11238 19156 11244 19168
rect 9272 19128 11244 19156
rect 9272 19116 9278 19128
rect 11238 19116 11244 19128
rect 11296 19116 11302 19168
rect 11514 19116 11520 19168
rect 11572 19156 11578 19168
rect 13998 19156 14004 19168
rect 11572 19128 14004 19156
rect 11572 19116 11578 19128
rect 13998 19116 14004 19128
rect 14056 19156 14062 19168
rect 14274 19156 14280 19168
rect 14056 19128 14280 19156
rect 14056 19116 14062 19128
rect 14274 19116 14280 19128
rect 14332 19116 14338 19168
rect 14461 19159 14519 19165
rect 14461 19125 14473 19159
rect 14507 19156 14519 19159
rect 14826 19156 14832 19168
rect 14507 19128 14832 19156
rect 14507 19125 14519 19128
rect 14461 19119 14519 19125
rect 14826 19116 14832 19128
rect 14884 19116 14890 19168
rect 14918 19116 14924 19168
rect 14976 19116 14982 19168
rect 15102 19116 15108 19168
rect 15160 19156 15166 19168
rect 15933 19159 15991 19165
rect 15933 19156 15945 19159
rect 15160 19128 15945 19156
rect 15160 19116 15166 19128
rect 15933 19125 15945 19128
rect 15979 19125 15991 19159
rect 15933 19119 15991 19125
rect 16390 19116 16396 19168
rect 16448 19156 16454 19168
rect 16758 19156 16764 19168
rect 16448 19128 16764 19156
rect 16448 19116 16454 19128
rect 16758 19116 16764 19128
rect 16816 19116 16822 19168
rect 18322 19116 18328 19168
rect 18380 19156 18386 19168
rect 20254 19156 20260 19168
rect 18380 19128 20260 19156
rect 18380 19116 18386 19128
rect 20254 19116 20260 19128
rect 20312 19156 20318 19168
rect 20438 19156 20444 19168
rect 20312 19128 20444 19156
rect 20312 19116 20318 19128
rect 20438 19116 20444 19128
rect 20496 19116 20502 19168
rect 22066 19156 22094 19264
rect 22646 19252 22652 19304
rect 22704 19252 22710 19304
rect 23492 19264 24440 19292
rect 22462 19184 22468 19236
rect 22520 19184 22526 19236
rect 23492 19156 23520 19264
rect 23658 19184 23664 19236
rect 23716 19224 23722 19236
rect 23937 19227 23995 19233
rect 23937 19224 23949 19227
rect 23716 19196 23949 19224
rect 23716 19184 23722 19196
rect 23937 19193 23949 19196
rect 23983 19193 23995 19227
rect 24412 19224 24440 19264
rect 24486 19252 24492 19304
rect 24544 19252 24550 19304
rect 25130 19292 25136 19304
rect 24596 19264 25136 19292
rect 24596 19224 24624 19264
rect 25130 19252 25136 19264
rect 25188 19252 25194 19304
rect 25225 19295 25283 19301
rect 25225 19261 25237 19295
rect 25271 19292 25283 19295
rect 25498 19292 25504 19304
rect 25271 19264 25504 19292
rect 25271 19261 25283 19264
rect 25225 19255 25283 19261
rect 25498 19252 25504 19264
rect 25556 19252 25562 19304
rect 26694 19252 26700 19304
rect 26752 19252 26758 19304
rect 27024 19295 27082 19301
rect 27024 19261 27036 19295
rect 27070 19292 27082 19295
rect 27522 19292 27528 19304
rect 27070 19264 27528 19292
rect 27070 19261 27082 19264
rect 27024 19255 27082 19261
rect 27522 19252 27528 19264
rect 27580 19292 27586 19304
rect 28997 19295 29055 19301
rect 27580 19264 28856 19292
rect 27580 19252 27586 19264
rect 28828 19236 28856 19264
rect 28997 19261 29009 19295
rect 29043 19292 29055 19295
rect 29178 19292 29184 19304
rect 29043 19264 29184 19292
rect 29043 19261 29055 19264
rect 28997 19255 29055 19261
rect 29178 19252 29184 19264
rect 29236 19252 29242 19304
rect 29273 19295 29331 19301
rect 29273 19261 29285 19295
rect 29319 19292 29331 19295
rect 29564 19292 29592 19332
rect 29822 19320 29828 19332
rect 29880 19320 29886 19372
rect 29319 19264 29592 19292
rect 29319 19261 29331 19264
rect 29273 19255 29331 19261
rect 29638 19252 29644 19304
rect 29696 19292 29702 19304
rect 30193 19295 30251 19301
rect 30193 19292 30205 19295
rect 29696 19264 30205 19292
rect 29696 19252 29702 19264
rect 30193 19261 30205 19264
rect 30239 19261 30251 19295
rect 30193 19255 30251 19261
rect 24412 19196 24624 19224
rect 26252 19196 26832 19224
rect 23937 19187 23995 19193
rect 22066 19128 23520 19156
rect 24486 19116 24492 19168
rect 24544 19156 24550 19168
rect 24955 19159 25013 19165
rect 24955 19156 24967 19159
rect 24544 19128 24967 19156
rect 24544 19116 24550 19128
rect 24955 19125 24967 19128
rect 25001 19156 25013 19159
rect 26252 19156 26280 19196
rect 26804 19168 26832 19196
rect 28166 19184 28172 19236
rect 28224 19224 28230 19236
rect 28224 19196 28672 19224
rect 28224 19184 28230 19196
rect 25001 19128 26280 19156
rect 25001 19125 25013 19128
rect 24955 19119 25013 19125
rect 26326 19116 26332 19168
rect 26384 19116 26390 19168
rect 26786 19116 26792 19168
rect 26844 19116 26850 19168
rect 26970 19116 26976 19168
rect 27028 19156 27034 19168
rect 28537 19159 28595 19165
rect 28537 19156 28549 19159
rect 27028 19128 28549 19156
rect 27028 19116 27034 19128
rect 28537 19125 28549 19128
rect 28583 19125 28595 19159
rect 28644 19156 28672 19196
rect 28810 19184 28816 19236
rect 28868 19184 28874 19236
rect 29288 19196 30144 19224
rect 29288 19156 29316 19196
rect 28644 19128 29316 19156
rect 28537 19119 28595 19125
rect 29362 19116 29368 19168
rect 29420 19156 29426 19168
rect 30116 19165 30144 19196
rect 29917 19159 29975 19165
rect 29917 19156 29929 19159
rect 29420 19128 29929 19156
rect 29420 19116 29426 19128
rect 29917 19125 29929 19128
rect 29963 19125 29975 19159
rect 29917 19119 29975 19125
rect 30101 19159 30159 19165
rect 30101 19125 30113 19159
rect 30147 19125 30159 19159
rect 30101 19119 30159 19125
rect 552 19066 31072 19088
rect 552 19014 7988 19066
rect 8040 19014 8052 19066
rect 8104 19014 8116 19066
rect 8168 19014 8180 19066
rect 8232 19014 8244 19066
rect 8296 19014 15578 19066
rect 15630 19014 15642 19066
rect 15694 19014 15706 19066
rect 15758 19014 15770 19066
rect 15822 19014 15834 19066
rect 15886 19014 23168 19066
rect 23220 19014 23232 19066
rect 23284 19014 23296 19066
rect 23348 19014 23360 19066
rect 23412 19014 23424 19066
rect 23476 19014 30758 19066
rect 30810 19014 30822 19066
rect 30874 19014 30886 19066
rect 30938 19014 30950 19066
rect 31002 19014 31014 19066
rect 31066 19014 31072 19066
rect 552 18992 31072 19014
rect 1578 18912 1584 18964
rect 1636 18952 1642 18964
rect 1771 18955 1829 18961
rect 1771 18952 1783 18955
rect 1636 18924 1783 18952
rect 1636 18912 1642 18924
rect 1771 18921 1783 18924
rect 1817 18921 1829 18955
rect 1771 18915 1829 18921
rect 3050 18912 3056 18964
rect 3108 18912 3114 18964
rect 3234 18912 3240 18964
rect 3292 18952 3298 18964
rect 7929 18955 7987 18961
rect 3292 18924 7328 18952
rect 3292 18912 3298 18924
rect 1210 18776 1216 18828
rect 1268 18776 1274 18828
rect 2866 18816 2872 18828
rect 1964 18788 2872 18816
rect 1801 18769 1859 18775
rect 1302 18708 1308 18760
rect 1360 18708 1366 18760
rect 1801 18735 1813 18769
rect 1847 18748 1859 18769
rect 1964 18748 1992 18788
rect 2866 18776 2872 18788
rect 2924 18776 2930 18828
rect 2958 18776 2964 18828
rect 3016 18776 3022 18828
rect 3068 18816 3096 18912
rect 3418 18844 3424 18896
rect 3476 18844 3482 18896
rect 5626 18844 5632 18896
rect 5684 18844 5690 18896
rect 5810 18844 5816 18896
rect 5868 18844 5874 18896
rect 5828 18816 5856 18844
rect 6178 18816 6184 18828
rect 3068 18788 4019 18816
rect 5828 18788 6184 18816
rect 1847 18735 1992 18748
rect 1801 18729 1992 18735
rect 1826 18720 1992 18729
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18748 2099 18751
rect 2498 18748 2504 18760
rect 2087 18720 2504 18748
rect 2087 18717 2099 18720
rect 2041 18711 2099 18717
rect 2498 18708 2504 18720
rect 2556 18708 2562 18760
rect 2976 18748 3004 18776
rect 3513 18751 3571 18757
rect 3513 18748 3525 18751
rect 2976 18720 3525 18748
rect 3513 18717 3525 18720
rect 3559 18717 3571 18751
rect 3513 18711 3571 18717
rect 1029 18615 1087 18621
rect 1029 18581 1041 18615
rect 1075 18612 1087 18615
rect 3418 18612 3424 18624
rect 1075 18584 3424 18612
rect 1075 18581 1087 18584
rect 1029 18575 1087 18581
rect 3418 18572 3424 18584
rect 3476 18572 3482 18624
rect 3528 18612 3556 18711
rect 3694 18708 3700 18760
rect 3752 18748 3758 18760
rect 3991 18759 4019 18788
rect 6178 18776 6184 18788
rect 6236 18825 6242 18828
rect 6236 18819 6290 18825
rect 6236 18785 6244 18819
rect 6278 18785 6290 18819
rect 6236 18779 6290 18785
rect 6236 18776 6242 18779
rect 3840 18751 3898 18757
rect 3840 18748 3852 18751
rect 3752 18720 3852 18748
rect 3752 18708 3758 18720
rect 3840 18717 3852 18720
rect 3886 18717 3898 18751
rect 3840 18711 3898 18717
rect 3976 18753 4034 18759
rect 3976 18719 3988 18753
rect 4022 18719 4034 18753
rect 3976 18713 4034 18719
rect 4249 18751 4307 18757
rect 4249 18717 4261 18751
rect 4295 18748 4307 18751
rect 4982 18748 4988 18760
rect 4295 18720 4988 18748
rect 4295 18717 4307 18720
rect 4249 18711 4307 18717
rect 4982 18708 4988 18720
rect 5040 18708 5046 18760
rect 5905 18751 5963 18757
rect 5905 18717 5917 18751
rect 5951 18748 5963 18751
rect 6086 18748 6092 18760
rect 5951 18720 6092 18748
rect 5951 18717 5963 18720
rect 5905 18711 5963 18717
rect 6086 18708 6092 18720
rect 6144 18708 6150 18760
rect 6362 18708 6368 18760
rect 6420 18708 6426 18760
rect 6638 18708 6644 18760
rect 6696 18708 6702 18760
rect 5534 18680 5540 18692
rect 5092 18652 5540 18680
rect 5092 18612 5120 18652
rect 5534 18640 5540 18652
rect 5592 18640 5598 18692
rect 7300 18680 7328 18924
rect 7929 18921 7941 18955
rect 7975 18952 7987 18955
rect 8478 18952 8484 18964
rect 7975 18924 8484 18952
rect 7975 18921 7987 18924
rect 7929 18915 7987 18921
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 9030 18952 9036 18964
rect 8588 18924 9036 18952
rect 7466 18844 7472 18896
rect 7524 18884 7530 18896
rect 8389 18887 8447 18893
rect 8389 18884 8401 18887
rect 7524 18856 8401 18884
rect 7524 18844 7530 18856
rect 8389 18853 8401 18856
rect 8435 18884 8447 18887
rect 8588 18884 8616 18924
rect 9030 18912 9036 18924
rect 9088 18912 9094 18964
rect 9122 18912 9128 18964
rect 9180 18961 9186 18964
rect 9180 18952 9189 18961
rect 11054 18952 11060 18964
rect 9180 18924 11060 18952
rect 9180 18915 9189 18924
rect 9180 18912 9186 18915
rect 11054 18912 11060 18924
rect 11112 18912 11118 18964
rect 11422 18912 11428 18964
rect 11480 18952 11486 18964
rect 14007 18955 14065 18961
rect 14007 18952 14019 18955
rect 11480 18924 14019 18952
rect 11480 18912 11486 18924
rect 14007 18921 14019 18924
rect 14053 18921 14065 18955
rect 14007 18915 14065 18921
rect 14918 18912 14924 18964
rect 14976 18912 14982 18964
rect 15010 18912 15016 18964
rect 15068 18952 15074 18964
rect 15381 18955 15439 18961
rect 15381 18952 15393 18955
rect 15068 18924 15393 18952
rect 15068 18912 15074 18924
rect 15381 18921 15393 18924
rect 15427 18921 15439 18955
rect 15381 18915 15439 18921
rect 15930 18912 15936 18964
rect 15988 18952 15994 18964
rect 15988 18924 16160 18952
rect 15988 18912 15994 18924
rect 8435 18856 8616 18884
rect 13372 18856 13676 18884
rect 8435 18853 8447 18856
rect 8389 18847 8447 18853
rect 7374 18776 7380 18828
rect 7432 18816 7438 18828
rect 7742 18816 7748 18828
rect 7432 18788 7748 18816
rect 7432 18776 7438 18788
rect 7742 18776 7748 18788
rect 7800 18816 7806 18828
rect 8113 18819 8171 18825
rect 8113 18816 8125 18819
rect 7800 18788 8125 18816
rect 7800 18776 7806 18788
rect 8113 18785 8125 18788
rect 8159 18785 8171 18819
rect 8499 18816 8708 18820
rect 10781 18819 10839 18825
rect 8113 18779 8171 18785
rect 8266 18792 9444 18816
rect 8266 18788 8527 18792
rect 8680 18788 9444 18792
rect 8266 18680 8294 18788
rect 8478 18708 8484 18760
rect 8536 18748 8542 18760
rect 8665 18751 8723 18757
rect 8665 18748 8677 18751
rect 8536 18720 8677 18748
rect 8536 18708 8542 18720
rect 8665 18717 8677 18720
rect 8711 18717 8723 18751
rect 8665 18711 8723 18717
rect 8938 18708 8944 18760
rect 8996 18748 9002 18760
rect 9416 18757 9444 18788
rect 10781 18785 10793 18819
rect 10827 18816 10839 18819
rect 13372 18816 13400 18856
rect 10827 18788 13400 18816
rect 10827 18785 10839 18788
rect 10781 18779 10839 18785
rect 13446 18776 13452 18828
rect 13504 18776 13510 18828
rect 13648 18816 13676 18856
rect 14277 18819 14335 18825
rect 13648 18800 13955 18816
rect 13648 18788 14047 18800
rect 13927 18775 14047 18788
rect 14277 18785 14289 18819
rect 14323 18816 14335 18819
rect 14936 18816 14964 18912
rect 14323 18788 14964 18816
rect 14323 18785 14335 18788
rect 14277 18779 14335 18785
rect 15930 18776 15936 18828
rect 15988 18776 15994 18828
rect 16132 18825 16160 18924
rect 16482 18912 16488 18964
rect 16540 18952 16546 18964
rect 16540 18924 17724 18952
rect 16540 18912 16546 18924
rect 16117 18819 16175 18825
rect 16117 18785 16129 18819
rect 16163 18785 16175 18819
rect 17696 18816 17724 18924
rect 17770 18912 17776 18964
rect 17828 18952 17834 18964
rect 20622 18952 20628 18964
rect 17828 18924 20628 18952
rect 17828 18912 17834 18924
rect 20622 18912 20628 18924
rect 20680 18912 20686 18964
rect 21284 18924 22968 18952
rect 21284 18896 21312 18924
rect 19794 18844 19800 18896
rect 19852 18844 19858 18896
rect 21266 18844 21272 18896
rect 21324 18844 21330 18896
rect 22940 18884 22968 18924
rect 23014 18912 23020 18964
rect 23072 18952 23078 18964
rect 23385 18955 23443 18961
rect 23385 18952 23397 18955
rect 23072 18924 23397 18952
rect 23072 18912 23078 18924
rect 23385 18921 23397 18924
rect 23431 18921 23443 18955
rect 23385 18915 23443 18921
rect 23477 18955 23535 18961
rect 23477 18921 23489 18955
rect 23523 18952 23535 18955
rect 25682 18952 25688 18964
rect 23523 18924 25688 18952
rect 23523 18921 23535 18924
rect 23477 18915 23535 18921
rect 25682 18912 25688 18924
rect 25740 18912 25746 18964
rect 26970 18912 26976 18964
rect 27028 18912 27034 18964
rect 28810 18912 28816 18964
rect 28868 18961 28874 18964
rect 28868 18952 28877 18961
rect 28868 18924 28913 18952
rect 28868 18915 28877 18924
rect 28868 18912 28874 18915
rect 29086 18912 29092 18964
rect 29144 18952 29150 18964
rect 29362 18952 29368 18964
rect 29144 18924 29368 18952
rect 29144 18912 29150 18924
rect 29362 18912 29368 18924
rect 29420 18912 29426 18964
rect 30190 18912 30196 18964
rect 30248 18912 30254 18964
rect 24210 18884 24216 18896
rect 22940 18856 24216 18884
rect 24210 18844 24216 18856
rect 24268 18844 24274 18896
rect 26988 18884 27016 18912
rect 25516 18856 27016 18884
rect 18601 18819 18659 18825
rect 17696 18788 18276 18816
rect 16117 18779 16175 18785
rect 13927 18772 14062 18775
rect 14004 18769 14062 18772
rect 9128 18751 9186 18757
rect 9128 18748 9140 18751
rect 8996 18720 9140 18748
rect 8996 18708 9002 18720
rect 9128 18717 9140 18720
rect 9174 18717 9186 18751
rect 9128 18711 9186 18717
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18717 9459 18751
rect 9401 18711 9459 18717
rect 10962 18708 10968 18760
rect 11020 18708 11026 18760
rect 11244 18708 11250 18760
rect 11302 18757 11308 18760
rect 11514 18759 11520 18760
rect 11302 18751 11350 18757
rect 11302 18717 11304 18751
rect 11338 18717 11350 18751
rect 11302 18711 11350 18717
rect 11471 18753 11520 18759
rect 11471 18719 11483 18753
rect 11517 18719 11520 18753
rect 11471 18713 11520 18719
rect 11302 18708 11308 18711
rect 11514 18708 11520 18713
rect 11572 18708 11578 18760
rect 11698 18708 11704 18760
rect 11756 18708 11762 18760
rect 11790 18708 11796 18760
rect 11848 18748 11854 18760
rect 13541 18751 13599 18757
rect 13541 18748 13553 18751
rect 11848 18720 13553 18748
rect 11848 18708 11854 18720
rect 13541 18717 13553 18720
rect 13587 18717 13599 18751
rect 14004 18735 14016 18769
rect 14050 18735 14062 18769
rect 14004 18729 14062 18735
rect 13541 18711 13599 18717
rect 7300 18652 8294 18680
rect 12710 18640 12716 18692
rect 12768 18680 12774 18692
rect 12805 18683 12863 18689
rect 12805 18680 12817 18683
rect 12768 18652 12817 18680
rect 12768 18640 12774 18652
rect 12805 18649 12817 18652
rect 12851 18649 12863 18683
rect 12805 18643 12863 18649
rect 3528 18584 5120 18612
rect 5166 18572 5172 18624
rect 5224 18612 5230 18624
rect 13078 18612 13084 18624
rect 5224 18584 13084 18612
rect 5224 18572 5230 18584
rect 13078 18572 13084 18584
rect 13136 18572 13142 18624
rect 13262 18572 13268 18624
rect 13320 18572 13326 18624
rect 13556 18612 13584 18711
rect 14366 18708 14372 18760
rect 14424 18748 14430 18760
rect 16444 18751 16502 18757
rect 16444 18748 16456 18751
rect 14424 18720 16456 18748
rect 14424 18708 14430 18720
rect 16444 18717 16456 18720
rect 16490 18717 16502 18751
rect 16444 18711 16502 18717
rect 16580 18751 16638 18757
rect 16580 18717 16592 18751
rect 16626 18748 16638 18751
rect 16758 18748 16764 18760
rect 16626 18720 16764 18748
rect 16626 18717 16638 18720
rect 16580 18711 16638 18717
rect 16758 18708 16764 18720
rect 16816 18708 16822 18760
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18748 16911 18751
rect 17678 18748 17684 18760
rect 16899 18720 17684 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 17678 18708 17684 18720
rect 17736 18708 17742 18760
rect 14734 18612 14740 18624
rect 13556 18584 14740 18612
rect 14734 18572 14740 18584
rect 14792 18572 14798 18624
rect 15749 18615 15807 18621
rect 15749 18581 15761 18615
rect 15795 18612 15807 18615
rect 16482 18612 16488 18624
rect 15795 18584 16488 18612
rect 15795 18581 15807 18584
rect 15749 18575 15807 18581
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 18138 18572 18144 18624
rect 18196 18572 18202 18624
rect 18248 18612 18276 18788
rect 18601 18785 18613 18819
rect 18647 18816 18659 18819
rect 18966 18816 18972 18828
rect 18647 18788 18972 18816
rect 18647 18785 18659 18788
rect 18601 18779 18659 18785
rect 18966 18776 18972 18788
rect 19024 18776 19030 18828
rect 19812 18816 19840 18844
rect 20165 18819 20223 18825
rect 20165 18816 20177 18819
rect 19812 18788 20177 18816
rect 20165 18785 20177 18788
rect 20211 18785 20223 18819
rect 20165 18779 20223 18785
rect 20438 18776 20444 18828
rect 20496 18816 20502 18828
rect 20533 18819 20591 18825
rect 20533 18816 20545 18819
rect 20496 18788 20545 18816
rect 20496 18776 20502 18788
rect 20533 18785 20545 18788
rect 20579 18785 20591 18819
rect 21545 18819 21603 18825
rect 21545 18816 21557 18819
rect 20533 18779 20591 18785
rect 20640 18788 21557 18816
rect 18325 18751 18383 18757
rect 18325 18717 18337 18751
rect 18371 18748 18383 18751
rect 18690 18748 18696 18760
rect 18371 18720 18696 18748
rect 18371 18717 18383 18720
rect 18325 18711 18383 18717
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 18782 18708 18788 18760
rect 18840 18748 18846 18760
rect 19981 18751 20039 18757
rect 18840 18720 19334 18748
rect 18840 18708 18846 18720
rect 19306 18680 19334 18720
rect 19981 18717 19993 18751
rect 20027 18748 20039 18751
rect 20640 18748 20668 18788
rect 21545 18785 21557 18788
rect 21591 18785 21603 18819
rect 21545 18779 21603 18785
rect 22278 18776 22284 18828
rect 22336 18816 22342 18828
rect 22336 18788 23060 18816
rect 22336 18776 22342 18788
rect 20027 18720 20668 18748
rect 20027 18717 20039 18720
rect 19981 18711 20039 18717
rect 20806 18708 20812 18760
rect 20864 18748 20870 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20864 18720 20913 18748
rect 20864 18708 20870 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 21276 18751 21334 18757
rect 21276 18748 21288 18751
rect 20901 18711 20959 18717
rect 21008 18720 21288 18748
rect 21008 18680 21036 18720
rect 21276 18717 21288 18720
rect 21322 18748 21334 18751
rect 21450 18748 21456 18760
rect 21322 18720 21456 18748
rect 21322 18717 21334 18720
rect 21276 18711 21334 18717
rect 21450 18708 21456 18720
rect 21508 18708 21514 18760
rect 22002 18708 22008 18760
rect 22060 18748 22066 18760
rect 22646 18748 22652 18760
rect 22060 18720 22652 18748
rect 22060 18708 22066 18720
rect 22646 18708 22652 18720
rect 22704 18708 22710 18760
rect 22922 18708 22928 18760
rect 22980 18708 22986 18760
rect 23032 18748 23060 18788
rect 23842 18776 23848 18828
rect 23900 18816 23906 18828
rect 24486 18825 24492 18828
rect 24029 18819 24087 18825
rect 24029 18816 24041 18819
rect 23900 18788 24041 18816
rect 23900 18776 23906 18788
rect 24029 18785 24041 18788
rect 24075 18785 24087 18819
rect 24029 18779 24087 18785
rect 24448 18819 24492 18825
rect 24448 18785 24460 18819
rect 24448 18779 24492 18785
rect 24486 18776 24492 18779
rect 24544 18776 24550 18828
rect 25516 18816 25544 18856
rect 27890 18844 27896 18896
rect 27948 18884 27954 18896
rect 27948 18856 28488 18884
rect 27948 18844 27954 18856
rect 24780 18788 25544 18816
rect 23569 18751 23627 18757
rect 23569 18748 23581 18751
rect 23032 18720 23581 18748
rect 23569 18717 23581 18720
rect 23615 18717 23627 18751
rect 23569 18711 23627 18717
rect 24121 18751 24179 18757
rect 24121 18717 24133 18751
rect 24167 18717 24179 18751
rect 24121 18711 24179 18717
rect 24627 18751 24685 18757
rect 24627 18717 24639 18751
rect 24673 18748 24685 18751
rect 24780 18748 24808 18788
rect 25866 18776 25872 18828
rect 25924 18816 25930 18828
rect 26697 18819 26755 18825
rect 26697 18816 26709 18819
rect 25924 18788 26709 18816
rect 25924 18776 25930 18788
rect 26697 18785 26709 18788
rect 26743 18816 26755 18819
rect 26878 18816 26884 18828
rect 26743 18788 26884 18816
rect 26743 18785 26755 18788
rect 26697 18779 26755 18785
rect 26878 18776 26884 18788
rect 26936 18776 26942 18828
rect 28258 18776 28264 18828
rect 28316 18816 28322 18828
rect 28353 18819 28411 18825
rect 28353 18816 28365 18819
rect 28316 18788 28365 18816
rect 28316 18776 28322 18788
rect 28353 18785 28365 18788
rect 28399 18785 28411 18819
rect 28460 18816 28488 18856
rect 29362 18816 29368 18828
rect 28460 18788 29368 18816
rect 28353 18779 28411 18785
rect 24673 18720 24808 18748
rect 24857 18751 24915 18757
rect 24673 18717 24685 18720
rect 24627 18711 24685 18717
rect 24857 18717 24869 18751
rect 24903 18748 24915 18751
rect 26050 18748 26056 18760
rect 24903 18720 26056 18748
rect 24903 18717 24915 18720
rect 24857 18711 24915 18717
rect 19306 18652 21036 18680
rect 22940 18680 22968 18708
rect 23017 18683 23075 18689
rect 23017 18680 23029 18683
rect 22940 18652 23029 18680
rect 23017 18649 23029 18652
rect 23063 18649 23075 18683
rect 23017 18643 23075 18649
rect 20993 18615 21051 18621
rect 20993 18612 21005 18615
rect 18248 18584 21005 18612
rect 20993 18581 21005 18584
rect 21039 18581 21051 18615
rect 20993 18575 21051 18581
rect 22833 18615 22891 18621
rect 22833 18581 22845 18615
rect 22879 18612 22891 18615
rect 23750 18612 23756 18624
rect 22879 18584 23756 18612
rect 22879 18581 22891 18584
rect 22833 18575 22891 18581
rect 23750 18572 23756 18584
rect 23808 18572 23814 18624
rect 23842 18572 23848 18624
rect 23900 18572 23906 18624
rect 24136 18612 24164 18711
rect 26050 18708 26056 18720
rect 26108 18708 26114 18760
rect 26142 18708 26148 18760
rect 26200 18748 26206 18760
rect 26421 18751 26479 18757
rect 26421 18748 26433 18751
rect 26200 18720 26433 18748
rect 26200 18708 26206 18720
rect 26421 18717 26433 18720
rect 26467 18717 26479 18751
rect 26421 18711 26479 18717
rect 25516 18652 26096 18680
rect 24394 18612 24400 18624
rect 24136 18584 24400 18612
rect 24394 18572 24400 18584
rect 24452 18612 24458 18624
rect 25516 18612 25544 18652
rect 24452 18584 25544 18612
rect 24452 18572 24458 18584
rect 25590 18572 25596 18624
rect 25648 18612 25654 18624
rect 25961 18615 26019 18621
rect 25961 18612 25973 18615
rect 25648 18584 25973 18612
rect 25648 18572 25654 18584
rect 25961 18581 25973 18584
rect 26007 18581 26019 18615
rect 26068 18612 26096 18652
rect 27890 18640 27896 18692
rect 27948 18680 27954 18692
rect 27985 18683 28043 18689
rect 27985 18680 27997 18683
rect 27948 18652 27997 18680
rect 27948 18640 27954 18652
rect 27985 18649 27997 18652
rect 28031 18649 28043 18683
rect 28276 18680 28304 18776
rect 28966 18760 28994 18788
rect 29362 18776 29368 18788
rect 29420 18776 29426 18828
rect 28810 18708 28816 18760
rect 28868 18708 28874 18760
rect 28966 18720 29000 18760
rect 28994 18708 29000 18720
rect 29052 18708 29058 18760
rect 29086 18708 29092 18760
rect 29144 18708 29150 18760
rect 27985 18643 28043 18649
rect 28092 18652 28304 18680
rect 26418 18612 26424 18624
rect 26068 18584 26424 18612
rect 25961 18575 26019 18581
rect 26418 18572 26424 18584
rect 26476 18572 26482 18624
rect 26694 18572 26700 18624
rect 26752 18612 26758 18624
rect 28092 18612 28120 18652
rect 26752 18584 28120 18612
rect 26752 18572 26758 18584
rect 28166 18572 28172 18624
rect 28224 18612 28230 18624
rect 28261 18615 28319 18621
rect 28261 18612 28273 18615
rect 28224 18584 28273 18612
rect 28224 18572 28230 18584
rect 28261 18581 28273 18584
rect 28307 18581 28319 18615
rect 28261 18575 28319 18581
rect 28534 18572 28540 18624
rect 28592 18612 28598 18624
rect 31294 18612 31300 18624
rect 28592 18584 31300 18612
rect 28592 18572 28598 18584
rect 31294 18572 31300 18584
rect 31352 18572 31358 18624
rect 552 18522 30912 18544
rect 552 18470 4193 18522
rect 4245 18470 4257 18522
rect 4309 18470 4321 18522
rect 4373 18470 4385 18522
rect 4437 18470 4449 18522
rect 4501 18470 11783 18522
rect 11835 18470 11847 18522
rect 11899 18470 11911 18522
rect 11963 18470 11975 18522
rect 12027 18470 12039 18522
rect 12091 18470 19373 18522
rect 19425 18470 19437 18522
rect 19489 18470 19501 18522
rect 19553 18470 19565 18522
rect 19617 18470 19629 18522
rect 19681 18470 26963 18522
rect 27015 18470 27027 18522
rect 27079 18470 27091 18522
rect 27143 18470 27155 18522
rect 27207 18470 27219 18522
rect 27271 18470 30912 18522
rect 552 18448 30912 18470
rect 1210 18368 1216 18420
rect 1268 18408 1274 18420
rect 3602 18408 3608 18420
rect 1268 18380 3608 18408
rect 1268 18368 1274 18380
rect 3602 18368 3608 18380
rect 3660 18368 3666 18420
rect 3694 18368 3700 18420
rect 3752 18408 3758 18420
rect 5718 18408 5724 18420
rect 3752 18380 5724 18408
rect 3752 18368 3758 18380
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 5905 18411 5963 18417
rect 5905 18377 5917 18411
rect 5951 18408 5963 18411
rect 6362 18408 6368 18420
rect 5951 18380 6368 18408
rect 5951 18377 5963 18380
rect 5905 18371 5963 18377
rect 6362 18368 6368 18380
rect 6420 18368 6426 18420
rect 6914 18368 6920 18420
rect 6972 18408 6978 18420
rect 13630 18408 13636 18420
rect 6972 18380 13636 18408
rect 6972 18368 6978 18380
rect 13630 18368 13636 18380
rect 13688 18368 13694 18420
rect 17862 18408 17868 18420
rect 13832 18380 17868 18408
rect 2961 18343 3019 18349
rect 2961 18309 2973 18343
rect 3007 18340 3019 18343
rect 13832 18340 13860 18380
rect 17862 18368 17868 18380
rect 17920 18368 17926 18420
rect 18046 18368 18052 18420
rect 18104 18408 18110 18420
rect 21266 18408 21272 18420
rect 18104 18380 21272 18408
rect 18104 18368 18110 18380
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 21450 18368 21456 18420
rect 21508 18408 21514 18420
rect 22741 18411 22799 18417
rect 22741 18408 22753 18411
rect 21508 18380 22753 18408
rect 21508 18368 21514 18380
rect 22741 18377 22753 18380
rect 22787 18377 22799 18411
rect 22741 18371 22799 18377
rect 23750 18368 23756 18420
rect 23808 18408 23814 18420
rect 28445 18411 28503 18417
rect 23808 18380 26096 18408
rect 23808 18368 23814 18380
rect 3007 18312 3924 18340
rect 3007 18309 3019 18312
rect 2961 18303 3019 18309
rect 1443 18275 1501 18281
rect 1443 18241 1455 18275
rect 1489 18272 1501 18275
rect 3050 18272 3056 18284
rect 1489 18244 3056 18272
rect 1489 18241 1501 18244
rect 1443 18235 1501 18241
rect 3050 18232 3056 18244
rect 3108 18232 3114 18284
rect 3896 18272 3924 18312
rect 12176 18312 13860 18340
rect 4246 18272 4252 18284
rect 3896 18244 4252 18272
rect 4246 18232 4252 18244
rect 4304 18232 4310 18284
rect 4387 18275 4445 18281
rect 4387 18241 4399 18275
rect 4433 18272 4445 18275
rect 5534 18272 5540 18284
rect 4433 18244 5540 18272
rect 4433 18241 4445 18244
rect 4387 18235 4445 18241
rect 5534 18232 5540 18244
rect 5592 18232 5598 18284
rect 5626 18232 5632 18284
rect 5684 18272 5690 18284
rect 6552 18275 6610 18281
rect 6552 18272 6564 18275
rect 5684 18244 6564 18272
rect 5684 18232 5690 18244
rect 6552 18241 6564 18244
rect 6598 18241 6610 18275
rect 8386 18272 8392 18284
rect 6552 18235 6610 18241
rect 6748 18244 8392 18272
rect 937 18207 995 18213
rect 937 18173 949 18207
rect 983 18173 995 18207
rect 937 18167 995 18173
rect 952 18068 980 18167
rect 1670 18164 1676 18216
rect 1728 18164 1734 18216
rect 3237 18207 3295 18213
rect 3237 18173 3249 18207
rect 3283 18173 3295 18207
rect 3237 18167 3295 18173
rect 1210 18068 1216 18080
rect 952 18040 1216 18068
rect 1210 18028 1216 18040
rect 1268 18028 1274 18080
rect 1403 18071 1461 18077
rect 1403 18037 1415 18071
rect 1449 18068 1461 18071
rect 1578 18068 1584 18080
rect 1449 18040 1584 18068
rect 1449 18037 1461 18040
rect 1403 18031 1461 18037
rect 1578 18028 1584 18040
rect 1636 18068 1642 18080
rect 1762 18068 1768 18080
rect 1636 18040 1768 18068
rect 1636 18028 1642 18040
rect 1762 18028 1768 18040
rect 1820 18028 1826 18080
rect 3252 18068 3280 18167
rect 3602 18164 3608 18216
rect 3660 18204 3666 18216
rect 3881 18207 3939 18213
rect 3881 18204 3893 18207
rect 3660 18176 3893 18204
rect 3660 18164 3666 18176
rect 3881 18173 3893 18176
rect 3927 18204 3939 18207
rect 4522 18204 4528 18216
rect 3927 18176 4528 18204
rect 3927 18173 3939 18176
rect 3881 18167 3939 18173
rect 4522 18164 4528 18176
rect 4580 18164 4586 18216
rect 4617 18207 4675 18213
rect 4617 18173 4629 18207
rect 4663 18204 4675 18207
rect 4706 18204 4712 18216
rect 4663 18176 4712 18204
rect 4663 18173 4675 18176
rect 4617 18167 4675 18173
rect 4706 18164 4712 18176
rect 4764 18164 4770 18216
rect 5442 18164 5448 18216
rect 5500 18164 5506 18216
rect 6086 18164 6092 18216
rect 6144 18164 6150 18216
rect 6748 18204 6776 18244
rect 8386 18232 8392 18244
rect 8444 18272 8450 18284
rect 8573 18275 8631 18281
rect 8573 18272 8585 18275
rect 8444 18244 8585 18272
rect 8444 18232 8450 18244
rect 8573 18241 8585 18244
rect 8619 18272 8631 18275
rect 8938 18272 8944 18284
rect 8619 18244 8944 18272
rect 8619 18241 8631 18244
rect 8573 18235 8631 18241
rect 8938 18232 8944 18244
rect 8996 18232 9002 18284
rect 9122 18279 9128 18284
rect 9079 18273 9128 18279
rect 9079 18239 9091 18273
rect 9125 18239 9128 18273
rect 9079 18233 9128 18239
rect 9122 18232 9128 18233
rect 9180 18232 9186 18284
rect 9306 18232 9312 18284
rect 9364 18232 9370 18284
rect 10689 18275 10747 18281
rect 10689 18241 10701 18275
rect 10735 18272 10747 18275
rect 11244 18275 11302 18281
rect 11244 18272 11256 18275
rect 10735 18244 11256 18272
rect 10735 18241 10747 18244
rect 10689 18235 10747 18241
rect 11244 18241 11256 18244
rect 11290 18241 11302 18275
rect 11244 18235 11302 18241
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18272 11575 18275
rect 12176 18272 12204 18312
rect 15930 18300 15936 18352
rect 15988 18340 15994 18352
rect 16206 18340 16212 18352
rect 15988 18312 16212 18340
rect 15988 18300 15994 18312
rect 16206 18300 16212 18312
rect 16264 18300 16270 18352
rect 19242 18300 19248 18352
rect 19300 18340 19306 18352
rect 19300 18312 19840 18340
rect 19300 18300 19306 18312
rect 11563 18244 12204 18272
rect 11563 18241 11575 18244
rect 11517 18235 11575 18241
rect 12250 18232 12256 18284
rect 12308 18272 12314 18284
rect 14182 18281 14188 18284
rect 14144 18275 14188 18281
rect 12308 18244 13952 18272
rect 12308 18232 12314 18244
rect 6196 18176 6776 18204
rect 6825 18207 6883 18213
rect 3513 18139 3571 18145
rect 3513 18105 3525 18139
rect 3559 18136 3571 18139
rect 5460 18136 5488 18164
rect 6196 18136 6224 18176
rect 6825 18173 6837 18207
rect 6871 18204 6883 18207
rect 7466 18204 7472 18216
rect 6871 18176 7472 18204
rect 6871 18173 6883 18176
rect 6825 18167 6883 18173
rect 7466 18164 7472 18176
rect 7524 18164 7530 18216
rect 8478 18164 8484 18216
rect 8536 18204 8542 18216
rect 10781 18207 10839 18213
rect 10781 18204 10793 18207
rect 8536 18176 10793 18204
rect 8536 18164 8542 18176
rect 10781 18173 10793 18176
rect 10827 18173 10839 18207
rect 10781 18167 10839 18173
rect 13357 18207 13415 18213
rect 13357 18173 13369 18207
rect 13403 18204 13415 18207
rect 13538 18204 13544 18216
rect 13403 18176 13544 18204
rect 13403 18173 13415 18176
rect 13357 18167 13415 18173
rect 3559 18108 3924 18136
rect 5460 18108 6224 18136
rect 8036 18108 8616 18136
rect 3559 18105 3571 18108
rect 3513 18099 3571 18105
rect 3896 18080 3924 18108
rect 3694 18068 3700 18080
rect 3252 18040 3700 18068
rect 3694 18028 3700 18040
rect 3752 18028 3758 18080
rect 3878 18028 3884 18080
rect 3936 18068 3942 18080
rect 4347 18071 4405 18077
rect 4347 18068 4359 18071
rect 3936 18040 4359 18068
rect 3936 18028 3942 18040
rect 4347 18037 4359 18040
rect 4393 18037 4405 18071
rect 4347 18031 4405 18037
rect 5074 18028 5080 18080
rect 5132 18068 5138 18080
rect 5902 18068 5908 18080
rect 5132 18040 5908 18068
rect 5132 18028 5138 18040
rect 5902 18028 5908 18040
rect 5960 18028 5966 18080
rect 6178 18028 6184 18080
rect 6236 18068 6242 18080
rect 6555 18071 6613 18077
rect 6555 18068 6567 18071
rect 6236 18040 6567 18068
rect 6236 18028 6242 18040
rect 6555 18037 6567 18040
rect 6601 18068 6613 18071
rect 6730 18068 6736 18080
rect 6601 18040 6736 18068
rect 6601 18037 6613 18040
rect 6555 18031 6613 18037
rect 6730 18028 6736 18040
rect 6788 18028 6794 18080
rect 6822 18028 6828 18080
rect 6880 18068 6886 18080
rect 8036 18068 8064 18108
rect 6880 18040 8064 18068
rect 8113 18071 8171 18077
rect 6880 18028 6886 18040
rect 8113 18037 8125 18071
rect 8159 18068 8171 18071
rect 8478 18068 8484 18080
rect 8159 18040 8484 18068
rect 8159 18037 8171 18040
rect 8113 18031 8171 18037
rect 8478 18028 8484 18040
rect 8536 18028 8542 18080
rect 8588 18068 8616 18108
rect 10686 18096 10692 18148
rect 10744 18136 10750 18148
rect 10796 18136 10824 18167
rect 13538 18164 13544 18176
rect 13596 18204 13602 18216
rect 13722 18204 13728 18216
rect 13596 18176 13728 18204
rect 13596 18164 13602 18176
rect 13722 18164 13728 18176
rect 13780 18164 13786 18216
rect 13814 18164 13820 18216
rect 13872 18164 13878 18216
rect 13924 18204 13952 18244
rect 14144 18241 14156 18275
rect 14144 18235 14188 18241
rect 14182 18232 14188 18235
rect 14240 18232 14246 18284
rect 14323 18275 14381 18281
rect 14323 18241 14335 18275
rect 14369 18272 14381 18275
rect 17034 18272 17040 18284
rect 14369 18244 16252 18272
rect 14369 18241 14381 18244
rect 14323 18235 14381 18241
rect 14553 18207 14611 18213
rect 14553 18204 14565 18207
rect 13924 18176 14565 18204
rect 14553 18173 14565 18176
rect 14599 18173 14611 18207
rect 14553 18167 14611 18173
rect 10744 18108 10824 18136
rect 16224 18136 16252 18244
rect 16776 18244 17040 18272
rect 16776 18213 16804 18244
rect 17034 18232 17040 18244
rect 17092 18232 17098 18284
rect 17126 18232 17132 18284
rect 17184 18232 17190 18284
rect 17310 18232 17316 18284
rect 17368 18272 17374 18284
rect 17368 18244 17908 18272
rect 17368 18232 17374 18244
rect 16301 18207 16359 18213
rect 16301 18173 16313 18207
rect 16347 18204 16359 18207
rect 16761 18207 16819 18213
rect 16761 18204 16773 18207
rect 16347 18176 16773 18204
rect 16347 18173 16359 18176
rect 16301 18167 16359 18173
rect 16761 18173 16773 18176
rect 16807 18173 16819 18207
rect 16761 18167 16819 18173
rect 16850 18164 16856 18216
rect 16908 18164 16914 18216
rect 17880 18204 17908 18244
rect 18322 18232 18328 18284
rect 18380 18272 18386 18284
rect 18693 18275 18751 18281
rect 18693 18272 18705 18275
rect 18380 18244 18705 18272
rect 18380 18232 18386 18244
rect 18693 18241 18705 18244
rect 18739 18241 18751 18275
rect 19812 18272 19840 18312
rect 19886 18300 19892 18352
rect 19944 18340 19950 18352
rect 20073 18343 20131 18349
rect 20073 18340 20085 18343
rect 19944 18312 20085 18340
rect 19944 18300 19950 18312
rect 20073 18309 20085 18312
rect 20119 18309 20131 18343
rect 20073 18303 20131 18309
rect 24394 18300 24400 18352
rect 24452 18300 24458 18352
rect 20349 18275 20407 18281
rect 19812 18244 20300 18272
rect 18693 18235 18751 18241
rect 18969 18207 19027 18213
rect 18969 18204 18981 18207
rect 16960 18176 17816 18204
rect 17880 18176 18981 18204
rect 16960 18136 16988 18176
rect 16224 18108 16988 18136
rect 10744 18096 10750 18108
rect 9030 18068 9036 18080
rect 9088 18077 9094 18080
rect 8588 18040 9036 18068
rect 9030 18028 9036 18040
rect 9088 18068 9097 18077
rect 9088 18040 9133 18068
rect 9088 18031 9097 18040
rect 9088 18028 9094 18031
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11247 18071 11305 18077
rect 11247 18068 11259 18071
rect 11112 18040 11259 18068
rect 11112 18028 11118 18040
rect 11247 18037 11259 18040
rect 11293 18037 11305 18071
rect 11247 18031 11305 18037
rect 12621 18071 12679 18077
rect 12621 18037 12633 18071
rect 12667 18068 12679 18071
rect 12986 18068 12992 18080
rect 12667 18040 12992 18068
rect 12667 18037 12679 18040
rect 12621 18031 12679 18037
rect 12986 18028 12992 18040
rect 13044 18028 13050 18080
rect 13170 18028 13176 18080
rect 13228 18028 13234 18080
rect 13906 18028 13912 18080
rect 13964 18068 13970 18080
rect 15657 18071 15715 18077
rect 15657 18068 15669 18071
rect 13964 18040 15669 18068
rect 13964 18028 13970 18040
rect 15657 18037 15669 18040
rect 15703 18037 15715 18071
rect 15657 18031 15715 18037
rect 15838 18028 15844 18080
rect 15896 18068 15902 18080
rect 16390 18068 16396 18080
rect 15896 18040 16396 18068
rect 15896 18028 15902 18040
rect 16390 18028 16396 18040
rect 16448 18028 16454 18080
rect 16577 18071 16635 18077
rect 16577 18037 16589 18071
rect 16623 18068 16635 18071
rect 17126 18068 17132 18080
rect 16623 18040 17132 18068
rect 16623 18037 16635 18040
rect 16577 18031 16635 18037
rect 17126 18028 17132 18040
rect 17184 18028 17190 18080
rect 17788 18068 17816 18176
rect 18969 18173 18981 18176
rect 19015 18204 19027 18207
rect 20162 18204 20168 18216
rect 19015 18176 20168 18204
rect 19015 18173 19027 18176
rect 18969 18167 19027 18173
rect 20162 18164 20168 18176
rect 20220 18164 20226 18216
rect 20272 18213 20300 18244
rect 20349 18241 20361 18275
rect 20395 18272 20407 18275
rect 20530 18272 20536 18284
rect 20395 18244 20536 18272
rect 20395 18241 20407 18244
rect 20349 18235 20407 18241
rect 20530 18232 20536 18244
rect 20588 18232 20594 18284
rect 20855 18275 20913 18281
rect 20855 18241 20867 18275
rect 20901 18272 20913 18275
rect 24026 18272 24032 18284
rect 20901 18244 24032 18272
rect 20901 18241 20913 18244
rect 20855 18235 20913 18241
rect 24026 18232 24032 18244
rect 24084 18232 24090 18284
rect 24210 18232 24216 18284
rect 24268 18272 24274 18284
rect 24673 18275 24731 18281
rect 24673 18272 24685 18275
rect 24268 18244 24685 18272
rect 24268 18232 24274 18244
rect 24673 18241 24685 18244
rect 24719 18241 24731 18275
rect 24673 18235 24731 18241
rect 24854 18232 24860 18284
rect 24912 18232 24918 18284
rect 25179 18275 25237 18281
rect 25179 18241 25191 18275
rect 25225 18272 25237 18275
rect 25590 18272 25596 18284
rect 25225 18244 25596 18272
rect 25225 18241 25237 18244
rect 25179 18235 25237 18241
rect 25590 18232 25596 18244
rect 25648 18232 25654 18284
rect 26068 18272 26096 18380
rect 26160 18380 28396 18408
rect 26160 18352 26188 18380
rect 26142 18300 26148 18352
rect 26200 18300 26206 18352
rect 28368 18340 28396 18380
rect 28445 18377 28457 18411
rect 28491 18408 28503 18411
rect 30098 18408 30104 18420
rect 28491 18380 30104 18408
rect 28491 18377 28503 18380
rect 28445 18371 28503 18377
rect 30098 18368 30104 18380
rect 30156 18368 30162 18420
rect 30282 18368 30288 18420
rect 30340 18368 30346 18420
rect 28718 18340 28724 18352
rect 28368 18312 28724 18340
rect 28718 18300 28724 18312
rect 28776 18300 28782 18352
rect 29730 18300 29736 18352
rect 29788 18340 29794 18352
rect 30374 18340 30380 18352
rect 29788 18312 30380 18340
rect 29788 18300 29794 18312
rect 30374 18300 30380 18312
rect 30432 18340 30438 18352
rect 30432 18312 30604 18340
rect 30432 18300 30438 18312
rect 27157 18275 27215 18281
rect 27157 18272 27169 18275
rect 26068 18244 27169 18272
rect 27157 18241 27169 18244
rect 27203 18241 27215 18275
rect 28736 18270 28764 18300
rect 28997 18275 29055 18281
rect 28997 18272 29009 18275
rect 28920 18270 29009 18272
rect 28736 18244 29009 18270
rect 28736 18242 28948 18244
rect 27157 18235 27215 18241
rect 28997 18241 29009 18244
rect 29043 18241 29055 18275
rect 28997 18235 29055 18241
rect 20257 18207 20315 18213
rect 20257 18173 20269 18207
rect 20303 18173 20315 18207
rect 20257 18167 20315 18173
rect 21085 18207 21143 18213
rect 21085 18173 21097 18207
rect 21131 18204 21143 18207
rect 21726 18204 21732 18216
rect 21131 18176 21732 18204
rect 21131 18173 21143 18176
rect 21085 18167 21143 18173
rect 21726 18164 21732 18176
rect 21784 18164 21790 18216
rect 22066 18176 23244 18204
rect 18509 18139 18567 18145
rect 18509 18105 18521 18139
rect 18555 18136 18567 18139
rect 19610 18136 19616 18148
rect 18555 18108 19616 18136
rect 18555 18105 18567 18108
rect 18509 18099 18567 18105
rect 19610 18096 19616 18108
rect 19668 18096 19674 18148
rect 19794 18096 19800 18148
rect 19852 18096 19858 18148
rect 17954 18068 17960 18080
rect 17788 18040 17960 18068
rect 17954 18028 17960 18040
rect 18012 18028 18018 18080
rect 19978 18028 19984 18080
rect 20036 18028 20042 18080
rect 20806 18028 20812 18080
rect 20864 18077 20870 18080
rect 20864 18068 20873 18077
rect 20864 18040 20909 18068
rect 20864 18031 20873 18040
rect 20864 18028 20870 18031
rect 20990 18028 20996 18080
rect 21048 18068 21054 18080
rect 22066 18068 22094 18176
rect 22462 18096 22468 18148
rect 22520 18136 22526 18148
rect 22649 18139 22707 18145
rect 22649 18136 22661 18139
rect 22520 18108 22661 18136
rect 22520 18096 22526 18108
rect 22649 18105 22661 18108
rect 22695 18136 22707 18139
rect 22830 18136 22836 18148
rect 22695 18108 22836 18136
rect 22695 18105 22707 18108
rect 22649 18099 22707 18105
rect 22830 18096 22836 18108
rect 22888 18096 22894 18148
rect 23216 18145 23244 18176
rect 24578 18164 24584 18216
rect 24636 18164 24642 18216
rect 24872 18204 24900 18232
rect 25409 18207 25467 18213
rect 25409 18204 25421 18207
rect 24872 18176 25421 18204
rect 25409 18173 25421 18176
rect 25455 18173 25467 18207
rect 25409 18167 25467 18173
rect 26050 18164 26056 18216
rect 26108 18164 26114 18216
rect 26510 18164 26516 18216
rect 26568 18204 26574 18216
rect 26881 18207 26939 18213
rect 26881 18204 26893 18207
rect 26568 18176 26893 18204
rect 26568 18164 26574 18176
rect 26881 18173 26893 18176
rect 26927 18173 26939 18207
rect 28534 18204 28540 18216
rect 26881 18167 26939 18173
rect 26988 18176 28540 18204
rect 23201 18139 23259 18145
rect 23201 18105 23213 18139
rect 23247 18136 23259 18139
rect 23247 18108 23428 18136
rect 23247 18105 23259 18108
rect 23201 18099 23259 18105
rect 21048 18040 22094 18068
rect 21048 18028 21054 18040
rect 22186 18028 22192 18080
rect 22244 18028 22250 18080
rect 23400 18068 23428 18108
rect 23566 18096 23572 18148
rect 23624 18096 23630 18148
rect 23750 18096 23756 18148
rect 23808 18136 23814 18148
rect 23937 18139 23995 18145
rect 23937 18136 23949 18139
rect 23808 18108 23949 18136
rect 23808 18096 23814 18108
rect 23937 18105 23949 18108
rect 23983 18136 23995 18139
rect 24118 18136 24124 18148
rect 23983 18108 24124 18136
rect 23983 18105 23995 18108
rect 23937 18099 23995 18105
rect 24118 18096 24124 18108
rect 24176 18096 24182 18148
rect 26068 18136 26096 18164
rect 26988 18136 27016 18176
rect 28534 18164 28540 18176
rect 28592 18164 28598 18216
rect 28813 18207 28871 18213
rect 28813 18173 28825 18207
rect 28859 18204 28871 18207
rect 29273 18207 29331 18213
rect 28859 18176 28948 18204
rect 28859 18173 28871 18176
rect 28813 18167 28871 18173
rect 28920 18148 28948 18176
rect 29273 18173 29285 18207
rect 29319 18204 29331 18207
rect 29730 18204 29736 18216
rect 29319 18201 29408 18204
rect 29656 18201 29736 18204
rect 29319 18176 29736 18201
rect 29319 18173 29331 18176
rect 29380 18173 29684 18176
rect 29273 18167 29331 18173
rect 29730 18164 29736 18176
rect 29788 18164 29794 18216
rect 30576 18213 30604 18312
rect 30101 18207 30159 18213
rect 30101 18173 30113 18207
rect 30147 18204 30159 18207
rect 30561 18207 30619 18213
rect 30147 18176 30512 18204
rect 30147 18173 30159 18176
rect 30101 18167 30159 18173
rect 26068 18108 27016 18136
rect 27890 18096 27896 18148
rect 27948 18136 27954 18148
rect 27948 18108 28764 18136
rect 27948 18096 27954 18108
rect 24029 18071 24087 18077
rect 24029 18068 24041 18071
rect 23400 18040 24041 18068
rect 24029 18037 24041 18040
rect 24075 18037 24087 18071
rect 24029 18031 24087 18037
rect 24946 18028 24952 18080
rect 25004 18068 25010 18080
rect 25139 18071 25197 18077
rect 25139 18068 25151 18071
rect 25004 18040 25151 18068
rect 25004 18028 25010 18040
rect 25139 18037 25151 18040
rect 25185 18037 25197 18071
rect 25139 18031 25197 18037
rect 25314 18028 25320 18080
rect 25372 18068 25378 18080
rect 26513 18071 26571 18077
rect 26513 18068 26525 18071
rect 25372 18040 26525 18068
rect 25372 18028 25378 18040
rect 26513 18037 26525 18040
rect 26559 18037 26571 18071
rect 26513 18031 26571 18037
rect 28350 18028 28356 18080
rect 28408 18068 28414 18080
rect 28629 18071 28687 18077
rect 28629 18068 28641 18071
rect 28408 18040 28641 18068
rect 28408 18028 28414 18040
rect 28629 18037 28641 18040
rect 28675 18037 28687 18071
rect 28736 18068 28764 18108
rect 28902 18096 28908 18148
rect 28960 18096 28966 18148
rect 29104 18108 30420 18136
rect 29104 18068 29132 18108
rect 28736 18040 29132 18068
rect 28629 18031 28687 18037
rect 29822 18028 29828 18080
rect 29880 18068 29886 18080
rect 30006 18068 30012 18080
rect 29880 18040 30012 18068
rect 29880 18028 29886 18040
rect 30006 18028 30012 18040
rect 30064 18028 30070 18080
rect 30392 18077 30420 18108
rect 30377 18071 30435 18077
rect 30377 18037 30389 18071
rect 30423 18037 30435 18071
rect 30484 18068 30512 18176
rect 30561 18173 30573 18207
rect 30607 18173 30619 18207
rect 30561 18167 30619 18173
rect 30484 18040 31156 18068
rect 30377 18031 30435 18037
rect 552 17978 31072 18000
rect 552 17926 7988 17978
rect 8040 17926 8052 17978
rect 8104 17926 8116 17978
rect 8168 17926 8180 17978
rect 8232 17926 8244 17978
rect 8296 17926 15578 17978
rect 15630 17926 15642 17978
rect 15694 17926 15706 17978
rect 15758 17926 15770 17978
rect 15822 17926 15834 17978
rect 15886 17926 23168 17978
rect 23220 17926 23232 17978
rect 23284 17926 23296 17978
rect 23348 17926 23360 17978
rect 23412 17926 23424 17978
rect 23476 17926 30758 17978
rect 30810 17926 30822 17978
rect 30874 17926 30886 17978
rect 30938 17926 30950 17978
rect 31002 17926 31014 17978
rect 31066 17926 31072 17978
rect 552 17904 31072 17926
rect 937 17867 995 17873
rect 937 17833 949 17867
rect 983 17864 995 17867
rect 1302 17864 1308 17876
rect 983 17836 1308 17864
rect 983 17833 995 17836
rect 937 17827 995 17833
rect 1302 17824 1308 17836
rect 1360 17824 1366 17876
rect 1762 17824 1768 17876
rect 1820 17873 1826 17876
rect 1820 17864 1829 17873
rect 1820 17836 3096 17864
rect 1820 17827 1829 17836
rect 1820 17824 1826 17827
rect 3068 17796 3096 17836
rect 3142 17824 3148 17876
rect 3200 17824 3206 17876
rect 3418 17824 3424 17876
rect 3476 17864 3482 17876
rect 8754 17864 8760 17876
rect 3476 17836 8760 17864
rect 3476 17824 3482 17836
rect 8754 17824 8760 17836
rect 8812 17824 8818 17876
rect 8938 17824 8944 17876
rect 8996 17864 9002 17876
rect 9131 17867 9189 17873
rect 9131 17864 9143 17867
rect 8996 17836 9143 17864
rect 8996 17824 9002 17836
rect 9131 17833 9143 17836
rect 9177 17864 9189 17867
rect 9674 17864 9680 17876
rect 9177 17836 9680 17864
rect 9177 17833 9189 17836
rect 9131 17827 9189 17833
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 10686 17824 10692 17876
rect 10744 17864 10750 17876
rect 11146 17864 11152 17876
rect 10744 17836 11152 17864
rect 10744 17824 10750 17836
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 11983 17867 12041 17873
rect 11983 17833 11995 17867
rect 12029 17864 12041 17867
rect 12158 17864 12164 17876
rect 12029 17836 12164 17864
rect 12029 17833 12041 17836
rect 11983 17827 12041 17833
rect 12158 17824 12164 17836
rect 12216 17824 12222 17876
rect 13556 17836 15240 17864
rect 13556 17808 13584 17836
rect 3068 17768 3648 17796
rect 1121 17731 1179 17737
rect 1121 17697 1133 17731
rect 1167 17728 1179 17731
rect 3142 17728 3148 17740
rect 1167 17700 1716 17728
rect 1167 17697 1179 17700
rect 1121 17691 1179 17697
rect 1688 17672 1716 17700
rect 1964 17700 3148 17728
rect 1305 17663 1363 17669
rect 1305 17629 1317 17663
rect 1351 17629 1363 17663
rect 1305 17623 1363 17629
rect 1210 17484 1216 17536
rect 1268 17524 1274 17536
rect 1320 17524 1348 17623
rect 1670 17620 1676 17672
rect 1728 17620 1734 17672
rect 1811 17665 1869 17671
rect 1811 17631 1823 17665
rect 1857 17660 1869 17665
rect 1964 17660 1992 17700
rect 3142 17688 3148 17700
rect 3200 17688 3206 17740
rect 3510 17688 3516 17740
rect 3568 17688 3574 17740
rect 3620 17728 3648 17768
rect 5626 17756 5632 17808
rect 5684 17756 5690 17808
rect 5718 17756 5724 17808
rect 5776 17796 5782 17808
rect 6089 17799 6147 17805
rect 6089 17796 6101 17799
rect 5776 17768 6101 17796
rect 5776 17756 5782 17768
rect 6089 17765 6101 17768
rect 6135 17765 6147 17799
rect 6089 17759 6147 17765
rect 3620 17700 3883 17728
rect 1857 17632 1992 17660
rect 2041 17663 2099 17669
rect 1857 17631 1869 17632
rect 1811 17625 1869 17631
rect 2041 17629 2053 17663
rect 2087 17660 2099 17663
rect 3234 17660 3240 17672
rect 2087 17632 3240 17660
rect 2087 17629 2099 17632
rect 2041 17623 2099 17629
rect 3234 17620 3240 17632
rect 3292 17620 3298 17672
rect 3528 17524 3556 17688
rect 3855 17672 3883 17700
rect 4172 17700 5672 17728
rect 4009 17681 4067 17687
rect 4009 17678 4021 17681
rect 3855 17669 3884 17672
rect 3840 17663 3884 17669
rect 3840 17629 3852 17663
rect 3840 17623 3884 17629
rect 3878 17620 3884 17623
rect 3936 17620 3942 17672
rect 4007 17647 4021 17678
rect 4055 17660 4067 17681
rect 4172 17660 4200 17700
rect 5644 17672 5672 17700
rect 5810 17688 5816 17740
rect 5868 17688 5874 17740
rect 6104 17728 6132 17759
rect 8570 17756 8576 17808
rect 8628 17756 8634 17808
rect 8662 17756 8668 17808
rect 8720 17756 8726 17808
rect 10778 17756 10784 17808
rect 10836 17756 10842 17808
rect 11330 17796 11336 17808
rect 11164 17768 11336 17796
rect 6104 17700 6684 17728
rect 6656 17672 6684 17700
rect 6730 17688 6736 17740
rect 6788 17737 6794 17740
rect 6788 17731 6842 17737
rect 6788 17697 6796 17731
rect 6830 17697 6842 17731
rect 6788 17691 6842 17697
rect 7193 17731 7251 17737
rect 7193 17697 7205 17731
rect 7239 17697 7251 17731
rect 8680 17728 8708 17756
rect 11164 17740 11192 17768
rect 11330 17756 11336 17768
rect 11388 17756 11394 17808
rect 13538 17756 13544 17808
rect 13596 17756 13602 17808
rect 9214 17728 9220 17740
rect 8680 17700 9220 17728
rect 7193 17691 7251 17697
rect 6788 17688 6794 17691
rect 4055 17647 4200 17660
rect 4007 17632 4200 17647
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 5442 17660 5448 17672
rect 4295 17632 5448 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 5442 17620 5448 17632
rect 5500 17620 5506 17672
rect 5626 17620 5632 17672
rect 5684 17620 5690 17672
rect 6086 17620 6092 17672
rect 6144 17660 6150 17672
rect 6457 17663 6515 17669
rect 6457 17660 6469 17663
rect 6144 17632 6469 17660
rect 6144 17620 6150 17632
rect 6457 17629 6469 17632
rect 6503 17629 6515 17663
rect 6457 17623 6515 17629
rect 6638 17620 6644 17672
rect 6696 17620 6702 17672
rect 6920 17665 6978 17671
rect 6920 17631 6932 17665
rect 6966 17660 6978 17665
rect 7006 17660 7012 17672
rect 6966 17632 7012 17660
rect 6966 17631 6978 17632
rect 6920 17625 6978 17631
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 7208 17660 7236 17691
rect 9214 17688 9220 17700
rect 9272 17688 9278 17740
rect 9401 17731 9459 17737
rect 9401 17697 9413 17731
rect 9447 17728 9459 17731
rect 9490 17728 9496 17740
rect 9447 17700 9496 17728
rect 9447 17697 9459 17700
rect 9401 17691 9459 17697
rect 9490 17688 9496 17700
rect 9548 17688 9554 17740
rect 11057 17731 11115 17737
rect 11057 17697 11069 17731
rect 11103 17728 11115 17731
rect 11146 17728 11152 17740
rect 11103 17700 11152 17728
rect 11103 17697 11115 17700
rect 11057 17691 11115 17697
rect 11146 17688 11152 17700
rect 11204 17688 11210 17740
rect 11238 17688 11244 17740
rect 11296 17728 11302 17740
rect 11517 17731 11575 17737
rect 11517 17728 11529 17731
rect 11296 17700 11529 17728
rect 11296 17688 11302 17700
rect 11517 17697 11529 17700
rect 11563 17728 11575 17731
rect 11606 17728 11612 17740
rect 11563 17700 11612 17728
rect 11563 17697 11575 17700
rect 11517 17691 11575 17697
rect 11606 17688 11612 17700
rect 11664 17688 11670 17740
rect 12176 17700 12434 17728
rect 8202 17660 8208 17672
rect 7208 17632 8208 17660
rect 8202 17620 8208 17632
rect 8260 17620 8266 17672
rect 8665 17663 8723 17669
rect 8665 17629 8677 17663
rect 8711 17629 8723 17663
rect 8665 17623 8723 17629
rect 8386 17552 8392 17604
rect 8444 17592 8450 17604
rect 8680 17592 8708 17623
rect 8846 17620 8852 17672
rect 8904 17660 8910 17672
rect 9128 17663 9186 17669
rect 9128 17660 9140 17663
rect 8904 17632 9140 17660
rect 8904 17620 8910 17632
rect 9128 17629 9140 17632
rect 9174 17629 9186 17663
rect 9128 17623 9186 17629
rect 12023 17663 12081 17669
rect 12023 17629 12035 17663
rect 12069 17660 12081 17663
rect 12176 17660 12204 17700
rect 12069 17632 12204 17660
rect 12069 17629 12081 17632
rect 12023 17623 12081 17629
rect 12250 17620 12256 17672
rect 12308 17620 12314 17672
rect 12406 17660 12434 17700
rect 13170 17688 13176 17740
rect 13228 17728 13234 17740
rect 14553 17731 14611 17737
rect 14553 17728 14565 17731
rect 13228 17700 14565 17728
rect 13228 17688 13234 17700
rect 14553 17697 14565 17700
rect 14599 17697 14611 17731
rect 15212 17728 15240 17836
rect 15286 17824 15292 17876
rect 15344 17864 15350 17876
rect 15657 17867 15715 17873
rect 15657 17864 15669 17867
rect 15344 17836 15669 17864
rect 15344 17824 15350 17836
rect 15657 17833 15669 17836
rect 15703 17833 15715 17867
rect 15657 17827 15715 17833
rect 16206 17824 16212 17876
rect 16264 17864 16270 17876
rect 16574 17864 16580 17876
rect 16264 17836 16580 17864
rect 16264 17824 16270 17836
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 16666 17824 16672 17876
rect 16724 17864 16730 17876
rect 16761 17867 16819 17873
rect 16761 17864 16773 17867
rect 16724 17836 16773 17864
rect 16724 17824 16730 17836
rect 16761 17833 16773 17836
rect 16807 17833 16819 17867
rect 17310 17864 17316 17876
rect 16761 17827 16819 17833
rect 17052 17836 17316 17864
rect 15562 17756 15568 17808
rect 15620 17796 15626 17808
rect 16022 17796 16028 17808
rect 15620 17768 16028 17796
rect 15620 17756 15626 17768
rect 16022 17756 16028 17768
rect 16080 17796 16086 17808
rect 17052 17796 17080 17836
rect 17310 17824 17316 17836
rect 17368 17824 17374 17876
rect 23109 17867 23167 17873
rect 23109 17864 23121 17867
rect 18432 17836 23121 17864
rect 16080 17768 17080 17796
rect 16080 17756 16086 17768
rect 16298 17728 16304 17740
rect 15212 17700 16304 17728
rect 14553 17691 14611 17697
rect 16298 17688 16304 17700
rect 16356 17688 16362 17740
rect 16500 17737 16528 17768
rect 16485 17731 16543 17737
rect 16485 17697 16497 17731
rect 16531 17728 16543 17731
rect 17272 17731 17330 17737
rect 17272 17728 17284 17731
rect 16531 17700 16565 17728
rect 16868 17700 17284 17728
rect 16531 17697 16543 17700
rect 16485 17691 16543 17697
rect 12406 17632 13768 17660
rect 8444 17564 8708 17592
rect 10060 17564 11284 17592
rect 8444 17552 8450 17564
rect 1268 17496 3556 17524
rect 1268 17484 1274 17496
rect 5810 17484 5816 17536
rect 5868 17524 5874 17536
rect 10060 17524 10088 17564
rect 5868 17496 10088 17524
rect 5868 17484 5874 17496
rect 10410 17484 10416 17536
rect 10468 17524 10474 17536
rect 11149 17527 11207 17533
rect 11149 17524 11161 17527
rect 10468 17496 11161 17524
rect 10468 17484 10474 17496
rect 11149 17493 11161 17496
rect 11195 17493 11207 17527
rect 11256 17524 11284 17564
rect 12250 17524 12256 17536
rect 11256 17496 12256 17524
rect 11149 17487 11207 17493
rect 12250 17484 12256 17496
rect 12308 17484 12314 17536
rect 12710 17484 12716 17536
rect 12768 17524 12774 17536
rect 13357 17527 13415 17533
rect 13357 17524 13369 17527
rect 12768 17496 13369 17524
rect 12768 17484 12774 17496
rect 13357 17493 13369 17496
rect 13403 17493 13415 17527
rect 13740 17524 13768 17632
rect 13814 17620 13820 17672
rect 13872 17620 13878 17672
rect 14182 17669 14188 17672
rect 14144 17663 14188 17669
rect 14144 17629 14156 17663
rect 14144 17623 14188 17629
rect 14182 17620 14188 17623
rect 14240 17620 14246 17672
rect 14323 17663 14381 17669
rect 14323 17629 14335 17663
rect 14369 17660 14381 17663
rect 14369 17632 16160 17660
rect 14369 17629 14381 17632
rect 14323 17623 14381 17629
rect 16132 17592 16160 17632
rect 16206 17620 16212 17672
rect 16264 17620 16270 17672
rect 16316 17660 16344 17688
rect 16868 17672 16896 17700
rect 17272 17697 17284 17700
rect 17318 17697 17330 17731
rect 18432 17728 18460 17836
rect 23109 17833 23121 17836
rect 23155 17833 23167 17867
rect 23934 17864 23940 17876
rect 23109 17827 23167 17833
rect 23676 17836 23940 17864
rect 17272 17691 17330 17697
rect 17610 17700 18460 17728
rect 17441 17681 17499 17687
rect 16316 17632 16620 17660
rect 16298 17592 16304 17604
rect 16132 17564 16304 17592
rect 16298 17552 16304 17564
rect 16356 17552 16362 17604
rect 15378 17524 15384 17536
rect 13740 17496 15384 17524
rect 13357 17487 13415 17493
rect 15378 17484 15384 17496
rect 15436 17484 15442 17536
rect 16592 17524 16620 17632
rect 16666 17620 16672 17672
rect 16724 17620 16730 17672
rect 16850 17620 16856 17672
rect 16908 17620 16914 17672
rect 16945 17663 17003 17669
rect 16945 17629 16957 17663
rect 16991 17629 17003 17663
rect 17441 17647 17453 17681
rect 17487 17660 17499 17681
rect 17610 17660 17638 17700
rect 18782 17688 18788 17740
rect 18840 17728 18846 17740
rect 19153 17731 19211 17737
rect 19153 17728 19165 17731
rect 18840 17700 19165 17728
rect 18840 17688 18846 17700
rect 19153 17697 19165 17700
rect 19199 17697 19211 17731
rect 19153 17691 19211 17697
rect 19429 17731 19487 17737
rect 19429 17697 19441 17731
rect 19475 17728 19487 17731
rect 20070 17728 20076 17740
rect 19475 17700 20076 17728
rect 19475 17697 19487 17700
rect 19429 17691 19487 17697
rect 20070 17688 20076 17700
rect 20128 17688 20134 17740
rect 20254 17688 20260 17740
rect 20312 17728 20318 17740
rect 21085 17731 21143 17737
rect 21085 17728 21097 17731
rect 20312 17700 21097 17728
rect 20312 17688 20318 17700
rect 21085 17697 21097 17700
rect 21131 17728 21143 17731
rect 22005 17731 22063 17737
rect 21131 17700 21220 17728
rect 21131 17697 21143 17700
rect 21085 17691 21143 17697
rect 17487 17647 17638 17660
rect 17441 17641 17638 17647
rect 17456 17632 17638 17641
rect 17681 17663 17739 17669
rect 16945 17623 17003 17629
rect 17681 17629 17693 17663
rect 17727 17660 17739 17663
rect 19518 17660 19524 17672
rect 17727 17632 19524 17660
rect 17727 17629 17739 17632
rect 17681 17623 17739 17629
rect 16684 17592 16712 17620
rect 16960 17592 16988 17623
rect 19518 17620 19524 17632
rect 19576 17620 19582 17672
rect 21192 17604 21220 17700
rect 22005 17697 22017 17731
rect 22051 17728 22063 17731
rect 22051 17700 22968 17728
rect 22051 17697 22063 17700
rect 22005 17691 22063 17697
rect 21266 17620 21272 17672
rect 21324 17620 21330 17672
rect 21450 17620 21456 17672
rect 21508 17660 21514 17672
rect 21596 17663 21654 17669
rect 21596 17660 21608 17663
rect 21508 17632 21608 17660
rect 21508 17620 21514 17632
rect 21596 17629 21608 17632
rect 21642 17629 21654 17663
rect 21596 17623 21654 17629
rect 21775 17663 21833 17669
rect 21775 17629 21787 17663
rect 21821 17660 21833 17663
rect 22940 17660 22968 17700
rect 23014 17688 23020 17740
rect 23072 17728 23078 17740
rect 23676 17737 23704 17836
rect 23934 17824 23940 17836
rect 23992 17824 23998 17876
rect 24026 17824 24032 17876
rect 24084 17864 24090 17876
rect 25961 17867 26019 17873
rect 25961 17864 25973 17867
rect 24084 17836 25973 17864
rect 24084 17824 24090 17836
rect 25961 17833 25973 17836
rect 26007 17833 26019 17867
rect 25961 17827 26019 17833
rect 26786 17824 26792 17876
rect 26844 17864 26850 17876
rect 26887 17867 26945 17873
rect 26887 17864 26899 17867
rect 26844 17836 26899 17864
rect 26844 17824 26850 17836
rect 26887 17833 26899 17836
rect 26933 17833 26945 17867
rect 26887 17827 26945 17833
rect 27062 17824 27068 17876
rect 27120 17864 27126 17876
rect 28534 17864 28540 17876
rect 27120 17836 28540 17864
rect 27120 17824 27126 17836
rect 28534 17824 28540 17836
rect 28592 17824 28598 17876
rect 28718 17824 28724 17876
rect 28776 17864 28782 17876
rect 29270 17864 29276 17876
rect 28776 17836 29276 17864
rect 28776 17824 28782 17836
rect 29270 17824 29276 17836
rect 29328 17864 29334 17876
rect 29638 17864 29644 17876
rect 29328 17836 29644 17864
rect 29328 17824 29334 17836
rect 29638 17824 29644 17836
rect 29696 17824 29702 17876
rect 28258 17756 28264 17808
rect 28316 17796 28322 17808
rect 28736 17796 28764 17824
rect 28316 17768 28396 17796
rect 28316 17756 28322 17768
rect 23661 17731 23719 17737
rect 23661 17728 23673 17731
rect 23072 17700 23673 17728
rect 23072 17688 23078 17700
rect 23661 17697 23673 17700
rect 23707 17697 23719 17731
rect 23661 17691 23719 17697
rect 23842 17688 23848 17740
rect 23900 17688 23906 17740
rect 24121 17731 24179 17737
rect 24121 17697 24133 17731
rect 24167 17728 24179 17731
rect 24210 17728 24216 17740
rect 24167 17700 24216 17728
rect 24167 17697 24179 17700
rect 24121 17691 24179 17697
rect 24210 17688 24216 17700
rect 24268 17688 24274 17740
rect 24394 17688 24400 17740
rect 24452 17737 24458 17740
rect 24452 17731 24506 17737
rect 24452 17697 24460 17731
rect 24494 17728 24506 17731
rect 24946 17728 24952 17740
rect 24494 17700 24952 17728
rect 24494 17697 24506 17700
rect 24452 17691 24506 17697
rect 24452 17688 24458 17691
rect 24946 17688 24952 17700
rect 25004 17688 25010 17740
rect 25222 17688 25228 17740
rect 25280 17728 25286 17740
rect 25866 17728 25872 17740
rect 25280 17700 25872 17728
rect 25280 17688 25286 17700
rect 25866 17688 25872 17700
rect 25924 17688 25930 17740
rect 23860 17660 23888 17688
rect 21821 17632 22876 17660
rect 22940 17632 23888 17660
rect 24627 17663 24685 17669
rect 21821 17629 21833 17632
rect 21775 17623 21833 17629
rect 20901 17595 20959 17601
rect 20901 17592 20913 17595
rect 16684 17564 16988 17592
rect 20088 17564 20913 17592
rect 18322 17524 18328 17536
rect 16592 17496 18328 17524
rect 18322 17484 18328 17496
rect 18380 17484 18386 17536
rect 18782 17484 18788 17536
rect 18840 17484 18846 17536
rect 19150 17484 19156 17536
rect 19208 17524 19214 17536
rect 20088 17524 20116 17564
rect 20901 17561 20913 17564
rect 20947 17561 20959 17595
rect 20901 17555 20959 17561
rect 21174 17552 21180 17604
rect 21232 17552 21238 17604
rect 22848 17592 22876 17632
rect 24627 17629 24639 17663
rect 24673 17660 24685 17663
rect 24762 17660 24768 17672
rect 24673 17632 24768 17660
rect 24673 17629 24685 17632
rect 24627 17623 24685 17629
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 24857 17663 24915 17669
rect 24857 17629 24869 17663
rect 24903 17660 24915 17663
rect 25590 17660 25596 17672
rect 24903 17632 25596 17660
rect 24903 17629 24915 17632
rect 24857 17623 24915 17629
rect 25590 17620 25596 17632
rect 25648 17620 25654 17672
rect 26142 17620 26148 17672
rect 26200 17660 26206 17672
rect 26418 17660 26424 17672
rect 26200 17632 26424 17660
rect 26200 17620 26206 17632
rect 26418 17620 26424 17632
rect 26476 17620 26482 17672
rect 26878 17620 26884 17672
rect 26936 17660 26942 17672
rect 27157 17663 27215 17669
rect 26936 17632 26981 17660
rect 26936 17620 26942 17632
rect 27157 17629 27169 17663
rect 27203 17660 27215 17663
rect 28368 17660 28396 17768
rect 28644 17768 28764 17796
rect 28644 17737 28672 17768
rect 28629 17731 28687 17737
rect 28629 17697 28641 17731
rect 28675 17697 28687 17731
rect 31128 17728 31156 18040
rect 30038 17714 31156 17728
rect 28629 17691 28687 17697
rect 30024 17700 31156 17714
rect 28460 17660 28491 17662
rect 27203 17632 28304 17660
rect 28368 17632 28494 17660
rect 27203 17629 27215 17632
rect 27157 17623 27215 17629
rect 22848 17564 23888 17592
rect 19208 17496 20116 17524
rect 20717 17527 20775 17533
rect 19208 17484 19214 17496
rect 20717 17493 20729 17527
rect 20763 17524 20775 17527
rect 21542 17524 21548 17536
rect 20763 17496 21548 17524
rect 20763 17493 20775 17496
rect 20717 17487 20775 17493
rect 21542 17484 21548 17496
rect 21600 17484 21606 17536
rect 23860 17524 23888 17564
rect 23934 17552 23940 17604
rect 23992 17552 23998 17604
rect 25774 17524 25780 17536
rect 23860 17496 25780 17524
rect 25774 17484 25780 17496
rect 25832 17484 25838 17536
rect 28276 17524 28304 17632
rect 28466 17601 28494 17632
rect 28534 17620 28540 17672
rect 28592 17660 28598 17672
rect 28905 17663 28963 17669
rect 28905 17660 28917 17663
rect 28592 17632 28917 17660
rect 28592 17620 28598 17632
rect 28905 17629 28917 17632
rect 28951 17629 28963 17663
rect 28905 17623 28963 17629
rect 28994 17620 29000 17672
rect 29052 17660 29058 17672
rect 29270 17660 29276 17672
rect 29052 17632 29276 17660
rect 29052 17620 29058 17632
rect 29270 17620 29276 17632
rect 29328 17660 29334 17672
rect 30024 17660 30052 17700
rect 29328 17632 30052 17660
rect 29328 17620 29334 17632
rect 28445 17595 28503 17601
rect 28445 17561 28457 17595
rect 28491 17561 28503 17595
rect 28445 17555 28503 17561
rect 30374 17552 30380 17604
rect 30432 17552 30438 17604
rect 30650 17524 30656 17536
rect 28276 17496 30656 17524
rect 30650 17484 30656 17496
rect 30708 17484 30714 17536
rect 552 17434 30912 17456
rect 552 17382 4193 17434
rect 4245 17382 4257 17434
rect 4309 17382 4321 17434
rect 4373 17382 4385 17434
rect 4437 17382 4449 17434
rect 4501 17382 11783 17434
rect 11835 17382 11847 17434
rect 11899 17382 11911 17434
rect 11963 17382 11975 17434
rect 12027 17382 12039 17434
rect 12091 17382 19373 17434
rect 19425 17382 19437 17434
rect 19489 17382 19501 17434
rect 19553 17382 19565 17434
rect 19617 17382 19629 17434
rect 19681 17382 26963 17434
rect 27015 17382 27027 17434
rect 27079 17382 27091 17434
rect 27143 17382 27155 17434
rect 27207 17382 27219 17434
rect 27271 17382 30912 17434
rect 552 17360 30912 17382
rect 2961 17323 3019 17329
rect 2961 17289 2973 17323
rect 3007 17320 3019 17323
rect 5718 17320 5724 17332
rect 3007 17292 5724 17320
rect 3007 17289 3019 17292
rect 2961 17283 3019 17289
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 5810 17280 5816 17332
rect 5868 17280 5874 17332
rect 9214 17320 9220 17332
rect 6104 17292 9220 17320
rect 6104 17252 6132 17292
rect 9214 17280 9220 17292
rect 9272 17280 9278 17332
rect 9306 17280 9312 17332
rect 9364 17320 9370 17332
rect 10505 17323 10563 17329
rect 10505 17320 10517 17323
rect 9364 17292 10517 17320
rect 9364 17280 9370 17292
rect 10505 17289 10517 17292
rect 10551 17289 10563 17323
rect 12158 17320 12164 17332
rect 10505 17283 10563 17289
rect 11262 17292 12164 17320
rect 5276 17224 6132 17252
rect 8389 17255 8447 17261
rect 5276 17196 5304 17224
rect 8389 17221 8401 17255
rect 8435 17221 8447 17255
rect 8389 17215 8447 17221
rect 937 17187 995 17193
rect 937 17153 949 17187
rect 983 17184 995 17187
rect 1210 17184 1216 17196
rect 983 17156 1216 17184
rect 983 17153 995 17156
rect 937 17147 995 17153
rect 1210 17144 1216 17156
rect 1268 17144 1274 17196
rect 1673 17187 1731 17193
rect 1418 17169 1624 17184
rect 1418 17138 1445 17169
rect 1433 17135 1445 17138
rect 1479 17156 1624 17169
rect 1479 17135 1491 17156
rect 1433 17129 1491 17135
rect 1596 17116 1624 17156
rect 1673 17153 1685 17187
rect 1719 17184 1731 17187
rect 2130 17184 2136 17196
rect 1719 17156 2136 17184
rect 1719 17153 1731 17156
rect 1673 17147 1731 17153
rect 2130 17144 2136 17156
rect 2188 17144 2194 17196
rect 3326 17144 3332 17196
rect 3384 17184 3390 17196
rect 3510 17184 3516 17196
rect 3384 17156 3516 17184
rect 3384 17144 3390 17156
rect 3510 17144 3516 17156
rect 3568 17144 3574 17196
rect 3835 17187 3893 17193
rect 3835 17153 3847 17187
rect 3881 17184 3893 17187
rect 3881 17156 4660 17184
rect 3881 17153 3893 17156
rect 3835 17147 3893 17153
rect 2958 17116 2964 17128
rect 1596 17088 2964 17116
rect 2958 17076 2964 17088
rect 3016 17076 3022 17128
rect 3656 17119 3714 17125
rect 3656 17085 3668 17119
rect 3702 17116 3714 17119
rect 3970 17116 3976 17128
rect 3702 17088 3976 17116
rect 3702 17085 3714 17088
rect 3656 17079 3714 17085
rect 3970 17076 3976 17088
rect 4028 17076 4034 17128
rect 4065 17119 4123 17125
rect 4065 17085 4077 17119
rect 4111 17116 4123 17119
rect 4522 17116 4528 17128
rect 4111 17088 4528 17116
rect 4111 17085 4123 17088
rect 4065 17079 4123 17085
rect 4522 17076 4528 17088
rect 4580 17076 4586 17128
rect 4632 17116 4660 17156
rect 5258 17144 5264 17196
rect 5316 17144 5322 17196
rect 5445 17187 5503 17193
rect 5445 17153 5457 17187
rect 5491 17184 5503 17187
rect 6552 17187 6610 17193
rect 6552 17184 6564 17187
rect 5491 17156 6564 17184
rect 5491 17153 5503 17156
rect 5445 17147 5503 17153
rect 6552 17153 6564 17156
rect 6598 17153 6610 17187
rect 6552 17147 6610 17153
rect 6822 17144 6828 17196
rect 6880 17144 6886 17196
rect 8404 17128 8432 17215
rect 8478 17212 8484 17264
rect 8536 17212 8542 17264
rect 10594 17212 10600 17264
rect 10652 17252 10658 17264
rect 10870 17252 10876 17264
rect 10652 17224 10876 17252
rect 10652 17212 10658 17224
rect 10870 17212 10876 17224
rect 10928 17252 10934 17264
rect 11057 17255 11115 17261
rect 11057 17252 11069 17255
rect 10928 17224 11069 17252
rect 10928 17212 10934 17224
rect 11057 17221 11069 17224
rect 11103 17221 11115 17255
rect 11057 17215 11115 17221
rect 8496 17184 8524 17212
rect 8665 17187 8723 17193
rect 8665 17184 8677 17187
rect 8496 17156 8677 17184
rect 8665 17153 8677 17156
rect 8711 17153 8723 17187
rect 9128 17187 9186 17193
rect 9128 17184 9140 17187
rect 8665 17147 8723 17153
rect 8772 17156 9140 17184
rect 5997 17119 6055 17125
rect 4632 17088 5764 17116
rect 5736 16992 5764 17088
rect 5997 17085 6009 17119
rect 6043 17085 6055 17119
rect 5997 17079 6055 17085
rect 1403 16983 1461 16989
rect 1403 16949 1415 16983
rect 1449 16980 1461 16983
rect 1762 16980 1768 16992
rect 1449 16952 1768 16980
rect 1449 16949 1461 16952
rect 1403 16943 1461 16949
rect 1762 16940 1768 16952
rect 1820 16940 1826 16992
rect 3878 16940 3884 16992
rect 3936 16980 3942 16992
rect 5074 16980 5080 16992
rect 3936 16952 5080 16980
rect 3936 16940 3942 16952
rect 5074 16940 5080 16952
rect 5132 16940 5138 16992
rect 5718 16940 5724 16992
rect 5776 16940 5782 16992
rect 6012 16980 6040 17079
rect 6086 17076 6092 17128
rect 6144 17076 6150 17128
rect 6178 17076 6184 17128
rect 6236 17116 6242 17128
rect 6416 17119 6474 17125
rect 6416 17116 6428 17119
rect 6236 17088 6428 17116
rect 6236 17076 6242 17088
rect 6416 17085 6428 17088
rect 6462 17116 6474 17119
rect 7098 17116 7104 17128
rect 6462 17088 7104 17116
rect 6462 17085 6474 17088
rect 6416 17079 6474 17085
rect 7098 17076 7104 17088
rect 7156 17076 7162 17128
rect 8386 17076 8392 17128
rect 8444 17076 8450 17128
rect 8570 17076 8576 17128
rect 8628 17076 8634 17128
rect 8205 17051 8263 17057
rect 8205 17017 8217 17051
rect 8251 17048 8263 17051
rect 8251 17020 8432 17048
rect 8251 17017 8263 17020
rect 8205 17011 8263 17017
rect 6914 16980 6920 16992
rect 6012 16952 6920 16980
rect 6914 16940 6920 16952
rect 6972 16940 6978 16992
rect 8404 16980 8432 17020
rect 8772 16980 8800 17156
rect 9128 17153 9140 17156
rect 9174 17153 9186 17187
rect 9128 17147 9186 17153
rect 9214 17144 9220 17196
rect 9272 17184 9278 17196
rect 9401 17187 9459 17193
rect 9401 17184 9413 17187
rect 9272 17156 9413 17184
rect 9272 17144 9278 17156
rect 9401 17153 9413 17156
rect 9447 17153 9459 17187
rect 11262 17184 11290 17292
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 12342 17280 12348 17332
rect 12400 17320 12406 17332
rect 14090 17320 14096 17332
rect 12400 17292 14096 17320
rect 12400 17280 12406 17292
rect 14090 17280 14096 17292
rect 14148 17280 14154 17332
rect 14185 17323 14243 17329
rect 14185 17289 14197 17323
rect 14231 17320 14243 17323
rect 15010 17320 15016 17332
rect 14231 17292 15016 17320
rect 14231 17289 14243 17292
rect 14185 17283 14243 17289
rect 15010 17280 15016 17292
rect 15068 17280 15074 17332
rect 16117 17323 16175 17329
rect 16117 17289 16129 17323
rect 16163 17320 16175 17323
rect 18046 17320 18052 17332
rect 16163 17292 18052 17320
rect 16163 17289 16175 17292
rect 16117 17283 16175 17289
rect 18046 17280 18052 17292
rect 18104 17280 18110 17332
rect 18598 17280 18604 17332
rect 18656 17320 18662 17332
rect 20254 17320 20260 17332
rect 18656 17292 20260 17320
rect 18656 17280 18662 17292
rect 20254 17280 20260 17292
rect 20312 17280 20318 17332
rect 20364 17292 21864 17320
rect 13538 17252 13544 17264
rect 13004 17224 13544 17252
rect 11568 17187 11626 17193
rect 11568 17184 11580 17187
rect 11262 17156 11580 17184
rect 9401 17147 9459 17153
rect 11568 17153 11580 17156
rect 11614 17153 11626 17187
rect 11568 17147 11626 17153
rect 11747 17187 11805 17193
rect 11747 17153 11759 17187
rect 11793 17184 11805 17187
rect 12802 17184 12808 17196
rect 11793 17156 12808 17184
rect 11793 17153 11805 17156
rect 11747 17147 11805 17153
rect 12802 17144 12808 17156
rect 12860 17144 12866 17196
rect 9030 17076 9036 17128
rect 9088 17116 9094 17128
rect 9306 17116 9312 17128
rect 9088 17088 9312 17116
rect 9088 17076 9094 17088
rect 9306 17076 9312 17088
rect 9364 17076 9370 17128
rect 9490 17076 9496 17128
rect 9548 17116 9554 17128
rect 10502 17116 10508 17128
rect 9548 17088 10508 17116
rect 9548 17076 9554 17088
rect 10502 17076 10508 17088
rect 10560 17076 10566 17128
rect 10870 17076 10876 17128
rect 10928 17076 10934 17128
rect 11238 17076 11244 17128
rect 11296 17076 11302 17128
rect 11977 17119 12035 17125
rect 11977 17116 11989 17119
rect 11348 17088 11989 17116
rect 10962 17008 10968 17060
rect 11020 17048 11026 17060
rect 11348 17048 11376 17088
rect 11977 17085 11989 17088
rect 12023 17085 12035 17119
rect 11977 17079 12035 17085
rect 12250 17076 12256 17128
rect 12308 17116 12314 17128
rect 13004 17116 13032 17224
rect 13538 17212 13544 17224
rect 13596 17252 13602 17264
rect 13596 17224 13768 17252
rect 13596 17212 13602 17224
rect 13078 17144 13084 17196
rect 13136 17144 13142 17196
rect 12308 17088 13032 17116
rect 12308 17076 12314 17088
rect 11020 17020 11376 17048
rect 13096 17048 13124 17144
rect 13740 17125 13768 17224
rect 16206 17212 16212 17264
rect 16264 17212 16270 17264
rect 20364 17252 20392 17292
rect 20272 17224 20392 17252
rect 21836 17252 21864 17292
rect 22370 17280 22376 17332
rect 22428 17280 22434 17332
rect 23198 17280 23204 17332
rect 23256 17320 23262 17332
rect 23256 17292 25728 17320
rect 23256 17280 23262 17292
rect 22002 17252 22008 17264
rect 21836 17224 22008 17252
rect 15562 17184 15568 17196
rect 13924 17156 15568 17184
rect 13924 17125 13952 17156
rect 15562 17144 15568 17156
rect 15620 17144 15626 17196
rect 13725 17119 13783 17125
rect 13725 17085 13737 17119
rect 13771 17085 13783 17119
rect 13725 17079 13783 17085
rect 13909 17119 13967 17125
rect 13909 17085 13921 17119
rect 13955 17085 13967 17119
rect 13909 17079 13967 17085
rect 14001 17119 14059 17125
rect 14001 17085 14013 17119
rect 14047 17116 14059 17119
rect 14553 17119 14611 17125
rect 14047 17088 14504 17116
rect 14047 17085 14059 17088
rect 14001 17079 14059 17085
rect 13924 17048 13952 17079
rect 13096 17020 13952 17048
rect 11020 17008 11026 17020
rect 8404 16952 8800 16980
rect 9131 16983 9189 16989
rect 9131 16949 9143 16983
rect 9177 16980 9189 16983
rect 9674 16980 9680 16992
rect 9177 16952 9680 16980
rect 9177 16949 9189 16952
rect 9131 16943 9189 16949
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 11330 16980 11336 16992
rect 10192 16952 11336 16980
rect 10192 16940 10198 16952
rect 11330 16940 11336 16952
rect 11388 16940 11394 16992
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 13081 16983 13139 16989
rect 13081 16980 13093 16983
rect 11940 16952 13093 16980
rect 11940 16940 11946 16952
rect 13081 16949 13093 16952
rect 13127 16949 13139 16983
rect 13081 16943 13139 16949
rect 13630 16940 13636 16992
rect 13688 16980 13694 16992
rect 14016 16980 14044 17079
rect 13688 16952 14044 16980
rect 14476 16980 14504 17088
rect 14553 17085 14565 17119
rect 14599 17116 14611 17119
rect 14829 17119 14887 17125
rect 14599 17088 14688 17116
rect 14599 17085 14611 17088
rect 14553 17079 14611 17085
rect 14660 17060 14688 17088
rect 14829 17085 14841 17119
rect 14875 17116 14887 17119
rect 14918 17116 14924 17128
rect 14875 17088 14924 17116
rect 14875 17085 14887 17088
rect 14829 17079 14887 17085
rect 14918 17076 14924 17088
rect 14976 17076 14982 17128
rect 14642 17008 14648 17060
rect 14700 17008 14706 17060
rect 16224 16980 16252 17212
rect 16899 17187 16957 17193
rect 16899 17153 16911 17187
rect 16945 17153 16957 17187
rect 16899 17147 16957 17153
rect 16393 17119 16451 17125
rect 16393 17085 16405 17119
rect 16439 17116 16451 17119
rect 16666 17116 16672 17128
rect 16439 17088 16672 17116
rect 16439 17085 16451 17088
rect 16393 17079 16451 17085
rect 16666 17076 16672 17088
rect 16724 17076 16730 17128
rect 16914 17116 16942 17147
rect 17126 17144 17132 17196
rect 17184 17144 17190 17196
rect 19978 17184 19984 17196
rect 18156 17156 19984 17184
rect 18156 17116 18184 17156
rect 19978 17144 19984 17156
rect 20036 17144 20042 17196
rect 16914 17088 18184 17116
rect 18690 17076 18696 17128
rect 18748 17076 18754 17128
rect 18969 17119 19027 17125
rect 18969 17085 18981 17119
rect 19015 17116 19027 17119
rect 20272 17116 20300 17224
rect 22002 17212 22008 17224
rect 22060 17212 22066 17264
rect 22388 17252 22416 17280
rect 25700 17252 25728 17292
rect 25774 17280 25780 17332
rect 25832 17280 25838 17332
rect 25958 17280 25964 17332
rect 26016 17320 26022 17332
rect 27985 17323 28043 17329
rect 27985 17320 27997 17323
rect 26016 17292 27997 17320
rect 26016 17280 26022 17292
rect 27985 17289 27997 17292
rect 28031 17289 28043 17323
rect 27985 17283 28043 17289
rect 28442 17280 28448 17332
rect 28500 17320 28506 17332
rect 28718 17320 28724 17332
rect 28500 17292 28724 17320
rect 28500 17280 28506 17292
rect 28718 17280 28724 17292
rect 28776 17280 28782 17332
rect 29822 17280 29828 17332
rect 29880 17320 29886 17332
rect 29917 17323 29975 17329
rect 29917 17320 29929 17323
rect 29880 17292 29929 17320
rect 29880 17280 29886 17292
rect 29917 17289 29929 17292
rect 29963 17289 29975 17323
rect 29917 17283 29975 17289
rect 25866 17252 25872 17264
rect 22388 17224 23428 17252
rect 25700 17224 25872 17252
rect 20947 17187 21005 17193
rect 20947 17153 20959 17187
rect 20993 17184 21005 17187
rect 21082 17184 21088 17196
rect 20993 17156 21088 17184
rect 20993 17153 21005 17156
rect 20947 17147 21005 17153
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 21174 17144 21180 17196
rect 21232 17144 21238 17196
rect 22833 17187 22891 17193
rect 22833 17184 22845 17187
rect 21468 17156 22845 17184
rect 21468 17128 21496 17156
rect 22833 17153 22845 17156
rect 22879 17153 22891 17187
rect 22833 17147 22891 17153
rect 19015 17088 20300 17116
rect 20441 17119 20499 17125
rect 19015 17085 19027 17088
rect 18969 17079 19027 17085
rect 20441 17085 20453 17119
rect 20487 17116 20499 17119
rect 20530 17116 20536 17128
rect 20487 17088 20536 17116
rect 20487 17085 20499 17088
rect 20441 17079 20499 17085
rect 20530 17076 20536 17088
rect 20588 17076 20594 17128
rect 20806 17125 20812 17128
rect 20768 17119 20812 17125
rect 20768 17085 20780 17119
rect 20864 17116 20870 17128
rect 21450 17116 21456 17128
rect 20864 17088 21456 17116
rect 20768 17079 20812 17085
rect 20806 17076 20812 17079
rect 20864 17076 20870 17088
rect 21450 17076 21456 17088
rect 21508 17076 21514 17128
rect 22554 17076 22560 17128
rect 22612 17116 22618 17128
rect 22649 17119 22707 17125
rect 22649 17116 22661 17119
rect 22612 17088 22661 17116
rect 22612 17076 22618 17088
rect 22649 17085 22661 17088
rect 22695 17116 22707 17119
rect 23198 17116 23204 17128
rect 22695 17088 23204 17116
rect 22695 17085 22707 17088
rect 22649 17079 22707 17085
rect 23198 17076 23204 17088
rect 23256 17076 23262 17128
rect 23400 17116 23428 17224
rect 25866 17212 25872 17224
rect 25924 17212 25930 17264
rect 27706 17212 27712 17264
rect 27764 17252 27770 17264
rect 30285 17255 30343 17261
rect 30285 17252 30297 17255
rect 27764 17224 30297 17252
rect 27764 17212 27770 17224
rect 30285 17221 30297 17224
rect 30331 17221 30343 17255
rect 30285 17215 30343 17221
rect 30377 17255 30435 17261
rect 30377 17221 30389 17255
rect 30423 17221 30435 17255
rect 30377 17215 30435 17221
rect 23937 17187 23995 17193
rect 23937 17153 23949 17187
rect 23983 17184 23995 17187
rect 24210 17184 24216 17196
rect 23983 17156 24216 17184
rect 23983 17153 23995 17156
rect 23937 17147 23995 17153
rect 24210 17144 24216 17156
rect 24268 17144 24274 17196
rect 24443 17187 24501 17193
rect 24443 17153 24455 17187
rect 24489 17184 24501 17187
rect 26326 17184 26332 17196
rect 24489 17156 26332 17184
rect 24489 17153 24501 17156
rect 24443 17147 24501 17153
rect 26326 17144 26332 17156
rect 26384 17144 26390 17196
rect 26608 17187 26666 17193
rect 26608 17184 26620 17187
rect 26528 17156 26620 17184
rect 26528 17128 26556 17156
rect 26608 17153 26620 17156
rect 26654 17153 26666 17187
rect 26608 17147 26666 17153
rect 26881 17187 26939 17193
rect 26881 17153 26893 17187
rect 26927 17184 26939 17187
rect 30392 17184 30420 17215
rect 26927 17156 30420 17184
rect 26927 17153 26939 17156
rect 26881 17147 26939 17153
rect 24673 17119 24731 17125
rect 24673 17116 24685 17119
rect 23400 17088 24685 17116
rect 24673 17085 24685 17088
rect 24719 17085 24731 17119
rect 24673 17079 24731 17085
rect 26142 17076 26148 17128
rect 26200 17076 26206 17128
rect 26510 17076 26516 17128
rect 26568 17076 26574 17128
rect 28074 17076 28080 17128
rect 28132 17116 28138 17128
rect 28445 17119 28503 17125
rect 28445 17116 28457 17119
rect 28132 17088 28457 17116
rect 28132 17076 28138 17088
rect 28445 17085 28457 17088
rect 28491 17085 28503 17119
rect 28445 17079 28503 17085
rect 29089 17119 29147 17125
rect 29089 17085 29101 17119
rect 29135 17116 29147 17119
rect 29270 17116 29276 17128
rect 29135 17088 29276 17116
rect 29135 17085 29147 17088
rect 29089 17079 29147 17085
rect 29270 17076 29276 17088
rect 29328 17076 29334 17128
rect 29638 17076 29644 17128
rect 29696 17076 29702 17128
rect 29825 17119 29883 17125
rect 29825 17085 29837 17119
rect 29871 17116 29883 17119
rect 30006 17116 30012 17128
rect 29871 17088 30012 17116
rect 29871 17085 29883 17088
rect 29825 17079 29883 17085
rect 23477 17051 23535 17057
rect 19996 17020 20208 17048
rect 14476 16952 16252 16980
rect 13688 16940 13694 16952
rect 16850 16940 16856 16992
rect 16908 16989 16914 16992
rect 16908 16943 16917 16989
rect 16908 16940 16914 16943
rect 17034 16940 17040 16992
rect 17092 16980 17098 16992
rect 18233 16983 18291 16989
rect 18233 16980 18245 16983
rect 17092 16952 18245 16980
rect 17092 16940 17098 16952
rect 18233 16949 18245 16952
rect 18279 16949 18291 16983
rect 18233 16943 18291 16949
rect 18414 16940 18420 16992
rect 18472 16980 18478 16992
rect 19996 16980 20024 17020
rect 18472 16952 20024 16980
rect 18472 16940 18478 16952
rect 20070 16940 20076 16992
rect 20128 16940 20134 16992
rect 20180 16980 20208 17020
rect 23477 17017 23489 17051
rect 23523 17017 23535 17051
rect 23477 17011 23535 17017
rect 22281 16983 22339 16989
rect 22281 16980 22293 16983
rect 20180 16952 22293 16980
rect 22281 16949 22293 16952
rect 22327 16949 22339 16983
rect 23492 16980 23520 17011
rect 24394 16980 24400 16992
rect 24452 16989 24458 16992
rect 23492 16952 24400 16980
rect 22281 16943 22339 16949
rect 24394 16940 24400 16952
rect 24452 16980 24461 16989
rect 24452 16952 24497 16980
rect 24452 16943 24461 16952
rect 24452 16940 24458 16943
rect 26418 16940 26424 16992
rect 26476 16980 26482 16992
rect 26611 16983 26669 16989
rect 26611 16980 26623 16983
rect 26476 16952 26623 16980
rect 26476 16940 26482 16952
rect 26611 16949 26623 16952
rect 26657 16980 26669 16983
rect 26786 16980 26792 16992
rect 26657 16952 26792 16980
rect 26657 16949 26669 16952
rect 26611 16943 26669 16949
rect 26786 16940 26792 16952
rect 26844 16940 26850 16992
rect 28534 16940 28540 16992
rect 28592 16980 28598 16992
rect 29454 16980 29460 16992
rect 28592 16952 29460 16980
rect 28592 16940 28598 16952
rect 29454 16940 29460 16952
rect 29512 16980 29518 16992
rect 29840 16980 29868 17079
rect 30006 17076 30012 17088
rect 30064 17076 30070 17128
rect 30561 17119 30619 17125
rect 30561 17085 30573 17119
rect 30607 17116 30619 17119
rect 31110 17116 31116 17128
rect 30607 17088 31116 17116
rect 30607 17085 30619 17088
rect 30561 17079 30619 17085
rect 31110 17076 31116 17088
rect 31168 17076 31174 17128
rect 30101 17051 30159 17057
rect 30101 17017 30113 17051
rect 30147 17017 30159 17051
rect 30101 17011 30159 17017
rect 29512 16952 29868 16980
rect 29512 16940 29518 16952
rect 30006 16940 30012 16992
rect 30064 16980 30070 16992
rect 30116 16980 30144 17011
rect 30064 16952 30144 16980
rect 30064 16940 30070 16952
rect 31018 16940 31024 16992
rect 31076 16980 31082 16992
rect 31076 16952 31156 16980
rect 31076 16940 31082 16952
rect 552 16890 31072 16912
rect 552 16838 7988 16890
rect 8040 16838 8052 16890
rect 8104 16838 8116 16890
rect 8168 16838 8180 16890
rect 8232 16838 8244 16890
rect 8296 16838 15578 16890
rect 15630 16838 15642 16890
rect 15694 16838 15706 16890
rect 15758 16838 15770 16890
rect 15822 16838 15834 16890
rect 15886 16838 23168 16890
rect 23220 16838 23232 16890
rect 23284 16838 23296 16890
rect 23348 16838 23360 16890
rect 23412 16838 23424 16890
rect 23476 16838 30758 16890
rect 30810 16838 30822 16890
rect 30874 16838 30886 16890
rect 30938 16838 30950 16890
rect 31002 16838 31014 16890
rect 31066 16838 31072 16890
rect 552 16816 31072 16838
rect 1210 16736 1216 16788
rect 1268 16776 1274 16788
rect 2314 16776 2320 16788
rect 1268 16748 2320 16776
rect 1268 16736 1274 16748
rect 2314 16736 2320 16748
rect 2372 16736 2378 16788
rect 3050 16736 3056 16788
rect 3108 16736 3114 16788
rect 3326 16736 3332 16788
rect 3384 16776 3390 16788
rect 3384 16748 4936 16776
rect 3384 16736 3390 16748
rect 1121 16643 1179 16649
rect 1121 16609 1133 16643
rect 1167 16640 1179 16643
rect 3602 16640 3608 16652
rect 1167 16612 3608 16640
rect 1167 16609 1179 16612
rect 1121 16603 1179 16609
rect 3602 16600 3608 16612
rect 3660 16600 3666 16652
rect 4249 16643 4307 16649
rect 4249 16609 4261 16643
rect 4295 16640 4307 16643
rect 4522 16640 4528 16652
rect 4295 16612 4528 16640
rect 4295 16609 4307 16612
rect 4249 16603 4307 16609
rect 4522 16600 4528 16612
rect 4580 16600 4586 16652
rect 4908 16640 4936 16748
rect 5534 16736 5540 16788
rect 5592 16736 5598 16788
rect 6279 16779 6337 16785
rect 6279 16776 6291 16779
rect 5644 16748 6291 16776
rect 5074 16668 5080 16720
rect 5132 16708 5138 16720
rect 5644 16708 5672 16748
rect 6279 16745 6291 16748
rect 6325 16745 6337 16779
rect 6279 16739 6337 16745
rect 7006 16736 7012 16788
rect 7064 16776 7070 16788
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 7064 16748 7665 16776
rect 7064 16736 7070 16748
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 7653 16739 7711 16745
rect 8481 16779 8539 16785
rect 8481 16745 8493 16779
rect 8527 16776 8539 16779
rect 8662 16776 8668 16788
rect 8527 16748 8668 16776
rect 8527 16745 8539 16748
rect 8481 16739 8539 16745
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 8938 16736 8944 16788
rect 8996 16776 9002 16788
rect 9131 16779 9189 16785
rect 9131 16776 9143 16779
rect 8996 16748 9143 16776
rect 8996 16736 9002 16748
rect 9131 16745 9143 16748
rect 9177 16745 9189 16779
rect 9131 16739 9189 16745
rect 10502 16736 10508 16788
rect 10560 16736 10566 16788
rect 11882 16776 11888 16788
rect 11164 16748 11888 16776
rect 5132 16680 5672 16708
rect 5132 16668 5138 16680
rect 7282 16668 7288 16720
rect 7340 16708 7346 16720
rect 8205 16711 8263 16717
rect 8205 16708 8217 16711
rect 7340 16680 8217 16708
rect 7340 16668 7346 16680
rect 8205 16677 8217 16680
rect 8251 16677 8263 16711
rect 11164 16708 11192 16748
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12802 16736 12808 16788
rect 12860 16776 12866 16788
rect 15657 16779 15715 16785
rect 15657 16776 15669 16779
rect 12860 16748 15669 16776
rect 12860 16736 12866 16748
rect 15657 16745 15669 16748
rect 15703 16745 15715 16779
rect 15657 16739 15715 16745
rect 16114 16736 16120 16788
rect 16172 16736 16178 16788
rect 17034 16736 17040 16788
rect 17092 16736 17098 16788
rect 17954 16736 17960 16788
rect 18012 16776 18018 16788
rect 18785 16779 18843 16785
rect 18785 16776 18797 16779
rect 18012 16748 18797 16776
rect 18012 16736 18018 16748
rect 18785 16745 18797 16748
rect 18831 16745 18843 16779
rect 18785 16739 18843 16745
rect 19150 16736 19156 16788
rect 19208 16736 19214 16788
rect 21174 16776 21180 16788
rect 19444 16748 21180 16776
rect 8205 16671 8263 16677
rect 10888 16680 11192 16708
rect 5813 16643 5871 16649
rect 5813 16640 5825 16643
rect 4908 16612 5825 16640
rect 5813 16609 5825 16612
rect 5859 16609 5871 16643
rect 5813 16603 5871 16609
rect 5902 16600 5908 16652
rect 5960 16640 5966 16652
rect 5960 16612 6040 16640
rect 5960 16600 5966 16612
rect 1026 16532 1032 16584
rect 1084 16572 1090 16584
rect 1578 16581 1584 16584
rect 1213 16575 1271 16581
rect 1213 16572 1225 16575
rect 1084 16544 1225 16572
rect 1084 16532 1090 16544
rect 1213 16541 1225 16544
rect 1259 16541 1271 16575
rect 1213 16535 1271 16541
rect 1540 16575 1584 16581
rect 1540 16541 1552 16575
rect 1540 16535 1584 16541
rect 1578 16532 1584 16535
rect 1636 16532 1642 16584
rect 1762 16583 1768 16584
rect 1719 16577 1768 16583
rect 1719 16543 1731 16577
rect 1765 16543 1768 16577
rect 1719 16537 1768 16543
rect 1762 16532 1768 16537
rect 1820 16532 1826 16584
rect 1949 16575 2007 16581
rect 1949 16541 1961 16575
rect 1995 16572 2007 16575
rect 3513 16575 3571 16581
rect 1995 16544 3464 16572
rect 1995 16541 2007 16544
rect 1949 16535 2007 16541
rect 934 16396 940 16448
rect 992 16396 998 16448
rect 3436 16436 3464 16544
rect 3513 16541 3525 16575
rect 3559 16572 3571 16575
rect 3694 16572 3700 16584
rect 3559 16544 3700 16572
rect 3559 16541 3571 16544
rect 3513 16535 3571 16541
rect 3694 16532 3700 16544
rect 3752 16532 3758 16584
rect 3878 16581 3884 16584
rect 3840 16575 3884 16581
rect 3840 16541 3852 16575
rect 3840 16535 3884 16541
rect 3878 16532 3884 16535
rect 3936 16532 3942 16584
rect 4062 16583 4068 16584
rect 4019 16577 4068 16583
rect 4019 16543 4031 16577
rect 4065 16543 4068 16577
rect 4019 16537 4068 16543
rect 4062 16532 4068 16537
rect 4120 16532 4126 16584
rect 6012 16572 6040 16612
rect 6546 16600 6552 16652
rect 6604 16600 6610 16652
rect 9398 16600 9404 16652
rect 9456 16600 9462 16652
rect 10888 16640 10916 16680
rect 13906 16668 13912 16720
rect 13964 16668 13970 16720
rect 17052 16708 17080 16736
rect 15396 16680 17080 16708
rect 9508 16612 10916 16640
rect 9161 16593 9219 16599
rect 6276 16575 6334 16581
rect 6276 16572 6288 16575
rect 6012 16544 6288 16572
rect 6276 16541 6288 16544
rect 6322 16541 6334 16575
rect 6276 16535 6334 16541
rect 8662 16532 8668 16584
rect 8720 16532 8726 16584
rect 9161 16559 9173 16593
rect 9207 16572 9219 16593
rect 9508 16572 9536 16612
rect 11054 16600 11060 16652
rect 11112 16600 11118 16652
rect 12345 16643 12403 16649
rect 12345 16640 12357 16643
rect 11164 16612 12357 16640
rect 9207 16559 9536 16572
rect 9161 16553 9536 16559
rect 9186 16544 9536 16553
rect 10318 16532 10324 16584
rect 10376 16572 10382 16584
rect 11164 16572 11192 16612
rect 12345 16609 12357 16612
rect 12391 16609 12403 16643
rect 13924 16640 13952 16668
rect 14182 16649 14188 16652
rect 12345 16603 12403 16609
rect 13740 16612 13952 16640
rect 14144 16643 14188 16649
rect 10376 16544 11192 16572
rect 10376 16532 10382 16544
rect 11238 16532 11244 16584
rect 11296 16572 11302 16584
rect 11609 16575 11667 16581
rect 11609 16572 11621 16575
rect 11296 16544 11621 16572
rect 11296 16532 11302 16544
rect 11609 16541 11621 16544
rect 11655 16541 11667 16575
rect 11609 16535 11667 16541
rect 11790 16532 11796 16584
rect 11848 16572 11854 16584
rect 11974 16581 11980 16584
rect 11936 16575 11980 16581
rect 11936 16572 11948 16575
rect 11848 16544 11948 16572
rect 11848 16532 11854 16544
rect 11936 16541 11948 16544
rect 11936 16535 11980 16541
rect 11974 16532 11980 16535
rect 12032 16532 12038 16584
rect 12115 16575 12173 16581
rect 12115 16541 12127 16575
rect 12161 16572 12173 16575
rect 13740 16572 13768 16612
rect 14144 16609 14156 16643
rect 14144 16603 14188 16609
rect 14182 16600 14188 16603
rect 14240 16600 14246 16652
rect 14384 16640 14596 16644
rect 15396 16640 15424 16680
rect 14328 16616 15424 16640
rect 14328 16612 14412 16616
rect 14568 16612 15424 16616
rect 12161 16544 13768 16572
rect 12161 16541 12173 16544
rect 12115 16535 12173 16541
rect 13814 16532 13820 16584
rect 13872 16532 13878 16584
rect 14328 16583 14356 16612
rect 15470 16600 15476 16652
rect 15528 16600 15534 16652
rect 16206 16600 16212 16652
rect 16264 16640 16270 16652
rect 16301 16643 16359 16649
rect 16301 16640 16313 16643
rect 16264 16612 16313 16640
rect 16264 16600 16270 16612
rect 16301 16609 16313 16612
rect 16347 16609 16359 16643
rect 16853 16643 16911 16649
rect 16853 16640 16865 16643
rect 16301 16603 16359 16609
rect 16408 16612 16865 16640
rect 14323 16577 14381 16583
rect 14323 16543 14335 16577
rect 14369 16543 14381 16577
rect 14323 16537 14381 16543
rect 14458 16534 14464 16586
rect 14516 16574 14522 16586
rect 14553 16575 14611 16581
rect 14553 16574 14565 16575
rect 14516 16546 14565 16574
rect 14516 16534 14522 16546
rect 14553 16541 14565 16546
rect 14599 16541 14611 16575
rect 15488 16572 15516 16600
rect 16408 16572 16436 16612
rect 16853 16609 16865 16612
rect 16899 16609 16911 16643
rect 16853 16603 16911 16609
rect 17034 16600 17040 16652
rect 17092 16640 17098 16652
rect 17272 16643 17330 16649
rect 17272 16640 17284 16643
rect 17092 16612 17284 16640
rect 17092 16600 17098 16612
rect 17272 16609 17284 16612
rect 17318 16609 17330 16643
rect 17272 16603 17330 16609
rect 17681 16643 17739 16649
rect 17681 16609 17693 16643
rect 17727 16640 17739 16643
rect 19168 16640 19196 16736
rect 19444 16649 19472 16748
rect 21174 16736 21180 16748
rect 21232 16736 21238 16788
rect 21284 16748 23612 16776
rect 17727 16612 19196 16640
rect 19337 16643 19395 16649
rect 17727 16609 17739 16612
rect 17681 16603 17739 16609
rect 19337 16609 19349 16643
rect 19383 16609 19395 16643
rect 19337 16603 19395 16609
rect 19429 16643 19487 16649
rect 19429 16609 19441 16643
rect 19475 16609 19487 16643
rect 19429 16603 19487 16609
rect 19705 16643 19763 16649
rect 19705 16609 19717 16643
rect 19751 16640 19763 16643
rect 20070 16640 20076 16652
rect 19751 16612 20076 16640
rect 19751 16609 19763 16612
rect 19705 16603 19763 16609
rect 17441 16593 17499 16599
rect 15488 16544 16436 16572
rect 14553 16535 14611 16541
rect 16666 16532 16672 16584
rect 16724 16572 16730 16584
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 16724 16544 16957 16572
rect 16724 16532 16730 16544
rect 16945 16541 16957 16544
rect 16991 16572 17003 16575
rect 17126 16572 17132 16584
rect 16991 16544 17132 16572
rect 16991 16541 17003 16544
rect 16945 16535 17003 16541
rect 17126 16532 17132 16544
rect 17184 16532 17190 16584
rect 17441 16559 17453 16593
rect 17487 16572 17499 16593
rect 18414 16572 18420 16584
rect 17487 16559 18420 16572
rect 17441 16553 18420 16559
rect 17456 16544 18420 16553
rect 18414 16532 18420 16544
rect 18472 16532 18478 16584
rect 19352 16572 19380 16603
rect 20070 16600 20076 16612
rect 20128 16600 20134 16652
rect 21082 16600 21088 16652
rect 21140 16600 21146 16652
rect 21284 16584 21312 16748
rect 23584 16717 23612 16748
rect 23842 16736 23848 16788
rect 23900 16776 23906 16788
rect 24210 16776 24216 16788
rect 23900 16748 24216 16776
rect 23900 16736 23906 16748
rect 23569 16711 23627 16717
rect 23569 16677 23581 16711
rect 23615 16677 23627 16711
rect 23569 16671 23627 16677
rect 21358 16600 21364 16652
rect 21416 16640 21422 16652
rect 22005 16643 22063 16649
rect 22005 16640 22017 16643
rect 21416 16612 22017 16640
rect 21416 16600 21422 16612
rect 22005 16609 22017 16612
rect 22051 16609 22063 16643
rect 22005 16603 22063 16609
rect 22370 16600 22376 16652
rect 22428 16640 22434 16652
rect 23934 16640 23940 16652
rect 22428 16612 23940 16640
rect 22428 16600 22434 16612
rect 23934 16600 23940 16612
rect 23992 16600 23998 16652
rect 24136 16649 24164 16748
rect 24210 16736 24216 16748
rect 24268 16736 24274 16788
rect 24394 16736 24400 16788
rect 24452 16776 24458 16788
rect 24587 16779 24645 16785
rect 24587 16776 24599 16779
rect 24452 16748 24599 16776
rect 24452 16736 24458 16748
rect 24587 16745 24599 16748
rect 24633 16745 24645 16779
rect 27890 16776 27896 16788
rect 24587 16739 24645 16745
rect 25976 16748 27896 16776
rect 24121 16643 24179 16649
rect 24121 16609 24133 16643
rect 24167 16609 24179 16643
rect 24121 16603 24179 16609
rect 24857 16643 24915 16649
rect 24857 16609 24869 16643
rect 24903 16640 24915 16643
rect 25976 16640 26004 16748
rect 27890 16736 27896 16748
rect 27948 16736 27954 16788
rect 28350 16736 28356 16788
rect 28408 16776 28414 16788
rect 29914 16776 29920 16788
rect 28408 16748 29920 16776
rect 28408 16736 28414 16748
rect 29914 16736 29920 16748
rect 29972 16736 29978 16788
rect 30374 16736 30380 16788
rect 30432 16736 30438 16788
rect 31018 16736 31024 16788
rect 31076 16776 31082 16788
rect 31128 16776 31156 16952
rect 31076 16748 31156 16776
rect 31076 16736 31082 16748
rect 27982 16668 27988 16720
rect 28040 16708 28046 16720
rect 28040 16680 28764 16708
rect 28040 16668 28046 16680
rect 24903 16612 26004 16640
rect 24903 16609 24915 16612
rect 24857 16603 24915 16609
rect 26050 16600 26056 16652
rect 26108 16640 26114 16652
rect 27157 16643 27215 16649
rect 27157 16640 27169 16643
rect 26108 16612 27169 16640
rect 26108 16600 26114 16612
rect 27157 16609 27169 16612
rect 27203 16609 27215 16643
rect 27157 16603 27215 16609
rect 27246 16600 27252 16652
rect 27304 16600 27310 16652
rect 27614 16600 27620 16652
rect 27672 16640 27678 16652
rect 28629 16643 28687 16649
rect 28629 16640 28641 16643
rect 27672 16612 28641 16640
rect 27672 16600 27678 16612
rect 28629 16609 28641 16612
rect 28675 16609 28687 16643
rect 28736 16640 28764 16680
rect 28905 16643 28963 16649
rect 28905 16640 28917 16643
rect 28736 16612 28917 16640
rect 28629 16603 28687 16609
rect 28905 16609 28917 16612
rect 28951 16609 28963 16643
rect 30561 16643 30619 16649
rect 30561 16640 30573 16643
rect 28905 16603 28963 16609
rect 29104 16612 30573 16640
rect 24584 16593 24642 16599
rect 19352 16544 20392 16572
rect 10778 16464 10784 16516
rect 10836 16504 10842 16516
rect 10836 16476 11284 16504
rect 10836 16464 10842 16476
rect 5258 16436 5264 16448
rect 3436 16408 5264 16436
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 5534 16396 5540 16448
rect 5592 16436 5598 16448
rect 10134 16436 10140 16448
rect 5592 16408 10140 16436
rect 5592 16396 5598 16408
rect 10134 16396 10140 16408
rect 10192 16396 10198 16448
rect 11256 16436 11284 16476
rect 11330 16464 11336 16516
rect 11388 16464 11394 16516
rect 15470 16504 15476 16516
rect 15212 16476 15476 16504
rect 12710 16436 12716 16448
rect 11256 16408 12716 16436
rect 12710 16396 12716 16408
rect 12768 16396 12774 16448
rect 13446 16396 13452 16448
rect 13504 16396 13510 16448
rect 14274 16396 14280 16448
rect 14332 16436 14338 16448
rect 15212 16436 15240 16476
rect 15470 16464 15476 16476
rect 15528 16504 15534 16516
rect 19426 16504 19432 16516
rect 15528 16476 16804 16504
rect 15528 16464 15534 16476
rect 14332 16408 15240 16436
rect 14332 16396 14338 16408
rect 15930 16396 15936 16448
rect 15988 16436 15994 16448
rect 16669 16439 16727 16445
rect 16669 16436 16681 16439
rect 15988 16408 16681 16436
rect 15988 16396 15994 16408
rect 16669 16405 16681 16408
rect 16715 16405 16727 16439
rect 16776 16436 16804 16476
rect 19306 16476 19432 16504
rect 19306 16448 19334 16476
rect 19426 16464 19432 16476
rect 19484 16464 19490 16516
rect 20364 16504 20392 16544
rect 20530 16532 20536 16584
rect 20588 16572 20594 16584
rect 20898 16572 20904 16584
rect 20588 16544 20904 16572
rect 20588 16532 20594 16544
rect 20898 16532 20904 16544
rect 20956 16572 20962 16584
rect 21266 16572 21272 16584
rect 20956 16544 21272 16572
rect 20956 16532 20962 16544
rect 21266 16532 21272 16544
rect 21324 16532 21330 16584
rect 21450 16532 21456 16584
rect 21508 16572 21514 16584
rect 21596 16575 21654 16581
rect 21596 16572 21608 16575
rect 21508 16544 21608 16572
rect 21508 16532 21514 16544
rect 21596 16541 21608 16544
rect 21642 16541 21654 16575
rect 21596 16535 21654 16541
rect 21775 16575 21833 16581
rect 21775 16541 21787 16575
rect 21821 16572 21833 16575
rect 21821 16544 24072 16572
rect 24584 16559 24596 16593
rect 24630 16572 24642 16593
rect 25038 16572 25044 16584
rect 24630 16559 25044 16572
rect 24584 16553 25044 16559
rect 24596 16544 25044 16553
rect 21821 16541 21833 16544
rect 21775 16535 21833 16541
rect 20364 16476 21128 16504
rect 21100 16448 21128 16476
rect 22738 16464 22744 16516
rect 22796 16504 22802 16516
rect 23109 16507 23167 16513
rect 23109 16504 23121 16507
rect 22796 16476 23121 16504
rect 22796 16464 22802 16476
rect 23109 16473 23121 16476
rect 23155 16473 23167 16507
rect 23109 16467 23167 16473
rect 18414 16436 18420 16448
rect 16776 16408 18420 16436
rect 16669 16399 16727 16405
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 19150 16396 19156 16448
rect 19208 16396 19214 16448
rect 19242 16396 19248 16448
rect 19300 16408 19334 16448
rect 19300 16396 19306 16408
rect 21082 16396 21088 16448
rect 21140 16396 21146 16448
rect 21174 16396 21180 16448
rect 21232 16436 21238 16448
rect 22462 16436 22468 16448
rect 21232 16408 22468 16436
rect 21232 16396 21238 16408
rect 22462 16396 22468 16408
rect 22520 16396 22526 16448
rect 24044 16436 24072 16544
rect 25038 16532 25044 16544
rect 25096 16532 25102 16584
rect 26142 16532 26148 16584
rect 26200 16572 26206 16584
rect 26786 16581 26792 16584
rect 26421 16575 26479 16581
rect 26421 16572 26433 16575
rect 26200 16544 26433 16572
rect 26200 16532 26206 16544
rect 26421 16541 26433 16544
rect 26467 16541 26479 16575
rect 26421 16535 26479 16541
rect 26748 16575 26792 16581
rect 26748 16541 26760 16575
rect 26748 16535 26792 16541
rect 26786 16532 26792 16535
rect 26844 16532 26850 16584
rect 26884 16577 26942 16583
rect 26884 16543 26896 16577
rect 26930 16572 26942 16577
rect 27264 16572 27292 16600
rect 26930 16544 27292 16572
rect 26930 16543 26942 16544
rect 26884 16537 26942 16543
rect 27890 16532 27896 16584
rect 27948 16572 27954 16584
rect 28166 16572 28172 16584
rect 27948 16544 28172 16572
rect 27948 16532 27954 16544
rect 28166 16532 28172 16544
rect 28224 16532 28230 16584
rect 28442 16532 28448 16584
rect 28500 16572 28506 16584
rect 29104 16574 29132 16612
rect 30561 16609 30573 16612
rect 30607 16609 30619 16643
rect 30561 16603 30619 16609
rect 29012 16572 29132 16574
rect 28500 16546 29132 16572
rect 28500 16544 29040 16546
rect 28500 16532 28506 16544
rect 29270 16532 29276 16584
rect 29328 16572 29334 16584
rect 29546 16572 29552 16584
rect 29328 16544 29552 16572
rect 29328 16532 29334 16544
rect 29546 16532 29552 16544
rect 29604 16532 29610 16584
rect 29638 16532 29644 16584
rect 29696 16572 29702 16584
rect 30009 16575 30067 16581
rect 30009 16572 30021 16575
rect 29696 16544 30021 16572
rect 29696 16532 29702 16544
rect 30009 16541 30021 16544
rect 30055 16541 30067 16575
rect 30009 16535 30067 16541
rect 25961 16507 26019 16513
rect 25961 16473 25973 16507
rect 26007 16473 26019 16507
rect 25961 16467 26019 16473
rect 27816 16476 28396 16504
rect 25976 16436 26004 16467
rect 24044 16408 26004 16436
rect 26786 16396 26792 16448
rect 26844 16436 26850 16448
rect 27816 16436 27844 16476
rect 26844 16408 27844 16436
rect 26844 16396 26850 16408
rect 28258 16396 28264 16448
rect 28316 16396 28322 16448
rect 28368 16436 28396 16476
rect 29362 16436 29368 16448
rect 28368 16408 29368 16436
rect 29362 16396 29368 16408
rect 29420 16396 29426 16448
rect 552 16346 30912 16368
rect 552 16294 4193 16346
rect 4245 16294 4257 16346
rect 4309 16294 4321 16346
rect 4373 16294 4385 16346
rect 4437 16294 4449 16346
rect 4501 16294 11783 16346
rect 11835 16294 11847 16346
rect 11899 16294 11911 16346
rect 11963 16294 11975 16346
rect 12027 16294 12039 16346
rect 12091 16294 19373 16346
rect 19425 16294 19437 16346
rect 19489 16294 19501 16346
rect 19553 16294 19565 16346
rect 19617 16294 19629 16346
rect 19681 16294 26963 16346
rect 27015 16294 27027 16346
rect 27079 16294 27091 16346
rect 27143 16294 27155 16346
rect 27207 16294 27219 16346
rect 27271 16294 30912 16346
rect 552 16272 30912 16294
rect 2958 16192 2964 16244
rect 3016 16192 3022 16244
rect 5534 16232 5540 16244
rect 3804 16204 5540 16232
rect 1443 16099 1501 16105
rect 1443 16065 1455 16099
rect 1489 16096 1501 16099
rect 3804 16096 3832 16204
rect 5534 16192 5540 16204
rect 5592 16192 5598 16244
rect 5626 16192 5632 16244
rect 5684 16192 5690 16244
rect 7929 16235 7987 16241
rect 7929 16232 7941 16235
rect 6104 16204 7941 16232
rect 1489 16068 3832 16096
rect 4295 16099 4353 16105
rect 1489 16065 1501 16068
rect 1443 16059 1501 16065
rect 4295 16065 4307 16099
rect 4341 16096 4353 16099
rect 6104 16096 6132 16204
rect 7929 16201 7941 16204
rect 7975 16201 7987 16235
rect 7929 16195 7987 16201
rect 8389 16235 8447 16241
rect 8389 16201 8401 16235
rect 8435 16232 8447 16235
rect 10318 16232 10324 16244
rect 8435 16204 10324 16232
rect 8435 16201 8447 16204
rect 8389 16195 8447 16201
rect 10318 16192 10324 16204
rect 10376 16192 10382 16244
rect 13446 16232 13452 16244
rect 10796 16204 13452 16232
rect 10134 16124 10140 16176
rect 10192 16164 10198 16176
rect 10505 16167 10563 16173
rect 10505 16164 10517 16167
rect 10192 16136 10517 16164
rect 10192 16124 10198 16136
rect 10505 16133 10517 16136
rect 10551 16133 10563 16167
rect 10505 16127 10563 16133
rect 8294 16096 8300 16108
rect 4341 16068 6132 16096
rect 6564 16081 8300 16096
rect 4341 16065 4353 16068
rect 4295 16059 4353 16065
rect 6564 16050 6597 16081
rect 6585 16047 6597 16050
rect 6631 16068 8300 16081
rect 6631 16047 6643 16068
rect 8294 16056 8300 16068
rect 8352 16056 8358 16108
rect 8386 16056 8392 16108
rect 8444 16096 8450 16108
rect 9171 16099 9229 16105
rect 8444 16068 8943 16096
rect 8444 16056 8450 16068
rect 6585 16041 6643 16047
rect 937 16031 995 16037
rect 937 15997 949 16031
rect 983 16028 995 16031
rect 1026 16028 1032 16040
rect 983 16000 1032 16028
rect 983 15997 995 16000
rect 937 15991 995 15997
rect 1026 15988 1032 16000
rect 1084 15988 1090 16040
rect 1673 16031 1731 16037
rect 1673 15997 1685 16031
rect 1719 16028 1731 16031
rect 1719 16000 3556 16028
rect 1719 15997 1731 16000
rect 1673 15991 1731 15997
rect 3326 15920 3332 15972
rect 3384 15920 3390 15972
rect 3528 15960 3556 16000
rect 3694 15988 3700 16040
rect 3752 16028 3758 16040
rect 3789 16031 3847 16037
rect 3789 16028 3801 16031
rect 3752 16000 3801 16028
rect 3752 15988 3758 16000
rect 3789 15997 3801 16000
rect 3835 15997 3847 16031
rect 4430 16028 4436 16040
rect 3789 15991 3847 15997
rect 3896 16000 4436 16028
rect 3896 15960 3924 16000
rect 4430 15988 4436 16000
rect 4488 15988 4494 16040
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 16028 4583 16031
rect 4890 16028 4896 16040
rect 4571 16000 4896 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 4890 15988 4896 16000
rect 4948 15988 4954 16040
rect 6089 16031 6147 16037
rect 6089 15997 6101 16031
rect 6135 16028 6147 16031
rect 6178 16028 6184 16040
rect 6135 16000 6184 16028
rect 6135 15997 6147 16000
rect 6089 15991 6147 15997
rect 6178 15988 6184 16000
rect 6236 15988 6242 16040
rect 6822 15988 6828 16040
rect 6880 15988 6886 16040
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 8478 16028 8484 16040
rect 7156 16000 8484 16028
rect 7156 15988 7162 16000
rect 8478 15988 8484 16000
rect 8536 15988 8542 16040
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 15997 8631 16031
rect 8573 15991 8631 15997
rect 3528 15932 3924 15960
rect 8588 15904 8616 15991
rect 8662 15988 8668 16040
rect 8720 15988 8726 16040
rect 8915 16028 8943 16068
rect 9171 16065 9183 16099
rect 9217 16096 9229 16099
rect 10796 16096 10824 16204
rect 13446 16192 13452 16204
rect 13504 16192 13510 16244
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 13817 16235 13875 16241
rect 13817 16232 13829 16235
rect 13780 16204 13829 16232
rect 13780 16192 13786 16204
rect 13817 16201 13829 16204
rect 13863 16201 13875 16235
rect 16393 16235 16451 16241
rect 16393 16232 16405 16235
rect 13817 16195 13875 16201
rect 14062 16204 16405 16232
rect 10965 16167 11023 16173
rect 10965 16133 10977 16167
rect 11011 16133 11023 16167
rect 10965 16127 11023 16133
rect 9217 16068 10824 16096
rect 9217 16065 9229 16068
rect 9171 16059 9229 16065
rect 9401 16031 9459 16037
rect 9401 16028 9413 16031
rect 8915 16000 9413 16028
rect 9401 15997 9413 16000
rect 9447 15997 9459 16031
rect 9401 15991 9459 15997
rect 9674 15988 9680 16040
rect 9732 16028 9738 16040
rect 10980 16028 11008 16127
rect 11238 16056 11244 16108
rect 11296 16056 11302 16108
rect 11422 16056 11428 16108
rect 11480 16056 11486 16108
rect 11747 16099 11805 16105
rect 11747 16065 11759 16099
rect 11793 16096 11805 16099
rect 14062 16096 14090 16204
rect 16393 16201 16405 16204
rect 16439 16201 16451 16235
rect 16393 16195 16451 16201
rect 16482 16192 16488 16244
rect 16540 16232 16546 16244
rect 16540 16204 18368 16232
rect 16540 16192 16546 16204
rect 14458 16124 14464 16176
rect 14516 16124 14522 16176
rect 14734 16096 14740 16108
rect 11793 16068 14090 16096
rect 14568 16068 14740 16096
rect 11793 16065 11805 16068
rect 11747 16059 11805 16065
rect 9732 16000 11008 16028
rect 11149 16031 11207 16037
rect 9732 15988 9738 16000
rect 11149 15997 11161 16031
rect 11195 16028 11207 16031
rect 11440 16028 11468 16056
rect 11195 16000 11468 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 11606 15988 11612 16040
rect 11664 16028 11670 16040
rect 14568 16037 14596 16068
rect 14734 16056 14740 16068
rect 14792 16056 14798 16108
rect 15016 16099 15074 16105
rect 15016 16096 15028 16099
rect 14844 16068 15028 16096
rect 14844 16040 14872 16068
rect 15016 16065 15028 16068
rect 15062 16065 15074 16099
rect 18233 16099 18291 16105
rect 18233 16096 18245 16099
rect 15016 16059 15074 16065
rect 15212 16068 18245 16096
rect 11977 16031 12035 16037
rect 11977 16028 11989 16031
rect 11664 16000 11989 16028
rect 11664 15988 11670 16000
rect 11977 15997 11989 16000
rect 12023 15997 12035 16031
rect 14553 16031 14611 16037
rect 14553 16028 14565 16031
rect 11977 15991 12035 15997
rect 13464 16000 14565 16028
rect 13464 15972 13492 16000
rect 14553 15997 14565 16000
rect 14599 15997 14611 16031
rect 14553 15991 14611 15997
rect 14826 15988 14832 16040
rect 14884 15988 14890 16040
rect 14918 15988 14924 16040
rect 14976 16028 14982 16040
rect 15212 16028 15240 16068
rect 18233 16065 18245 16068
rect 18279 16065 18291 16099
rect 18340 16096 18368 16204
rect 18414 16192 18420 16244
rect 18472 16232 18478 16244
rect 20530 16232 20536 16244
rect 18472 16204 20536 16232
rect 18472 16192 18478 16204
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 22094 16232 22100 16244
rect 20640 16204 22100 16232
rect 19199 16099 19257 16105
rect 18340 16068 18828 16096
rect 18233 16059 18291 16065
rect 14976 16000 15240 16028
rect 14976 15988 14982 16000
rect 15286 15988 15292 16040
rect 15344 15988 15350 16040
rect 16850 15988 16856 16040
rect 16908 15988 16914 16040
rect 17129 16031 17187 16037
rect 17129 15997 17141 16031
rect 17175 16028 17187 16031
rect 17494 16028 17500 16040
rect 17175 16000 17500 16028
rect 17175 15997 17187 16000
rect 17129 15991 17187 15997
rect 17494 15988 17500 16000
rect 17552 15988 17558 16040
rect 18693 16031 18751 16037
rect 18693 15997 18705 16031
rect 18739 15997 18751 16031
rect 18800 16028 18828 16068
rect 19199 16065 19211 16099
rect 19245 16096 19257 16099
rect 20640 16096 20668 16204
rect 22094 16192 22100 16204
rect 22152 16192 22158 16244
rect 22830 16192 22836 16244
rect 22888 16232 22894 16244
rect 25685 16235 25743 16241
rect 25685 16232 25697 16235
rect 22888 16204 25697 16232
rect 22888 16192 22894 16204
rect 25685 16201 25697 16204
rect 25731 16201 25743 16235
rect 27154 16232 27160 16244
rect 25685 16195 25743 16201
rect 26068 16204 27160 16232
rect 20714 16124 20720 16176
rect 20772 16124 20778 16176
rect 22646 16124 22652 16176
rect 22704 16164 22710 16176
rect 23201 16167 23259 16173
rect 23201 16164 23213 16167
rect 22704 16136 23213 16164
rect 22704 16124 22710 16136
rect 23201 16133 23213 16136
rect 23247 16133 23259 16167
rect 23201 16127 23259 16133
rect 25314 16124 25320 16176
rect 25372 16164 25378 16176
rect 26068 16164 26096 16204
rect 27154 16192 27160 16204
rect 27212 16192 27218 16244
rect 28350 16232 28356 16244
rect 27632 16204 28356 16232
rect 27632 16176 27660 16204
rect 28350 16192 28356 16204
rect 28408 16192 28414 16244
rect 28442 16192 28448 16244
rect 28500 16192 28506 16244
rect 28902 16192 28908 16244
rect 28960 16232 28966 16244
rect 30285 16235 30343 16241
rect 30285 16232 30297 16235
rect 28960 16204 30297 16232
rect 28960 16192 28966 16204
rect 30285 16201 30297 16204
rect 30331 16232 30343 16235
rect 30331 16204 30512 16232
rect 30331 16201 30343 16204
rect 30285 16195 30343 16201
rect 25372 16136 26096 16164
rect 25372 16124 25378 16136
rect 27614 16124 27620 16176
rect 27672 16124 27678 16176
rect 28994 16164 29000 16176
rect 28966 16124 29000 16164
rect 29052 16124 29058 16176
rect 29546 16124 29552 16176
rect 29604 16124 29610 16176
rect 29641 16167 29699 16173
rect 29641 16133 29653 16167
rect 29687 16133 29699 16167
rect 29641 16127 29699 16133
rect 21266 16105 21272 16108
rect 21228 16099 21272 16105
rect 21228 16096 21240 16099
rect 19245 16068 20668 16096
rect 20824 16068 21240 16096
rect 19245 16065 19257 16068
rect 19199 16059 19257 16065
rect 20824 16040 20852 16068
rect 21228 16065 21240 16068
rect 21228 16059 21272 16065
rect 21266 16056 21272 16059
rect 21324 16056 21330 16108
rect 21407 16099 21465 16105
rect 21407 16065 21419 16099
rect 21453 16096 21465 16099
rect 21453 16068 23704 16096
rect 21453 16065 21465 16068
rect 21407 16059 21465 16065
rect 19429 16031 19487 16037
rect 19429 16028 19441 16031
rect 18800 16000 19441 16028
rect 18693 15991 18751 15997
rect 19429 15997 19441 16000
rect 19475 15997 19487 16031
rect 19429 15991 19487 15997
rect 13446 15960 13452 15972
rect 13004 15932 13452 15960
rect 1403 15895 1461 15901
rect 1403 15861 1415 15895
rect 1449 15892 1461 15895
rect 1670 15892 1676 15904
rect 1449 15864 1676 15892
rect 1449 15861 1461 15864
rect 1403 15855 1461 15861
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 3510 15852 3516 15904
rect 3568 15892 3574 15904
rect 3605 15895 3663 15901
rect 3605 15892 3617 15895
rect 3568 15864 3617 15892
rect 3568 15852 3574 15864
rect 3605 15861 3617 15864
rect 3651 15892 3663 15895
rect 3694 15892 3700 15904
rect 3651 15864 3700 15892
rect 3651 15861 3663 15864
rect 3605 15855 3663 15861
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 3878 15852 3884 15904
rect 3936 15892 3942 15904
rect 4255 15895 4313 15901
rect 4255 15892 4267 15895
rect 3936 15864 4267 15892
rect 3936 15852 3942 15864
rect 4255 15861 4267 15864
rect 4301 15861 4313 15895
rect 4255 15855 4313 15861
rect 4430 15852 4436 15904
rect 4488 15892 4494 15904
rect 6086 15892 6092 15904
rect 4488 15864 6092 15892
rect 4488 15852 4494 15864
rect 6086 15852 6092 15864
rect 6144 15852 6150 15904
rect 6454 15852 6460 15904
rect 6512 15892 6518 15904
rect 6555 15895 6613 15901
rect 6555 15892 6567 15895
rect 6512 15864 6567 15892
rect 6512 15852 6518 15864
rect 6555 15861 6567 15864
rect 6601 15861 6613 15895
rect 6555 15855 6613 15861
rect 8570 15852 8576 15904
rect 8628 15852 8634 15904
rect 8938 15852 8944 15904
rect 8996 15892 9002 15904
rect 9131 15895 9189 15901
rect 9131 15892 9143 15895
rect 8996 15864 9143 15892
rect 8996 15852 9002 15864
rect 9131 15861 9143 15864
rect 9177 15861 9189 15895
rect 9131 15855 9189 15861
rect 11698 15852 11704 15904
rect 11756 15901 11762 15904
rect 11756 15892 11765 15901
rect 11756 15864 11801 15892
rect 11756 15855 11765 15864
rect 11756 15852 11762 15855
rect 11882 15852 11888 15904
rect 11940 15892 11946 15904
rect 13004 15892 13032 15932
rect 13446 15920 13452 15932
rect 13504 15920 13510 15972
rect 13538 15920 13544 15972
rect 13596 15960 13602 15972
rect 13725 15963 13783 15969
rect 13725 15960 13737 15963
rect 13596 15932 13737 15960
rect 13596 15920 13602 15932
rect 13725 15929 13737 15932
rect 13771 15960 13783 15963
rect 13998 15960 14004 15972
rect 13771 15932 14004 15960
rect 13771 15929 13783 15932
rect 13725 15923 13783 15929
rect 13998 15920 14004 15932
rect 14056 15920 14062 15972
rect 14274 15920 14280 15972
rect 14332 15920 14338 15972
rect 11940 15864 13032 15892
rect 11940 15852 11946 15864
rect 13078 15852 13084 15904
rect 13136 15852 13142 15904
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 15010 15892 15016 15904
rect 15068 15901 15074 15904
rect 14240 15864 15016 15892
rect 14240 15852 14246 15864
rect 15010 15852 15016 15864
rect 15068 15855 15077 15901
rect 15068 15852 15074 15855
rect 17126 15852 17132 15904
rect 17184 15892 17190 15904
rect 18708 15892 18736 15991
rect 20806 15988 20812 16040
rect 20864 15988 20870 16040
rect 20898 15988 20904 16040
rect 20956 15988 20962 16040
rect 21637 16031 21695 16037
rect 21637 16028 21649 16031
rect 21008 16000 21649 16028
rect 20162 15920 20168 15972
rect 20220 15960 20226 15972
rect 21008 15960 21036 16000
rect 21637 15997 21649 16000
rect 21683 15997 21695 16031
rect 21637 15991 21695 15997
rect 22922 15988 22928 16040
rect 22980 16028 22986 16040
rect 23109 16031 23167 16037
rect 23109 16028 23121 16031
rect 22980 16000 23121 16028
rect 22980 15988 22986 16000
rect 23109 15997 23121 16000
rect 23155 15997 23167 16031
rect 23109 15991 23167 15997
rect 20220 15932 21036 15960
rect 20220 15920 20226 15932
rect 17184 15864 18736 15892
rect 17184 15852 17190 15864
rect 19058 15852 19064 15904
rect 19116 15892 19122 15904
rect 19159 15895 19217 15901
rect 19159 15892 19171 15895
rect 19116 15864 19171 15892
rect 19116 15852 19122 15864
rect 19159 15861 19171 15864
rect 19205 15861 19217 15895
rect 19159 15855 19217 15861
rect 22738 15852 22744 15904
rect 22796 15852 22802 15904
rect 23676 15892 23704 16068
rect 23842 16056 23848 16108
rect 23900 16056 23906 16108
rect 24210 16105 24216 16108
rect 24172 16099 24216 16105
rect 24172 16065 24184 16099
rect 24172 16059 24216 16065
rect 24210 16056 24216 16059
rect 24268 16056 24274 16108
rect 24351 16099 24409 16105
rect 24351 16065 24363 16099
rect 24397 16096 24409 16099
rect 25958 16096 25964 16108
rect 24397 16068 25964 16096
rect 24397 16065 24409 16068
rect 24351 16059 24409 16065
rect 25958 16056 25964 16068
rect 26016 16056 26022 16108
rect 26418 16105 26424 16108
rect 26380 16099 26424 16105
rect 26380 16065 26392 16099
rect 26380 16059 26424 16065
rect 26418 16056 26424 16059
rect 26476 16056 26482 16108
rect 26516 16097 26574 16103
rect 26516 16063 26528 16097
rect 26562 16096 26574 16097
rect 26789 16099 26847 16105
rect 26562 16068 26648 16096
rect 26562 16063 26574 16068
rect 26516 16057 26574 16063
rect 26620 16040 26648 16068
rect 26789 16065 26801 16099
rect 26835 16096 26847 16099
rect 28966 16096 28994 16124
rect 26835 16068 28994 16096
rect 26835 16065 26847 16068
rect 26789 16059 26847 16065
rect 29270 16056 29276 16108
rect 29328 16056 29334 16108
rect 29457 16099 29515 16105
rect 29457 16065 29469 16099
rect 29503 16096 29515 16099
rect 29564 16096 29592 16124
rect 29503 16068 29592 16096
rect 29656 16096 29684 16127
rect 30006 16124 30012 16176
rect 30064 16124 30070 16176
rect 30024 16096 30052 16124
rect 29656 16068 30052 16096
rect 29503 16065 29515 16068
rect 29457 16059 29515 16065
rect 23934 15988 23940 16040
rect 23992 16028 23998 16040
rect 24581 16031 24639 16037
rect 24581 16028 24593 16031
rect 23992 16000 24593 16028
rect 23992 15988 23998 16000
rect 24581 15997 24593 16000
rect 24627 15997 24639 16031
rect 24581 15991 24639 15997
rect 26053 16031 26111 16037
rect 26053 15997 26065 16031
rect 26099 16028 26111 16031
rect 26142 16028 26148 16040
rect 26099 16000 26148 16028
rect 26099 15997 26111 16000
rect 26053 15991 26111 15997
rect 26142 15988 26148 16000
rect 26200 15988 26206 16040
rect 26602 15988 26608 16040
rect 26660 15988 26666 16040
rect 27154 15988 27160 16040
rect 27212 16028 27218 16040
rect 28166 16028 28172 16040
rect 27212 16000 28172 16028
rect 27212 15988 27218 16000
rect 28166 15988 28172 16000
rect 28224 16028 28230 16040
rect 28261 16031 28319 16037
rect 28261 16028 28273 16031
rect 28224 16000 28273 16028
rect 28224 15988 28230 16000
rect 28261 15997 28273 16000
rect 28307 15997 28319 16031
rect 28261 15991 28319 15997
rect 28718 15988 28724 16040
rect 28776 15988 28782 16040
rect 28813 16031 28871 16037
rect 28813 15997 28825 16031
rect 28859 16028 28871 16031
rect 28902 16028 28908 16040
rect 28859 16000 28908 16028
rect 28859 15997 28871 16000
rect 28813 15991 28871 15997
rect 28902 15988 28908 16000
rect 28960 15988 28966 16040
rect 28994 15988 29000 16040
rect 29052 16028 29058 16040
rect 29181 16031 29239 16037
rect 29052 16024 29132 16028
rect 29181 16024 29193 16031
rect 29052 16000 29193 16024
rect 29052 15988 29058 16000
rect 29104 15997 29193 16000
rect 29227 15997 29239 16031
rect 29104 15996 29239 15997
rect 29288 16024 29316 16056
rect 30009 16031 30067 16037
rect 30009 16028 30021 16031
rect 29288 16015 29390 16024
rect 29656 16022 30021 16028
rect 29288 16009 29405 16015
rect 29288 15996 29359 16009
rect 29181 15991 29239 15996
rect 27522 15920 27528 15972
rect 27580 15960 27586 15972
rect 28736 15960 28764 15988
rect 29347 15975 29359 15996
rect 29393 15975 29405 16009
rect 29564 16004 30021 16022
rect 29347 15969 29405 15975
rect 29472 16000 30021 16004
rect 29472 15994 29684 16000
rect 30009 15997 30021 16000
rect 30055 15997 30067 16031
rect 29472 15976 29592 15994
rect 30009 15991 30067 15997
rect 30193 16031 30251 16037
rect 30193 15997 30205 16031
rect 30239 15997 30251 16031
rect 30193 15991 30251 15997
rect 27580 15932 28672 15960
rect 28736 15932 29224 15960
rect 27580 15920 27586 15932
rect 24118 15892 24124 15904
rect 23676 15864 24124 15892
rect 24118 15852 24124 15864
rect 24176 15852 24182 15904
rect 24302 15852 24308 15904
rect 24360 15892 24366 15904
rect 28644 15901 28672 15932
rect 27893 15895 27951 15901
rect 27893 15892 27905 15895
rect 24360 15864 27905 15892
rect 24360 15852 24366 15864
rect 27893 15861 27905 15864
rect 27939 15861 27951 15895
rect 27893 15855 27951 15861
rect 28629 15895 28687 15901
rect 28629 15861 28641 15895
rect 28675 15861 28687 15895
rect 29196 15892 29224 15932
rect 29270 15892 29276 15904
rect 29196 15864 29276 15892
rect 28629 15855 28687 15861
rect 29270 15852 29276 15864
rect 29328 15892 29334 15904
rect 29472 15892 29500 15976
rect 29328 15864 29500 15892
rect 29328 15852 29334 15864
rect 29546 15852 29552 15904
rect 29604 15892 29610 15904
rect 29825 15895 29883 15901
rect 29825 15892 29837 15895
rect 29604 15864 29837 15892
rect 29604 15852 29610 15864
rect 29825 15861 29837 15864
rect 29871 15861 29883 15895
rect 29825 15855 29883 15861
rect 30006 15852 30012 15904
rect 30064 15892 30070 15904
rect 30208 15892 30236 15991
rect 30374 15920 30380 15972
rect 30432 15960 30438 15972
rect 30484 15960 30512 16204
rect 30432 15932 30512 15960
rect 30432 15920 30438 15932
rect 30064 15864 30236 15892
rect 30064 15852 30070 15864
rect 31018 15852 31024 15904
rect 31076 15892 31082 15904
rect 31076 15864 31340 15892
rect 31076 15852 31082 15864
rect 552 15802 31072 15824
rect 552 15750 7988 15802
rect 8040 15750 8052 15802
rect 8104 15750 8116 15802
rect 8168 15750 8180 15802
rect 8232 15750 8244 15802
rect 8296 15750 15578 15802
rect 15630 15750 15642 15802
rect 15694 15750 15706 15802
rect 15758 15750 15770 15802
rect 15822 15750 15834 15802
rect 15886 15750 23168 15802
rect 23220 15750 23232 15802
rect 23284 15750 23296 15802
rect 23348 15750 23360 15802
rect 23412 15750 23424 15802
rect 23476 15750 30758 15802
rect 30810 15750 30822 15802
rect 30874 15750 30886 15802
rect 30938 15750 30950 15802
rect 31002 15750 31014 15802
rect 31066 15750 31072 15802
rect 552 15728 31072 15750
rect 1044 15660 3096 15688
rect 1044 15561 1072 15660
rect 3068 15620 3096 15660
rect 3142 15648 3148 15700
rect 3200 15648 3206 15700
rect 4982 15688 4988 15700
rect 3620 15660 4988 15688
rect 3620 15620 3648 15660
rect 4982 15648 4988 15660
rect 5040 15648 5046 15700
rect 10505 15691 10563 15697
rect 10505 15688 10517 15691
rect 5736 15660 10517 15688
rect 3068 15592 3648 15620
rect 1029 15555 1087 15561
rect 1029 15521 1041 15555
rect 1075 15521 1087 15555
rect 5736 15552 5764 15660
rect 10505 15657 10517 15660
rect 10551 15657 10563 15691
rect 10505 15651 10563 15657
rect 11425 15691 11483 15697
rect 11425 15657 11437 15691
rect 11471 15688 11483 15691
rect 11882 15688 11888 15700
rect 11471 15660 11888 15688
rect 11471 15657 11483 15660
rect 11425 15651 11483 15657
rect 11882 15648 11888 15660
rect 11940 15648 11946 15700
rect 11974 15648 11980 15700
rect 12032 15688 12038 15700
rect 13078 15688 13084 15700
rect 12032 15660 13084 15688
rect 12032 15648 12038 15660
rect 13078 15648 13084 15660
rect 13136 15648 13142 15700
rect 14182 15648 14188 15700
rect 14240 15688 14246 15700
rect 14283 15691 14341 15697
rect 14283 15688 14295 15691
rect 14240 15660 14295 15688
rect 14240 15648 14246 15660
rect 14283 15657 14295 15660
rect 14329 15657 14341 15691
rect 14283 15651 14341 15657
rect 14826 15648 14832 15700
rect 14884 15688 14890 15700
rect 18230 15688 18236 15700
rect 14884 15660 18236 15688
rect 14884 15648 14890 15660
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 23750 15688 23756 15700
rect 19352 15660 23756 15688
rect 6454 15580 6460 15632
rect 6512 15580 6518 15632
rect 11698 15580 11704 15632
rect 11756 15580 11762 15632
rect 16942 15580 16948 15632
rect 17000 15620 17006 15632
rect 17000 15592 17264 15620
rect 17000 15580 17006 15592
rect 1029 15515 1087 15521
rect 1970 15524 5764 15552
rect 5905 15555 5963 15561
rect 1801 15505 1859 15511
rect 1670 15493 1676 15496
rect 1305 15487 1363 15493
rect 1305 15453 1317 15487
rect 1351 15453 1363 15487
rect 1305 15447 1363 15453
rect 1632 15487 1676 15493
rect 1632 15453 1644 15487
rect 1632 15447 1676 15453
rect 842 15308 848 15360
rect 900 15308 906 15360
rect 1118 15308 1124 15360
rect 1176 15348 1182 15360
rect 1320 15348 1348 15447
rect 1670 15444 1676 15447
rect 1728 15444 1734 15496
rect 1801 15471 1813 15505
rect 1847 15484 1859 15505
rect 1970 15484 1998 15524
rect 5905 15521 5917 15555
rect 5951 15521 5963 15555
rect 6472 15552 6500 15580
rect 6784 15555 6842 15561
rect 6784 15552 6796 15555
rect 6472 15524 6796 15552
rect 5905 15515 5963 15521
rect 6784 15521 6796 15524
rect 6830 15521 6842 15555
rect 11149 15555 11207 15561
rect 6784 15515 6842 15521
rect 7116 15524 11100 15552
rect 1847 15471 1998 15484
rect 1801 15465 1998 15471
rect 1816 15456 1998 15465
rect 2038 15444 2044 15496
rect 2096 15444 2102 15496
rect 3510 15444 3516 15496
rect 3568 15444 3574 15496
rect 3878 15493 3884 15496
rect 3840 15487 3884 15493
rect 3840 15453 3852 15487
rect 3840 15447 3884 15453
rect 3878 15444 3884 15447
rect 3936 15444 3942 15496
rect 3970 15444 3976 15496
rect 4028 15484 4034 15496
rect 4249 15487 4307 15493
rect 4028 15456 4073 15484
rect 4028 15444 4034 15456
rect 4249 15453 4261 15487
rect 4295 15484 4307 15487
rect 4614 15484 4620 15496
rect 4295 15456 4620 15484
rect 4295 15453 4307 15456
rect 4249 15447 4307 15453
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 5629 15487 5687 15493
rect 5629 15453 5641 15487
rect 5675 15484 5687 15487
rect 5718 15484 5724 15496
rect 5675 15456 5724 15484
rect 5675 15453 5687 15456
rect 5629 15447 5687 15453
rect 5718 15444 5724 15456
rect 5776 15444 5782 15496
rect 3528 15348 3556 15444
rect 3786 15348 3792 15360
rect 1176 15320 3792 15348
rect 1176 15308 1182 15320
rect 3786 15308 3792 15320
rect 3844 15348 3850 15360
rect 5920 15348 5948 15515
rect 6953 15505 7011 15511
rect 6953 15502 6965 15505
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15453 6515 15487
rect 6938 15471 6965 15502
rect 6999 15484 7011 15505
rect 7116 15484 7144 15524
rect 6999 15471 7144 15484
rect 6938 15456 7144 15471
rect 6457 15447 6515 15453
rect 3844 15320 5948 15348
rect 3844 15308 3850 15320
rect 6178 15308 6184 15360
rect 6236 15348 6242 15360
rect 6472 15348 6500 15447
rect 7190 15444 7196 15496
rect 7248 15444 7254 15496
rect 7650 15444 7656 15496
rect 7708 15484 7714 15496
rect 7834 15484 7840 15496
rect 7708 15456 7840 15484
rect 7708 15444 7714 15456
rect 7834 15444 7840 15456
rect 7892 15444 7898 15496
rect 8662 15484 8668 15496
rect 8266 15456 8668 15484
rect 8266 15416 8294 15456
rect 8662 15444 8668 15456
rect 8720 15444 8726 15496
rect 8846 15444 8852 15496
rect 8904 15484 8910 15496
rect 8992 15487 9050 15493
rect 8992 15484 9004 15487
rect 8904 15456 9004 15484
rect 8904 15444 8910 15456
rect 8992 15453 9004 15456
rect 9038 15453 9050 15487
rect 8992 15447 9050 15453
rect 9122 15444 9128 15496
rect 9180 15484 9186 15496
rect 9180 15456 9225 15484
rect 9180 15444 9186 15456
rect 9306 15444 9312 15496
rect 9364 15484 9370 15496
rect 9401 15487 9459 15493
rect 9401 15484 9413 15487
rect 9364 15456 9413 15484
rect 9364 15444 9370 15456
rect 9401 15453 9413 15456
rect 9447 15453 9459 15487
rect 9401 15447 9459 15453
rect 7852 15388 8294 15416
rect 7852 15348 7880 15388
rect 6236 15320 7880 15348
rect 6236 15308 6242 15320
rect 8294 15308 8300 15360
rect 8352 15308 8358 15360
rect 11072 15348 11100 15524
rect 11149 15521 11161 15555
rect 11195 15552 11207 15555
rect 11238 15552 11244 15564
rect 11195 15524 11244 15552
rect 11195 15521 11207 15524
rect 11149 15515 11207 15521
rect 11238 15512 11244 15524
rect 11296 15552 11302 15564
rect 11609 15555 11667 15561
rect 11609 15552 11621 15555
rect 11296 15524 11621 15552
rect 11296 15512 11302 15524
rect 11609 15521 11621 15524
rect 11655 15521 11667 15555
rect 11716 15552 11744 15580
rect 11936 15555 11994 15561
rect 11936 15552 11948 15555
rect 11716 15524 11948 15552
rect 11609 15515 11667 15521
rect 11936 15521 11948 15524
rect 11982 15521 11994 15555
rect 11936 15515 11994 15521
rect 12268 15524 12848 15552
rect 12115 15487 12173 15493
rect 12115 15453 12127 15487
rect 12161 15484 12173 15487
rect 12268 15484 12296 15524
rect 12161 15456 12296 15484
rect 12345 15487 12403 15493
rect 12161 15453 12173 15456
rect 12115 15447 12173 15453
rect 12345 15453 12357 15487
rect 12391 15484 12403 15487
rect 12710 15484 12716 15496
rect 12391 15456 12716 15484
rect 12391 15453 12403 15456
rect 12345 15447 12403 15453
rect 12710 15444 12716 15456
rect 12768 15444 12774 15496
rect 12820 15484 12848 15524
rect 13446 15512 13452 15564
rect 13504 15552 13510 15564
rect 13814 15552 13820 15564
rect 13504 15524 13820 15552
rect 13504 15512 13510 15524
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 14458 15512 14464 15564
rect 14516 15512 14522 15564
rect 14553 15555 14611 15561
rect 14553 15521 14565 15555
rect 14599 15552 14611 15555
rect 15930 15552 15936 15564
rect 14599 15524 15936 15552
rect 14599 15521 14611 15524
rect 14553 15515 14611 15521
rect 15930 15512 15936 15524
rect 15988 15512 15994 15564
rect 16209 15555 16267 15561
rect 16209 15521 16221 15555
rect 16255 15521 16267 15555
rect 16209 15515 16267 15521
rect 14323 15487 14381 15493
rect 12820 15456 13860 15484
rect 11974 15348 11980 15360
rect 11072 15320 11980 15348
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 13446 15308 13452 15360
rect 13504 15308 13510 15360
rect 13832 15348 13860 15456
rect 14323 15453 14335 15487
rect 14369 15484 14381 15487
rect 14476 15484 14504 15512
rect 14369 15456 14504 15484
rect 14369 15453 14381 15456
rect 14323 15447 14381 15453
rect 14734 15444 14740 15496
rect 14792 15484 14798 15496
rect 16224 15484 16252 15515
rect 17034 15512 17040 15564
rect 17092 15512 17098 15564
rect 17236 15552 17264 15592
rect 17456 15555 17514 15561
rect 17456 15552 17468 15555
rect 17236 15524 17468 15552
rect 17328 15496 17356 15524
rect 17456 15521 17468 15524
rect 17502 15521 17514 15555
rect 17456 15515 17514 15521
rect 17865 15555 17923 15561
rect 17865 15521 17877 15555
rect 17911 15552 17923 15555
rect 19150 15552 19156 15564
rect 17911 15524 19156 15552
rect 17911 15521 17923 15524
rect 17865 15515 17923 15521
rect 19150 15512 19156 15524
rect 19208 15512 19214 15564
rect 17625 15505 17683 15511
rect 17625 15502 17637 15505
rect 17126 15484 17132 15496
rect 14792 15456 16252 15484
rect 16684 15456 17132 15484
rect 14792 15444 14798 15456
rect 15212 15388 16068 15416
rect 15212 15348 15240 15388
rect 16040 15360 16068 15388
rect 16684 15360 16712 15456
rect 17126 15444 17132 15456
rect 17184 15444 17190 15496
rect 17310 15444 17316 15496
rect 17368 15444 17374 15496
rect 17604 15471 17637 15502
rect 17671 15484 17683 15505
rect 19352 15484 19380 15660
rect 23750 15648 23756 15660
rect 23808 15648 23814 15700
rect 23943 15691 24001 15697
rect 23943 15657 23955 15691
rect 23989 15688 24001 15691
rect 24210 15688 24216 15700
rect 23989 15660 24216 15688
rect 23989 15657 24001 15660
rect 23943 15651 24001 15657
rect 24210 15648 24216 15660
rect 24268 15648 24274 15700
rect 27522 15688 27528 15700
rect 24872 15660 27528 15688
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15552 19763 15555
rect 21358 15552 21364 15564
rect 19751 15524 21364 15552
rect 19751 15521 19763 15524
rect 19705 15515 19763 15521
rect 21358 15512 21364 15524
rect 21416 15512 21422 15564
rect 21542 15512 21548 15564
rect 21600 15561 21606 15564
rect 21600 15555 21654 15561
rect 21600 15521 21608 15555
rect 21642 15521 21654 15555
rect 21600 15515 21654 15521
rect 21600 15512 21606 15515
rect 23842 15512 23848 15564
rect 23900 15512 23906 15564
rect 24213 15555 24271 15561
rect 24213 15521 24225 15555
rect 24259 15552 24271 15555
rect 24872 15552 24900 15660
rect 27522 15648 27528 15660
rect 27580 15648 27586 15700
rect 28258 15648 28264 15700
rect 28316 15688 28322 15700
rect 28451 15691 28509 15697
rect 28451 15688 28463 15691
rect 28316 15660 28463 15688
rect 28316 15648 28322 15660
rect 28451 15657 28463 15660
rect 28497 15657 28509 15691
rect 28451 15651 28509 15657
rect 28994 15648 29000 15700
rect 29052 15688 29058 15700
rect 29052 15660 29408 15688
rect 29052 15648 29058 15660
rect 26418 15580 26424 15632
rect 26476 15620 26482 15632
rect 27157 15623 27215 15629
rect 27157 15620 27169 15623
rect 26476 15592 27169 15620
rect 26476 15580 26482 15592
rect 27157 15589 27169 15592
rect 27203 15589 27215 15623
rect 29380 15620 29408 15660
rect 29638 15648 29644 15700
rect 29696 15688 29702 15700
rect 29825 15691 29883 15697
rect 29825 15688 29837 15691
rect 29696 15660 29837 15688
rect 29696 15648 29702 15660
rect 29825 15657 29837 15660
rect 29871 15657 29883 15691
rect 29825 15651 29883 15657
rect 31018 15648 31024 15700
rect 31076 15688 31082 15700
rect 31202 15688 31208 15700
rect 31076 15660 31208 15688
rect 31076 15648 31082 15660
rect 31202 15648 31208 15660
rect 31260 15648 31266 15700
rect 29730 15620 29736 15632
rect 29380 15592 29736 15620
rect 27157 15583 27215 15589
rect 29730 15580 29736 15592
rect 29788 15580 29794 15632
rect 30926 15580 30932 15632
rect 30984 15620 30990 15632
rect 31312 15620 31340 15864
rect 30984 15592 31340 15620
rect 30984 15580 30990 15592
rect 24259 15524 24900 15552
rect 25777 15555 25835 15561
rect 24259 15521 24271 15524
rect 24213 15515 24271 15521
rect 25777 15521 25789 15555
rect 25823 15521 25835 15555
rect 25777 15515 25835 15521
rect 17671 15471 19380 15484
rect 17604 15456 19380 15471
rect 19429 15487 19487 15493
rect 19429 15453 19441 15487
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 18598 15376 18604 15428
rect 18656 15416 18662 15428
rect 19242 15416 19248 15428
rect 18656 15388 19248 15416
rect 18656 15376 18662 15388
rect 19242 15376 19248 15388
rect 19300 15416 19306 15428
rect 19444 15416 19472 15447
rect 19794 15444 19800 15496
rect 19852 15484 19858 15496
rect 20898 15484 20904 15496
rect 19852 15456 20904 15484
rect 19852 15444 19858 15456
rect 20898 15444 20904 15456
rect 20956 15484 20962 15496
rect 21266 15484 21272 15496
rect 20956 15456 21272 15484
rect 20956 15444 20962 15456
rect 21266 15444 21272 15456
rect 21324 15444 21330 15496
rect 21818 15495 21824 15496
rect 21775 15489 21824 15495
rect 21775 15455 21787 15489
rect 21821 15455 21824 15489
rect 21775 15449 21824 15455
rect 21818 15444 21824 15449
rect 21876 15444 21882 15496
rect 22002 15444 22008 15496
rect 22060 15444 22066 15496
rect 23477 15487 23535 15493
rect 23477 15453 23489 15487
rect 23523 15484 23535 15487
rect 23658 15484 23664 15496
rect 23523 15456 23664 15484
rect 23523 15453 23535 15456
rect 23477 15447 23535 15453
rect 23658 15444 23664 15456
rect 23716 15484 23722 15496
rect 23860 15484 23888 15512
rect 23973 15505 24031 15511
rect 23973 15502 23985 15505
rect 23716 15456 23888 15484
rect 23971 15471 23985 15502
rect 24019 15498 24031 15505
rect 24019 15471 24032 15498
rect 23971 15456 24032 15471
rect 23716 15444 23722 15456
rect 24026 15446 24032 15456
rect 24084 15446 24090 15498
rect 24118 15444 24124 15496
rect 24176 15484 24182 15496
rect 24176 15456 25360 15484
rect 24176 15444 24182 15456
rect 25332 15425 25360 15456
rect 25317 15419 25375 15425
rect 19300 15388 19472 15416
rect 20364 15388 21128 15416
rect 19300 15376 19306 15388
rect 13832 15320 15240 15348
rect 15378 15308 15384 15360
rect 15436 15348 15442 15360
rect 15657 15351 15715 15357
rect 15657 15348 15669 15351
rect 15436 15320 15669 15348
rect 15436 15308 15442 15320
rect 15657 15317 15669 15320
rect 15703 15317 15715 15351
rect 15657 15311 15715 15317
rect 16022 15308 16028 15360
rect 16080 15308 16086 15360
rect 16485 15351 16543 15357
rect 16485 15317 16497 15351
rect 16531 15348 16543 15351
rect 16666 15348 16672 15360
rect 16531 15320 16672 15348
rect 16531 15317 16543 15320
rect 16485 15311 16543 15317
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 16850 15308 16856 15360
rect 16908 15308 16914 15360
rect 18966 15308 18972 15360
rect 19024 15308 19030 15360
rect 19794 15308 19800 15360
rect 19852 15348 19858 15360
rect 20364 15348 20392 15388
rect 19852 15320 20392 15348
rect 19852 15308 19858 15320
rect 20990 15308 20996 15360
rect 21048 15308 21054 15360
rect 21100 15348 21128 15388
rect 25317 15385 25329 15419
rect 25363 15385 25375 15419
rect 25317 15379 25375 15385
rect 22002 15348 22008 15360
rect 21100 15320 22008 15348
rect 22002 15308 22008 15320
rect 22060 15308 22066 15360
rect 22646 15308 22652 15360
rect 22704 15348 22710 15360
rect 23109 15351 23167 15357
rect 23109 15348 23121 15351
rect 22704 15320 23121 15348
rect 22704 15308 22710 15320
rect 23109 15317 23121 15320
rect 23155 15317 23167 15351
rect 23109 15311 23167 15317
rect 24026 15308 24032 15360
rect 24084 15348 24090 15360
rect 25792 15348 25820 15515
rect 26326 15512 26332 15564
rect 26384 15552 26390 15564
rect 26513 15555 26571 15561
rect 26513 15552 26525 15555
rect 26384 15524 26525 15552
rect 26384 15512 26390 15524
rect 26513 15521 26525 15524
rect 26559 15552 26571 15555
rect 26786 15552 26792 15564
rect 26559 15524 26792 15552
rect 26559 15521 26571 15524
rect 26513 15515 26571 15521
rect 26786 15512 26792 15524
rect 26844 15512 26850 15564
rect 26881 15555 26939 15561
rect 26881 15521 26893 15555
rect 26927 15552 26939 15555
rect 26970 15552 26976 15564
rect 26927 15524 26976 15552
rect 26927 15521 26939 15524
rect 26881 15515 26939 15521
rect 26970 15512 26976 15524
rect 27028 15512 27034 15564
rect 27614 15512 27620 15564
rect 27672 15512 27678 15564
rect 28368 15524 28994 15552
rect 26053 15487 26111 15493
rect 26053 15453 26065 15487
rect 26099 15484 26111 15487
rect 26142 15484 26148 15496
rect 26099 15456 26148 15484
rect 26099 15453 26111 15456
rect 26053 15447 26111 15453
rect 26142 15444 26148 15456
rect 26200 15484 26206 15496
rect 26200 15456 27936 15484
rect 26200 15444 26206 15456
rect 27801 15419 27859 15425
rect 27801 15416 27813 15419
rect 26344 15388 27813 15416
rect 26344 15360 26372 15388
rect 27801 15385 27813 15388
rect 27847 15385 27859 15419
rect 27801 15379 27859 15385
rect 24084 15320 25820 15348
rect 24084 15308 24090 15320
rect 26326 15308 26332 15360
rect 26384 15308 26390 15360
rect 26418 15308 26424 15360
rect 26476 15348 26482 15360
rect 26697 15351 26755 15357
rect 26697 15348 26709 15351
rect 26476 15320 26709 15348
rect 26476 15308 26482 15320
rect 26697 15317 26709 15320
rect 26743 15317 26755 15351
rect 26697 15311 26755 15317
rect 26786 15308 26792 15360
rect 26844 15348 26850 15360
rect 26970 15348 26976 15360
rect 26844 15320 26976 15348
rect 26844 15308 26850 15320
rect 26970 15308 26976 15320
rect 27028 15308 27034 15360
rect 27908 15348 27936 15456
rect 27982 15444 27988 15496
rect 28040 15444 28046 15496
rect 28166 15444 28172 15496
rect 28224 15484 28230 15496
rect 28368 15484 28396 15524
rect 28534 15493 28540 15496
rect 28224 15456 28396 15484
rect 28491 15487 28540 15493
rect 28224 15444 28230 15456
rect 28491 15453 28503 15487
rect 28537 15453 28540 15487
rect 28491 15447 28540 15453
rect 28534 15444 28540 15447
rect 28592 15444 28598 15496
rect 28718 15444 28724 15496
rect 28776 15444 28782 15496
rect 28966 15484 28994 15524
rect 30006 15512 30012 15564
rect 30064 15552 30070 15564
rect 30193 15555 30251 15561
rect 30193 15552 30205 15555
rect 30064 15524 30205 15552
rect 30064 15512 30070 15524
rect 30193 15521 30205 15524
rect 30239 15521 30251 15555
rect 30193 15515 30251 15521
rect 28966 15456 30420 15484
rect 30392 15425 30420 15456
rect 30377 15419 30435 15425
rect 30377 15385 30389 15419
rect 30423 15416 30435 15419
rect 31202 15416 31208 15428
rect 30423 15388 31208 15416
rect 30423 15385 30435 15388
rect 30377 15379 30435 15385
rect 31202 15376 31208 15388
rect 31260 15376 31266 15428
rect 28350 15348 28356 15360
rect 27908 15320 28356 15348
rect 28350 15308 28356 15320
rect 28408 15308 28414 15360
rect 552 15258 30912 15280
rect 552 15206 4193 15258
rect 4245 15206 4257 15258
rect 4309 15206 4321 15258
rect 4373 15206 4385 15258
rect 4437 15206 4449 15258
rect 4501 15206 11783 15258
rect 11835 15206 11847 15258
rect 11899 15206 11911 15258
rect 11963 15206 11975 15258
rect 12027 15206 12039 15258
rect 12091 15206 19373 15258
rect 19425 15206 19437 15258
rect 19489 15206 19501 15258
rect 19553 15206 19565 15258
rect 19617 15206 19629 15258
rect 19681 15206 26963 15258
rect 27015 15206 27027 15258
rect 27079 15206 27091 15258
rect 27143 15206 27155 15258
rect 27207 15206 27219 15258
rect 27271 15206 30912 15258
rect 552 15184 30912 15206
rect 1394 15104 1400 15156
rect 1452 15144 1458 15156
rect 2777 15147 2835 15153
rect 1452 15116 2360 15144
rect 1452 15104 1458 15116
rect 2332 15076 2360 15116
rect 2777 15113 2789 15147
rect 2823 15144 2835 15147
rect 2866 15144 2872 15156
rect 2823 15116 2872 15144
rect 2823 15113 2835 15116
rect 2777 15107 2835 15113
rect 2866 15104 2872 15116
rect 2924 15104 2930 15156
rect 5718 15144 5724 15156
rect 3252 15116 5724 15144
rect 3252 15076 3280 15116
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 5813 15147 5871 15153
rect 5813 15113 5825 15147
rect 5859 15144 5871 15147
rect 5902 15144 5908 15156
rect 5859 15116 5908 15144
rect 5859 15113 5871 15116
rect 5813 15107 5871 15113
rect 5902 15104 5908 15116
rect 5960 15104 5966 15156
rect 8294 15144 8300 15156
rect 6104 15116 8300 15144
rect 2332 15048 3280 15076
rect 937 15011 995 15017
rect 937 14977 949 15011
rect 983 15008 995 15011
rect 1118 15008 1124 15020
rect 983 14980 1124 15008
rect 983 14977 995 14980
rect 937 14971 995 14977
rect 1118 14968 1124 14980
rect 1176 14968 1182 15020
rect 1302 14968 1308 15020
rect 1360 14968 1366 15020
rect 1443 15011 1501 15017
rect 1443 14977 1455 15011
rect 1489 15008 1501 15011
rect 3050 15008 3056 15020
rect 1489 14980 3056 15008
rect 1489 14977 1501 14980
rect 1443 14971 1501 14977
rect 3050 14968 3056 14980
rect 3108 14968 3114 15020
rect 1320 14940 1348 14968
rect 3252 14949 3280 15048
rect 3786 14968 3792 15020
rect 3844 14968 3850 15020
rect 4295 15011 4353 15017
rect 4295 14977 4307 15011
rect 4341 15008 4353 15011
rect 6104 15008 6132 15116
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 13081 15147 13139 15153
rect 13081 15144 13093 15147
rect 8680 15116 13093 15144
rect 4341 14980 6132 15008
rect 6595 15011 6653 15017
rect 4341 14977 4353 14980
rect 4295 14971 4353 14977
rect 6595 14977 6607 15011
rect 6641 15008 6653 15011
rect 8680 15008 8708 15116
rect 13081 15113 13093 15116
rect 13127 15113 13139 15147
rect 13081 15107 13139 15113
rect 13262 15104 13268 15156
rect 13320 15144 13326 15156
rect 14277 15147 14335 15153
rect 14277 15144 14289 15147
rect 13320 15116 14289 15144
rect 13320 15104 13326 15116
rect 14277 15113 14289 15116
rect 14323 15144 14335 15147
rect 14458 15144 14464 15156
rect 14323 15116 14464 15144
rect 14323 15113 14335 15116
rect 14277 15107 14335 15113
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 15838 15144 15844 15156
rect 14568 15116 15844 15144
rect 10962 15036 10968 15088
rect 11020 15036 11026 15088
rect 13998 15036 14004 15088
rect 14056 15076 14062 15088
rect 14568 15076 14596 15116
rect 15838 15104 15844 15116
rect 15896 15104 15902 15156
rect 18432 15116 21128 15144
rect 18432 15085 18460 15116
rect 14056 15048 14596 15076
rect 18417 15079 18475 15085
rect 14056 15036 14062 15048
rect 18417 15045 18429 15079
rect 18463 15045 18475 15079
rect 18417 15039 18475 15045
rect 6641 14980 8708 15008
rect 6641 14977 6653 14980
rect 6595 14971 6653 14977
rect 8846 14968 8852 15020
rect 8904 15008 8910 15020
rect 8992 15011 9050 15017
rect 8992 15008 9004 15011
rect 8904 14980 9004 15008
rect 8904 14968 8910 14980
rect 8992 14977 9004 14980
rect 9038 14977 9050 15011
rect 8992 14971 9050 14977
rect 9171 15011 9229 15017
rect 9171 14977 9183 15011
rect 9217 15008 9229 15011
rect 10778 15008 10784 15020
rect 9217 14980 10784 15008
rect 9217 14977 9229 14980
rect 9171 14971 9229 14977
rect 10778 14968 10784 14980
rect 10836 14968 10842 15020
rect 11238 14968 11244 15020
rect 11296 14968 11302 15020
rect 11747 15011 11805 15017
rect 11747 14977 11759 15011
rect 11793 15008 11805 15011
rect 11793 14980 13492 15008
rect 11793 14977 11805 14980
rect 11747 14971 11805 14977
rect 1673 14943 1731 14949
rect 1673 14940 1685 14943
rect 1320 14912 1685 14940
rect 1673 14909 1685 14912
rect 1719 14909 1731 14943
rect 1673 14903 1731 14909
rect 3237 14943 3295 14949
rect 3237 14909 3249 14943
rect 3283 14909 3295 14943
rect 3237 14903 3295 14909
rect 3878 14900 3884 14952
rect 3936 14940 3942 14952
rect 4116 14943 4174 14949
rect 4116 14940 4128 14943
rect 3936 14912 4128 14940
rect 3936 14900 3942 14912
rect 4116 14909 4128 14912
rect 4162 14909 4174 14943
rect 4116 14903 4174 14909
rect 4522 14900 4528 14952
rect 4580 14900 4586 14952
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 6089 14943 6147 14949
rect 6089 14940 6101 14943
rect 5684 14912 6101 14940
rect 5684 14900 5690 14912
rect 6089 14909 6101 14912
rect 6135 14940 6147 14943
rect 6178 14940 6184 14952
rect 6135 14912 6184 14940
rect 6135 14909 6147 14912
rect 6089 14903 6147 14909
rect 6178 14900 6184 14912
rect 6236 14900 6242 14952
rect 6454 14949 6460 14952
rect 6416 14943 6460 14949
rect 6416 14909 6428 14943
rect 6512 14940 6518 14952
rect 6730 14940 6736 14952
rect 6512 14912 6736 14940
rect 6416 14903 6460 14909
rect 6454 14900 6460 14903
rect 6512 14900 6518 14912
rect 6730 14900 6736 14912
rect 6788 14900 6794 14952
rect 6822 14900 6828 14952
rect 6880 14900 6886 14952
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 8386 14940 8392 14952
rect 6972 14912 8392 14940
rect 6972 14900 6978 14912
rect 8386 14900 8392 14912
rect 8444 14940 8450 14952
rect 8573 14943 8631 14949
rect 8573 14940 8585 14943
rect 8444 14912 8585 14940
rect 8444 14900 8450 14912
rect 8573 14909 8585 14912
rect 8619 14909 8631 14943
rect 8573 14903 8631 14909
rect 8662 14900 8668 14952
rect 8720 14900 8726 14952
rect 9401 14943 9459 14949
rect 9401 14940 9413 14943
rect 8772 14912 9413 14940
rect 3513 14875 3571 14881
rect 3513 14872 3525 14875
rect 2746 14844 3525 14872
rect 1403 14807 1461 14813
rect 1403 14773 1415 14807
rect 1449 14804 1461 14807
rect 1670 14804 1676 14816
rect 1449 14776 1676 14804
rect 1449 14773 1461 14776
rect 1403 14767 1461 14773
rect 1670 14764 1676 14776
rect 1728 14804 1734 14816
rect 2746 14804 2774 14844
rect 3513 14841 3525 14844
rect 3559 14872 3571 14875
rect 3896 14872 3924 14900
rect 3559 14844 3924 14872
rect 3559 14841 3571 14844
rect 3513 14835 3571 14841
rect 7558 14832 7564 14884
rect 7616 14872 7622 14884
rect 8478 14872 8484 14884
rect 7616 14844 8484 14872
rect 7616 14832 7622 14844
rect 8478 14832 8484 14844
rect 8536 14832 8542 14884
rect 1728 14776 2774 14804
rect 1728 14764 1734 14776
rect 4062 14764 4068 14816
rect 4120 14804 4126 14816
rect 7929 14807 7987 14813
rect 7929 14804 7941 14807
rect 4120 14776 7941 14804
rect 4120 14764 4126 14776
rect 7929 14773 7941 14776
rect 7975 14773 7987 14807
rect 7929 14767 7987 14773
rect 8389 14807 8447 14813
rect 8389 14773 8401 14807
rect 8435 14804 8447 14807
rect 8772 14804 8800 14912
rect 9401 14909 9413 14912
rect 9447 14909 9459 14943
rect 11149 14943 11207 14949
rect 11149 14940 11161 14943
rect 9401 14903 9459 14909
rect 10980 14912 11161 14940
rect 10980 14816 11008 14912
rect 11149 14909 11161 14912
rect 11195 14940 11207 14943
rect 11330 14940 11336 14952
rect 11195 14912 11336 14940
rect 11195 14909 11207 14912
rect 11149 14903 11207 14909
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 11974 14900 11980 14952
rect 12032 14900 12038 14952
rect 12802 14900 12808 14952
rect 12860 14900 12866 14952
rect 13464 14940 13492 14980
rect 13538 14968 13544 15020
rect 13596 14968 13602 15020
rect 15010 15017 15016 15020
rect 14972 15011 15016 15017
rect 13740 14980 14780 15008
rect 13740 14940 13768 14980
rect 13464 14912 13768 14940
rect 14001 14943 14059 14949
rect 14001 14909 14013 14943
rect 14047 14909 14059 14943
rect 14001 14903 14059 14909
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14909 14703 14943
rect 14752 14940 14780 14980
rect 14972 14977 14984 15011
rect 14972 14971 15016 14977
rect 15010 14968 15016 14971
rect 15068 14968 15074 15020
rect 15151 15011 15209 15017
rect 15151 14977 15163 15011
rect 15197 15008 15209 15011
rect 15197 14980 16804 15008
rect 15197 14977 15209 14980
rect 15151 14971 15209 14977
rect 15286 14940 15292 14952
rect 14752 14912 15292 14940
rect 14645 14903 14703 14909
rect 12820 14872 12848 14900
rect 14016 14872 14044 14903
rect 12820 14844 14044 14872
rect 14185 14875 14243 14881
rect 14185 14841 14197 14875
rect 14231 14872 14243 14875
rect 14458 14872 14464 14884
rect 14231 14844 14464 14872
rect 14231 14841 14243 14844
rect 14185 14835 14243 14841
rect 14458 14832 14464 14844
rect 14516 14832 14522 14884
rect 14660 14872 14688 14903
rect 15286 14900 15292 14912
rect 15344 14900 15350 14952
rect 15378 14900 15384 14952
rect 15436 14900 15442 14952
rect 14734 14872 14740 14884
rect 14660 14844 14740 14872
rect 14734 14832 14740 14844
rect 14792 14832 14798 14884
rect 16776 14816 16804 14980
rect 17126 14968 17132 15020
rect 17184 14968 17190 15020
rect 17310 14968 17316 15020
rect 17368 15008 17374 15020
rect 18877 15011 18935 15017
rect 18877 15008 18889 15011
rect 17368 14980 18889 15008
rect 17368 14968 17374 14980
rect 18877 14977 18889 14980
rect 18923 15008 18935 15011
rect 19058 15008 19064 15020
rect 18923 14980 19064 15008
rect 18923 14977 18935 14980
rect 18877 14971 18935 14977
rect 19058 14968 19064 14980
rect 19116 14968 19122 15020
rect 19702 15008 19708 15020
rect 19306 14980 19708 15008
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14940 16911 14943
rect 16942 14940 16948 14952
rect 16899 14912 16948 14940
rect 16899 14909 16911 14912
rect 16853 14903 16911 14909
rect 16942 14900 16948 14912
rect 17000 14940 17006 14952
rect 17586 14940 17592 14952
rect 17000 14912 17592 14940
rect 17000 14900 17006 14912
rect 17586 14900 17592 14912
rect 17644 14900 17650 14952
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14940 18751 14943
rect 18782 14940 18788 14952
rect 18739 14912 18788 14940
rect 18739 14909 18751 14912
rect 18693 14903 18751 14909
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 19306 14940 19334 14980
rect 19702 14968 19708 14980
rect 19760 14968 19766 15020
rect 20211 15011 20269 15017
rect 20211 14977 20223 15011
rect 20257 15008 20269 15011
rect 20898 15008 20904 15020
rect 20257 14980 20904 15008
rect 20257 14977 20269 14980
rect 20211 14971 20269 14977
rect 20898 14968 20904 14980
rect 20956 14968 20962 15020
rect 21100 15008 21128 15116
rect 21358 15104 21364 15156
rect 21416 15144 21422 15156
rect 23385 15147 23443 15153
rect 23385 15144 23397 15147
rect 21416 15116 23397 15144
rect 21416 15104 21422 15116
rect 23385 15113 23397 15116
rect 23431 15113 23443 15147
rect 23385 15107 23443 15113
rect 23842 15104 23848 15156
rect 23900 15144 23906 15156
rect 25685 15147 25743 15153
rect 25685 15144 25697 15147
rect 23900 15116 25697 15144
rect 23900 15104 23906 15116
rect 25685 15113 25697 15116
rect 25731 15113 25743 15147
rect 25685 15107 25743 15113
rect 26050 15104 26056 15156
rect 26108 15104 26114 15156
rect 27062 15104 27068 15156
rect 27120 15144 27126 15156
rect 27430 15144 27436 15156
rect 27120 15116 27436 15144
rect 27120 15104 27126 15116
rect 27430 15104 27436 15116
rect 27488 15104 27494 15156
rect 28074 15104 28080 15156
rect 28132 15104 28138 15156
rect 28537 15147 28595 15153
rect 28537 15113 28549 15147
rect 28583 15144 28595 15147
rect 28626 15144 28632 15156
rect 28583 15116 28632 15144
rect 28583 15113 28595 15116
rect 28537 15107 28595 15113
rect 28626 15104 28632 15116
rect 28684 15104 28690 15156
rect 29638 15104 29644 15156
rect 29696 15144 29702 15156
rect 30374 15144 30380 15156
rect 29696 15116 30380 15144
rect 29696 15104 29702 15116
rect 30374 15104 30380 15116
rect 30432 15104 30438 15156
rect 31110 15104 31116 15156
rect 31168 15104 31174 15156
rect 26513 15079 26571 15085
rect 26513 15045 26525 15079
rect 26559 15045 26571 15079
rect 28092 15076 28120 15104
rect 29825 15079 29883 15085
rect 29825 15076 29837 15079
rect 28092 15048 29837 15076
rect 26513 15039 26571 15045
rect 29825 15045 29837 15048
rect 29871 15076 29883 15079
rect 29914 15076 29920 15088
rect 29871 15048 29920 15076
rect 29871 15045 29883 15048
rect 29825 15039 29883 15045
rect 22281 15011 22339 15017
rect 22281 15008 22293 15011
rect 21100 14980 22293 15008
rect 22281 14977 22293 14980
rect 22327 14977 22339 15011
rect 22281 14971 22339 14977
rect 23658 14968 23664 15020
rect 23716 15008 23722 15020
rect 23845 15011 23903 15017
rect 23845 15008 23857 15011
rect 23716 14980 23857 15008
rect 23716 14968 23722 14980
rect 23845 14977 23857 14980
rect 23891 15008 23903 15011
rect 24026 15008 24032 15020
rect 23891 14980 24032 15008
rect 23891 14977 23903 14980
rect 23845 14971 23903 14977
rect 24026 14968 24032 14980
rect 24084 14968 24090 15020
rect 24210 15017 24216 15020
rect 24172 15011 24216 15017
rect 24172 14977 24184 15011
rect 24172 14971 24216 14977
rect 24210 14968 24216 14971
rect 24268 14968 24274 15020
rect 24351 15011 24409 15017
rect 24351 14977 24363 15011
rect 24397 15008 24409 15011
rect 24762 15008 24768 15020
rect 24397 14980 24768 15008
rect 24397 14977 24409 14980
rect 24351 14971 24409 14977
rect 24762 14968 24768 14980
rect 24820 14968 24826 15020
rect 26418 15008 26424 15020
rect 26252 14980 26424 15008
rect 19076 14912 19334 14940
rect 19429 14943 19487 14949
rect 19076 14816 19104 14912
rect 19429 14909 19441 14943
rect 19475 14909 19487 14943
rect 19429 14903 19487 14909
rect 20441 14943 20499 14949
rect 20441 14909 20453 14943
rect 20487 14940 20499 14943
rect 21450 14940 21456 14952
rect 20487 14912 21456 14940
rect 20487 14909 20499 14912
rect 20441 14903 20499 14909
rect 8435 14776 8800 14804
rect 8435 14773 8447 14776
rect 8389 14767 8447 14773
rect 9766 14764 9772 14816
rect 9824 14804 9830 14816
rect 10410 14804 10416 14816
rect 9824 14776 10416 14804
rect 9824 14764 9830 14776
rect 10410 14764 10416 14776
rect 10468 14764 10474 14816
rect 10502 14764 10508 14816
rect 10560 14764 10566 14816
rect 10962 14764 10968 14816
rect 11020 14764 11026 14816
rect 11698 14764 11704 14816
rect 11756 14813 11762 14816
rect 11756 14804 11765 14813
rect 11756 14776 11801 14804
rect 11756 14767 11765 14776
rect 11756 14764 11762 14767
rect 13814 14764 13820 14816
rect 13872 14764 13878 14816
rect 16482 14764 16488 14816
rect 16540 14764 16546 14816
rect 16758 14764 16764 14816
rect 16816 14764 16822 14816
rect 19058 14764 19064 14816
rect 19116 14764 19122 14816
rect 19242 14764 19248 14816
rect 19300 14764 19306 14816
rect 19444 14804 19472 14903
rect 21450 14900 21456 14912
rect 21508 14900 21514 14952
rect 22005 14943 22063 14949
rect 22005 14909 22017 14943
rect 22051 14940 22063 14943
rect 22370 14940 22376 14952
rect 22051 14912 22376 14940
rect 22051 14909 22063 14912
rect 22005 14903 22063 14909
rect 22370 14900 22376 14912
rect 22428 14900 22434 14952
rect 24581 14943 24639 14949
rect 24581 14940 24593 14943
rect 23584 14912 24593 14940
rect 23014 14832 23020 14884
rect 23072 14872 23078 14884
rect 23584 14872 23612 14912
rect 24581 14909 24593 14912
rect 24627 14909 24639 14943
rect 24581 14903 24639 14909
rect 25038 14900 25044 14952
rect 25096 14940 25102 14952
rect 26252 14949 26280 14980
rect 26418 14968 26424 14980
rect 26476 14968 26482 15020
rect 26528 15008 26556 15039
rect 29914 15036 29920 15048
rect 29972 15036 29978 15088
rect 27062 15017 27068 15020
rect 27024 15011 27068 15017
rect 26528 14980 26832 15008
rect 26237 14943 26295 14949
rect 26237 14940 26249 14943
rect 25096 14912 26249 14940
rect 25096 14900 25102 14912
rect 26237 14909 26249 14912
rect 26283 14909 26295 14943
rect 26237 14903 26295 14909
rect 26326 14900 26332 14952
rect 26384 14900 26390 14952
rect 23072 14844 23612 14872
rect 23072 14832 23078 14844
rect 25498 14832 25504 14884
rect 25556 14872 25562 14884
rect 26142 14872 26148 14884
rect 25556 14844 26148 14872
rect 25556 14832 25562 14844
rect 26142 14832 26148 14844
rect 26200 14832 26206 14884
rect 26528 14872 26556 14980
rect 26694 14900 26700 14952
rect 26752 14900 26758 14952
rect 26804 14940 26832 14980
rect 27024 14977 27036 15011
rect 27024 14971 27068 14977
rect 27062 14968 27068 14971
rect 27120 14968 27126 15020
rect 27246 15015 27252 15020
rect 27203 15009 27252 15015
rect 27203 14975 27215 15009
rect 27249 14975 27252 15009
rect 27203 14969 27252 14975
rect 27246 14968 27252 14969
rect 27304 14968 27310 15020
rect 27433 15011 27491 15017
rect 27433 14977 27445 15011
rect 27479 15008 27491 15011
rect 27614 15008 27620 15020
rect 27479 14980 27620 15008
rect 27479 14977 27491 14980
rect 27433 14971 27491 14977
rect 27614 14968 27620 14980
rect 27672 14968 27678 15020
rect 31128 15008 31156 15104
rect 27724 14980 31156 15008
rect 27724 14940 27752 14980
rect 26804 14912 27752 14940
rect 27890 14900 27896 14952
rect 27948 14940 27954 14952
rect 27948 14912 28120 14940
rect 27948 14900 27954 14912
rect 26252 14844 26556 14872
rect 26252 14816 26280 14844
rect 20070 14804 20076 14816
rect 19444 14776 20076 14804
rect 20070 14764 20076 14776
rect 20128 14764 20134 14816
rect 20171 14807 20229 14813
rect 20171 14773 20183 14807
rect 20217 14804 20229 14807
rect 20806 14804 20812 14816
rect 20217 14776 20812 14804
rect 20217 14773 20229 14776
rect 20171 14767 20229 14773
rect 20806 14764 20812 14776
rect 20864 14764 20870 14816
rect 20898 14764 20904 14816
rect 20956 14804 20962 14816
rect 21545 14807 21603 14813
rect 21545 14804 21557 14807
rect 20956 14776 21557 14804
rect 20956 14764 20962 14776
rect 21545 14773 21557 14776
rect 21591 14773 21603 14807
rect 21545 14767 21603 14773
rect 21818 14764 21824 14816
rect 21876 14804 21882 14816
rect 22278 14804 22284 14816
rect 21876 14776 22284 14804
rect 21876 14764 21882 14776
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 26234 14764 26240 14816
rect 26292 14764 26298 14816
rect 26418 14764 26424 14816
rect 26476 14804 26482 14816
rect 26712 14804 26740 14900
rect 28092 14872 28120 14912
rect 28350 14900 28356 14952
rect 28408 14940 28414 14952
rect 29089 14943 29147 14949
rect 29089 14940 29101 14943
rect 28408 14912 29101 14940
rect 28408 14900 28414 14912
rect 29089 14909 29101 14912
rect 29135 14909 29147 14943
rect 29089 14903 29147 14909
rect 29454 14900 29460 14952
rect 29512 14940 29518 14952
rect 29641 14943 29699 14949
rect 29641 14940 29653 14943
rect 29512 14912 29653 14940
rect 29512 14900 29518 14912
rect 29641 14909 29653 14912
rect 29687 14909 29699 14943
rect 29641 14903 29699 14909
rect 30193 14943 30251 14949
rect 30193 14909 30205 14943
rect 30239 14940 30251 14943
rect 30282 14940 30288 14952
rect 30239 14912 30288 14940
rect 30239 14909 30251 14912
rect 30193 14903 30251 14909
rect 30282 14900 30288 14912
rect 30340 14900 30346 14952
rect 30377 14943 30435 14949
rect 30377 14909 30389 14943
rect 30423 14940 30435 14943
rect 30742 14940 30748 14952
rect 30423 14912 30748 14940
rect 30423 14909 30435 14912
rect 30377 14903 30435 14909
rect 28902 14872 28908 14884
rect 28092 14844 28908 14872
rect 28902 14832 28908 14844
rect 28960 14832 28966 14884
rect 28994 14804 29000 14816
rect 26476 14776 29000 14804
rect 26476 14764 26482 14776
rect 28994 14764 29000 14776
rect 29052 14804 29058 14816
rect 29181 14807 29239 14813
rect 29181 14804 29193 14807
rect 29052 14776 29193 14804
rect 29052 14764 29058 14776
rect 29181 14773 29193 14776
rect 29227 14773 29239 14807
rect 29181 14767 29239 14773
rect 30282 14764 30288 14816
rect 30340 14804 30346 14816
rect 30392 14804 30420 14903
rect 30742 14900 30748 14912
rect 30800 14900 30806 14952
rect 30340 14776 30420 14804
rect 30340 14764 30346 14776
rect 30926 14764 30932 14816
rect 30984 14804 30990 14816
rect 30984 14776 31156 14804
rect 30984 14764 30990 14776
rect 552 14714 31072 14736
rect 552 14662 7988 14714
rect 8040 14662 8052 14714
rect 8104 14662 8116 14714
rect 8168 14662 8180 14714
rect 8232 14662 8244 14714
rect 8296 14662 15578 14714
rect 15630 14662 15642 14714
rect 15694 14662 15706 14714
rect 15758 14662 15770 14714
rect 15822 14662 15834 14714
rect 15886 14662 23168 14714
rect 23220 14662 23232 14714
rect 23284 14662 23296 14714
rect 23348 14662 23360 14714
rect 23412 14662 23424 14714
rect 23476 14662 30758 14714
rect 30810 14662 30822 14714
rect 30874 14662 30886 14714
rect 30938 14662 30950 14714
rect 31002 14662 31014 14714
rect 31066 14662 31072 14714
rect 552 14640 31072 14662
rect 934 14560 940 14612
rect 992 14600 998 14612
rect 992 14572 1624 14600
rect 992 14560 998 14572
rect 1210 14492 1216 14544
rect 1268 14492 1274 14544
rect 1394 14492 1400 14544
rect 1452 14492 1458 14544
rect 937 14467 995 14473
rect 937 14433 949 14467
rect 983 14464 995 14467
rect 1412 14464 1440 14492
rect 983 14436 1440 14464
rect 1596 14464 1624 14572
rect 2222 14560 2228 14612
rect 2280 14600 2286 14612
rect 3786 14600 3792 14612
rect 2280 14572 3792 14600
rect 2280 14560 2286 14572
rect 3786 14560 3792 14572
rect 3844 14600 3850 14612
rect 4065 14603 4123 14609
rect 3844 14572 4035 14600
rect 3844 14560 3850 14572
rect 3602 14492 3608 14544
rect 3660 14492 3666 14544
rect 4007 14532 4035 14572
rect 4065 14569 4077 14603
rect 4111 14600 4123 14603
rect 4430 14600 4436 14612
rect 4111 14572 4436 14600
rect 4111 14569 4123 14572
rect 4065 14563 4123 14569
rect 4430 14560 4436 14572
rect 4488 14560 4494 14612
rect 4522 14560 4528 14612
rect 4580 14600 4586 14612
rect 4617 14603 4675 14609
rect 4617 14600 4629 14603
rect 4580 14572 4629 14600
rect 4580 14560 4586 14572
rect 4617 14569 4629 14572
rect 4663 14569 4675 14603
rect 4617 14563 4675 14569
rect 4706 14560 4712 14612
rect 4764 14600 4770 14612
rect 5169 14603 5227 14609
rect 5169 14600 5181 14603
rect 4764 14572 5181 14600
rect 4764 14560 4770 14572
rect 5169 14569 5181 14572
rect 5215 14569 5227 14603
rect 5169 14563 5227 14569
rect 5442 14560 5448 14612
rect 5500 14560 5506 14612
rect 6178 14560 6184 14612
rect 6236 14600 6242 14612
rect 6273 14603 6331 14609
rect 6273 14600 6285 14603
rect 6236 14572 6285 14600
rect 6236 14560 6242 14572
rect 6273 14569 6285 14572
rect 6319 14569 6331 14603
rect 6273 14563 6331 14569
rect 6549 14603 6607 14609
rect 6549 14569 6561 14603
rect 6595 14600 6607 14603
rect 6822 14600 6828 14612
rect 6595 14572 6828 14600
rect 6595 14569 6607 14572
rect 6549 14563 6607 14569
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 7374 14560 7380 14612
rect 7432 14600 7438 14612
rect 8294 14600 8300 14612
rect 7432 14572 8300 14600
rect 7432 14560 7438 14572
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 9125 14603 9183 14609
rect 9125 14569 9137 14603
rect 9171 14600 9183 14603
rect 9306 14600 9312 14612
rect 9171 14572 9312 14600
rect 9171 14569 9183 14572
rect 9125 14563 9183 14569
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 9398 14560 9404 14612
rect 9456 14560 9462 14612
rect 10410 14560 10416 14612
rect 10468 14600 10474 14612
rect 10505 14603 10563 14609
rect 10505 14600 10517 14603
rect 10468 14572 10517 14600
rect 10468 14560 10474 14572
rect 10505 14569 10517 14572
rect 10551 14569 10563 14603
rect 10505 14563 10563 14569
rect 11057 14603 11115 14609
rect 11057 14569 11069 14603
rect 11103 14600 11115 14603
rect 11333 14603 11391 14609
rect 11103 14572 11284 14600
rect 11103 14569 11115 14572
rect 11057 14563 11115 14569
rect 5534 14532 5540 14544
rect 4007 14504 5540 14532
rect 2225 14467 2283 14473
rect 2225 14464 2237 14467
rect 1596 14436 2237 14464
rect 983 14433 995 14436
rect 937 14427 995 14433
rect 2225 14433 2237 14436
rect 2271 14433 2283 14467
rect 3620 14464 3648 14492
rect 4540 14473 4568 14504
rect 3973 14467 4031 14473
rect 3973 14464 3985 14467
rect 3620 14436 3985 14464
rect 2225 14427 2283 14433
rect 3973 14433 3985 14436
rect 4019 14464 4031 14467
rect 4249 14467 4307 14473
rect 4249 14464 4261 14467
rect 4019 14436 4261 14464
rect 4019 14433 4031 14436
rect 3973 14427 4031 14433
rect 4249 14433 4261 14436
rect 4295 14433 4307 14467
rect 4249 14427 4307 14433
rect 4525 14467 4583 14473
rect 4525 14433 4537 14467
rect 4571 14433 4583 14467
rect 4525 14427 4583 14433
rect 4801 14467 4859 14473
rect 4801 14433 4813 14467
rect 4847 14464 4859 14467
rect 4982 14464 4988 14476
rect 4847 14436 4988 14464
rect 4847 14433 4859 14436
rect 4801 14427 4859 14433
rect 1394 14356 1400 14408
rect 1452 14396 1458 14408
rect 1489 14399 1547 14405
rect 1489 14396 1501 14399
rect 1452 14368 1501 14396
rect 1452 14356 1458 14368
rect 1489 14365 1501 14368
rect 1535 14365 1547 14399
rect 1489 14359 1547 14365
rect 1670 14356 1676 14408
rect 1728 14396 1734 14408
rect 1816 14399 1874 14405
rect 1816 14396 1828 14399
rect 1728 14368 1828 14396
rect 1728 14356 1734 14368
rect 1816 14365 1828 14368
rect 1862 14365 1874 14399
rect 1816 14359 1874 14365
rect 1946 14356 1952 14408
rect 2004 14407 2010 14408
rect 2004 14401 2053 14407
rect 2004 14367 2007 14401
rect 2041 14367 2053 14401
rect 2004 14361 2053 14367
rect 2004 14356 2010 14361
rect 2130 14356 2136 14408
rect 2188 14396 2194 14408
rect 2590 14396 2596 14408
rect 2188 14368 2596 14396
rect 2188 14356 2194 14368
rect 2590 14356 2596 14368
rect 2648 14356 2654 14408
rect 4264 14396 4292 14427
rect 4982 14424 4988 14436
rect 5040 14424 5046 14476
rect 5368 14473 5396 14504
rect 5534 14492 5540 14504
rect 5592 14532 5598 14544
rect 5592 14504 6224 14532
rect 5592 14492 5598 14504
rect 5077 14467 5135 14473
rect 5077 14433 5089 14467
rect 5123 14433 5135 14467
rect 5077 14427 5135 14433
rect 5353 14467 5411 14473
rect 5353 14433 5365 14467
rect 5399 14433 5411 14467
rect 5353 14427 5411 14433
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 5902 14464 5908 14476
rect 5675 14436 5908 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 5092 14396 5120 14427
rect 5644 14396 5672 14427
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 6196 14473 6224 14504
rect 6291 14504 6598 14532
rect 6291 14476 6319 14504
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14433 6239 14467
rect 6181 14427 6239 14433
rect 6273 14424 6279 14476
rect 6331 14424 6337 14476
rect 6457 14467 6515 14473
rect 6457 14433 6469 14467
rect 6503 14433 6515 14467
rect 6570 14464 6598 14504
rect 6638 14492 6644 14544
rect 6696 14532 6702 14544
rect 9766 14532 9772 14544
rect 6696 14504 6966 14532
rect 6696 14492 6702 14504
rect 6733 14467 6791 14473
rect 6733 14464 6745 14467
rect 6570 14436 6745 14464
rect 6457 14427 6515 14433
rect 6733 14433 6745 14436
rect 6779 14433 6791 14467
rect 6938 14464 6966 14504
rect 9600 14504 9772 14532
rect 6938 14436 8156 14464
rect 6733 14427 6791 14433
rect 6291 14396 6319 14424
rect 4264 14368 5028 14396
rect 5092 14368 5672 14396
rect 5920 14368 6319 14396
rect 3789 14331 3847 14337
rect 3789 14297 3801 14331
rect 3835 14328 3847 14331
rect 4798 14328 4804 14340
rect 3835 14300 4804 14328
rect 3835 14297 3847 14300
rect 3789 14291 3847 14297
rect 4798 14288 4804 14300
rect 4856 14288 4862 14340
rect 4890 14288 4896 14340
rect 4948 14288 4954 14340
rect 5000 14328 5028 14368
rect 5920 14328 5948 14368
rect 5000 14300 5948 14328
rect 5997 14331 6055 14337
rect 5997 14297 6009 14331
rect 6043 14328 6055 14331
rect 6270 14328 6276 14340
rect 6043 14300 6276 14328
rect 6043 14297 6055 14300
rect 5997 14291 6055 14297
rect 6270 14288 6276 14300
rect 6328 14288 6334 14340
rect 1762 14220 1768 14272
rect 1820 14260 1826 14272
rect 3326 14260 3332 14272
rect 1820 14232 3332 14260
rect 1820 14220 1826 14232
rect 3326 14220 3332 14232
rect 3384 14220 3390 14272
rect 3510 14220 3516 14272
rect 3568 14220 3574 14272
rect 4341 14263 4399 14269
rect 4341 14229 4353 14263
rect 4387 14260 4399 14263
rect 4614 14260 4620 14272
rect 4387 14232 4620 14260
rect 4387 14229 4399 14232
rect 4341 14223 4399 14229
rect 4614 14220 4620 14232
rect 4672 14220 4678 14272
rect 4982 14220 4988 14272
rect 5040 14260 5046 14272
rect 5718 14260 5724 14272
rect 5040 14232 5724 14260
rect 5040 14220 5046 14232
rect 5718 14220 5724 14232
rect 5776 14260 5782 14272
rect 6472 14260 6500 14427
rect 6822 14356 6828 14408
rect 6880 14356 6886 14408
rect 7190 14405 7196 14408
rect 7152 14399 7196 14405
rect 7152 14365 7164 14399
rect 7152 14359 7196 14365
rect 7190 14356 7196 14359
rect 7248 14356 7254 14408
rect 7282 14356 7288 14408
rect 7340 14356 7346 14408
rect 7558 14356 7564 14408
rect 7616 14356 7622 14408
rect 8128 14396 8156 14436
rect 8570 14424 8576 14476
rect 8628 14464 8634 14476
rect 9600 14473 9628 14504
rect 9766 14492 9772 14504
rect 9824 14532 9830 14544
rect 9824 14504 9996 14532
rect 9824 14492 9830 14504
rect 9309 14467 9367 14473
rect 9309 14464 9321 14467
rect 8628 14436 9321 14464
rect 8628 14424 8634 14436
rect 9309 14433 9321 14436
rect 9355 14433 9367 14467
rect 9309 14427 9367 14433
rect 9585 14467 9643 14473
rect 9585 14433 9597 14467
rect 9631 14433 9643 14467
rect 9585 14427 9643 14433
rect 9861 14467 9919 14473
rect 9861 14433 9873 14467
rect 9907 14433 9919 14467
rect 9968 14464 9996 14504
rect 10042 14492 10048 14544
rect 10100 14492 10106 14544
rect 11146 14492 11152 14544
rect 11204 14492 11210 14544
rect 11256 14532 11284 14572
rect 11333 14569 11345 14603
rect 11379 14600 11391 14603
rect 11974 14600 11980 14612
rect 11379 14572 11980 14600
rect 11379 14569 11391 14572
rect 11333 14563 11391 14569
rect 11974 14560 11980 14572
rect 12032 14560 12038 14612
rect 12066 14560 12072 14612
rect 12124 14609 12130 14612
rect 12124 14600 12133 14609
rect 12124 14572 12169 14600
rect 12124 14563 12133 14572
rect 12124 14560 12130 14563
rect 12986 14560 12992 14612
rect 13044 14600 13050 14612
rect 13449 14603 13507 14609
rect 13449 14600 13461 14603
rect 13044 14572 13461 14600
rect 13044 14560 13050 14572
rect 13449 14569 13461 14572
rect 13495 14569 13507 14603
rect 16482 14600 16488 14612
rect 13449 14563 13507 14569
rect 13556 14572 16488 14600
rect 11606 14532 11612 14544
rect 11256 14504 11612 14532
rect 11606 14492 11612 14504
rect 11664 14492 11670 14544
rect 10689 14467 10747 14473
rect 10689 14464 10701 14467
rect 9968 14436 10701 14464
rect 9861 14427 9919 14433
rect 10689 14433 10701 14436
rect 10735 14464 10747 14467
rect 10962 14464 10968 14476
rect 10735 14436 10968 14464
rect 10735 14433 10747 14436
rect 10689 14427 10747 14433
rect 9324 14396 9352 14427
rect 9876 14396 9904 14427
rect 10962 14424 10968 14436
rect 11020 14424 11026 14476
rect 11164 14464 11192 14492
rect 11241 14467 11299 14473
rect 11241 14464 11253 14467
rect 11164 14436 11253 14464
rect 11241 14433 11253 14436
rect 11287 14433 11299 14467
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 11241 14427 11299 14433
rect 11348 14436 11529 14464
rect 11348 14408 11376 14436
rect 11517 14433 11529 14436
rect 11563 14433 11575 14467
rect 13556 14464 13584 14572
rect 16482 14560 16488 14572
rect 16540 14560 16546 14612
rect 16758 14560 16764 14612
rect 16816 14600 16822 14612
rect 18509 14603 18567 14609
rect 18509 14600 18521 14603
rect 16816 14572 18521 14600
rect 16816 14560 16822 14572
rect 18509 14569 18521 14572
rect 18555 14569 18567 14603
rect 18509 14563 18567 14569
rect 19242 14560 19248 14612
rect 19300 14560 19306 14612
rect 20806 14560 20812 14612
rect 20864 14600 20870 14612
rect 22103 14603 22161 14609
rect 22103 14600 22115 14603
rect 20864 14572 22115 14600
rect 20864 14560 20870 14572
rect 22103 14569 22115 14572
rect 22149 14569 22161 14603
rect 22103 14563 22161 14569
rect 22278 14560 22284 14612
rect 22336 14600 22342 14612
rect 25685 14603 25743 14609
rect 25685 14600 25697 14603
rect 22336 14572 25697 14600
rect 22336 14560 22342 14572
rect 25685 14569 25697 14572
rect 25731 14569 25743 14603
rect 25685 14563 25743 14569
rect 26142 14560 26148 14612
rect 26200 14600 26206 14612
rect 26200 14572 28120 14600
rect 26200 14560 26206 14572
rect 15286 14492 15292 14544
rect 15344 14532 15350 14544
rect 15933 14535 15991 14541
rect 15933 14532 15945 14535
rect 15344 14504 15945 14532
rect 15344 14492 15350 14504
rect 15933 14501 15945 14504
rect 15979 14501 15991 14535
rect 15933 14495 15991 14501
rect 18322 14492 18328 14544
rect 18380 14532 18386 14544
rect 19061 14535 19119 14541
rect 19061 14532 19073 14535
rect 18380 14504 19073 14532
rect 18380 14492 18386 14504
rect 19061 14501 19073 14504
rect 19107 14532 19119 14535
rect 19150 14532 19156 14544
rect 19107 14504 19156 14532
rect 19107 14501 19119 14504
rect 19061 14495 19119 14501
rect 19150 14492 19156 14504
rect 19208 14492 19214 14544
rect 11517 14427 11575 14433
rect 12268 14436 13584 14464
rect 13817 14467 13875 14473
rect 8128 14368 9204 14396
rect 9324 14368 9904 14396
rect 6638 14260 6644 14272
rect 5776 14232 6644 14260
rect 5776 14220 5782 14232
rect 6638 14220 6644 14232
rect 6696 14260 6702 14272
rect 7006 14260 7012 14272
rect 6696 14232 7012 14260
rect 6696 14220 6702 14232
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 8202 14220 8208 14272
rect 8260 14260 8266 14272
rect 8754 14260 8760 14272
rect 8260 14232 8760 14260
rect 8260 14220 8266 14232
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 8846 14220 8852 14272
rect 8904 14220 8910 14272
rect 9176 14260 9204 14368
rect 9677 14331 9735 14337
rect 9677 14328 9689 14331
rect 9508 14300 9689 14328
rect 9508 14260 9536 14300
rect 9677 14297 9689 14300
rect 9723 14297 9735 14331
rect 9876 14328 9904 14368
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 10367 14368 11284 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 11256 14340 11284 14368
rect 11330 14356 11336 14408
rect 11388 14356 11394 14408
rect 11609 14399 11667 14405
rect 11609 14365 11621 14399
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 12115 14399 12173 14405
rect 12115 14365 12127 14399
rect 12161 14396 12173 14399
rect 12268 14396 12296 14436
rect 13817 14433 13829 14467
rect 13863 14464 13875 14467
rect 13906 14464 13912 14476
rect 13863 14436 13912 14464
rect 13863 14433 13875 14436
rect 13817 14427 13875 14433
rect 13906 14424 13912 14436
rect 13964 14424 13970 14476
rect 15194 14464 15200 14476
rect 14016 14436 15200 14464
rect 14016 14408 14044 14436
rect 15194 14424 15200 14436
rect 15252 14424 15258 14476
rect 16114 14424 16120 14476
rect 16172 14424 16178 14476
rect 16758 14424 16764 14476
rect 16816 14464 16822 14476
rect 16996 14467 17054 14473
rect 16996 14464 17008 14467
rect 16816 14436 17008 14464
rect 16816 14424 16822 14436
rect 16996 14433 17008 14436
rect 17042 14464 17054 14467
rect 17310 14464 17316 14476
rect 17042 14436 17316 14464
rect 17042 14433 17054 14436
rect 16996 14427 17054 14433
rect 17310 14424 17316 14436
rect 17368 14424 17374 14476
rect 17405 14467 17463 14473
rect 17405 14433 17417 14467
rect 17451 14464 17463 14467
rect 19260 14464 19288 14560
rect 21085 14535 21143 14541
rect 21085 14501 21097 14535
rect 21131 14532 21143 14535
rect 21634 14532 21640 14544
rect 21131 14504 21640 14532
rect 21131 14501 21143 14504
rect 21085 14495 21143 14501
rect 21634 14492 21640 14504
rect 21692 14492 21698 14544
rect 23750 14492 23756 14544
rect 23808 14492 23814 14544
rect 26786 14532 26792 14544
rect 26712 14504 26792 14532
rect 17451 14436 19288 14464
rect 19352 14436 21036 14464
rect 17451 14433 17463 14436
rect 17405 14427 17463 14433
rect 12161 14368 12296 14396
rect 12161 14365 12173 14368
rect 12115 14359 12173 14365
rect 11146 14328 11152 14340
rect 9876 14300 11152 14328
rect 9677 14291 9735 14297
rect 11146 14288 11152 14300
rect 11204 14288 11210 14340
rect 11238 14288 11244 14340
rect 11296 14328 11302 14340
rect 11624 14328 11652 14359
rect 12342 14356 12348 14408
rect 12400 14356 12406 14408
rect 13446 14356 13452 14408
rect 13504 14356 13510 14408
rect 13998 14356 14004 14408
rect 14056 14356 14062 14408
rect 14182 14405 14188 14408
rect 14144 14399 14188 14405
rect 14144 14365 14156 14399
rect 14144 14359 14188 14365
rect 14182 14356 14188 14359
rect 14240 14356 14246 14408
rect 14323 14399 14381 14405
rect 14323 14365 14335 14399
rect 14369 14396 14381 14399
rect 14458 14396 14464 14408
rect 14369 14368 14464 14396
rect 14369 14365 14381 14368
rect 14323 14359 14381 14365
rect 14458 14356 14464 14368
rect 14516 14356 14522 14408
rect 14550 14356 14556 14408
rect 14608 14356 14614 14408
rect 16666 14356 16672 14408
rect 16724 14356 16730 14408
rect 17175 14399 17233 14405
rect 17175 14365 17187 14399
rect 17221 14396 17233 14399
rect 19352 14396 19380 14436
rect 17221 14368 19380 14396
rect 19429 14399 19487 14405
rect 17221 14365 17233 14368
rect 17175 14359 17233 14365
rect 19429 14365 19441 14399
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 11296 14300 11652 14328
rect 11296 14288 11302 14300
rect 9176 14232 9536 14260
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 13464 14260 13492 14356
rect 15212 14300 16436 14328
rect 9916 14232 13492 14260
rect 9916 14220 9922 14232
rect 14090 14220 14096 14272
rect 14148 14260 14154 14272
rect 14642 14260 14648 14272
rect 14148 14232 14648 14260
rect 14148 14220 14154 14232
rect 14642 14220 14648 14232
rect 14700 14220 14706 14272
rect 14734 14220 14740 14272
rect 14792 14260 14798 14272
rect 15212 14260 15240 14300
rect 14792 14232 15240 14260
rect 14792 14220 14798 14232
rect 16298 14220 16304 14272
rect 16356 14220 16362 14272
rect 16408 14260 16436 14300
rect 18966 14288 18972 14340
rect 19024 14288 19030 14340
rect 19150 14288 19156 14340
rect 19208 14328 19214 14340
rect 19444 14328 19472 14359
rect 19702 14356 19708 14408
rect 19760 14356 19766 14408
rect 19208 14300 19472 14328
rect 21008 14328 21036 14436
rect 21266 14424 21272 14476
rect 21324 14424 21330 14476
rect 22830 14464 22836 14476
rect 22204 14436 22836 14464
rect 21284 14396 21312 14424
rect 21637 14399 21695 14405
rect 21637 14396 21649 14399
rect 21284 14368 21649 14396
rect 21637 14365 21649 14368
rect 21683 14365 21695 14399
rect 21637 14359 21695 14365
rect 22116 14399 22174 14405
rect 22116 14365 22128 14399
rect 22162 14396 22174 14399
rect 22204 14396 22232 14436
rect 22830 14424 22836 14436
rect 22888 14424 22894 14476
rect 23658 14424 23664 14476
rect 23716 14464 23722 14476
rect 24210 14473 24216 14476
rect 23845 14467 23903 14473
rect 23845 14464 23857 14467
rect 23716 14436 23857 14464
rect 23716 14424 23722 14436
rect 23845 14433 23857 14436
rect 23891 14433 23903 14467
rect 23845 14427 23903 14433
rect 24172 14467 24216 14473
rect 24172 14433 24184 14467
rect 24172 14427 24216 14433
rect 24210 14424 24216 14427
rect 24268 14424 24274 14476
rect 24670 14424 24676 14476
rect 24728 14464 24734 14476
rect 26234 14473 26240 14476
rect 26229 14464 26240 14473
rect 24728 14436 26240 14464
rect 24728 14424 24734 14436
rect 26229 14427 26240 14436
rect 26234 14424 26240 14427
rect 26292 14424 26298 14476
rect 26712 14473 26740 14504
rect 26786 14492 26792 14504
rect 26844 14492 26850 14544
rect 26973 14535 27031 14541
rect 26973 14501 26985 14535
rect 27019 14532 27031 14535
rect 27062 14532 27068 14544
rect 27019 14504 27068 14532
rect 27019 14501 27031 14504
rect 26973 14495 27031 14501
rect 27062 14492 27068 14504
rect 27120 14492 27126 14544
rect 27246 14492 27252 14544
rect 27304 14532 27310 14544
rect 27341 14535 27399 14541
rect 27341 14532 27353 14535
rect 27304 14504 27353 14532
rect 27304 14492 27310 14504
rect 27341 14501 27353 14504
rect 27387 14501 27399 14535
rect 27341 14495 27399 14501
rect 27709 14535 27767 14541
rect 27709 14501 27721 14535
rect 27755 14532 27767 14535
rect 27890 14532 27896 14544
rect 27755 14504 27896 14532
rect 27755 14501 27767 14504
rect 27709 14495 27767 14501
rect 27890 14492 27896 14504
rect 27948 14492 27954 14544
rect 26605 14467 26663 14473
rect 26605 14433 26617 14467
rect 26651 14433 26663 14467
rect 26605 14427 26663 14433
rect 26707 14467 26765 14473
rect 26707 14433 26719 14467
rect 26753 14433 26765 14467
rect 26707 14427 26765 14433
rect 24341 14417 24399 14423
rect 24341 14408 24353 14417
rect 22162 14368 22232 14396
rect 22162 14365 22174 14368
rect 22116 14359 22174 14365
rect 22278 14356 22284 14408
rect 22336 14396 22342 14408
rect 22373 14399 22431 14405
rect 22373 14396 22385 14399
rect 22336 14368 22385 14396
rect 22336 14356 22342 14368
rect 22373 14365 22385 14368
rect 22419 14365 22431 14399
rect 22373 14359 22431 14365
rect 24302 14356 24308 14408
rect 24387 14383 24399 14417
rect 24360 14377 24399 14383
rect 24360 14368 24394 14377
rect 24360 14356 24366 14368
rect 24486 14356 24492 14408
rect 24544 14396 24550 14408
rect 24581 14399 24639 14405
rect 24581 14396 24593 14399
rect 24544 14368 24593 14396
rect 24544 14356 24550 14368
rect 24581 14365 24593 14368
rect 24627 14365 24639 14399
rect 24581 14359 24639 14365
rect 24946 14356 24952 14408
rect 25004 14396 25010 14408
rect 26620 14396 26648 14427
rect 27982 14424 27988 14476
rect 28040 14424 28046 14476
rect 28092 14464 28120 14572
rect 28258 14560 28264 14612
rect 28316 14600 28322 14612
rect 28451 14603 28509 14609
rect 28451 14600 28463 14603
rect 28316 14572 28463 14600
rect 28316 14560 28322 14572
rect 28451 14569 28463 14572
rect 28497 14569 28509 14603
rect 28451 14563 28509 14569
rect 29178 14560 29184 14612
rect 29236 14600 29242 14612
rect 29825 14603 29883 14609
rect 29825 14600 29837 14603
rect 29236 14572 29837 14600
rect 29236 14560 29242 14572
rect 29825 14569 29837 14572
rect 29871 14569 29883 14603
rect 29825 14563 29883 14569
rect 29914 14560 29920 14612
rect 29972 14560 29978 14612
rect 30742 14560 30748 14612
rect 30800 14600 30806 14612
rect 31128 14600 31156 14776
rect 30800 14572 31156 14600
rect 30800 14560 30806 14572
rect 29454 14492 29460 14544
rect 29512 14532 29518 14544
rect 29932 14532 29960 14560
rect 29512 14504 30420 14532
rect 29512 14492 29518 14504
rect 30392 14473 30420 14504
rect 30377 14467 30435 14473
rect 28092 14436 30052 14464
rect 25004 14368 26648 14396
rect 25004 14356 25010 14368
rect 26620 14328 26648 14368
rect 28350 14356 28356 14408
rect 28408 14396 28414 14408
rect 28448 14399 28506 14405
rect 28448 14396 28460 14399
rect 28408 14368 28460 14396
rect 28408 14356 28414 14368
rect 28448 14365 28460 14368
rect 28494 14365 28506 14399
rect 28448 14359 28506 14365
rect 28721 14399 28779 14405
rect 28721 14365 28733 14399
rect 28767 14396 28779 14399
rect 29914 14396 29920 14408
rect 28767 14368 29920 14396
rect 28767 14365 28779 14368
rect 28721 14359 28779 14365
rect 29914 14356 29920 14368
rect 29972 14356 29978 14408
rect 27890 14328 27896 14340
rect 21008 14300 21670 14328
rect 26620 14300 27896 14328
rect 19208 14288 19214 14300
rect 18984 14260 19012 14288
rect 16408 14232 19012 14260
rect 19444 14260 19472 14300
rect 21453 14263 21511 14269
rect 21453 14260 21465 14263
rect 19444 14232 21465 14260
rect 21453 14229 21465 14232
rect 21499 14260 21511 14263
rect 21542 14260 21548 14272
rect 21499 14232 21548 14260
rect 21499 14229 21511 14232
rect 21453 14223 21511 14229
rect 21542 14220 21548 14232
rect 21600 14220 21606 14272
rect 21642 14260 21670 14300
rect 27890 14288 27896 14300
rect 27948 14288 27954 14340
rect 30024 14328 30052 14436
rect 30377 14433 30389 14467
rect 30423 14433 30435 14467
rect 30377 14427 30435 14433
rect 30193 14331 30251 14337
rect 30193 14328 30205 14331
rect 30024 14300 30205 14328
rect 30193 14297 30205 14300
rect 30239 14297 30251 14331
rect 30193 14291 30251 14297
rect 22738 14260 22744 14272
rect 21642 14232 22744 14260
rect 22738 14220 22744 14232
rect 22796 14220 22802 14272
rect 23290 14220 23296 14272
rect 23348 14260 23354 14272
rect 25038 14260 25044 14272
rect 23348 14232 25044 14260
rect 23348 14220 23354 14232
rect 25038 14220 25044 14232
rect 25096 14220 25102 14272
rect 26050 14220 26056 14272
rect 26108 14220 26114 14272
rect 26421 14263 26479 14269
rect 26421 14229 26433 14263
rect 26467 14260 26479 14263
rect 26694 14260 26700 14272
rect 26467 14232 26700 14260
rect 26467 14229 26479 14232
rect 26421 14223 26479 14229
rect 26694 14220 26700 14232
rect 26752 14220 26758 14272
rect 26786 14220 26792 14272
rect 26844 14260 26850 14272
rect 27062 14260 27068 14272
rect 26844 14232 27068 14260
rect 26844 14220 26850 14232
rect 27062 14220 27068 14232
rect 27120 14220 27126 14272
rect 27154 14220 27160 14272
rect 27212 14260 27218 14272
rect 27614 14260 27620 14272
rect 27212 14232 27620 14260
rect 27212 14220 27218 14232
rect 27614 14220 27620 14232
rect 27672 14220 27678 14272
rect 552 14170 30912 14192
rect 552 14118 4193 14170
rect 4245 14118 4257 14170
rect 4309 14118 4321 14170
rect 4373 14118 4385 14170
rect 4437 14118 4449 14170
rect 4501 14118 11783 14170
rect 11835 14118 11847 14170
rect 11899 14118 11911 14170
rect 11963 14118 11975 14170
rect 12027 14118 12039 14170
rect 12091 14118 19373 14170
rect 19425 14118 19437 14170
rect 19489 14118 19501 14170
rect 19553 14118 19565 14170
rect 19617 14118 19629 14170
rect 19681 14118 26963 14170
rect 27015 14118 27027 14170
rect 27079 14118 27091 14170
rect 27143 14118 27155 14170
rect 27207 14118 27219 14170
rect 27271 14118 30912 14170
rect 552 14096 30912 14118
rect 3510 14016 3516 14068
rect 3568 14056 3574 14068
rect 4154 14056 4160 14068
rect 3568 14028 4160 14056
rect 3568 14016 3574 14028
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 5905 14059 5963 14065
rect 5905 14025 5917 14059
rect 5951 14056 5963 14059
rect 7282 14056 7288 14068
rect 5951 14028 7288 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 9858 14056 9864 14068
rect 8220 14028 9864 14056
rect 750 13880 756 13932
rect 808 13920 814 13932
rect 937 13923 995 13929
rect 937 13920 949 13923
rect 808 13892 949 13920
rect 808 13880 814 13892
rect 937 13889 949 13892
rect 983 13889 995 13923
rect 937 13883 995 13889
rect 1443 13923 1501 13929
rect 1443 13889 1455 13923
rect 1489 13920 1501 13923
rect 2774 13920 2780 13932
rect 1489 13892 2780 13920
rect 1489 13889 1501 13892
rect 1443 13883 1501 13889
rect 2774 13880 2780 13892
rect 2832 13880 2838 13932
rect 3881 13923 3939 13929
rect 3436 13918 3832 13920
rect 3881 13918 3893 13923
rect 3436 13892 3893 13918
rect 3436 13864 3464 13892
rect 3804 13890 3893 13892
rect 3881 13889 3893 13890
rect 3927 13889 3939 13923
rect 3881 13883 3939 13889
rect 4154 13880 4160 13932
rect 4212 13920 4218 13932
rect 4344 13923 4402 13929
rect 4344 13920 4356 13923
rect 4212 13892 4356 13920
rect 4212 13880 4218 13892
rect 4344 13889 4356 13892
rect 4390 13889 4402 13923
rect 4344 13883 4402 13889
rect 5626 13880 5632 13932
rect 5684 13920 5690 13932
rect 5684 13892 6132 13920
rect 5684 13880 5690 13892
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 2590 13852 2596 13864
rect 1719 13824 2596 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 3050 13812 3056 13864
rect 3108 13812 3114 13864
rect 3418 13812 3424 13864
rect 3476 13812 3482 13864
rect 3510 13812 3516 13864
rect 3568 13812 3574 13864
rect 4617 13855 4675 13861
rect 3789 13831 3847 13837
rect 3789 13797 3801 13831
rect 3835 13797 3847 13831
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 5810 13852 5816 13864
rect 4663 13824 5816 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 5810 13812 5816 13824
rect 5868 13812 5874 13864
rect 6104 13861 6132 13892
rect 6270 13880 6276 13932
rect 6328 13880 6334 13932
rect 6454 13929 6460 13932
rect 6416 13923 6460 13929
rect 6416 13889 6428 13923
rect 6416 13883 6460 13889
rect 6454 13880 6460 13883
rect 6512 13880 6518 13932
rect 6595 13923 6653 13929
rect 6595 13889 6607 13923
rect 6641 13920 6653 13923
rect 8220 13920 8248 14028
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 9950 14016 9956 14068
rect 10008 14056 10014 14068
rect 11606 14056 11612 14068
rect 10008 14028 11612 14056
rect 10008 14016 10014 14028
rect 11606 14016 11612 14028
rect 11664 14016 11670 14068
rect 12342 14016 12348 14068
rect 12400 14056 12406 14068
rect 12437 14059 12495 14065
rect 12437 14056 12449 14059
rect 12400 14028 12449 14056
rect 12400 14016 12406 14028
rect 12437 14025 12449 14028
rect 12483 14025 12495 14059
rect 12437 14019 12495 14025
rect 12526 14016 12532 14068
rect 12584 14056 12590 14068
rect 12989 14059 13047 14065
rect 12989 14056 13001 14059
rect 12584 14028 13001 14056
rect 12584 14016 12590 14028
rect 12989 14025 13001 14028
rect 13035 14025 13047 14059
rect 12989 14019 13047 14025
rect 13262 14016 13268 14068
rect 13320 14016 13326 14068
rect 13909 14059 13967 14065
rect 13909 14025 13921 14059
rect 13955 14056 13967 14059
rect 14550 14056 14556 14068
rect 13955 14028 14556 14056
rect 13955 14025 13967 14028
rect 13909 14019 13967 14025
rect 14550 14016 14556 14028
rect 14608 14016 14614 14068
rect 16850 14056 16856 14068
rect 15856 14028 16856 14056
rect 8386 13948 8392 14000
rect 8444 13988 8450 14000
rect 8941 13991 8999 13997
rect 8444 13960 8708 13988
rect 8444 13948 8450 13960
rect 8573 13923 8631 13929
rect 8573 13920 8585 13923
rect 6641 13892 8248 13920
rect 8312 13892 8585 13920
rect 6641 13889 6653 13892
rect 6595 13883 6653 13889
rect 6089 13855 6147 13861
rect 6089 13821 6101 13855
rect 6135 13821 6147 13855
rect 6288 13852 6316 13880
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6288 13824 6837 13852
rect 6089 13815 6147 13821
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 8202 13852 8208 13864
rect 6972 13824 8208 13852
rect 6972 13812 6978 13824
rect 8202 13812 8208 13824
rect 8260 13852 8266 13864
rect 8312 13852 8340 13892
rect 8573 13889 8585 13892
rect 8619 13889 8631 13923
rect 8573 13883 8631 13889
rect 8260 13824 8340 13852
rect 8260 13812 8266 13824
rect 8386 13812 8392 13864
rect 8444 13812 8450 13864
rect 8680 13852 8708 13960
rect 8941 13957 8953 13991
rect 8987 13988 8999 13991
rect 9122 13988 9128 14000
rect 8987 13960 9128 13988
rect 8987 13957 8999 13960
rect 8941 13951 8999 13957
rect 9122 13948 9128 13960
rect 9180 13948 9186 14000
rect 11146 13948 11152 14000
rect 11204 13988 11210 14000
rect 11204 13960 12204 13988
rect 11204 13948 11210 13960
rect 10140 13923 10198 13929
rect 10140 13920 10152 13923
rect 9416 13892 10152 13920
rect 9416 13864 9444 13892
rect 10140 13889 10152 13892
rect 10186 13889 10198 13923
rect 11330 13920 11336 13932
rect 10140 13883 10198 13889
rect 10520 13892 11336 13920
rect 10520 13864 10548 13892
rect 11330 13880 11336 13892
rect 11388 13880 11394 13932
rect 11698 13880 11704 13932
rect 11756 13920 11762 13932
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 11756 13892 12081 13920
rect 11756 13880 11762 13892
rect 12069 13889 12081 13892
rect 12115 13889 12127 13923
rect 12176 13920 12204 13960
rect 12710 13948 12716 14000
rect 12768 13948 12774 14000
rect 13280 13920 13308 14016
rect 13633 13991 13691 13997
rect 13633 13957 13645 13991
rect 13679 13988 13691 13991
rect 13998 13988 14004 14000
rect 13679 13960 14004 13988
rect 13679 13957 13691 13960
rect 13633 13951 13691 13957
rect 13998 13948 14004 13960
rect 14056 13948 14062 14000
rect 13446 13920 13452 13932
rect 12176 13892 12756 13920
rect 12069 13883 12127 13889
rect 9125 13855 9183 13861
rect 9125 13852 9137 13855
rect 8680 13824 9137 13852
rect 9125 13821 9137 13824
rect 9171 13852 9183 13855
rect 9306 13852 9312 13864
rect 9171 13824 9312 13852
rect 9171 13821 9183 13824
rect 9125 13815 9183 13821
rect 9306 13812 9312 13824
rect 9364 13812 9370 13864
rect 9398 13812 9404 13864
rect 9456 13812 9462 13864
rect 9490 13812 9496 13864
rect 9548 13852 9554 13864
rect 10042 13861 10048 13864
rect 9677 13855 9735 13861
rect 9677 13852 9689 13855
rect 9548 13824 9689 13852
rect 9548 13812 9554 13824
rect 9677 13821 9689 13824
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 10004 13855 10048 13861
rect 10004 13821 10016 13855
rect 10004 13815 10048 13821
rect 10042 13812 10048 13815
rect 10100 13812 10106 13864
rect 10410 13812 10416 13864
rect 10468 13812 10474 13864
rect 10502 13812 10508 13864
rect 10560 13812 10566 13864
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 11882 13852 11888 13864
rect 11112 13824 11888 13852
rect 11112 13812 11118 13824
rect 11882 13812 11888 13824
rect 11940 13812 11946 13864
rect 12621 13855 12679 13861
rect 12621 13821 12633 13855
rect 12667 13821 12679 13855
rect 12621 13815 12679 13821
rect 3789 13791 3847 13797
rect 3804 13728 3832 13791
rect 5534 13744 5540 13796
rect 5592 13744 5598 13796
rect 7834 13744 7840 13796
rect 7892 13784 7898 13796
rect 9217 13787 9275 13793
rect 9217 13784 9229 13787
rect 7892 13756 9229 13784
rect 7892 13744 7898 13756
rect 9217 13753 9229 13756
rect 9263 13753 9275 13787
rect 9217 13747 9275 13753
rect 11422 13744 11428 13796
rect 11480 13744 11486 13796
rect 11790 13744 11796 13796
rect 11848 13744 11854 13796
rect 1403 13719 1461 13725
rect 1403 13685 1415 13719
rect 1449 13716 1461 13719
rect 1946 13716 1952 13728
rect 1449 13688 1952 13716
rect 1449 13685 1461 13688
rect 1403 13679 1461 13685
rect 1946 13676 1952 13688
rect 2004 13676 2010 13728
rect 3326 13676 3332 13728
rect 3384 13676 3390 13728
rect 3605 13719 3663 13725
rect 3605 13685 3617 13719
rect 3651 13716 3663 13719
rect 3694 13716 3700 13728
rect 3651 13688 3700 13716
rect 3651 13685 3663 13688
rect 3605 13679 3663 13685
rect 3694 13676 3700 13688
rect 3752 13676 3758 13728
rect 3786 13676 3792 13728
rect 3844 13676 3850 13728
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 4347 13719 4405 13725
rect 4347 13716 4359 13719
rect 4028 13688 4359 13716
rect 4028 13676 4034 13688
rect 4347 13685 4359 13688
rect 4393 13716 4405 13719
rect 4522 13716 4528 13728
rect 4393 13688 4528 13716
rect 4393 13685 4405 13688
rect 4347 13679 4405 13685
rect 4522 13676 4528 13688
rect 4580 13676 4586 13728
rect 5552 13716 5580 13744
rect 6454 13716 6460 13728
rect 5552 13688 6460 13716
rect 6454 13676 6460 13688
rect 6512 13676 6518 13728
rect 6638 13676 6644 13728
rect 6696 13716 6702 13728
rect 7929 13719 7987 13725
rect 7929 13716 7941 13719
rect 6696 13688 7941 13716
rect 6696 13676 6702 13688
rect 7929 13685 7941 13688
rect 7975 13685 7987 13719
rect 7929 13679 7987 13685
rect 8662 13676 8668 13728
rect 8720 13716 8726 13728
rect 11440 13716 11468 13744
rect 12250 13716 12256 13728
rect 8720 13688 12256 13716
rect 8720 13676 8726 13688
rect 12250 13676 12256 13688
rect 12308 13716 12314 13728
rect 12636 13716 12664 13815
rect 12728 13784 12756 13892
rect 12912 13892 13452 13920
rect 12912 13861 12940 13892
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 13722 13880 13728 13932
rect 13780 13880 13786 13932
rect 13906 13880 13912 13932
rect 13964 13880 13970 13932
rect 14648 13921 14706 13927
rect 14108 13892 14596 13920
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13852 13231 13855
rect 13740 13852 13768 13880
rect 13219 13824 13768 13852
rect 13817 13855 13875 13861
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 13817 13821 13829 13855
rect 13863 13821 13875 13855
rect 13817 13815 13875 13821
rect 13188 13784 13216 13815
rect 12728 13756 13216 13784
rect 13722 13744 13728 13796
rect 13780 13784 13786 13796
rect 13832 13784 13860 13815
rect 13780 13756 13860 13784
rect 13924 13784 13952 13880
rect 14108 13861 14136 13892
rect 14093 13855 14151 13861
rect 14093 13821 14105 13855
rect 14139 13821 14151 13855
rect 14093 13815 14151 13821
rect 14185 13855 14243 13861
rect 14185 13821 14197 13855
rect 14231 13821 14243 13855
rect 14568 13852 14596 13892
rect 14648 13887 14660 13921
rect 14694 13920 14706 13921
rect 14734 13920 14740 13932
rect 14694 13892 14740 13920
rect 14694 13887 14706 13892
rect 14648 13881 14706 13887
rect 14734 13880 14740 13892
rect 14792 13880 14798 13932
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13920 14979 13923
rect 15856 13920 15884 14028
rect 16850 14016 16856 14028
rect 16908 14016 16914 14068
rect 18230 14016 18236 14068
rect 18288 14016 18294 14068
rect 19058 14016 19064 14068
rect 19116 14016 19122 14068
rect 21910 14056 21916 14068
rect 19996 14028 21916 14056
rect 16022 13948 16028 14000
rect 16080 13948 16086 14000
rect 18690 13948 18696 14000
rect 18748 13988 18754 14000
rect 19521 13991 19579 13997
rect 19521 13988 19533 13991
rect 18748 13960 19533 13988
rect 18748 13948 18754 13960
rect 19521 13957 19533 13960
rect 19567 13957 19579 13991
rect 19521 13951 19579 13957
rect 16758 13929 16764 13932
rect 14967 13892 15884 13920
rect 16720 13923 16764 13929
rect 14967 13889 14979 13892
rect 14921 13883 14979 13889
rect 16720 13889 16732 13923
rect 16720 13883 16764 13889
rect 16758 13880 16764 13883
rect 16816 13880 16822 13932
rect 16899 13923 16957 13929
rect 16899 13889 16911 13923
rect 16945 13920 16957 13923
rect 19996 13920 20024 14028
rect 21910 14016 21916 14028
rect 21968 14016 21974 14068
rect 22465 14059 22523 14065
rect 22465 14025 22477 14059
rect 22511 14056 22523 14059
rect 24854 14056 24860 14068
rect 22511 14028 24860 14056
rect 22511 14025 22523 14028
rect 22465 14019 22523 14025
rect 24854 14016 24860 14028
rect 24912 14016 24918 14068
rect 26050 14016 26056 14068
rect 26108 14016 26114 14068
rect 26510 14016 26516 14068
rect 26568 14016 26574 14068
rect 26602 14016 26608 14068
rect 26660 14056 26666 14068
rect 27430 14056 27436 14068
rect 26660 14028 27436 14056
rect 26660 14016 26666 14028
rect 27430 14016 27436 14028
rect 27488 14016 27494 14068
rect 27522 14016 27528 14068
rect 27580 14056 27586 14068
rect 28997 14059 29055 14065
rect 28997 14056 29009 14059
rect 27580 14028 29009 14056
rect 27580 14016 27586 14028
rect 28997 14025 29009 14028
rect 29043 14025 29055 14059
rect 28997 14019 29055 14025
rect 29086 14016 29092 14068
rect 29144 14056 29150 14068
rect 29273 14059 29331 14065
rect 29273 14056 29285 14059
rect 29144 14028 29285 14056
rect 29144 14016 29150 14028
rect 29273 14025 29285 14028
rect 29319 14025 29331 14059
rect 29273 14019 29331 14025
rect 29546 14016 29552 14068
rect 29604 14016 29610 14068
rect 29822 14016 29828 14068
rect 29880 14016 29886 14068
rect 30285 14059 30343 14065
rect 30285 14025 30297 14059
rect 30331 14056 30343 14059
rect 31110 14056 31116 14068
rect 30331 14028 31116 14056
rect 30331 14025 30343 14028
rect 30285 14019 30343 14025
rect 31110 14016 31116 14028
rect 31168 14016 31174 14068
rect 21450 13948 21456 14000
rect 21508 13988 21514 14000
rect 22189 13991 22247 13997
rect 22189 13988 22201 13991
rect 21508 13960 22201 13988
rect 21508 13948 21514 13960
rect 22189 13957 22201 13960
rect 22235 13957 22247 13991
rect 22189 13951 22247 13957
rect 22741 13991 22799 13997
rect 22741 13957 22753 13991
rect 22787 13988 22799 13991
rect 24486 13988 24492 14000
rect 22787 13960 24492 13988
rect 22787 13957 22799 13960
rect 22741 13951 22799 13957
rect 24486 13948 24492 13960
rect 24544 13948 24550 14000
rect 20530 13927 20536 13932
rect 16945 13892 20024 13920
rect 20487 13921 20536 13927
rect 16945 13889 16957 13892
rect 16899 13883 16957 13889
rect 20487 13887 20499 13921
rect 20533 13887 20536 13921
rect 20487 13881 20536 13887
rect 20530 13880 20536 13881
rect 20588 13880 20594 13932
rect 22097 13923 22155 13929
rect 22097 13889 22109 13923
rect 22143 13920 22155 13923
rect 24210 13920 24216 13932
rect 22143 13892 24216 13920
rect 22143 13889 22155 13892
rect 22097 13883 22155 13889
rect 24210 13880 24216 13892
rect 24268 13880 24274 13932
rect 24394 13920 24400 13932
rect 24320 13892 24400 13920
rect 14826 13852 14832 13864
rect 14568 13824 14832 13852
rect 14185 13815 14243 13821
rect 14200 13784 14228 13815
rect 14826 13812 14832 13824
rect 14884 13812 14890 13864
rect 16393 13855 16451 13861
rect 16393 13821 16405 13855
rect 16439 13852 16451 13855
rect 17129 13855 17187 13861
rect 16439 13824 16528 13852
rect 16439 13821 16451 13824
rect 16393 13815 16451 13821
rect 13924 13756 14228 13784
rect 13780 13744 13786 13756
rect 13078 13716 13084 13728
rect 12308 13688 13084 13716
rect 12308 13676 12314 13688
rect 13078 13676 13084 13688
rect 13136 13676 13142 13728
rect 14182 13676 14188 13728
rect 14240 13716 14246 13728
rect 14651 13719 14709 13725
rect 14651 13716 14663 13719
rect 14240 13688 14663 13716
rect 14240 13676 14246 13688
rect 14651 13685 14663 13688
rect 14697 13716 14709 13719
rect 14918 13716 14924 13728
rect 14697 13688 14924 13716
rect 14697 13685 14709 13688
rect 14651 13679 14709 13685
rect 14918 13676 14924 13688
rect 14976 13676 14982 13728
rect 16500 13716 16528 13824
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 19429 13855 19487 13861
rect 17175 13824 19288 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 18785 13787 18843 13793
rect 18785 13784 18797 13787
rect 17788 13756 18797 13784
rect 16666 13716 16672 13728
rect 16500 13688 16672 13716
rect 16666 13676 16672 13688
rect 16724 13716 16730 13728
rect 17126 13716 17132 13728
rect 16724 13688 17132 13716
rect 16724 13676 16730 13688
rect 17126 13676 17132 13688
rect 17184 13716 17190 13728
rect 17788 13716 17816 13756
rect 18785 13753 18797 13756
rect 18831 13753 18843 13787
rect 18785 13747 18843 13753
rect 19260 13725 19288 13824
rect 19429 13821 19441 13855
rect 19475 13821 19487 13855
rect 19429 13815 19487 13821
rect 19705 13855 19763 13861
rect 19705 13821 19717 13855
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 17184 13688 17816 13716
rect 19245 13719 19303 13725
rect 17184 13676 17190 13688
rect 19245 13685 19257 13719
rect 19291 13685 19303 13719
rect 19245 13679 19303 13685
rect 19334 13676 19340 13728
rect 19392 13716 19398 13728
rect 19444 13716 19472 13815
rect 19720 13784 19748 13815
rect 19978 13812 19984 13864
rect 20036 13812 20042 13864
rect 20622 13852 20628 13864
rect 20088 13824 20628 13852
rect 20088 13784 20116 13824
rect 20622 13812 20628 13824
rect 20680 13812 20686 13864
rect 20714 13812 20720 13864
rect 20772 13812 20778 13864
rect 22373 13855 22431 13861
rect 22373 13821 22385 13855
rect 22419 13852 22431 13855
rect 22649 13855 22707 13861
rect 22419 13824 22600 13852
rect 22419 13821 22431 13824
rect 22373 13815 22431 13821
rect 22572 13796 22600 13824
rect 22649 13821 22661 13855
rect 22695 13852 22707 13855
rect 22922 13852 22928 13864
rect 22695 13824 22928 13852
rect 22695 13821 22707 13824
rect 22649 13815 22707 13821
rect 19720 13756 20116 13784
rect 22554 13744 22560 13796
rect 22612 13744 22618 13796
rect 20346 13716 20352 13728
rect 19392 13688 20352 13716
rect 19392 13676 19398 13688
rect 20346 13676 20352 13688
rect 20404 13676 20410 13728
rect 20447 13719 20505 13725
rect 20447 13685 20459 13719
rect 20493 13716 20505 13719
rect 20806 13716 20812 13728
rect 20493 13688 20812 13716
rect 20493 13685 20505 13688
rect 20447 13679 20505 13685
rect 20806 13676 20812 13688
rect 20864 13676 20870 13728
rect 21910 13676 21916 13728
rect 21968 13716 21974 13728
rect 22664 13716 22692 13815
rect 22922 13812 22928 13824
rect 22980 13812 22986 13864
rect 23201 13855 23259 13861
rect 23201 13821 23213 13855
rect 23247 13852 23259 13855
rect 23290 13852 23296 13864
rect 23247 13824 23296 13852
rect 23247 13821 23259 13824
rect 23201 13815 23259 13821
rect 22738 13744 22744 13796
rect 22796 13784 22802 13796
rect 23216 13784 23244 13815
rect 23290 13812 23296 13824
rect 23348 13812 23354 13864
rect 23382 13812 23388 13864
rect 23440 13812 23446 13864
rect 23750 13852 23756 13864
rect 23584 13824 23756 13852
rect 22796 13756 23244 13784
rect 22796 13744 22802 13756
rect 21968 13688 22692 13716
rect 21968 13676 21974 13688
rect 23014 13676 23020 13728
rect 23072 13676 23078 13728
rect 23584 13725 23612 13824
rect 23750 13812 23756 13824
rect 23808 13812 23814 13864
rect 23934 13852 23940 13864
rect 23860 13824 23940 13852
rect 23860 13725 23888 13824
rect 23934 13812 23940 13824
rect 23992 13812 23998 13864
rect 24026 13812 24032 13864
rect 24084 13852 24090 13864
rect 24320 13861 24348 13892
rect 24394 13880 24400 13892
rect 24452 13880 24458 13932
rect 24995 13923 25053 13929
rect 24995 13889 25007 13923
rect 25041 13920 25053 13923
rect 25225 13923 25283 13929
rect 25041 13892 25176 13920
rect 25041 13889 25053 13892
rect 24995 13883 25053 13889
rect 24305 13855 24363 13861
rect 24084 13824 24164 13852
rect 24084 13812 24090 13824
rect 24136 13784 24164 13824
rect 24305 13821 24317 13855
rect 24351 13821 24363 13855
rect 24305 13815 24363 13821
rect 24489 13855 24547 13861
rect 24489 13821 24501 13855
rect 24535 13852 24547 13855
rect 24762 13852 24768 13864
rect 24535 13824 24768 13852
rect 24535 13821 24547 13824
rect 24489 13815 24547 13821
rect 24762 13812 24768 13824
rect 24820 13812 24826 13864
rect 25148 13852 25176 13892
rect 25225 13889 25237 13923
rect 25271 13920 25283 13923
rect 26068 13920 26096 14016
rect 28537 13991 28595 13997
rect 28537 13957 28549 13991
rect 28583 13957 28595 13991
rect 28537 13951 28595 13957
rect 25271 13892 26096 13920
rect 25271 13889 25283 13892
rect 25225 13883 25283 13889
rect 26418 13880 26424 13932
rect 26476 13920 26482 13932
rect 26697 13923 26755 13929
rect 26697 13920 26709 13923
rect 26476 13892 26709 13920
rect 26476 13880 26482 13892
rect 26697 13889 26709 13892
rect 26743 13889 26755 13923
rect 27160 13923 27218 13929
rect 27160 13920 27172 13923
rect 26697 13883 26755 13889
rect 26988 13892 27172 13920
rect 26988 13864 27016 13892
rect 27160 13889 27172 13892
rect 27206 13889 27218 13923
rect 27160 13883 27218 13889
rect 27338 13880 27344 13932
rect 27396 13920 27402 13932
rect 28552 13920 28580 13951
rect 29178 13948 29184 14000
rect 29236 13988 29242 14000
rect 30561 13991 30619 13997
rect 29236 13960 29684 13988
rect 29236 13948 29242 13960
rect 29656 13932 29684 13960
rect 30561 13957 30573 13991
rect 30607 13988 30619 13991
rect 30742 13988 30748 14000
rect 30607 13960 30748 13988
rect 30607 13957 30619 13960
rect 30561 13951 30619 13957
rect 30742 13948 30748 13960
rect 30800 13948 30806 14000
rect 27396 13892 28580 13920
rect 27396 13880 27402 13892
rect 29546 13880 29552 13932
rect 29604 13880 29610 13932
rect 29638 13880 29644 13932
rect 29696 13920 29702 13932
rect 31386 13920 31392 13932
rect 29696 13892 30052 13920
rect 29696 13880 29702 13892
rect 25682 13852 25688 13864
rect 25148 13824 25688 13852
rect 25682 13812 25688 13824
rect 25740 13812 25746 13864
rect 26970 13812 26976 13864
rect 27028 13812 27034 13864
rect 27433 13855 27491 13861
rect 27433 13821 27445 13855
rect 27479 13852 27491 13855
rect 27522 13852 27528 13864
rect 27479 13824 27528 13852
rect 27479 13821 27491 13824
rect 27433 13815 27491 13821
rect 27522 13812 27528 13824
rect 27580 13812 27586 13864
rect 28902 13812 28908 13864
rect 28960 13852 28966 13864
rect 29086 13852 29092 13864
rect 28960 13824 29092 13852
rect 28960 13812 28966 13824
rect 29086 13812 29092 13824
rect 29144 13812 29150 13864
rect 29181 13855 29239 13861
rect 29181 13821 29193 13855
rect 29227 13852 29239 13855
rect 29270 13852 29276 13864
rect 29227 13824 29276 13852
rect 29227 13821 29239 13824
rect 29181 13815 29239 13821
rect 24578 13784 24584 13796
rect 24136 13756 24584 13784
rect 24578 13744 24584 13756
rect 24636 13744 24642 13796
rect 23569 13719 23627 13725
rect 23569 13685 23581 13719
rect 23615 13685 23627 13719
rect 23569 13679 23627 13685
rect 23845 13719 23903 13725
rect 23845 13685 23857 13719
rect 23891 13685 23903 13719
rect 23845 13679 23903 13685
rect 24118 13676 24124 13728
rect 24176 13676 24182 13728
rect 24955 13719 25013 13725
rect 24955 13685 24967 13719
rect 25001 13716 25013 13719
rect 26510 13716 26516 13728
rect 25001 13688 26516 13716
rect 25001 13685 25013 13688
rect 24955 13679 25013 13685
rect 26510 13676 26516 13688
rect 26568 13676 26574 13728
rect 27154 13676 27160 13728
rect 27212 13725 27218 13728
rect 27212 13716 27221 13725
rect 29196 13716 29224 13815
rect 29270 13812 29276 13824
rect 29328 13812 29334 13864
rect 29457 13855 29515 13861
rect 29457 13821 29469 13855
rect 29503 13821 29515 13855
rect 29564 13852 29592 13880
rect 30024 13861 30052 13892
rect 30300 13892 31392 13920
rect 29733 13855 29791 13861
rect 29733 13852 29745 13855
rect 29564 13824 29745 13852
rect 29457 13815 29515 13821
rect 29733 13821 29745 13824
rect 29779 13821 29791 13855
rect 29733 13815 29791 13821
rect 30009 13855 30067 13861
rect 30009 13821 30021 13855
rect 30055 13821 30067 13855
rect 30009 13815 30067 13821
rect 30101 13855 30159 13861
rect 30101 13821 30113 13855
rect 30147 13852 30159 13855
rect 30300 13852 30328 13892
rect 31386 13880 31392 13892
rect 31444 13880 31450 13932
rect 30147 13824 30328 13852
rect 30147 13821 30159 13824
rect 30101 13815 30159 13821
rect 29472 13784 29500 13815
rect 30374 13812 30380 13864
rect 30432 13812 30438 13864
rect 29638 13784 29644 13796
rect 29472 13756 29644 13784
rect 29638 13744 29644 13756
rect 29696 13784 29702 13796
rect 30282 13784 30288 13796
rect 29696 13756 30288 13784
rect 29696 13744 29702 13756
rect 30282 13744 30288 13756
rect 30340 13744 30346 13796
rect 29822 13716 29828 13728
rect 27212 13688 27257 13716
rect 29196 13688 29828 13716
rect 27212 13679 27221 13688
rect 27212 13676 27218 13679
rect 29822 13676 29828 13688
rect 29880 13676 29886 13728
rect 552 13626 31072 13648
rect 552 13574 7988 13626
rect 8040 13574 8052 13626
rect 8104 13574 8116 13626
rect 8168 13574 8180 13626
rect 8232 13574 8244 13626
rect 8296 13574 15578 13626
rect 15630 13574 15642 13626
rect 15694 13574 15706 13626
rect 15758 13574 15770 13626
rect 15822 13574 15834 13626
rect 15886 13574 23168 13626
rect 23220 13574 23232 13626
rect 23284 13574 23296 13626
rect 23348 13574 23360 13626
rect 23412 13574 23424 13626
rect 23476 13574 30758 13626
rect 30810 13574 30822 13626
rect 30874 13574 30886 13626
rect 30938 13574 30950 13626
rect 31002 13574 31014 13626
rect 31066 13574 31072 13626
rect 552 13552 31072 13574
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 1771 13515 1829 13521
rect 1771 13512 1783 13515
rect 1728 13484 1783 13512
rect 1728 13472 1734 13484
rect 1771 13481 1783 13484
rect 1817 13481 1829 13515
rect 1771 13475 1829 13481
rect 3418 13472 3424 13524
rect 3476 13472 3482 13524
rect 3970 13472 3976 13524
rect 4028 13521 4034 13524
rect 4028 13512 4037 13521
rect 4028 13484 4073 13512
rect 4028 13475 4037 13484
rect 4028 13472 4034 13475
rect 5810 13472 5816 13524
rect 5868 13472 5874 13524
rect 6086 13472 6092 13524
rect 6144 13472 6150 13524
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7190 13512 7196 13524
rect 6972 13484 7196 13512
rect 6972 13472 6978 13484
rect 7190 13472 7196 13484
rect 7248 13512 7254 13524
rect 7291 13515 7349 13521
rect 7291 13512 7303 13515
rect 7248 13484 7303 13512
rect 7248 13472 7254 13484
rect 7291 13481 7303 13484
rect 7337 13481 7349 13515
rect 7291 13475 7349 13481
rect 7834 13472 7840 13524
rect 7892 13512 7898 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 7892 13484 9045 13512
rect 7892 13472 7898 13484
rect 9033 13481 9045 13484
rect 9079 13481 9091 13515
rect 9033 13475 9091 13481
rect 9214 13472 9220 13524
rect 9272 13512 9278 13524
rect 9493 13515 9551 13521
rect 9493 13512 9505 13515
rect 9272 13484 9505 13512
rect 9272 13472 9278 13484
rect 9493 13481 9505 13484
rect 9539 13481 9551 13515
rect 9493 13475 9551 13481
rect 9784 13484 10180 13512
rect 3436 13444 3464 13472
rect 3436 13416 3556 13444
rect 842 13336 848 13388
rect 900 13336 906 13388
rect 1210 13336 1216 13388
rect 1268 13336 1274 13388
rect 1302 13336 1308 13388
rect 1360 13336 1366 13388
rect 3528 13385 3556 13416
rect 5828 13416 6966 13444
rect 5828 13388 5856 13416
rect 2041 13379 2099 13385
rect 2041 13376 2053 13379
rect 1688 13348 2053 13376
rect 860 13308 888 13336
rect 1688 13308 1716 13348
rect 2041 13345 2053 13348
rect 2087 13345 2099 13379
rect 2041 13339 2099 13345
rect 3513 13379 3571 13385
rect 3513 13345 3525 13379
rect 3559 13345 3571 13379
rect 3513 13339 3571 13345
rect 5810 13336 5816 13388
rect 5868 13336 5874 13388
rect 5997 13379 6055 13385
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 6178 13376 6184 13388
rect 6043 13348 6184 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 6178 13336 6184 13348
rect 6236 13336 6242 13388
rect 6288 13385 6316 13416
rect 6273 13379 6331 13385
rect 6273 13345 6285 13379
rect 6319 13345 6331 13379
rect 6273 13339 6331 13345
rect 6454 13336 6460 13388
rect 6512 13376 6518 13388
rect 6733 13379 6791 13385
rect 6733 13376 6745 13379
rect 6512 13348 6745 13376
rect 6512 13336 6518 13348
rect 6733 13345 6745 13348
rect 6779 13345 6791 13379
rect 6733 13339 6791 13345
rect 6822 13336 6828 13388
rect 6880 13336 6886 13388
rect 6938 13376 6966 13416
rect 8478 13404 8484 13456
rect 8536 13444 8542 13456
rect 9122 13444 9128 13456
rect 8536 13416 9128 13444
rect 8536 13404 8542 13416
rect 9122 13404 9128 13416
rect 9180 13404 9186 13456
rect 9232 13416 9444 13444
rect 8846 13376 8852 13388
rect 6938 13348 8852 13376
rect 8846 13336 8852 13348
rect 8904 13376 8910 13388
rect 9232 13376 9260 13416
rect 8904 13348 9260 13376
rect 8904 13336 8910 13348
rect 9306 13336 9312 13388
rect 9364 13336 9370 13388
rect 9416 13376 9444 13416
rect 9582 13404 9588 13456
rect 9640 13404 9646 13456
rect 9784 13376 9812 13484
rect 10152 13444 10180 13484
rect 11146 13472 11152 13524
rect 11204 13472 11210 13524
rect 11790 13472 11796 13524
rect 11848 13512 11854 13524
rect 11848 13484 12572 13512
rect 11848 13472 11854 13484
rect 10152 13416 11744 13444
rect 9416 13348 9812 13376
rect 9858 13336 9864 13388
rect 9916 13336 9922 13388
rect 10152 13385 10180 13416
rect 11716 13388 11744 13416
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 10413 13363 10471 13369
rect 10413 13329 10425 13363
rect 10459 13329 10471 13363
rect 10962 13336 10968 13388
rect 11020 13376 11026 13388
rect 11422 13376 11428 13388
rect 11020 13348 11428 13376
rect 11020 13336 11026 13348
rect 11422 13336 11428 13348
rect 11480 13336 11486 13388
rect 11606 13336 11612 13388
rect 11664 13336 11670 13388
rect 11698 13336 11704 13388
rect 11756 13376 11762 13388
rect 11793 13379 11851 13385
rect 11793 13376 11805 13379
rect 11756 13348 11805 13376
rect 11756 13336 11762 13348
rect 11793 13345 11805 13348
rect 11839 13376 11851 13379
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 11839 13348 12081 13376
rect 11839 13345 11851 13348
rect 11793 13339 11851 13345
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 12544 13376 12572 13484
rect 14458 13472 14464 13524
rect 14516 13512 14522 13524
rect 14516 13484 15148 13512
rect 14516 13472 14522 13484
rect 14918 13404 14924 13456
rect 14976 13444 14982 13456
rect 15013 13447 15071 13453
rect 15013 13444 15025 13447
rect 14976 13416 15025 13444
rect 14976 13404 14982 13416
rect 15013 13413 15025 13416
rect 15059 13413 15071 13447
rect 15120 13444 15148 13484
rect 15378 13472 15384 13524
rect 15436 13512 15442 13524
rect 16117 13515 16175 13521
rect 16117 13512 16129 13515
rect 15436 13484 16129 13512
rect 15436 13472 15442 13484
rect 16117 13481 16129 13484
rect 16163 13481 16175 13515
rect 18969 13515 19027 13521
rect 18969 13512 18981 13515
rect 16117 13475 16175 13481
rect 16224 13484 18981 13512
rect 16224 13444 16252 13484
rect 18969 13481 18981 13484
rect 19015 13481 19027 13515
rect 18969 13475 19027 13481
rect 20346 13472 20352 13524
rect 20404 13472 20410 13524
rect 20714 13472 20720 13524
rect 20772 13512 20778 13524
rect 21545 13515 21603 13521
rect 21545 13512 21557 13515
rect 20772 13484 21557 13512
rect 20772 13472 20778 13484
rect 21545 13481 21557 13484
rect 21591 13481 21603 13515
rect 21545 13475 21603 13481
rect 21910 13472 21916 13524
rect 21968 13472 21974 13524
rect 22020 13484 23888 13512
rect 15120 13416 16252 13444
rect 15013 13407 15071 13413
rect 16758 13404 16764 13456
rect 16816 13404 16822 13456
rect 20364 13444 20392 13472
rect 21928 13444 21956 13472
rect 20364 13416 21956 13444
rect 12820 13376 12943 13380
rect 12544 13352 12943 13376
rect 12544 13348 12848 13352
rect 12069 13339 12127 13345
rect 10413 13323 10471 13329
rect 860 13280 1716 13308
rect 1811 13311 1869 13317
rect 1811 13277 1823 13311
rect 1857 13308 1869 13311
rect 2222 13308 2228 13320
rect 1857 13280 2228 13308
rect 1857 13277 1869 13280
rect 1811 13271 1869 13277
rect 2222 13268 2228 13280
rect 2280 13268 2286 13320
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13308 3479 13311
rect 3786 13310 3792 13320
rect 3718 13308 3792 13310
rect 3467 13282 3792 13308
rect 3467 13280 3746 13282
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 3786 13268 3792 13282
rect 3844 13268 3850 13320
rect 3970 13268 3976 13320
rect 4028 13308 4034 13320
rect 4249 13311 4307 13317
rect 4028 13280 4073 13308
rect 4028 13268 4034 13280
rect 4249 13277 4261 13311
rect 4295 13308 4307 13311
rect 5074 13308 5080 13320
rect 4295 13280 5080 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 5074 13268 5080 13280
rect 5132 13268 5138 13320
rect 5629 13311 5687 13317
rect 5629 13277 5641 13311
rect 5675 13308 5687 13311
rect 7190 13308 7196 13320
rect 5675 13280 7196 13308
rect 5675 13277 5687 13280
rect 5629 13271 5687 13277
rect 7190 13268 7196 13280
rect 7248 13268 7254 13320
rect 7282 13268 7288 13320
rect 7340 13268 7346 13320
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13308 7619 13311
rect 8754 13308 8760 13320
rect 7607 13280 8760 13308
rect 7607 13277 7619 13280
rect 7561 13271 7619 13277
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 9122 13268 9128 13320
rect 9180 13308 9186 13320
rect 9646 13308 9812 13310
rect 9180 13282 10364 13308
rect 9180 13280 9674 13282
rect 9784 13280 10364 13282
rect 9180 13268 9186 13280
rect 5350 13200 5356 13252
rect 5408 13240 5414 13252
rect 6270 13240 6276 13252
rect 5408 13212 6276 13240
rect 5408 13200 5414 13212
rect 6270 13200 6276 13212
rect 6328 13200 6334 13252
rect 6362 13200 6368 13252
rect 6420 13240 6426 13252
rect 6730 13240 6736 13252
rect 6420 13212 6736 13240
rect 6420 13200 6426 13212
rect 6730 13200 6736 13212
rect 6788 13200 6794 13252
rect 8849 13243 8907 13249
rect 8849 13209 8861 13243
rect 8895 13240 8907 13243
rect 9490 13240 9496 13252
rect 8895 13212 9496 13240
rect 8895 13209 8907 13212
rect 8849 13203 8907 13209
rect 9490 13200 9496 13212
rect 9548 13200 9554 13252
rect 10045 13243 10103 13249
rect 10045 13209 10057 13243
rect 10091 13240 10103 13243
rect 10134 13240 10140 13252
rect 10091 13212 10140 13240
rect 10091 13209 10103 13212
rect 10045 13203 10103 13209
rect 10134 13200 10140 13212
rect 10192 13200 10198 13252
rect 10336 13249 10364 13280
rect 10321 13243 10379 13249
rect 10321 13209 10333 13243
rect 10367 13209 10379 13243
rect 10321 13203 10379 13209
rect 10428 13240 10456 13323
rect 10686 13268 10692 13320
rect 10744 13268 10750 13320
rect 11054 13268 11060 13320
rect 11112 13268 11118 13320
rect 11238 13268 11244 13320
rect 11296 13268 11302 13320
rect 11330 13268 11336 13320
rect 11388 13308 11394 13320
rect 11517 13311 11575 13317
rect 11517 13308 11529 13311
rect 11388 13280 11529 13308
rect 11388 13268 11394 13280
rect 11517 13277 11529 13280
rect 11563 13277 11575 13311
rect 11624 13308 11652 13336
rect 12342 13308 12348 13320
rect 11624 13280 12348 13308
rect 11517 13271 11575 13277
rect 12342 13268 12348 13280
rect 12400 13268 12406 13320
rect 12434 13268 12440 13320
rect 12492 13268 12498 13320
rect 12802 13317 12808 13320
rect 12764 13311 12808 13317
rect 12764 13277 12776 13311
rect 12764 13271 12808 13277
rect 12802 13268 12808 13271
rect 12860 13268 12866 13320
rect 12915 13319 12943 13352
rect 13078 13336 13084 13388
rect 13136 13376 13142 13388
rect 14737 13379 14795 13385
rect 13136 13348 13768 13376
rect 13136 13336 13142 13348
rect 12900 13313 12958 13319
rect 12900 13279 12912 13313
rect 12946 13279 12958 13313
rect 12900 13273 12958 13279
rect 12986 13268 12992 13320
rect 13044 13308 13050 13320
rect 13173 13311 13231 13317
rect 13173 13308 13185 13311
rect 13044 13280 13185 13308
rect 13044 13268 13050 13280
rect 13173 13277 13185 13280
rect 13219 13277 13231 13311
rect 13740 13308 13768 13348
rect 14737 13345 14749 13379
rect 14783 13376 14795 13379
rect 15102 13376 15108 13388
rect 14783 13348 15108 13376
rect 14783 13345 14795 13348
rect 14737 13339 14795 13345
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 15381 13379 15439 13385
rect 15381 13345 15393 13379
rect 15427 13376 15439 13379
rect 15470 13376 15476 13388
rect 15427 13348 15476 13376
rect 15427 13345 15439 13348
rect 15381 13339 15439 13345
rect 15470 13336 15476 13348
rect 15528 13336 15534 13388
rect 16298 13376 16304 13388
rect 15580 13348 16304 13376
rect 15580 13308 15608 13348
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 16485 13379 16543 13385
rect 16485 13345 16497 13379
rect 16531 13376 16543 13379
rect 16574 13376 16580 13388
rect 16531 13348 16580 13376
rect 16531 13345 16543 13348
rect 16485 13339 16543 13345
rect 13740 13280 15608 13308
rect 13173 13271 13231 13277
rect 10704 13240 10732 13268
rect 10428 13212 10732 13240
rect 11072 13240 11100 13268
rect 11977 13243 12035 13249
rect 11977 13240 11989 13243
rect 11072 13212 11989 13240
rect 1029 13175 1087 13181
rect 1029 13141 1041 13175
rect 1075 13172 1087 13175
rect 1578 13172 1584 13184
rect 1075 13144 1584 13172
rect 1075 13141 1087 13144
rect 1029 13135 1087 13141
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 3142 13132 3148 13184
rect 3200 13172 3206 13184
rect 3510 13172 3516 13184
rect 3200 13144 3516 13172
rect 3200 13132 3206 13144
rect 3510 13132 3516 13144
rect 3568 13172 3574 13184
rect 6086 13172 6092 13184
rect 3568 13144 6092 13172
rect 3568 13132 3574 13144
rect 6086 13132 6092 13144
rect 6144 13132 6150 13184
rect 6549 13175 6607 13181
rect 6549 13141 6561 13175
rect 6595 13172 6607 13175
rect 7098 13172 7104 13184
rect 6595 13144 7104 13172
rect 6595 13141 6607 13144
rect 6549 13135 6607 13141
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 9214 13172 9220 13184
rect 7708 13144 9220 13172
rect 7708 13132 7714 13144
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 9306 13132 9312 13184
rect 9364 13172 9370 13184
rect 10428 13172 10456 13212
rect 11977 13209 11989 13212
rect 12023 13209 12035 13243
rect 11977 13203 12035 13209
rect 13832 13212 14412 13240
rect 13832 13184 13860 13212
rect 9364 13144 10456 13172
rect 9364 13132 9370 13144
rect 10594 13132 10600 13184
rect 10652 13132 10658 13184
rect 12253 13175 12311 13181
rect 12253 13141 12265 13175
rect 12299 13172 12311 13175
rect 13354 13172 13360 13184
rect 12299 13144 13360 13172
rect 12299 13141 12311 13144
rect 12253 13135 12311 13141
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 13814 13132 13820 13184
rect 13872 13132 13878 13184
rect 13998 13132 14004 13184
rect 14056 13172 14062 13184
rect 14277 13175 14335 13181
rect 14277 13172 14289 13175
rect 14056 13144 14289 13172
rect 14056 13132 14062 13144
rect 14277 13141 14289 13144
rect 14323 13141 14335 13175
rect 14384 13172 14412 13212
rect 14734 13200 14740 13252
rect 14792 13240 14798 13252
rect 16500 13240 16528 13339
rect 16574 13336 16580 13348
rect 16632 13336 16638 13388
rect 16776 13376 16804 13404
rect 17456 13379 17514 13385
rect 17456 13376 17468 13379
rect 16776 13348 17468 13376
rect 17456 13345 17468 13348
rect 17502 13345 17514 13379
rect 17456 13339 17514 13345
rect 17865 13379 17923 13385
rect 17865 13345 17877 13379
rect 17911 13376 17923 13379
rect 18690 13376 18696 13388
rect 17911 13348 18696 13376
rect 17911 13345 17923 13348
rect 17865 13339 17923 13345
rect 18690 13336 18696 13348
rect 18748 13336 18754 13388
rect 20898 13376 20904 13388
rect 19352 13348 20904 13376
rect 17126 13268 17132 13320
rect 17184 13268 17190 13320
rect 17635 13311 17693 13317
rect 17635 13277 17647 13311
rect 17681 13308 17693 13311
rect 19352 13308 19380 13348
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 21266 13336 21272 13388
rect 21324 13376 21330 13388
rect 21453 13379 21511 13385
rect 21453 13376 21465 13379
rect 21324 13348 21465 13376
rect 21324 13336 21330 13348
rect 21453 13345 21465 13348
rect 21499 13376 21511 13379
rect 21634 13376 21640 13388
rect 21499 13348 21640 13376
rect 21499 13345 21511 13348
rect 21453 13339 21511 13345
rect 21634 13336 21640 13348
rect 21692 13336 21698 13388
rect 21744 13385 21772 13416
rect 21729 13379 21787 13385
rect 21729 13345 21741 13379
rect 21775 13345 21787 13379
rect 21729 13339 21787 13345
rect 21913 13379 21971 13385
rect 21913 13345 21925 13379
rect 21959 13376 21971 13379
rect 22020 13376 22048 13484
rect 23860 13456 23888 13484
rect 23934 13472 23940 13524
rect 23992 13472 23998 13524
rect 24118 13472 24124 13524
rect 24176 13512 24182 13524
rect 26970 13512 26976 13524
rect 24176 13484 26976 13512
rect 24176 13472 24182 13484
rect 26970 13472 26976 13484
rect 27028 13472 27034 13524
rect 27430 13472 27436 13524
rect 27488 13512 27494 13524
rect 28261 13515 28319 13521
rect 28261 13512 28273 13515
rect 27488 13484 28273 13512
rect 27488 13472 27494 13484
rect 28261 13481 28273 13484
rect 28307 13481 28319 13515
rect 28261 13475 28319 13481
rect 29270 13472 29276 13524
rect 29328 13512 29334 13524
rect 29730 13512 29736 13524
rect 29328 13484 29736 13512
rect 29328 13472 29334 13484
rect 29730 13472 29736 13484
rect 29788 13472 29794 13524
rect 23842 13404 23848 13456
rect 23900 13444 23906 13456
rect 23900 13416 24164 13444
rect 23900 13404 23906 13416
rect 24136 13385 24164 13416
rect 24210 13404 24216 13456
rect 24268 13404 24274 13456
rect 21959 13348 22048 13376
rect 22240 13379 22298 13385
rect 21959 13345 21971 13348
rect 21913 13339 21971 13345
rect 22240 13345 22252 13379
rect 22286 13376 22298 13379
rect 24121 13379 24179 13385
rect 22286 13348 23888 13376
rect 22286 13345 22298 13348
rect 22240 13339 22298 13345
rect 17681 13280 19380 13308
rect 17681 13277 17693 13280
rect 17635 13271 17693 13277
rect 19426 13268 19432 13320
rect 19484 13268 19490 13320
rect 19705 13311 19763 13317
rect 19705 13277 19717 13311
rect 19751 13308 19763 13311
rect 19886 13308 19892 13320
rect 19751 13280 19892 13308
rect 19751 13277 19763 13280
rect 19705 13271 19763 13277
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13308 21143 13311
rect 22094 13308 22100 13320
rect 21131 13280 22100 13308
rect 21131 13277 21143 13280
rect 21085 13271 21143 13277
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 22370 13268 22376 13320
rect 22428 13268 22434 13320
rect 22646 13268 22652 13320
rect 22704 13268 22710 13320
rect 23860 13308 23888 13348
rect 24121 13345 24133 13379
rect 24167 13345 24179 13379
rect 24228 13376 24256 13404
rect 24504 13376 24627 13380
rect 24228 13352 24627 13376
rect 24228 13348 24532 13352
rect 24121 13339 24179 13345
rect 24302 13308 24308 13320
rect 23860 13280 24308 13308
rect 24302 13268 24308 13280
rect 24360 13308 24366 13320
rect 24599 13319 24627 13352
rect 24854 13336 24860 13388
rect 24912 13336 24918 13388
rect 26237 13379 26295 13385
rect 26237 13345 26249 13379
rect 26283 13376 26295 13379
rect 26283 13348 26927 13376
rect 26283 13345 26295 13348
rect 26237 13339 26295 13345
rect 24448 13311 24506 13317
rect 24448 13308 24460 13311
rect 24360 13280 24460 13308
rect 24360 13268 24366 13280
rect 24448 13277 24460 13280
rect 24494 13277 24506 13311
rect 24448 13271 24506 13277
rect 24584 13313 24642 13319
rect 24584 13279 24596 13313
rect 24630 13279 24642 13313
rect 24584 13273 24642 13279
rect 24762 13268 24768 13320
rect 24820 13308 24826 13320
rect 26418 13308 26424 13320
rect 24820 13280 26424 13308
rect 24820 13268 24826 13280
rect 26418 13268 26424 13280
rect 26476 13268 26482 13320
rect 26602 13268 26608 13320
rect 26660 13308 26666 13320
rect 26786 13317 26792 13320
rect 26748 13311 26792 13317
rect 26748 13308 26760 13311
rect 26660 13280 26760 13308
rect 26660 13268 26666 13280
rect 26748 13277 26760 13280
rect 26748 13271 26792 13277
rect 26786 13268 26792 13271
rect 26844 13268 26850 13320
rect 26899 13319 26927 13348
rect 26970 13336 26976 13388
rect 27028 13376 27034 13388
rect 27157 13379 27215 13385
rect 27157 13376 27169 13379
rect 27028 13348 27169 13376
rect 27028 13336 27034 13348
rect 27157 13345 27169 13348
rect 27203 13345 27215 13379
rect 30561 13379 30619 13385
rect 30561 13376 30573 13379
rect 27157 13339 27215 13345
rect 27816 13348 28948 13376
rect 26884 13313 26942 13319
rect 26884 13279 26896 13313
rect 26930 13279 26942 13313
rect 26884 13273 26942 13279
rect 14792 13212 16528 13240
rect 21284 13212 21680 13240
rect 14792 13200 14798 13212
rect 15473 13175 15531 13181
rect 15473 13172 15485 13175
rect 14384 13144 15485 13172
rect 14277 13135 14335 13141
rect 15473 13141 15485 13144
rect 15519 13172 15531 13175
rect 16206 13172 16212 13184
rect 15519 13144 16212 13172
rect 15519 13141 15531 13144
rect 15473 13135 15531 13141
rect 16206 13132 16212 13144
rect 16264 13132 16270 13184
rect 16666 13132 16672 13184
rect 16724 13172 16730 13184
rect 17402 13172 17408 13184
rect 16724 13144 17408 13172
rect 16724 13132 16730 13144
rect 17402 13132 17408 13144
rect 17460 13132 17466 13184
rect 19702 13132 19708 13184
rect 19760 13172 19766 13184
rect 20162 13172 20168 13184
rect 19760 13144 20168 13172
rect 19760 13132 19766 13144
rect 20162 13132 20168 13144
rect 20220 13132 20226 13184
rect 21284 13181 21312 13212
rect 21269 13175 21327 13181
rect 21269 13141 21281 13175
rect 21315 13141 21327 13175
rect 21652 13172 21680 13212
rect 24026 13200 24032 13252
rect 24084 13200 24090 13252
rect 22278 13172 22284 13184
rect 21652 13144 22284 13172
rect 21269 13135 21327 13141
rect 22278 13132 22284 13144
rect 22336 13132 22342 13184
rect 23014 13132 23020 13184
rect 23072 13172 23078 13184
rect 24044 13172 24072 13200
rect 23072 13144 24072 13172
rect 23072 13132 23078 13144
rect 26786 13132 26792 13184
rect 26844 13172 26850 13184
rect 27816 13172 27844 13348
rect 28626 13268 28632 13320
rect 28684 13268 28690 13320
rect 28920 13317 28948 13348
rect 29840 13348 30573 13376
rect 29840 13320 29868 13348
rect 30561 13345 30573 13348
rect 30607 13345 30619 13379
rect 30561 13339 30619 13345
rect 28905 13311 28963 13317
rect 28905 13277 28917 13311
rect 28951 13277 28963 13311
rect 28905 13271 28963 13277
rect 29822 13268 29828 13320
rect 29880 13268 29886 13320
rect 30377 13243 30435 13249
rect 30377 13240 30389 13243
rect 30300 13212 30389 13240
rect 30300 13184 30328 13212
rect 30377 13209 30389 13212
rect 30423 13209 30435 13243
rect 30377 13203 30435 13209
rect 26844 13144 27844 13172
rect 26844 13132 26850 13144
rect 28902 13132 28908 13184
rect 28960 13172 28966 13184
rect 30009 13175 30067 13181
rect 30009 13172 30021 13175
rect 28960 13144 30021 13172
rect 28960 13132 28966 13144
rect 30009 13141 30021 13144
rect 30055 13141 30067 13175
rect 30009 13135 30067 13141
rect 30282 13132 30288 13184
rect 30340 13132 30346 13184
rect 552 13082 30912 13104
rect 552 13030 4193 13082
rect 4245 13030 4257 13082
rect 4309 13030 4321 13082
rect 4373 13030 4385 13082
rect 4437 13030 4449 13082
rect 4501 13030 11783 13082
rect 11835 13030 11847 13082
rect 11899 13030 11911 13082
rect 11963 13030 11975 13082
rect 12027 13030 12039 13082
rect 12091 13030 19373 13082
rect 19425 13030 19437 13082
rect 19489 13030 19501 13082
rect 19553 13030 19565 13082
rect 19617 13030 19629 13082
rect 19681 13030 26963 13082
rect 27015 13030 27027 13082
rect 27079 13030 27091 13082
rect 27143 13030 27155 13082
rect 27207 13030 27219 13082
rect 27271 13030 30912 13082
rect 552 13008 30912 13030
rect 1210 12928 1216 12980
rect 1268 12968 1274 12980
rect 2961 12971 3019 12977
rect 1268 12940 2360 12968
rect 1268 12928 1274 12940
rect 937 12835 995 12841
rect 937 12801 949 12835
rect 983 12832 995 12835
rect 1302 12832 1308 12844
rect 983 12804 1308 12832
rect 983 12801 995 12804
rect 937 12795 995 12801
rect 1302 12792 1308 12804
rect 1360 12792 1366 12844
rect 1443 12833 1501 12839
rect 1443 12799 1455 12833
rect 1489 12799 1501 12833
rect 1443 12793 1501 12799
rect 1458 12764 1486 12793
rect 1578 12792 1584 12844
rect 1636 12832 1642 12844
rect 1673 12835 1731 12841
rect 1673 12832 1685 12835
rect 1636 12804 1685 12832
rect 1636 12792 1642 12804
rect 1673 12801 1685 12804
rect 1719 12801 1731 12835
rect 2332 12832 2360 12940
rect 2961 12937 2973 12971
rect 3007 12968 3019 12971
rect 4246 12968 4252 12980
rect 3007 12940 4252 12968
rect 3007 12937 3019 12940
rect 2961 12931 3019 12937
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 7282 12968 7288 12980
rect 5951 12940 7288 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 7282 12928 7288 12940
rect 7340 12928 7346 12980
rect 8754 12928 8760 12980
rect 8812 12928 8818 12980
rect 8956 12940 9168 12968
rect 3237 12903 3295 12909
rect 3237 12869 3249 12903
rect 3283 12900 3295 12903
rect 3418 12900 3424 12912
rect 3283 12872 3424 12900
rect 3283 12869 3295 12872
rect 3237 12863 3295 12869
rect 3418 12860 3424 12872
rect 3476 12860 3482 12912
rect 3605 12903 3663 12909
rect 3605 12869 3617 12903
rect 3651 12869 3663 12903
rect 3605 12863 3663 12869
rect 3620 12832 3648 12863
rect 8386 12860 8392 12912
rect 8444 12900 8450 12912
rect 8573 12903 8631 12909
rect 8573 12900 8585 12903
rect 8444 12872 8585 12900
rect 8444 12860 8450 12872
rect 8573 12869 8585 12872
rect 8619 12900 8631 12903
rect 8956 12900 8984 12940
rect 8619 12872 8984 12900
rect 9033 12903 9091 12909
rect 8619 12869 8631 12872
rect 8573 12863 8631 12869
rect 9033 12869 9045 12903
rect 9079 12869 9091 12903
rect 9033 12863 9091 12869
rect 2332 12804 3556 12832
rect 3620 12804 4200 12832
rect 1673 12795 1731 12801
rect 2314 12764 2320 12776
rect 1458 12736 2320 12764
rect 2314 12724 2320 12736
rect 2372 12764 2378 12776
rect 2958 12764 2964 12776
rect 2372 12736 2964 12764
rect 2372 12724 2378 12736
rect 2958 12724 2964 12736
rect 3016 12724 3022 12776
rect 3418 12724 3424 12776
rect 3476 12724 3482 12776
rect 3528 12764 3556 12804
rect 3602 12764 3608 12776
rect 3528 12736 3608 12764
rect 3602 12724 3608 12736
rect 3660 12764 3666 12776
rect 3789 12767 3847 12773
rect 3789 12764 3801 12767
rect 3660 12736 3801 12764
rect 3660 12724 3666 12736
rect 3789 12733 3801 12736
rect 3835 12733 3847 12767
rect 3789 12727 3847 12733
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12733 3939 12767
rect 4172 12764 4200 12804
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4344 12835 4402 12841
rect 4344 12832 4356 12835
rect 4304 12804 4356 12832
rect 4304 12792 4310 12804
rect 4344 12801 4356 12804
rect 4390 12801 4402 12835
rect 4344 12795 4402 12801
rect 5626 12792 5632 12844
rect 5684 12832 5690 12844
rect 6552 12835 6610 12841
rect 6552 12832 6564 12835
rect 5684 12804 6564 12832
rect 5684 12792 5690 12804
rect 6552 12801 6564 12804
rect 6598 12801 6610 12835
rect 6552 12795 6610 12801
rect 6730 12792 6736 12844
rect 6788 12792 6794 12844
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 9048 12832 9076 12863
rect 6871 12804 9076 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 4617 12767 4675 12773
rect 4617 12764 4629 12767
rect 4172 12736 4629 12764
rect 3881 12727 3939 12733
rect 4617 12733 4629 12736
rect 4663 12733 4675 12767
rect 4617 12727 4675 12733
rect 6089 12767 6147 12773
rect 6089 12733 6101 12767
rect 6135 12764 6147 12767
rect 6638 12764 6644 12776
rect 6135 12736 6644 12764
rect 6135 12733 6147 12736
rect 6089 12727 6147 12733
rect 3896 12696 3924 12727
rect 6638 12724 6644 12736
rect 6696 12724 6702 12776
rect 6748 12764 6776 12792
rect 6748 12736 7696 12764
rect 3528 12668 3924 12696
rect 3528 12640 3556 12668
rect 1403 12631 1461 12637
rect 1403 12597 1415 12631
rect 1449 12628 1461 12631
rect 1670 12628 1676 12640
rect 1449 12600 1676 12628
rect 1449 12597 1461 12600
rect 1403 12591 1461 12597
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 3510 12588 3516 12640
rect 3568 12588 3574 12640
rect 4347 12631 4405 12637
rect 4347 12597 4359 12631
rect 4393 12628 4405 12631
rect 4522 12628 4528 12640
rect 4393 12600 4528 12628
rect 4393 12597 4405 12600
rect 4347 12591 4405 12597
rect 4522 12588 4528 12600
rect 4580 12588 4586 12640
rect 6555 12631 6613 12637
rect 6555 12597 6567 12631
rect 6601 12628 6613 12631
rect 6914 12628 6920 12640
rect 6601 12600 6920 12628
rect 6601 12597 6613 12600
rect 6555 12591 6613 12597
rect 6914 12588 6920 12600
rect 6972 12588 6978 12640
rect 7668 12628 7696 12736
rect 7834 12724 7840 12776
rect 7892 12764 7898 12776
rect 8389 12767 8447 12773
rect 8389 12764 8401 12767
rect 7892 12736 8401 12764
rect 7892 12724 7898 12736
rect 8389 12733 8401 12736
rect 8435 12764 8447 12767
rect 8570 12764 8576 12776
rect 8435 12736 8576 12764
rect 8435 12733 8447 12736
rect 8389 12727 8447 12733
rect 8570 12724 8576 12736
rect 8628 12724 8634 12776
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 8812 12736 8953 12764
rect 8812 12724 8818 12736
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 9140 12764 9168 12940
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 11238 12968 11244 12980
rect 9272 12940 11244 12968
rect 9272 12928 9278 12940
rect 11238 12928 11244 12940
rect 11296 12928 11302 12980
rect 12066 12928 12072 12980
rect 12124 12928 12130 12980
rect 12161 12971 12219 12977
rect 12161 12937 12173 12971
rect 12207 12968 12219 12971
rect 12342 12968 12348 12980
rect 12207 12940 12348 12968
rect 12207 12937 12219 12940
rect 12161 12931 12219 12937
rect 12342 12928 12348 12940
rect 12400 12928 12406 12980
rect 12544 12940 14964 12968
rect 9398 12860 9404 12912
rect 9456 12900 9462 12912
rect 12544 12900 12572 12940
rect 9456 12872 9720 12900
rect 9456 12860 9462 12872
rect 9692 12841 9720 12872
rect 11072 12872 12572 12900
rect 12621 12903 12679 12909
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12801 9735 12835
rect 9677 12795 9735 12801
rect 9950 12792 9956 12844
rect 10008 12832 10014 12844
rect 10140 12835 10198 12841
rect 10140 12832 10152 12835
rect 10008 12804 10152 12832
rect 10008 12792 10014 12804
rect 10140 12801 10152 12804
rect 10186 12801 10198 12835
rect 10140 12795 10198 12801
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 11072 12832 11100 12872
rect 12621 12869 12633 12903
rect 12667 12869 12679 12903
rect 12621 12863 12679 12869
rect 13173 12903 13231 12909
rect 13173 12869 13185 12903
rect 13219 12900 13231 12903
rect 13354 12900 13360 12912
rect 13219 12872 13360 12900
rect 13219 12869 13231 12872
rect 13173 12863 13231 12869
rect 10928 12804 11100 12832
rect 10928 12792 10934 12804
rect 11698 12792 11704 12844
rect 11756 12832 11762 12844
rect 12636 12832 12664 12863
rect 13354 12860 13360 12872
rect 13412 12860 13418 12912
rect 11756 12804 12388 12832
rect 12636 12804 13676 12832
rect 11756 12792 11762 12804
rect 9217 12767 9275 12773
rect 9217 12764 9229 12767
rect 9140 12736 9229 12764
rect 8941 12727 8999 12733
rect 9217 12733 9229 12736
rect 9263 12733 9275 12767
rect 9217 12727 9275 12733
rect 10413 12767 10471 12773
rect 10413 12733 10425 12767
rect 10459 12764 10471 12767
rect 11238 12764 11244 12776
rect 10459 12736 11244 12764
rect 10459 12733 10471 12736
rect 10413 12727 10471 12733
rect 11238 12724 11244 12736
rect 11296 12724 11302 12776
rect 12360 12773 12388 12804
rect 11885 12767 11943 12773
rect 11885 12764 11897 12767
rect 11624 12736 11897 12764
rect 8205 12699 8263 12705
rect 8205 12665 8217 12699
rect 8251 12696 8263 12699
rect 8251 12668 9674 12696
rect 8251 12665 8263 12668
rect 8205 12659 8263 12665
rect 9646 12640 9674 12668
rect 9309 12631 9367 12637
rect 9309 12628 9321 12631
rect 7668 12600 9321 12628
rect 9309 12597 9321 12600
rect 9355 12597 9367 12631
rect 9646 12600 9680 12640
rect 9309 12591 9367 12597
rect 9674 12588 9680 12600
rect 9732 12588 9738 12640
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10143 12631 10201 12637
rect 10143 12628 10155 12631
rect 10008 12600 10155 12628
rect 10008 12588 10014 12600
rect 10143 12597 10155 12600
rect 10189 12597 10201 12631
rect 10143 12591 10201 12597
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 11330 12628 11336 12640
rect 10744 12600 11336 12628
rect 10744 12588 10750 12600
rect 11330 12588 11336 12600
rect 11388 12628 11394 12640
rect 11624 12628 11652 12736
rect 11885 12733 11897 12736
rect 11931 12733 11943 12767
rect 11885 12727 11943 12733
rect 12345 12767 12403 12773
rect 12345 12733 12357 12767
rect 12391 12733 12403 12767
rect 12345 12727 12403 12733
rect 12805 12767 12863 12773
rect 12805 12733 12817 12767
rect 12851 12764 12863 12767
rect 12894 12764 12900 12776
rect 12851 12736 12900 12764
rect 12851 12733 12863 12736
rect 12805 12727 12863 12733
rect 12894 12724 12900 12736
rect 12952 12724 12958 12776
rect 13081 12767 13139 12773
rect 13081 12733 13093 12767
rect 13127 12764 13139 12767
rect 13170 12764 13176 12776
rect 13127 12736 13176 12764
rect 13127 12733 13139 12736
rect 13081 12727 13139 12733
rect 11790 12656 11796 12708
rect 11848 12696 11854 12708
rect 13096 12696 13124 12727
rect 13170 12724 13176 12736
rect 13228 12724 13234 12776
rect 13357 12767 13415 12773
rect 13357 12733 13369 12767
rect 13403 12764 13415 12767
rect 13446 12764 13452 12776
rect 13403 12736 13452 12764
rect 13403 12733 13415 12736
rect 13357 12727 13415 12733
rect 13446 12724 13452 12736
rect 13504 12724 13510 12776
rect 13538 12724 13544 12776
rect 13596 12724 13602 12776
rect 13648 12764 13676 12804
rect 13814 12792 13820 12844
rect 13872 12830 13878 12844
rect 14047 12833 14105 12839
rect 14047 12832 14059 12833
rect 13924 12830 14059 12832
rect 13872 12804 14059 12830
rect 13872 12802 13952 12804
rect 13872 12792 13878 12802
rect 14047 12799 14059 12804
rect 14093 12799 14105 12833
rect 14936 12832 14964 12940
rect 15102 12928 15108 12980
rect 15160 12968 15166 12980
rect 17310 12968 17316 12980
rect 15160 12940 17316 12968
rect 15160 12928 15166 12940
rect 17310 12928 17316 12940
rect 17368 12928 17374 12980
rect 21634 12968 21640 12980
rect 18432 12940 21640 12968
rect 18432 12909 18460 12940
rect 21634 12928 21640 12940
rect 21692 12928 21698 12980
rect 22189 12971 22247 12977
rect 22189 12937 22201 12971
rect 22235 12968 22247 12971
rect 22646 12968 22652 12980
rect 22235 12940 22652 12968
rect 22235 12937 22247 12940
rect 22189 12931 22247 12937
rect 22646 12928 22652 12940
rect 22704 12928 22710 12980
rect 22741 12971 22799 12977
rect 22741 12937 22753 12971
rect 22787 12968 22799 12971
rect 22787 12940 23152 12968
rect 22787 12937 22799 12940
rect 22741 12931 22799 12937
rect 18417 12903 18475 12909
rect 18417 12869 18429 12903
rect 18463 12869 18475 12903
rect 18417 12863 18475 12869
rect 19334 12860 19340 12912
rect 19392 12860 19398 12912
rect 19702 12860 19708 12912
rect 19760 12860 19766 12912
rect 19886 12860 19892 12912
rect 19944 12860 19950 12912
rect 22005 12903 22063 12909
rect 22005 12869 22017 12903
rect 22051 12900 22063 12903
rect 22370 12900 22376 12912
rect 22051 12872 22376 12900
rect 22051 12869 22063 12872
rect 22005 12863 22063 12869
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 22554 12860 22560 12912
rect 22612 12860 22618 12912
rect 16856 12835 16914 12841
rect 16856 12832 16868 12835
rect 14936 12804 16868 12832
rect 14047 12793 14105 12799
rect 16856 12801 16868 12804
rect 16902 12801 16914 12835
rect 16856 12795 16914 12801
rect 14277 12767 14335 12773
rect 14277 12764 14289 12767
rect 13648 12760 13860 12764
rect 13924 12760 14289 12764
rect 13648 12736 14289 12760
rect 13832 12732 13952 12736
rect 14277 12733 14289 12736
rect 14323 12733 14335 12767
rect 14277 12727 14335 12733
rect 16390 12724 16396 12776
rect 16448 12724 16454 12776
rect 17129 12767 17187 12773
rect 17129 12764 17141 12767
rect 16500 12736 17141 12764
rect 11848 12668 13124 12696
rect 15657 12699 15715 12705
rect 11848 12656 11854 12668
rect 15657 12665 15669 12699
rect 15703 12696 15715 12699
rect 16022 12696 16028 12708
rect 15703 12668 16028 12696
rect 15703 12665 15715 12668
rect 15657 12659 15715 12665
rect 16022 12656 16028 12668
rect 16080 12656 16086 12708
rect 16301 12699 16359 12705
rect 16301 12665 16313 12699
rect 16347 12696 16359 12699
rect 16500 12696 16528 12736
rect 17129 12733 17141 12736
rect 17175 12764 17187 12767
rect 17175 12736 17816 12764
rect 17175 12733 17187 12736
rect 17129 12727 17187 12733
rect 16347 12668 16528 12696
rect 17788 12696 17816 12736
rect 19058 12724 19064 12776
rect 19116 12724 19122 12776
rect 19352 12773 19380 12860
rect 19904 12832 19932 12860
rect 19981 12835 20039 12841
rect 19981 12832 19993 12835
rect 19904 12804 19993 12832
rect 19981 12801 19993 12804
rect 20027 12801 20039 12835
rect 19981 12795 20039 12801
rect 20162 12792 20168 12844
rect 20220 12832 20226 12844
rect 20444 12835 20502 12841
rect 20444 12832 20456 12835
rect 20220 12804 20456 12832
rect 20220 12792 20226 12804
rect 20444 12801 20456 12804
rect 20490 12801 20502 12835
rect 20444 12795 20502 12801
rect 20622 12792 20628 12844
rect 20680 12832 20686 12844
rect 22572 12832 22600 12860
rect 20680 12804 22600 12832
rect 23124 12832 23152 12940
rect 23750 12928 23756 12980
rect 23808 12968 23814 12980
rect 24946 12968 24952 12980
rect 23808 12940 24952 12968
rect 23808 12928 23814 12940
rect 24946 12928 24952 12940
rect 25004 12928 25010 12980
rect 25590 12928 25596 12980
rect 25648 12928 25654 12980
rect 25682 12928 25688 12980
rect 25740 12928 25746 12980
rect 27154 12968 27160 12980
rect 26068 12940 27160 12968
rect 25608 12900 25636 12928
rect 26068 12900 26096 12940
rect 27154 12928 27160 12940
rect 27212 12928 27218 12980
rect 29914 12928 29920 12980
rect 29972 12928 29978 12980
rect 30374 12928 30380 12980
rect 30432 12928 30438 12980
rect 25608 12872 26096 12900
rect 27706 12860 27712 12912
rect 27764 12900 27770 12912
rect 27764 12872 30604 12900
rect 27764 12860 27770 12872
rect 23124 12804 23980 12832
rect 20680 12792 20686 12804
rect 19337 12767 19395 12773
rect 19337 12733 19349 12767
rect 19383 12764 19395 12767
rect 19426 12764 19432 12776
rect 19383 12736 19432 12764
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 19426 12724 19432 12736
rect 19484 12764 19490 12776
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 19484 12736 19625 12764
rect 19484 12724 19490 12736
rect 19613 12733 19625 12736
rect 19659 12733 19671 12767
rect 19613 12727 19671 12733
rect 19889 12767 19947 12773
rect 19889 12733 19901 12767
rect 19935 12764 19947 12767
rect 20070 12764 20076 12776
rect 19935 12736 20076 12764
rect 19935 12733 19947 12736
rect 19889 12727 19947 12733
rect 20070 12724 20076 12736
rect 20128 12724 20134 12776
rect 20254 12724 20260 12776
rect 20312 12764 20318 12776
rect 20717 12767 20775 12773
rect 20717 12764 20729 12767
rect 20312 12736 20729 12764
rect 20312 12724 20318 12736
rect 20717 12733 20729 12736
rect 20763 12733 20775 12767
rect 20717 12727 20775 12733
rect 22373 12767 22431 12773
rect 22373 12733 22385 12767
rect 22419 12764 22431 12767
rect 22572 12764 22600 12804
rect 22419 12736 22600 12764
rect 22419 12733 22431 12736
rect 22373 12727 22431 12733
rect 22572 12696 22600 12736
rect 22922 12724 22928 12776
rect 22980 12724 22986 12776
rect 23385 12767 23443 12773
rect 23385 12733 23397 12767
rect 23431 12733 23443 12767
rect 23385 12727 23443 12733
rect 23661 12767 23719 12773
rect 23661 12733 23673 12767
rect 23707 12764 23719 12767
rect 23750 12764 23756 12776
rect 23707 12736 23756 12764
rect 23707 12733 23719 12736
rect 23661 12727 23719 12733
rect 23400 12696 23428 12727
rect 23750 12724 23756 12736
rect 23808 12724 23814 12776
rect 23842 12724 23848 12776
rect 23900 12724 23906 12776
rect 23952 12764 23980 12804
rect 24026 12792 24032 12844
rect 24084 12832 24090 12844
rect 24308 12835 24366 12841
rect 24308 12832 24320 12835
rect 24084 12804 24320 12832
rect 24084 12792 24090 12804
rect 24308 12801 24320 12804
rect 24354 12801 24366 12835
rect 24308 12795 24366 12801
rect 25590 12792 25596 12844
rect 25648 12832 25654 12844
rect 26516 12835 26574 12841
rect 26516 12832 26528 12835
rect 25648 12804 26528 12832
rect 25648 12792 25654 12804
rect 26516 12801 26528 12804
rect 26562 12801 26574 12835
rect 26516 12795 26574 12801
rect 26694 12792 26700 12844
rect 26752 12832 26758 12844
rect 26789 12835 26847 12841
rect 26789 12832 26801 12835
rect 26752 12804 26801 12832
rect 26752 12792 26758 12804
rect 26789 12801 26801 12804
rect 26835 12801 26847 12835
rect 26789 12795 26847 12801
rect 27154 12792 27160 12844
rect 27212 12832 27218 12844
rect 30282 12832 30288 12844
rect 27212 12804 30288 12832
rect 27212 12792 27218 12804
rect 30282 12792 30288 12804
rect 30340 12792 30346 12844
rect 24581 12767 24639 12773
rect 24581 12764 24593 12767
rect 23952 12736 24593 12764
rect 24581 12733 24593 12736
rect 24627 12733 24639 12767
rect 24581 12727 24639 12733
rect 24854 12724 24860 12776
rect 24912 12764 24918 12776
rect 25866 12764 25872 12776
rect 24912 12736 25872 12764
rect 24912 12724 24918 12736
rect 25866 12724 25872 12736
rect 25924 12724 25930 12776
rect 26053 12767 26111 12773
rect 26053 12733 26065 12767
rect 26099 12764 26111 12767
rect 26418 12764 26424 12776
rect 26099 12736 26424 12764
rect 26099 12733 26111 12736
rect 26053 12727 26111 12733
rect 26418 12724 26424 12736
rect 26476 12724 26482 12776
rect 27982 12724 27988 12776
rect 28040 12764 28046 12776
rect 28353 12767 28411 12773
rect 28353 12764 28365 12767
rect 28040 12736 28365 12764
rect 28040 12724 28046 12736
rect 28353 12733 28365 12736
rect 28399 12764 28411 12767
rect 29457 12767 29515 12773
rect 29457 12764 29469 12767
rect 28399 12736 29469 12764
rect 28399 12733 28411 12736
rect 28353 12727 28411 12733
rect 29457 12733 29469 12736
rect 29503 12733 29515 12767
rect 30101 12767 30159 12773
rect 30101 12764 30113 12767
rect 29457 12727 29515 12733
rect 29564 12736 30113 12764
rect 17788 12668 20024 12696
rect 22572 12668 23428 12696
rect 16347 12665 16359 12668
rect 16301 12659 16359 12665
rect 19996 12640 20024 12668
rect 23566 12656 23572 12708
rect 23624 12696 23630 12708
rect 23934 12696 23940 12708
rect 23624 12668 23940 12696
rect 23624 12656 23630 12668
rect 23934 12656 23940 12668
rect 23992 12656 23998 12708
rect 25884 12696 25912 12724
rect 26142 12696 26148 12708
rect 25884 12668 26148 12696
rect 26142 12656 26148 12668
rect 26200 12656 26206 12708
rect 27522 12656 27528 12708
rect 27580 12696 27586 12708
rect 27580 12668 28488 12696
rect 27580 12656 27586 12668
rect 11388 12600 11652 12628
rect 11701 12631 11759 12637
rect 11388 12588 11394 12600
rect 11701 12597 11713 12631
rect 11747 12628 11759 12631
rect 11974 12628 11980 12640
rect 11747 12600 11980 12628
rect 11747 12597 11759 12600
rect 11701 12591 11759 12597
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13078 12628 13084 12640
rect 12943 12600 13084 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13078 12588 13084 12600
rect 13136 12588 13142 12640
rect 14007 12631 14065 12637
rect 14007 12597 14019 12631
rect 14053 12628 14065 12631
rect 14182 12628 14188 12640
rect 14053 12600 14188 12628
rect 14053 12597 14065 12600
rect 14007 12591 14065 12597
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 16850 12588 16856 12640
rect 16908 12637 16914 12640
rect 16908 12591 16917 12637
rect 16908 12588 16914 12591
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 18782 12628 18788 12640
rect 17460 12600 18788 12628
rect 17460 12588 17466 12600
rect 18782 12588 18788 12600
rect 18840 12588 18846 12640
rect 18874 12588 18880 12640
rect 18932 12588 18938 12640
rect 19153 12631 19211 12637
rect 19153 12597 19165 12631
rect 19199 12628 19211 12631
rect 19334 12628 19340 12640
rect 19199 12600 19340 12628
rect 19199 12597 19211 12600
rect 19153 12591 19211 12597
rect 19334 12588 19340 12600
rect 19392 12588 19398 12640
rect 19429 12631 19487 12637
rect 19429 12597 19441 12631
rect 19475 12628 19487 12631
rect 19794 12628 19800 12640
rect 19475 12600 19800 12628
rect 19475 12597 19487 12600
rect 19429 12591 19487 12597
rect 19794 12588 19800 12600
rect 19852 12588 19858 12640
rect 19978 12588 19984 12640
rect 20036 12588 20042 12640
rect 20447 12631 20505 12637
rect 20447 12597 20459 12631
rect 20493 12628 20505 12631
rect 20806 12628 20812 12640
rect 20493 12600 20812 12628
rect 20493 12597 20505 12600
rect 20447 12591 20505 12597
rect 20806 12588 20812 12600
rect 20864 12628 20870 12640
rect 22002 12628 22008 12640
rect 20864 12600 22008 12628
rect 20864 12588 20870 12600
rect 22002 12588 22008 12600
rect 22060 12588 22066 12640
rect 22830 12588 22836 12640
rect 22888 12628 22894 12640
rect 23201 12631 23259 12637
rect 23201 12628 23213 12631
rect 22888 12600 23213 12628
rect 22888 12588 22894 12600
rect 23201 12597 23213 12600
rect 23247 12597 23259 12631
rect 23201 12591 23259 12597
rect 23477 12631 23535 12637
rect 23477 12597 23489 12631
rect 23523 12628 23535 12631
rect 24118 12628 24124 12640
rect 23523 12600 24124 12628
rect 23523 12597 23535 12600
rect 23477 12591 23535 12597
rect 24118 12588 24124 12600
rect 24176 12588 24182 12640
rect 24302 12588 24308 12640
rect 24360 12637 24366 12640
rect 24360 12628 24369 12637
rect 26519 12631 26577 12637
rect 24360 12600 24405 12628
rect 24360 12591 24369 12600
rect 26519 12597 26531 12631
rect 26565 12628 26577 12631
rect 26878 12628 26884 12640
rect 26565 12600 26884 12628
rect 26565 12597 26577 12600
rect 26519 12591 26577 12597
rect 24360 12588 24366 12591
rect 26878 12588 26884 12600
rect 26936 12588 26942 12640
rect 27430 12588 27436 12640
rect 27488 12628 27494 12640
rect 28460 12637 28488 12668
rect 28994 12656 29000 12708
rect 29052 12696 29058 12708
rect 29089 12699 29147 12705
rect 29089 12696 29101 12699
rect 29052 12668 29101 12696
rect 29052 12656 29058 12668
rect 29089 12665 29101 12668
rect 29135 12665 29147 12699
rect 29089 12659 29147 12665
rect 29178 12656 29184 12708
rect 29236 12696 29242 12708
rect 29564 12696 29592 12736
rect 30101 12733 30113 12736
rect 30147 12764 30159 12767
rect 30374 12764 30380 12776
rect 30147 12736 30380 12764
rect 30147 12733 30159 12736
rect 30101 12727 30159 12733
rect 30374 12724 30380 12736
rect 30432 12724 30438 12776
rect 30576 12773 30604 12872
rect 30561 12767 30619 12773
rect 30561 12733 30573 12767
rect 30607 12733 30619 12767
rect 30561 12727 30619 12733
rect 29236 12668 29592 12696
rect 29236 12656 29242 12668
rect 29638 12656 29644 12708
rect 29696 12656 29702 12708
rect 27893 12631 27951 12637
rect 27893 12628 27905 12631
rect 27488 12600 27905 12628
rect 27488 12588 27494 12600
rect 27893 12597 27905 12600
rect 27939 12597 27951 12631
rect 27893 12591 27951 12597
rect 28445 12631 28503 12637
rect 28445 12597 28457 12631
rect 28491 12597 28503 12631
rect 28445 12591 28503 12597
rect 29454 12588 29460 12640
rect 29512 12628 29518 12640
rect 29656 12628 29684 12656
rect 29512 12600 29684 12628
rect 29512 12588 29518 12600
rect 29730 12588 29736 12640
rect 29788 12588 29794 12640
rect 552 12538 31072 12560
rect 552 12486 7988 12538
rect 8040 12486 8052 12538
rect 8104 12486 8116 12538
rect 8168 12486 8180 12538
rect 8232 12486 8244 12538
rect 8296 12486 15578 12538
rect 15630 12486 15642 12538
rect 15694 12486 15706 12538
rect 15758 12486 15770 12538
rect 15822 12486 15834 12538
rect 15886 12486 23168 12538
rect 23220 12486 23232 12538
rect 23284 12486 23296 12538
rect 23348 12486 23360 12538
rect 23412 12486 23424 12538
rect 23476 12486 30758 12538
rect 30810 12486 30822 12538
rect 30874 12486 30886 12538
rect 30938 12486 30950 12538
rect 31002 12486 31014 12538
rect 31066 12486 31072 12538
rect 552 12464 31072 12486
rect 3142 12424 3148 12436
rect 1228 12396 3148 12424
rect 1228 12297 1256 12396
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 3234 12384 3240 12436
rect 3292 12424 3298 12436
rect 3786 12424 3792 12436
rect 3292 12396 3792 12424
rect 3292 12384 3298 12396
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 3970 12384 3976 12436
rect 4028 12433 4034 12436
rect 4028 12424 4037 12433
rect 4522 12424 4528 12436
rect 4028 12396 4528 12424
rect 4028 12387 4037 12396
rect 4028 12384 4034 12387
rect 4522 12384 4528 12396
rect 4580 12384 4586 12436
rect 5537 12427 5595 12433
rect 5537 12393 5549 12427
rect 5583 12424 5595 12427
rect 5626 12424 5632 12436
rect 5583 12396 5632 12424
rect 5583 12393 5595 12396
rect 5537 12387 5595 12393
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 5718 12384 5724 12436
rect 5776 12384 5782 12436
rect 5902 12384 5908 12436
rect 5960 12384 5966 12436
rect 6270 12384 6276 12436
rect 6328 12424 6334 12436
rect 8294 12424 8300 12436
rect 6328 12396 8300 12424
rect 6328 12384 6334 12396
rect 8294 12384 8300 12396
rect 8352 12384 8358 12436
rect 8478 12384 8484 12436
rect 8536 12424 8542 12436
rect 8536 12396 10088 12424
rect 8536 12384 8542 12396
rect 1213 12291 1271 12297
rect 1213 12257 1225 12291
rect 1259 12257 1271 12291
rect 1213 12251 1271 12257
rect 1302 12248 1308 12300
rect 1360 12248 1366 12300
rect 1670 12297 1676 12300
rect 1632 12291 1676 12297
rect 1632 12257 1644 12291
rect 1632 12251 1676 12257
rect 1670 12248 1676 12251
rect 1728 12248 1734 12300
rect 3421 12291 3479 12297
rect 3421 12257 3433 12291
rect 3467 12288 3479 12291
rect 5736 12288 5764 12384
rect 5920 12356 5948 12384
rect 10060 12356 10088 12396
rect 11238 12384 11244 12436
rect 11296 12384 11302 12436
rect 12158 12424 12164 12436
rect 11348 12396 12164 12424
rect 11348 12356 11376 12396
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 12894 12424 12900 12436
rect 12268 12396 12900 12424
rect 12268 12356 12296 12396
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 13262 12384 13268 12436
rect 13320 12424 13326 12436
rect 14182 12424 14188 12436
rect 13320 12396 14188 12424
rect 13320 12384 13326 12396
rect 14182 12384 14188 12396
rect 14240 12424 14246 12436
rect 14240 12396 14964 12424
rect 14240 12384 14246 12396
rect 14936 12365 14964 12396
rect 15194 12384 15200 12436
rect 15252 12424 15258 12436
rect 15381 12427 15439 12433
rect 15381 12424 15393 12427
rect 15252 12396 15393 12424
rect 15252 12384 15258 12396
rect 15381 12393 15393 12396
rect 15427 12393 15439 12427
rect 15381 12387 15439 12393
rect 15930 12384 15936 12436
rect 15988 12424 15994 12436
rect 16301 12427 16359 12433
rect 16301 12424 16313 12427
rect 15988 12396 16313 12424
rect 15988 12384 15994 12396
rect 16301 12393 16313 12396
rect 16347 12393 16359 12427
rect 16301 12387 16359 12393
rect 16574 12384 16580 12436
rect 16632 12424 16638 12436
rect 16669 12427 16727 12433
rect 16669 12424 16681 12427
rect 16632 12396 16681 12424
rect 16632 12384 16638 12396
rect 16669 12393 16681 12396
rect 16715 12393 16727 12427
rect 19058 12424 19064 12436
rect 16669 12387 16727 12393
rect 17236 12396 19064 12424
rect 5920 12328 6598 12356
rect 10060 12328 11376 12356
rect 11440 12328 11928 12356
rect 5997 12291 6055 12297
rect 5997 12288 6009 12291
rect 3467 12260 4016 12288
rect 5736 12260 6009 12288
rect 3467 12257 3479 12260
rect 3421 12251 3479 12257
rect 1801 12241 1859 12247
rect 1801 12232 1813 12241
rect 1762 12180 1768 12232
rect 1847 12207 1859 12241
rect 1820 12201 1859 12207
rect 1820 12192 1844 12201
rect 1820 12180 1826 12192
rect 1946 12180 1952 12232
rect 2004 12220 2010 12232
rect 2041 12223 2099 12229
rect 2041 12220 2053 12223
rect 2004 12192 2053 12220
rect 2004 12180 2010 12192
rect 2041 12189 2053 12192
rect 2087 12189 2099 12223
rect 2041 12183 2099 12189
rect 3234 12180 3240 12232
rect 3292 12220 3298 12232
rect 3510 12220 3516 12232
rect 3292 12192 3516 12220
rect 3292 12180 3298 12192
rect 3510 12180 3516 12192
rect 3568 12220 3574 12232
rect 3878 12220 3884 12232
rect 3568 12192 3884 12220
rect 3568 12180 3574 12192
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 3988 12229 4016 12260
rect 5997 12257 6009 12260
rect 6043 12257 6055 12291
rect 5997 12251 6055 12257
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12288 6331 12291
rect 6362 12288 6368 12300
rect 6319 12260 6368 12288
rect 6319 12257 6331 12260
rect 6273 12251 6331 12257
rect 3976 12223 4034 12229
rect 3976 12189 3988 12223
rect 4022 12189 4034 12223
rect 3976 12183 4034 12189
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4249 12223 4307 12229
rect 4249 12220 4261 12223
rect 4120 12192 4261 12220
rect 4120 12180 4126 12192
rect 4249 12189 4261 12192
rect 4295 12189 4307 12223
rect 4249 12183 4307 12189
rect 5074 12180 5080 12232
rect 5132 12220 5138 12232
rect 6012 12220 6040 12251
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 6454 12248 6460 12300
rect 6512 12248 6518 12300
rect 6570 12288 6598 12328
rect 6570 12260 7052 12288
rect 6638 12220 6644 12232
rect 5132 12192 5856 12220
rect 6012 12192 6644 12220
rect 5132 12180 5138 12192
rect 3326 12112 3332 12164
rect 3384 12112 3390 12164
rect 5828 12161 5856 12192
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 6822 12229 6828 12232
rect 6784 12223 6828 12229
rect 6784 12189 6796 12223
rect 6784 12183 6828 12189
rect 6822 12180 6828 12183
rect 6880 12180 6886 12232
rect 6914 12180 6920 12232
rect 6972 12180 6978 12232
rect 7024 12220 7052 12260
rect 7098 12248 7104 12300
rect 7156 12288 7162 12300
rect 7193 12291 7251 12297
rect 7193 12288 7205 12291
rect 7156 12260 7205 12288
rect 7156 12248 7162 12260
rect 7193 12257 7205 12260
rect 7239 12257 7251 12291
rect 7193 12251 7251 12257
rect 7466 12248 7472 12300
rect 7524 12288 7530 12300
rect 8992 12291 9050 12297
rect 7524 12260 8892 12288
rect 7524 12248 7530 12260
rect 8864 12232 8892 12260
rect 8992 12257 9004 12291
rect 9038 12288 9050 12291
rect 9858 12288 9864 12300
rect 9038 12260 9864 12288
rect 9038 12257 9050 12260
rect 8992 12251 9050 12257
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 11146 12248 11152 12300
rect 11204 12248 11210 12300
rect 11440 12297 11468 12328
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12257 11483 12291
rect 11425 12251 11483 12257
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12288 11759 12291
rect 11790 12288 11796 12300
rect 11747 12260 11796 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 8570 12220 8576 12232
rect 7024 12192 8576 12220
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 8665 12223 8723 12229
rect 8665 12189 8677 12223
rect 8711 12189 8723 12223
rect 8665 12183 8723 12189
rect 5813 12155 5871 12161
rect 5813 12121 5825 12155
rect 5859 12121 5871 12155
rect 5813 12115 5871 12121
rect 6178 12112 6184 12164
rect 6236 12112 6242 12164
rect 1029 12087 1087 12093
rect 1029 12053 1041 12087
rect 1075 12084 1087 12087
rect 1946 12084 1952 12096
rect 1075 12056 1952 12084
rect 1075 12053 1087 12056
rect 1029 12047 1087 12053
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 3344 12084 3372 12112
rect 4062 12084 4068 12096
rect 3344 12056 4068 12084
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 6086 12044 6092 12096
rect 6144 12044 6150 12096
rect 6196 12084 6224 12112
rect 8018 12084 8024 12096
rect 6196 12056 8024 12084
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8478 12044 8484 12096
rect 8536 12044 8542 12096
rect 8680 12084 8708 12183
rect 8846 12180 8852 12232
rect 8904 12180 8910 12232
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12220 9459 12223
rect 11900 12220 11928 12328
rect 11992 12328 12296 12356
rect 14921 12359 14979 12365
rect 11992 12297 12020 12328
rect 14921 12325 14933 12359
rect 14967 12325 14979 12359
rect 14921 12319 14979 12325
rect 11977 12291 12035 12297
rect 11977 12257 11989 12291
rect 12023 12257 12035 12291
rect 11977 12251 12035 12257
rect 12066 12248 12072 12300
rect 12124 12248 12130 12300
rect 12345 12291 12403 12297
rect 12345 12257 12357 12291
rect 12391 12257 12403 12291
rect 12345 12251 12403 12257
rect 12084 12220 12112 12248
rect 12360 12220 12388 12251
rect 12434 12248 12440 12300
rect 12492 12248 12498 12300
rect 12802 12297 12808 12300
rect 12764 12291 12808 12297
rect 12764 12257 12776 12291
rect 12860 12288 12866 12300
rect 13173 12291 13231 12297
rect 12860 12260 13124 12288
rect 12764 12251 12808 12257
rect 12802 12248 12808 12251
rect 12860 12248 12866 12260
rect 9447 12192 11560 12220
rect 11900 12192 12388 12220
rect 9447 12189 9459 12192
rect 9401 12183 9459 12189
rect 10686 12112 10692 12164
rect 10744 12112 10750 12164
rect 11532 12161 11560 12192
rect 12618 12180 12624 12232
rect 12676 12220 12682 12232
rect 12900 12223 12958 12229
rect 12900 12220 12912 12223
rect 12676 12192 12912 12220
rect 12676 12180 12682 12192
rect 12900 12189 12912 12192
rect 12946 12189 12958 12223
rect 13096 12220 13124 12260
rect 13173 12257 13185 12291
rect 13219 12288 13231 12291
rect 13219 12260 13400 12288
rect 13219 12257 13231 12260
rect 13173 12251 13231 12257
rect 13372 12232 13400 12260
rect 13446 12248 13452 12300
rect 13504 12288 13510 12300
rect 14645 12291 14703 12297
rect 14645 12288 14657 12291
rect 13504 12260 14657 12288
rect 13504 12248 13510 12260
rect 14645 12257 14657 12260
rect 14691 12257 14703 12291
rect 14645 12251 14703 12257
rect 14826 12248 14832 12300
rect 14884 12288 14890 12300
rect 17236 12297 17264 12396
rect 19058 12384 19064 12396
rect 19116 12424 19122 12436
rect 19981 12427 20039 12433
rect 19116 12396 19932 12424
rect 19116 12384 19122 12396
rect 19904 12356 19932 12396
rect 19981 12393 19993 12427
rect 20027 12424 20039 12427
rect 20162 12424 20168 12436
rect 20027 12396 20168 12424
rect 20027 12393 20039 12396
rect 19981 12387 20039 12393
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 20254 12384 20260 12436
rect 20312 12384 20318 12436
rect 20622 12384 20628 12436
rect 20680 12384 20686 12436
rect 20717 12427 20775 12433
rect 20717 12393 20729 12427
rect 20763 12393 20775 12427
rect 20717 12387 20775 12393
rect 21735 12427 21793 12433
rect 21735 12393 21747 12427
rect 21781 12424 21793 12427
rect 22002 12424 22008 12436
rect 21781 12396 22008 12424
rect 21781 12393 21793 12396
rect 21735 12387 21793 12393
rect 20640 12356 20668 12384
rect 19904 12328 20668 12356
rect 20732 12356 20760 12387
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 23106 12384 23112 12436
rect 23164 12384 23170 12436
rect 23842 12424 23848 12436
rect 23492 12396 23848 12424
rect 20732 12328 21404 12356
rect 17221 12291 17279 12297
rect 17221 12288 17233 12291
rect 14884 12260 17233 12288
rect 14884 12248 14890 12260
rect 17221 12257 17233 12260
rect 17267 12257 17279 12291
rect 17221 12251 17279 12257
rect 17402 12248 17408 12300
rect 17460 12248 17466 12300
rect 17681 12291 17739 12297
rect 17681 12257 17693 12291
rect 17727 12288 17739 12291
rect 18284 12291 18342 12297
rect 18284 12288 18296 12291
rect 17727 12260 18296 12288
rect 17727 12257 17739 12260
rect 17681 12251 17739 12257
rect 18284 12257 18296 12260
rect 18330 12288 18342 12291
rect 18330 12260 18644 12288
rect 18330 12257 18342 12260
rect 18284 12251 18342 12257
rect 13262 12220 13268 12232
rect 13096 12192 13268 12220
rect 12900 12183 12958 12189
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 13354 12180 13360 12232
rect 13412 12180 13418 12232
rect 14274 12220 14280 12232
rect 14019 12192 14280 12220
rect 11517 12155 11575 12161
rect 11517 12121 11529 12155
rect 11563 12121 11575 12155
rect 11517 12115 11575 12121
rect 9398 12084 9404 12096
rect 8680 12056 9404 12084
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 10965 12087 11023 12093
rect 10965 12084 10977 12087
rect 10652 12056 10977 12084
rect 10652 12044 10658 12056
rect 10965 12053 10977 12056
rect 11011 12053 11023 12087
rect 10965 12047 11023 12053
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 11793 12087 11851 12093
rect 11793 12084 11805 12087
rect 11112 12056 11805 12084
rect 11112 12044 11118 12056
rect 11793 12053 11805 12056
rect 11839 12053 11851 12087
rect 11793 12047 11851 12053
rect 12161 12087 12219 12093
rect 12161 12053 12173 12087
rect 12207 12084 12219 12087
rect 14019 12084 14047 12192
rect 14274 12180 14280 12192
rect 14332 12180 14338 12232
rect 15838 12180 15844 12232
rect 15896 12180 15902 12232
rect 16574 12180 16580 12232
rect 16632 12220 16638 12232
rect 17862 12220 17868 12232
rect 16632 12192 17868 12220
rect 16632 12180 16638 12192
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 17954 12180 17960 12232
rect 18012 12180 18018 12232
rect 18414 12180 18420 12232
rect 18472 12180 18478 12232
rect 18616 12220 18644 12260
rect 18690 12248 18696 12300
rect 18748 12248 18754 12300
rect 20441 12291 20499 12297
rect 20441 12257 20453 12291
rect 20487 12288 20499 12291
rect 20640 12288 20668 12328
rect 20487 12260 20668 12288
rect 20901 12291 20959 12297
rect 20487 12257 20499 12260
rect 20441 12251 20499 12257
rect 20901 12257 20913 12291
rect 20947 12288 20959 12291
rect 21174 12288 21180 12300
rect 20947 12260 21180 12288
rect 20947 12257 20959 12260
rect 20901 12251 20959 12257
rect 21174 12248 21180 12260
rect 21232 12248 21238 12300
rect 21376 12288 21404 12328
rect 23492 12297 23520 12396
rect 23842 12384 23848 12396
rect 23900 12424 23906 12436
rect 25501 12427 25559 12433
rect 23900 12396 24900 12424
rect 23900 12384 23906 12396
rect 24872 12356 24900 12396
rect 25501 12393 25513 12427
rect 25547 12424 25559 12427
rect 25590 12424 25596 12436
rect 25547 12396 25596 12424
rect 25547 12393 25559 12396
rect 25501 12387 25559 12393
rect 25590 12384 25596 12396
rect 25648 12384 25654 12436
rect 25774 12384 25780 12436
rect 25832 12424 25838 12436
rect 27522 12424 27528 12436
rect 25832 12396 27528 12424
rect 25832 12384 25838 12396
rect 27522 12384 27528 12396
rect 27580 12384 27586 12436
rect 27614 12384 27620 12436
rect 27672 12424 27678 12436
rect 28261 12427 28319 12433
rect 28261 12424 28273 12427
rect 27672 12396 28273 12424
rect 27672 12384 27678 12396
rect 28261 12393 28273 12396
rect 28307 12393 28319 12427
rect 28261 12387 28319 12393
rect 28442 12384 28448 12436
rect 28500 12424 28506 12436
rect 30377 12427 30435 12433
rect 30377 12424 30389 12427
rect 28500 12396 30389 12424
rect 28500 12384 28506 12396
rect 30377 12393 30389 12396
rect 30423 12393 30435 12427
rect 30377 12387 30435 12393
rect 24872 12328 26464 12356
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 21376 12260 22017 12288
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 23477 12291 23535 12297
rect 23477 12257 23489 12291
rect 23523 12257 23535 12291
rect 23477 12251 23535 12257
rect 23804 12291 23862 12297
rect 23804 12257 23816 12291
rect 23850 12288 23862 12291
rect 23850 12260 24072 12288
rect 23850 12257 23862 12260
rect 23804 12251 23862 12257
rect 19058 12220 19064 12232
rect 18616 12192 19064 12220
rect 19058 12180 19064 12192
rect 19116 12180 19122 12232
rect 19886 12180 19892 12232
rect 19944 12220 19950 12232
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 19944 12192 21281 12220
rect 19944 12180 19950 12192
rect 21269 12189 21281 12192
rect 21315 12220 21327 12223
rect 21542 12220 21548 12232
rect 21315 12192 21548 12220
rect 21315 12189 21327 12192
rect 21269 12183 21327 12189
rect 21542 12180 21548 12192
rect 21600 12180 21606 12232
rect 21818 12229 21824 12232
rect 21775 12223 21824 12229
rect 21775 12189 21787 12223
rect 21821 12189 21824 12223
rect 21775 12183 21824 12189
rect 21818 12180 21824 12183
rect 21876 12180 21882 12232
rect 23934 12180 23940 12232
rect 23992 12180 23998 12232
rect 24044 12220 24072 12260
rect 24118 12248 24124 12300
rect 24176 12288 24182 12300
rect 24213 12291 24271 12297
rect 24213 12288 24225 12291
rect 24176 12260 24225 12288
rect 24176 12248 24182 12260
rect 24213 12257 24225 12260
rect 24259 12257 24271 12291
rect 24213 12251 24271 12257
rect 25774 12248 25780 12300
rect 25832 12248 25838 12300
rect 26436 12297 26464 12328
rect 26421 12291 26479 12297
rect 26421 12257 26433 12291
rect 26467 12288 26479 12291
rect 26510 12288 26516 12300
rect 26467 12260 26516 12288
rect 26467 12257 26479 12260
rect 26421 12251 26479 12257
rect 26510 12248 26516 12260
rect 26568 12288 26574 12300
rect 26568 12260 27016 12288
rect 26568 12248 26574 12260
rect 24302 12220 24308 12232
rect 24044 12192 24308 12220
rect 24302 12180 24308 12192
rect 24360 12220 24366 12232
rect 26748 12223 26806 12229
rect 26748 12220 26760 12223
rect 24360 12192 26760 12220
rect 24360 12180 24366 12192
rect 12207 12056 14047 12084
rect 12207 12053 12219 12056
rect 12161 12047 12219 12053
rect 14090 12044 14096 12096
rect 14148 12084 14154 12096
rect 14277 12087 14335 12093
rect 14277 12084 14289 12087
rect 14148 12056 14289 12084
rect 14148 12044 14154 12056
rect 14277 12053 14289 12056
rect 14323 12053 14335 12087
rect 14277 12047 14335 12053
rect 17034 12044 17040 12096
rect 17092 12044 17098 12096
rect 18322 12044 18328 12096
rect 18380 12084 18386 12096
rect 19426 12084 19432 12096
rect 18380 12056 19432 12084
rect 18380 12044 18386 12056
rect 19426 12044 19432 12056
rect 19484 12044 19490 12096
rect 20990 12044 20996 12096
rect 21048 12084 21054 12096
rect 25774 12084 25780 12096
rect 21048 12056 25780 12084
rect 21048 12044 21054 12056
rect 25774 12044 25780 12056
rect 25832 12044 25838 12096
rect 26053 12087 26111 12093
rect 26053 12053 26065 12087
rect 26099 12084 26111 12087
rect 26326 12084 26332 12096
rect 26099 12056 26332 12084
rect 26099 12053 26111 12056
rect 26053 12047 26111 12053
rect 26326 12044 26332 12056
rect 26384 12044 26390 12096
rect 26436 12084 26464 12192
rect 26748 12189 26760 12192
rect 26794 12189 26806 12223
rect 26748 12183 26806 12189
rect 26878 12180 26884 12232
rect 26936 12180 26942 12232
rect 26988 12220 27016 12260
rect 27154 12248 27160 12300
rect 27212 12248 27218 12300
rect 27982 12288 27988 12300
rect 27264 12260 27988 12288
rect 27264 12220 27292 12260
rect 27982 12248 27988 12260
rect 28040 12248 28046 12300
rect 28902 12248 28908 12300
rect 28960 12248 28966 12300
rect 29730 12248 29736 12300
rect 29788 12288 29794 12300
rect 30561 12291 30619 12297
rect 30561 12288 30573 12291
rect 29788 12260 30573 12288
rect 29788 12248 29794 12260
rect 30561 12257 30573 12260
rect 30607 12257 30619 12291
rect 30561 12251 30619 12257
rect 26988 12192 27292 12220
rect 27798 12180 27804 12232
rect 27856 12220 27862 12232
rect 28629 12223 28687 12229
rect 28629 12220 28641 12223
rect 27856 12192 28641 12220
rect 27856 12180 27862 12192
rect 28629 12189 28641 12192
rect 28675 12189 28687 12223
rect 28629 12183 28687 12189
rect 28258 12112 28264 12164
rect 28316 12112 28322 12164
rect 27614 12084 27620 12096
rect 26436 12056 27620 12084
rect 27614 12044 27620 12056
rect 27672 12084 27678 12096
rect 28276 12084 28304 12112
rect 27672 12056 28304 12084
rect 27672 12044 27678 12056
rect 28902 12044 28908 12096
rect 28960 12084 28966 12096
rect 30009 12087 30067 12093
rect 30009 12084 30021 12087
rect 28960 12056 30021 12084
rect 28960 12044 28966 12056
rect 30009 12053 30021 12056
rect 30055 12053 30067 12087
rect 30009 12047 30067 12053
rect 552 11994 30912 12016
rect 552 11942 4193 11994
rect 4245 11942 4257 11994
rect 4309 11942 4321 11994
rect 4373 11942 4385 11994
rect 4437 11942 4449 11994
rect 4501 11942 11783 11994
rect 11835 11942 11847 11994
rect 11899 11942 11911 11994
rect 11963 11942 11975 11994
rect 12027 11942 12039 11994
rect 12091 11942 19373 11994
rect 19425 11942 19437 11994
rect 19489 11942 19501 11994
rect 19553 11942 19565 11994
rect 19617 11942 19629 11994
rect 19681 11942 26963 11994
rect 27015 11942 27027 11994
rect 27079 11942 27091 11994
rect 27143 11942 27155 11994
rect 27207 11942 27219 11994
rect 27271 11942 30912 11994
rect 552 11920 30912 11942
rect 1394 11840 1400 11892
rect 1452 11880 1458 11892
rect 2866 11880 2872 11892
rect 1452 11852 2872 11880
rect 1452 11840 1458 11852
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 6086 11880 6092 11892
rect 5092 11852 6092 11880
rect 1443 11747 1501 11753
rect 1443 11713 1455 11747
rect 1489 11744 1501 11747
rect 2038 11744 2044 11756
rect 1489 11716 2044 11744
rect 1489 11713 1501 11716
rect 1443 11707 1501 11713
rect 2038 11704 2044 11716
rect 2096 11704 2102 11756
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11744 3111 11747
rect 3510 11744 3516 11756
rect 3099 11716 3516 11744
rect 3099 11713 3111 11716
rect 3053 11707 3111 11713
rect 3510 11704 3516 11716
rect 3568 11704 3574 11756
rect 3792 11747 3850 11753
rect 3792 11744 3804 11747
rect 3620 11716 3804 11744
rect 3620 11688 3648 11716
rect 3792 11713 3804 11716
rect 3838 11713 3850 11747
rect 3792 11707 3850 11713
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11744 4123 11747
rect 5092 11744 5120 11852
rect 6086 11840 6092 11852
rect 6144 11840 6150 11892
rect 6914 11840 6920 11892
rect 6972 11840 6978 11892
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 8021 11883 8079 11889
rect 8021 11880 8033 11883
rect 7616 11852 8033 11880
rect 7616 11840 7622 11852
rect 8021 11849 8033 11852
rect 8067 11849 8079 11883
rect 8021 11843 8079 11849
rect 8570 11840 8576 11892
rect 8628 11880 8634 11892
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 8628 11852 8861 11880
rect 8628 11840 8634 11852
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 8849 11843 8907 11849
rect 9030 11840 9036 11892
rect 9088 11880 9094 11892
rect 9125 11883 9183 11889
rect 9125 11880 9137 11883
rect 9088 11852 9137 11880
rect 9088 11840 9094 11852
rect 9125 11849 9137 11852
rect 9171 11849 9183 11883
rect 9125 11843 9183 11849
rect 9401 11883 9459 11889
rect 9401 11849 9413 11883
rect 9447 11880 9459 11883
rect 9447 11852 9674 11880
rect 9447 11849 9459 11852
rect 9401 11843 9459 11849
rect 4111 11716 5120 11744
rect 5445 11747 5503 11753
rect 4111 11713 4123 11716
rect 4065 11707 4123 11713
rect 5445 11713 5457 11747
rect 5491 11744 5503 11747
rect 6000 11745 6058 11751
rect 5491 11716 5948 11744
rect 5491 11713 5503 11716
rect 5445 11707 5503 11713
rect 934 11636 940 11688
rect 992 11636 998 11688
rect 1670 11636 1676 11688
rect 1728 11636 1734 11688
rect 3234 11636 3240 11688
rect 3292 11676 3298 11688
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 3292 11648 3341 11676
rect 3292 11636 3298 11648
rect 3329 11645 3341 11648
rect 3375 11645 3387 11679
rect 3329 11639 3387 11645
rect 3602 11636 3608 11688
rect 3660 11636 3666 11688
rect 4706 11636 4712 11688
rect 4764 11676 4770 11688
rect 5534 11676 5540 11688
rect 4764 11648 5540 11676
rect 4764 11636 4770 11648
rect 5534 11636 5540 11648
rect 5592 11636 5598 11688
rect 5920 11676 5948 11716
rect 6000 11711 6012 11745
rect 6046 11744 6058 11745
rect 6086 11744 6092 11756
rect 6046 11716 6092 11744
rect 6046 11711 6058 11716
rect 6000 11705 6058 11711
rect 6086 11704 6092 11716
rect 6144 11704 6150 11756
rect 6932 11744 6960 11840
rect 9646 11824 9674 11852
rect 11514 11840 11520 11892
rect 11572 11840 11578 11892
rect 12342 11840 12348 11892
rect 12400 11840 12406 11892
rect 12805 11883 12863 11889
rect 12805 11849 12817 11883
rect 12851 11880 12863 11883
rect 12986 11880 12992 11892
rect 12851 11852 12992 11880
rect 12851 11849 12863 11852
rect 12805 11843 12863 11849
rect 12986 11840 12992 11852
rect 13044 11840 13050 11892
rect 13078 11840 13084 11892
rect 13136 11840 13142 11892
rect 18322 11880 18328 11892
rect 16316 11852 18328 11880
rect 9646 11784 9680 11824
rect 9674 11772 9680 11784
rect 9732 11772 9738 11824
rect 11330 11772 11336 11824
rect 11388 11812 11394 11824
rect 12710 11812 12716 11824
rect 11388 11784 12716 11812
rect 11388 11772 11394 11784
rect 12710 11772 12716 11784
rect 12768 11772 12774 11824
rect 6196 11716 6960 11744
rect 6196 11676 6224 11716
rect 7834 11704 7840 11756
rect 7892 11744 7898 11756
rect 7892 11716 8432 11744
rect 7892 11704 7898 11716
rect 5920 11648 6224 11676
rect 6270 11636 6276 11688
rect 6328 11636 6334 11688
rect 6638 11636 6644 11688
rect 6696 11676 6702 11688
rect 7929 11679 7987 11685
rect 7929 11676 7941 11679
rect 6696 11648 7941 11676
rect 6696 11636 6702 11648
rect 7929 11645 7941 11648
rect 7975 11645 7987 11679
rect 7929 11639 7987 11645
rect 8018 11636 8024 11688
rect 8076 11676 8082 11688
rect 8205 11679 8263 11685
rect 8205 11676 8217 11679
rect 8076 11648 8217 11676
rect 8076 11636 8082 11648
rect 8205 11645 8217 11648
rect 8251 11645 8263 11679
rect 8205 11639 8263 11645
rect 1403 11543 1461 11549
rect 1403 11509 1415 11543
rect 1449 11540 1461 11543
rect 2866 11540 2872 11552
rect 1449 11512 2872 11540
rect 1449 11509 1461 11512
rect 1403 11503 1461 11509
rect 2866 11500 2872 11512
rect 2924 11500 2930 11552
rect 3795 11543 3853 11549
rect 3795 11509 3807 11543
rect 3841 11540 3853 11543
rect 3970 11540 3976 11552
rect 3841 11512 3976 11540
rect 3841 11509 3853 11512
rect 3795 11503 3853 11509
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 5626 11540 5632 11552
rect 4120 11512 5632 11540
rect 4120 11500 4126 11512
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 6003 11543 6061 11549
rect 6003 11509 6015 11543
rect 6049 11540 6061 11543
rect 6730 11540 6736 11552
rect 6049 11512 6736 11540
rect 6049 11509 6061 11512
rect 6003 11503 6061 11509
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 7006 11500 7012 11552
rect 7064 11540 7070 11552
rect 7377 11543 7435 11549
rect 7377 11540 7389 11543
rect 7064 11512 7389 11540
rect 7064 11500 7070 11512
rect 7377 11509 7389 11512
rect 7423 11509 7435 11543
rect 7377 11503 7435 11509
rect 7558 11500 7564 11552
rect 7616 11540 7622 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 7616 11512 7757 11540
rect 7616 11500 7622 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 8220 11540 8248 11639
rect 8294 11636 8300 11688
rect 8352 11636 8358 11688
rect 8404 11676 8432 11716
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 10140 11747 10198 11753
rect 10140 11744 10152 11747
rect 8536 11716 10152 11744
rect 8536 11704 8542 11716
rect 10140 11713 10152 11716
rect 10186 11713 10198 11747
rect 10140 11707 10198 11713
rect 10413 11747 10471 11753
rect 10413 11713 10425 11747
rect 10459 11744 10471 11747
rect 10594 11744 10600 11756
rect 10459 11716 10600 11744
rect 10459 11713 10471 11716
rect 10413 11707 10471 11713
rect 10594 11704 10600 11716
rect 10652 11704 10658 11756
rect 10704 11716 13032 11744
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 8404 11648 8677 11676
rect 8665 11645 8677 11648
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 8754 11636 8760 11688
rect 8812 11676 8818 11688
rect 8941 11679 8999 11685
rect 8941 11676 8953 11679
rect 8812 11648 8953 11676
rect 8812 11636 8818 11648
rect 8941 11645 8953 11648
rect 8987 11645 8999 11679
rect 8941 11639 8999 11645
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11676 9275 11679
rect 9306 11676 9312 11688
rect 9263 11648 9312 11676
rect 9263 11645 9275 11648
rect 9217 11639 9275 11645
rect 9306 11636 9312 11648
rect 9364 11636 9370 11688
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 9677 11679 9735 11685
rect 9677 11676 9689 11679
rect 9456 11648 9689 11676
rect 9456 11636 9462 11648
rect 9677 11645 9689 11648
rect 9723 11645 9735 11679
rect 10704 11676 10732 11716
rect 9677 11639 9735 11645
rect 9784 11648 10732 11676
rect 8312 11608 8340 11636
rect 8389 11611 8447 11617
rect 8389 11608 8401 11611
rect 8312 11580 8401 11608
rect 8389 11577 8401 11580
rect 8435 11577 8447 11611
rect 9784 11608 9812 11648
rect 10778 11636 10784 11688
rect 10836 11676 10842 11688
rect 12069 11679 12127 11685
rect 10836 11648 11100 11676
rect 10836 11636 10842 11648
rect 8389 11571 8447 11577
rect 8772 11580 9812 11608
rect 11072 11608 11100 11648
rect 12069 11645 12081 11679
rect 12115 11676 12127 11679
rect 12250 11676 12256 11688
rect 12115 11648 12256 11676
rect 12115 11645 12127 11648
rect 12069 11639 12127 11645
rect 12250 11636 12256 11648
rect 12308 11636 12314 11688
rect 13004 11685 13032 11716
rect 13096 11688 13124 11840
rect 13170 11772 13176 11824
rect 13228 11812 13234 11824
rect 13357 11815 13415 11821
rect 13357 11812 13369 11815
rect 13228 11784 13369 11812
rect 13228 11772 13234 11784
rect 13357 11781 13369 11784
rect 13403 11781 13415 11815
rect 13357 11775 13415 11781
rect 13262 11704 13268 11756
rect 13320 11744 13326 11756
rect 13868 11747 13926 11753
rect 13868 11744 13880 11747
rect 13320 11716 13880 11744
rect 13320 11704 13326 11716
rect 13868 11713 13880 11716
rect 13914 11713 13926 11747
rect 13868 11707 13926 11713
rect 14047 11747 14105 11753
rect 14047 11713 14059 11747
rect 14093 11744 14105 11747
rect 14182 11744 14188 11756
rect 14093 11716 14188 11744
rect 14093 11713 14105 11716
rect 14047 11707 14105 11713
rect 14182 11704 14188 11716
rect 14240 11704 14246 11756
rect 14274 11704 14280 11756
rect 14332 11704 14338 11756
rect 12989 11679 13047 11685
rect 12989 11645 13001 11679
rect 13035 11645 13047 11679
rect 12989 11639 13047 11645
rect 13078 11636 13084 11688
rect 13136 11636 13142 11688
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11676 13231 11679
rect 13219 11648 13400 11676
rect 13219 11645 13231 11648
rect 13173 11639 13231 11645
rect 13372 11608 13400 11648
rect 13538 11636 13544 11688
rect 13596 11636 13602 11688
rect 13630 11636 13636 11688
rect 13688 11636 13694 11688
rect 15838 11676 15844 11688
rect 14936 11648 15844 11676
rect 13648 11608 13676 11636
rect 11072 11580 13308 11608
rect 13372 11580 13676 11608
rect 8772 11540 8800 11580
rect 8220 11512 8800 11540
rect 7745 11503 7803 11509
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 9950 11540 9956 11552
rect 8904 11512 9956 11540
rect 8904 11500 8910 11512
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 10042 11500 10048 11552
rect 10100 11540 10106 11552
rect 10143 11543 10201 11549
rect 10143 11540 10155 11543
rect 10100 11512 10155 11540
rect 10100 11500 10106 11512
rect 10143 11509 10155 11512
rect 10189 11509 10201 11543
rect 10143 11503 10201 11509
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 11885 11543 11943 11549
rect 11885 11540 11897 11543
rect 10376 11512 11897 11540
rect 10376 11500 10382 11512
rect 11885 11509 11897 11512
rect 11931 11509 11943 11543
rect 13280 11540 13308 11580
rect 14936 11540 14964 11648
rect 15838 11636 15844 11648
rect 15896 11636 15902 11688
rect 16316 11685 16344 11852
rect 18322 11840 18328 11852
rect 18380 11840 18386 11892
rect 18414 11840 18420 11892
rect 18472 11840 18478 11892
rect 18708 11852 20490 11880
rect 17862 11772 17868 11824
rect 17920 11812 17926 11824
rect 18708 11812 18736 11852
rect 17920 11784 18736 11812
rect 20462 11812 20490 11852
rect 20530 11840 20536 11892
rect 20588 11840 20594 11892
rect 21542 11840 21548 11892
rect 21600 11880 21606 11892
rect 23569 11883 23627 11889
rect 21600 11852 22968 11880
rect 21600 11840 21606 11852
rect 20990 11812 20996 11824
rect 20462 11784 20996 11812
rect 17920 11772 17926 11784
rect 20990 11772 20996 11784
rect 21048 11772 21054 11824
rect 16899 11745 16957 11751
rect 16899 11711 16911 11745
rect 16945 11711 16957 11745
rect 16899 11705 16957 11711
rect 16301 11679 16359 11685
rect 16301 11645 16313 11679
rect 16347 11645 16359 11679
rect 16301 11639 16359 11645
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11676 16451 11679
rect 16666 11676 16672 11688
rect 16439 11648 16672 11676
rect 16439 11645 16451 11648
rect 16393 11639 16451 11645
rect 16666 11636 16672 11648
rect 16724 11636 16730 11688
rect 16914 11676 16942 11705
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 17092 11716 17141 11744
rect 17092 11704 17098 11716
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 18690 11744 18696 11756
rect 18012 11716 18696 11744
rect 18012 11704 18018 11716
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 19156 11747 19214 11753
rect 19156 11744 19168 11747
rect 18800 11716 19168 11744
rect 17862 11676 17868 11688
rect 16914 11648 17868 11676
rect 17862 11636 17868 11648
rect 17920 11636 17926 11688
rect 18800 11552 18828 11716
rect 19156 11713 19168 11716
rect 19202 11713 19214 11747
rect 19156 11707 19214 11713
rect 19334 11704 19340 11756
rect 19392 11744 19398 11756
rect 21560 11753 21588 11840
rect 22940 11812 22968 11852
rect 23569 11849 23581 11883
rect 23615 11880 23627 11883
rect 23934 11880 23940 11892
rect 23615 11852 23940 11880
rect 23615 11849 23627 11852
rect 23569 11843 23627 11849
rect 23934 11840 23940 11852
rect 23992 11840 23998 11892
rect 25682 11880 25688 11892
rect 24504 11852 25688 11880
rect 24504 11812 24532 11852
rect 25682 11840 25688 11852
rect 25740 11840 25746 11892
rect 26513 11883 26571 11889
rect 26513 11849 26525 11883
rect 26559 11880 26571 11883
rect 26878 11880 26884 11892
rect 26559 11852 26884 11880
rect 26559 11849 26571 11852
rect 26513 11843 26571 11849
rect 26878 11840 26884 11852
rect 26936 11840 26942 11892
rect 26970 11840 26976 11892
rect 27028 11880 27034 11892
rect 28721 11883 28779 11889
rect 27028 11852 28672 11880
rect 27028 11840 27034 11852
rect 22940 11784 24532 11812
rect 19429 11747 19487 11753
rect 19429 11744 19441 11747
rect 19392 11716 19441 11744
rect 19392 11704 19398 11716
rect 19429 11713 19441 11716
rect 19475 11713 19487 11747
rect 19429 11707 19487 11713
rect 21545 11747 21603 11753
rect 21545 11713 21557 11747
rect 21591 11713 21603 11747
rect 21545 11707 21603 11713
rect 22051 11747 22109 11753
rect 22051 11713 22063 11747
rect 22097 11744 22109 11747
rect 24213 11747 24271 11753
rect 22097 11716 22968 11744
rect 22097 11713 22109 11716
rect 22051 11707 22109 11713
rect 22940 11688 22968 11716
rect 24213 11713 24225 11747
rect 24259 11744 24271 11747
rect 24302 11744 24308 11756
rect 24259 11716 24308 11744
rect 24259 11713 24271 11716
rect 24213 11707 24271 11713
rect 24302 11704 24308 11716
rect 24360 11704 24366 11756
rect 24504 11753 24532 11784
rect 28442 11772 28448 11824
rect 28500 11772 28506 11824
rect 28644 11812 28672 11852
rect 28721 11849 28733 11883
rect 28767 11880 28779 11883
rect 28810 11880 28816 11892
rect 28767 11852 28816 11880
rect 28767 11849 28779 11852
rect 28721 11843 28779 11849
rect 28810 11840 28816 11852
rect 28868 11840 28874 11892
rect 29546 11812 29552 11824
rect 28644 11784 29552 11812
rect 29546 11772 29552 11784
rect 29604 11772 29610 11824
rect 30101 11815 30159 11821
rect 30101 11781 30113 11815
rect 30147 11781 30159 11815
rect 30101 11775 30159 11781
rect 24489 11747 24547 11753
rect 24489 11713 24501 11747
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 24995 11747 25053 11753
rect 24995 11713 25007 11747
rect 25041 11744 25053 11747
rect 25041 11716 25544 11744
rect 25041 11713 25053 11716
rect 24995 11707 25053 11713
rect 25516 11688 25544 11716
rect 26510 11704 26516 11756
rect 26568 11744 26574 11756
rect 26697 11747 26755 11753
rect 26697 11744 26709 11747
rect 26568 11716 26709 11744
rect 26568 11704 26574 11716
rect 26697 11713 26709 11716
rect 26743 11713 26755 11747
rect 26697 11707 26755 11713
rect 27203 11747 27261 11753
rect 27203 11713 27215 11747
rect 27249 11744 27261 11747
rect 27433 11747 27491 11753
rect 27249 11716 27384 11744
rect 27249 11713 27261 11716
rect 27203 11707 27261 11713
rect 19886 11636 19892 11688
rect 19944 11676 19950 11688
rect 21174 11676 21180 11688
rect 19944 11648 21180 11676
rect 19944 11636 19950 11648
rect 21174 11636 21180 11648
rect 21232 11636 21238 11688
rect 22278 11636 22284 11688
rect 22336 11636 22342 11688
rect 22922 11636 22928 11688
rect 22980 11636 22986 11688
rect 23934 11636 23940 11688
rect 23992 11676 23998 11688
rect 24854 11676 24860 11688
rect 23992 11648 24860 11676
rect 23992 11636 23998 11648
rect 24854 11636 24860 11648
rect 24912 11636 24918 11688
rect 25222 11636 25228 11688
rect 25280 11636 25286 11688
rect 25498 11636 25504 11688
rect 25556 11636 25562 11688
rect 27356 11676 27384 11716
rect 27433 11713 27445 11747
rect 27479 11744 27491 11747
rect 28460 11744 28488 11772
rect 27479 11716 28488 11744
rect 27479 11713 27491 11716
rect 27433 11707 27491 11713
rect 28718 11704 28724 11756
rect 28776 11744 28782 11756
rect 30116 11744 30144 11775
rect 28776 11716 30144 11744
rect 28776 11704 28782 11716
rect 29457 11679 29515 11685
rect 27356 11648 28580 11676
rect 28552 11620 28580 11648
rect 29457 11645 29469 11679
rect 29503 11676 29515 11679
rect 29549 11679 29607 11685
rect 29549 11676 29561 11679
rect 29503 11648 29561 11676
rect 29503 11645 29515 11648
rect 29457 11639 29515 11645
rect 29549 11645 29561 11648
rect 29595 11645 29607 11679
rect 29549 11639 29607 11645
rect 20088 11580 21680 11608
rect 13280 11512 14964 11540
rect 11885 11503 11943 11509
rect 15194 11500 15200 11552
rect 15252 11540 15258 11552
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 15252 11512 15393 11540
rect 15252 11500 15258 11512
rect 15381 11509 15393 11512
rect 15427 11509 15439 11543
rect 15381 11503 15439 11509
rect 15930 11500 15936 11552
rect 15988 11500 15994 11552
rect 16114 11500 16120 11552
rect 16172 11500 16178 11552
rect 16859 11543 16917 11549
rect 16859 11509 16871 11543
rect 16905 11540 16917 11543
rect 17126 11540 17132 11552
rect 16905 11512 17132 11540
rect 16905 11509 16917 11512
rect 16859 11503 16917 11509
rect 17126 11500 17132 11512
rect 17184 11500 17190 11552
rect 18782 11500 18788 11552
rect 18840 11500 18846 11552
rect 19058 11500 19064 11552
rect 19116 11540 19122 11552
rect 19159 11543 19217 11549
rect 19159 11540 19171 11543
rect 19116 11512 19171 11540
rect 19116 11500 19122 11512
rect 19159 11509 19171 11512
rect 19205 11540 19217 11543
rect 20088 11540 20116 11580
rect 21652 11552 21680 11580
rect 28534 11568 28540 11620
rect 28592 11568 28598 11620
rect 28994 11568 29000 11620
rect 29052 11608 29058 11620
rect 29089 11611 29147 11617
rect 29089 11608 29101 11611
rect 29052 11580 29101 11608
rect 29052 11568 29058 11580
rect 29089 11577 29101 11580
rect 29135 11577 29147 11611
rect 29089 11571 29147 11577
rect 19205 11512 20116 11540
rect 19205 11509 19217 11512
rect 19159 11503 19217 11509
rect 21082 11500 21088 11552
rect 21140 11500 21146 11552
rect 21634 11500 21640 11552
rect 21692 11500 21698 11552
rect 22002 11540 22008 11552
rect 22060 11549 22066 11552
rect 21969 11512 22008 11540
rect 22002 11500 22008 11512
rect 22060 11540 22069 11549
rect 24955 11543 25013 11549
rect 24955 11540 24967 11543
rect 22060 11512 24967 11540
rect 22060 11503 22069 11512
rect 24955 11509 24967 11512
rect 25001 11540 25013 11543
rect 26970 11540 26976 11552
rect 25001 11512 26976 11540
rect 25001 11509 25013 11512
rect 24955 11503 25013 11509
rect 22060 11500 22066 11503
rect 26970 11500 26976 11512
rect 27028 11500 27034 11552
rect 27163 11543 27221 11549
rect 27163 11509 27175 11543
rect 27209 11540 27221 11543
rect 27522 11540 27528 11552
rect 27209 11512 27528 11540
rect 27209 11509 27221 11512
rect 27163 11503 27221 11509
rect 27522 11500 27528 11512
rect 27580 11500 27586 11552
rect 27706 11500 27712 11552
rect 27764 11540 27770 11552
rect 29564 11540 29592 11639
rect 29638 11636 29644 11688
rect 29696 11676 29702 11688
rect 30285 11679 30343 11685
rect 30285 11676 30297 11679
rect 29696 11648 30297 11676
rect 29696 11636 29702 11648
rect 30285 11645 30297 11648
rect 30331 11645 30343 11679
rect 30285 11639 30343 11645
rect 29825 11611 29883 11617
rect 29825 11608 29837 11611
rect 29656 11580 29837 11608
rect 29656 11552 29684 11580
rect 29825 11577 29837 11580
rect 29871 11577 29883 11611
rect 29825 11571 29883 11577
rect 30300 11552 30328 11639
rect 30374 11636 30380 11688
rect 30432 11676 30438 11688
rect 30561 11679 30619 11685
rect 30561 11676 30573 11679
rect 30432 11648 30573 11676
rect 30432 11636 30438 11648
rect 30561 11645 30573 11648
rect 30607 11645 30619 11679
rect 30561 11639 30619 11645
rect 31294 11636 31300 11688
rect 31352 11636 31358 11688
rect 27764 11512 29592 11540
rect 27764 11500 27770 11512
rect 29638 11500 29644 11552
rect 29696 11500 29702 11552
rect 30282 11500 30288 11552
rect 30340 11500 30346 11552
rect 30377 11543 30435 11549
rect 30377 11509 30389 11543
rect 30423 11540 30435 11543
rect 31312 11540 31340 11636
rect 30423 11512 31340 11540
rect 30423 11509 30435 11512
rect 30377 11503 30435 11509
rect 552 11450 31072 11472
rect 552 11398 7988 11450
rect 8040 11398 8052 11450
rect 8104 11398 8116 11450
rect 8168 11398 8180 11450
rect 8232 11398 8244 11450
rect 8296 11398 15578 11450
rect 15630 11398 15642 11450
rect 15694 11398 15706 11450
rect 15758 11398 15770 11450
rect 15822 11398 15834 11450
rect 15886 11398 23168 11450
rect 23220 11398 23232 11450
rect 23284 11398 23296 11450
rect 23348 11398 23360 11450
rect 23412 11398 23424 11450
rect 23476 11398 30758 11450
rect 30810 11398 30822 11450
rect 30874 11398 30886 11450
rect 30938 11398 30950 11450
rect 31002 11398 31014 11450
rect 31066 11398 31072 11450
rect 552 11376 31072 11398
rect 1394 11296 1400 11348
rect 1452 11296 1458 11348
rect 1762 11296 1768 11348
rect 1820 11336 1826 11348
rect 1955 11339 2013 11345
rect 1955 11336 1967 11339
rect 1820 11308 1967 11336
rect 1820 11296 1826 11308
rect 1955 11305 1967 11308
rect 2001 11305 2013 11339
rect 1955 11299 2013 11305
rect 2130 11296 2136 11348
rect 2188 11336 2194 11348
rect 3513 11339 3571 11345
rect 2188 11308 3464 11336
rect 2188 11296 2194 11308
rect 658 11228 664 11280
rect 716 11268 722 11280
rect 3436 11268 3464 11308
rect 3513 11305 3525 11339
rect 3559 11336 3571 11339
rect 3602 11336 3608 11348
rect 3559 11308 3608 11336
rect 3559 11305 3571 11308
rect 3513 11299 3571 11305
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 3878 11296 3884 11348
rect 3936 11336 3942 11348
rect 4801 11339 4859 11345
rect 4801 11336 4813 11339
rect 3936 11308 4813 11336
rect 3936 11296 3942 11308
rect 4801 11305 4813 11308
rect 4847 11305 4859 11339
rect 4801 11299 4859 11305
rect 4982 11296 4988 11348
rect 5040 11336 5046 11348
rect 5445 11339 5503 11345
rect 5445 11336 5457 11339
rect 5040 11308 5457 11336
rect 5040 11296 5046 11308
rect 5445 11305 5457 11308
rect 5491 11305 5503 11339
rect 5445 11299 5503 11305
rect 5813 11339 5871 11345
rect 5813 11305 5825 11339
rect 5859 11336 5871 11339
rect 5994 11336 6000 11348
rect 5859 11308 6000 11336
rect 5859 11305 5871 11308
rect 5813 11299 5871 11305
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 6270 11296 6276 11348
rect 6328 11296 6334 11348
rect 8849 11339 8907 11345
rect 6932 11308 8248 11336
rect 716 11240 1624 11268
rect 3436 11240 3832 11268
rect 716 11228 722 11240
rect 1302 11160 1308 11212
rect 1360 11200 1366 11212
rect 1489 11203 1547 11209
rect 1489 11200 1501 11203
rect 1360 11172 1501 11200
rect 1360 11160 1366 11172
rect 1489 11169 1501 11172
rect 1535 11169 1547 11203
rect 1596 11200 1624 11240
rect 2130 11200 2136 11212
rect 1596 11172 2136 11200
rect 1489 11163 1547 11169
rect 2130 11160 2136 11172
rect 2188 11160 2194 11212
rect 2225 11203 2283 11209
rect 2225 11169 2237 11203
rect 2271 11200 2283 11203
rect 3697 11203 3755 11209
rect 2271 11172 3188 11200
rect 2271 11169 2283 11172
rect 2225 11163 2283 11169
rect 1946 11092 1952 11144
rect 2004 11141 2010 11144
rect 2004 11135 2053 11141
rect 2004 11101 2007 11135
rect 2041 11101 2053 11135
rect 2004 11095 2053 11101
rect 2004 11092 2010 11095
rect 3160 11064 3188 11172
rect 3697 11169 3709 11203
rect 3743 11169 3755 11203
rect 3804 11200 3832 11240
rect 3970 11228 3976 11280
rect 4028 11228 4034 11280
rect 6288 11268 6316 11296
rect 6730 11268 6736 11280
rect 4080 11240 5304 11268
rect 4080 11200 4108 11240
rect 3804 11172 4108 11200
rect 4433 11203 4491 11209
rect 3697 11163 3755 11169
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 4614 11200 4620 11212
rect 4479 11172 4620 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 3602 11064 3608 11076
rect 3160 11036 3608 11064
rect 3602 11024 3608 11036
rect 3660 11024 3666 11076
rect 3712 11064 3740 11163
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 4706 11160 4712 11212
rect 4764 11160 4770 11212
rect 3786 11092 3792 11144
rect 3844 11132 3850 11144
rect 3844 11104 5212 11132
rect 3844 11092 3850 11104
rect 4062 11064 4068 11076
rect 3712 11036 4068 11064
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 5184 11073 5212 11104
rect 5169 11067 5227 11073
rect 4172 11036 4660 11064
rect 1670 10956 1676 11008
rect 1728 10996 1734 11008
rect 4172 10996 4200 11036
rect 1728 10968 4200 10996
rect 4249 10999 4307 11005
rect 1728 10956 1734 10968
rect 4249 10965 4261 10999
rect 4295 10996 4307 10999
rect 4522 10996 4528 11008
rect 4295 10968 4528 10996
rect 4295 10965 4307 10968
rect 4249 10959 4307 10965
rect 4522 10956 4528 10968
rect 4580 10956 4586 11008
rect 4632 10996 4660 11036
rect 5169 11033 5181 11067
rect 5215 11033 5227 11067
rect 5276 11064 5304 11240
rect 5460 11240 6316 11268
rect 6380 11240 6736 11268
rect 5460 11212 5488 11240
rect 5353 11203 5411 11209
rect 5353 11169 5365 11203
rect 5399 11169 5411 11203
rect 5353 11163 5411 11169
rect 5368 11132 5396 11163
rect 5442 11160 5448 11212
rect 5500 11160 5506 11212
rect 5629 11203 5687 11209
rect 5629 11169 5641 11203
rect 5675 11200 5687 11203
rect 5718 11200 5724 11212
rect 5675 11172 5724 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 5644 11132 5672 11163
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 5810 11160 5816 11212
rect 5868 11200 5874 11212
rect 6380 11209 6408 11240
rect 6730 11228 6736 11240
rect 6788 11268 6794 11280
rect 6932 11268 6960 11308
rect 6788 11240 6960 11268
rect 8220 11268 8248 11308
rect 8849 11305 8861 11339
rect 8895 11336 8907 11339
rect 9122 11336 9128 11348
rect 8895 11308 9128 11336
rect 8895 11305 8907 11308
rect 8849 11299 8907 11305
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 9398 11296 9404 11348
rect 9456 11336 9462 11348
rect 9677 11339 9735 11345
rect 9677 11336 9689 11339
rect 9456 11308 9689 11336
rect 9456 11296 9462 11308
rect 9677 11305 9689 11308
rect 9723 11305 9735 11339
rect 9677 11299 9735 11305
rect 10229 11339 10287 11345
rect 10229 11305 10241 11339
rect 10275 11336 10287 11339
rect 10410 11336 10416 11348
rect 10275 11308 10416 11336
rect 10275 11305 10287 11308
rect 10229 11299 10287 11305
rect 10410 11296 10416 11308
rect 10468 11296 10474 11348
rect 10686 11296 10692 11348
rect 10744 11336 10750 11348
rect 10744 11308 12572 11336
rect 10744 11296 10750 11308
rect 9416 11268 9444 11296
rect 10778 11268 10784 11280
rect 8220 11240 9444 11268
rect 9876 11240 10784 11268
rect 6788 11228 6794 11240
rect 5997 11203 6055 11209
rect 5997 11200 6009 11203
rect 5868 11172 6009 11200
rect 5868 11160 5874 11172
rect 5997 11169 6009 11172
rect 6043 11169 6055 11203
rect 5997 11163 6055 11169
rect 6365 11203 6423 11209
rect 6365 11169 6377 11203
rect 6411 11169 6423 11203
rect 6365 11163 6423 11169
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 7152 11203 7210 11209
rect 7152 11200 7164 11203
rect 6972 11172 7164 11200
rect 6972 11160 6978 11172
rect 7152 11169 7164 11172
rect 7198 11169 7210 11203
rect 7152 11163 7210 11169
rect 7558 11160 7564 11212
rect 7616 11160 7622 11212
rect 7650 11160 7656 11212
rect 7708 11200 7714 11212
rect 9033 11203 9091 11209
rect 7708 11172 8800 11200
rect 7708 11160 7714 11172
rect 5368 11104 5672 11132
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 6825 11135 6883 11141
rect 6825 11132 6837 11135
rect 6696 11104 6837 11132
rect 6696 11092 6702 11104
rect 6825 11101 6837 11104
rect 6871 11101 6883 11135
rect 7282 11132 7288 11144
rect 7248 11104 7288 11132
rect 6825 11095 6883 11101
rect 7282 11092 7288 11104
rect 7340 11092 7346 11144
rect 8772 11132 8800 11172
rect 9033 11169 9045 11203
rect 9079 11200 9091 11203
rect 9306 11200 9312 11212
rect 9079 11172 9312 11200
rect 9079 11169 9091 11172
rect 9033 11163 9091 11169
rect 9306 11160 9312 11172
rect 9364 11160 9370 11212
rect 9490 11160 9496 11212
rect 9548 11200 9554 11212
rect 9585 11203 9643 11209
rect 9585 11200 9597 11203
rect 9548 11172 9597 11200
rect 9548 11160 9554 11172
rect 9585 11169 9597 11172
rect 9631 11169 9643 11203
rect 9585 11163 9643 11169
rect 9876 11132 9904 11240
rect 10778 11228 10784 11240
rect 10836 11228 10842 11280
rect 10962 11228 10968 11280
rect 11020 11268 11026 11280
rect 12253 11271 12311 11277
rect 12253 11268 12265 11271
rect 11020 11240 12265 11268
rect 11020 11228 11026 11240
rect 12253 11237 12265 11240
rect 12299 11237 12311 11271
rect 12253 11231 12311 11237
rect 10042 11160 10048 11212
rect 10100 11160 10106 11212
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 10594 11200 10600 11212
rect 10459 11172 10600 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 10594 11160 10600 11172
rect 10652 11160 10658 11212
rect 10686 11160 10692 11212
rect 10744 11160 10750 11212
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11200 11207 11203
rect 11425 11203 11483 11209
rect 11425 11200 11437 11203
rect 11195 11172 11437 11200
rect 11195 11169 11207 11172
rect 11149 11163 11207 11169
rect 11425 11169 11437 11172
rect 11471 11200 11483 11203
rect 11701 11203 11759 11209
rect 11701 11200 11713 11203
rect 11471 11172 11713 11200
rect 11471 11169 11483 11172
rect 11425 11163 11483 11169
rect 11701 11169 11713 11172
rect 11747 11200 11759 11203
rect 11977 11203 12035 11209
rect 11747 11172 11836 11200
rect 11747 11169 11759 11172
rect 11701 11163 11759 11169
rect 8772 11104 9904 11132
rect 5350 11064 5356 11076
rect 5276 11036 5356 11064
rect 5169 11027 5227 11033
rect 5350 11024 5356 11036
rect 5408 11024 5414 11076
rect 6386 11036 6598 11064
rect 6386 10996 6414 11036
rect 4632 10968 6414 10996
rect 6454 10956 6460 11008
rect 6512 10956 6518 11008
rect 6570 10996 6598 11036
rect 9122 11024 9128 11076
rect 9180 11064 9186 11076
rect 9217 11067 9275 11073
rect 9217 11064 9229 11067
rect 9180 11036 9229 11064
rect 9180 11024 9186 11036
rect 9217 11033 9229 11036
rect 9263 11033 9275 11067
rect 9217 11027 9275 11033
rect 9306 11024 9312 11076
rect 9364 11064 9370 11076
rect 10060 11064 10088 11160
rect 10134 11092 10140 11144
rect 10192 11132 10198 11144
rect 11808 11132 11836 11172
rect 11977 11169 11989 11203
rect 12023 11200 12035 11203
rect 12158 11200 12164 11212
rect 12023 11172 12164 11200
rect 12023 11169 12035 11172
rect 11977 11163 12035 11169
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 12544 11200 12572 11308
rect 14642 11296 14648 11348
rect 14700 11336 14706 11348
rect 15749 11339 15807 11345
rect 15749 11336 15761 11339
rect 14700 11308 15761 11336
rect 14700 11296 14706 11308
rect 15749 11305 15761 11308
rect 15795 11305 15807 11339
rect 15749 11299 15807 11305
rect 16114 11296 16120 11348
rect 16172 11296 16178 11348
rect 16669 11339 16727 11345
rect 16669 11305 16681 11339
rect 16715 11336 16727 11339
rect 18598 11336 18604 11348
rect 16715 11308 18604 11336
rect 16715 11305 16727 11308
rect 16669 11299 16727 11305
rect 18598 11296 18604 11308
rect 18656 11296 18662 11348
rect 18782 11296 18788 11348
rect 18840 11296 18846 11348
rect 20530 11336 20536 11348
rect 18892 11308 20536 11336
rect 12820 11200 12943 11204
rect 12544 11176 12943 11200
rect 12544 11172 12848 11176
rect 10192 11104 11744 11132
rect 11808 11104 12296 11132
rect 10192 11092 10198 11104
rect 9364 11036 10088 11064
rect 9364 11024 9370 11036
rect 10502 11024 10508 11076
rect 10560 11024 10566 11076
rect 10962 11024 10968 11076
rect 11020 11024 11026 11076
rect 11241 11067 11299 11073
rect 11241 11033 11253 11067
rect 11287 11064 11299 11067
rect 11606 11064 11612 11076
rect 11287 11036 11612 11064
rect 11287 11033 11299 11036
rect 11241 11027 11299 11033
rect 11606 11024 11612 11036
rect 11664 11024 11670 11076
rect 11146 10996 11152 11008
rect 6570 10968 11152 10996
rect 11146 10956 11152 10968
rect 11204 10956 11210 11008
rect 11517 10999 11575 11005
rect 11517 10965 11529 10999
rect 11563 10996 11575 10999
rect 11716 10996 11744 11104
rect 12268 11076 12296 11104
rect 12434 11092 12440 11144
rect 12492 11092 12498 11144
rect 12802 11141 12808 11144
rect 12764 11135 12808 11141
rect 12764 11101 12776 11135
rect 12764 11095 12808 11101
rect 12802 11092 12808 11095
rect 12860 11092 12866 11144
rect 12915 11143 12943 11176
rect 13078 11160 13084 11212
rect 13136 11200 13142 11212
rect 13173 11203 13231 11209
rect 13173 11200 13185 11203
rect 13136 11172 13185 11200
rect 13136 11160 13142 11172
rect 13173 11169 13185 11172
rect 13219 11169 13231 11203
rect 13173 11163 13231 11169
rect 14826 11160 14832 11212
rect 14884 11160 14890 11212
rect 15105 11203 15163 11209
rect 15105 11169 15117 11203
rect 15151 11200 15163 11203
rect 15470 11200 15476 11212
rect 15151 11172 15476 11200
rect 15151 11169 15163 11172
rect 15105 11163 15163 11169
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 16132 11200 16160 11296
rect 17497 11203 17555 11209
rect 17497 11200 17509 11203
rect 16132 11172 17509 11200
rect 17497 11169 17509 11172
rect 17543 11169 17555 11203
rect 17497 11163 17555 11169
rect 12900 11137 12958 11143
rect 12900 11103 12912 11137
rect 12946 11103 12958 11137
rect 14844 11132 14872 11160
rect 16574 11132 16580 11144
rect 14844 11104 16580 11132
rect 12900 11097 12958 11103
rect 16574 11092 16580 11104
rect 16632 11092 16638 11144
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 16761 11135 16819 11141
rect 16761 11132 16773 11135
rect 16724 11104 16773 11132
rect 16724 11092 16730 11104
rect 16761 11101 16773 11104
rect 16807 11132 16819 11135
rect 16942 11132 16948 11144
rect 16807 11104 16948 11132
rect 16807 11101 16819 11104
rect 16761 11095 16819 11101
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 17126 11141 17132 11144
rect 17088 11135 17132 11141
rect 17088 11101 17100 11135
rect 17088 11095 17132 11101
rect 17126 11092 17132 11095
rect 17184 11092 17190 11144
rect 17267 11135 17325 11141
rect 17267 11101 17279 11135
rect 17313 11132 17325 11135
rect 18892 11132 18920 11308
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 20993 11339 21051 11345
rect 20993 11305 21005 11339
rect 21039 11336 21051 11339
rect 21818 11336 21824 11348
rect 21039 11308 21824 11336
rect 21039 11305 21051 11308
rect 20993 11299 21051 11305
rect 21818 11296 21824 11308
rect 21876 11296 21882 11348
rect 22195 11339 22253 11345
rect 22195 11305 22207 11339
rect 22241 11336 22253 11339
rect 22922 11336 22928 11348
rect 22241 11308 22928 11336
rect 22241 11305 22253 11308
rect 22195 11299 22253 11305
rect 22922 11296 22928 11308
rect 22980 11296 22986 11348
rect 24403 11339 24461 11345
rect 24403 11336 24415 11339
rect 23584 11308 24415 11336
rect 19058 11228 19064 11280
rect 19116 11228 19122 11280
rect 19076 11200 19104 11228
rect 19296 11203 19354 11209
rect 19296 11200 19308 11203
rect 19076 11172 19308 11200
rect 19296 11169 19308 11172
rect 19342 11169 19354 11203
rect 19296 11163 19354 11169
rect 19518 11160 19524 11212
rect 19576 11200 19582 11212
rect 19705 11203 19763 11209
rect 19705 11200 19717 11203
rect 19576 11172 19717 11200
rect 19576 11160 19582 11172
rect 19705 11169 19717 11172
rect 19751 11169 19763 11203
rect 19705 11163 19763 11169
rect 20622 11160 20628 11212
rect 20680 11200 20686 11212
rect 21453 11203 21511 11209
rect 21453 11200 21465 11203
rect 20680 11172 21465 11200
rect 20680 11160 20686 11172
rect 21453 11169 21465 11172
rect 21499 11169 21511 11203
rect 23584 11200 23612 11308
rect 24403 11305 24415 11308
rect 24449 11336 24461 11339
rect 24449 11308 25360 11336
rect 24449 11305 24461 11308
rect 24403 11299 24461 11305
rect 21453 11163 21511 11169
rect 22112 11172 23612 11200
rect 23845 11203 23903 11209
rect 22112 11144 22140 11172
rect 23845 11169 23857 11203
rect 23891 11200 23903 11203
rect 25332 11200 25360 11308
rect 25498 11296 25504 11348
rect 25556 11336 25562 11348
rect 25777 11339 25835 11345
rect 25777 11336 25789 11339
rect 25556 11308 25789 11336
rect 25556 11296 25562 11308
rect 25777 11305 25789 11308
rect 25823 11305 25835 11339
rect 25777 11299 25835 11305
rect 26142 11296 26148 11348
rect 26200 11336 26206 11348
rect 28994 11336 29000 11348
rect 26200 11308 29000 11336
rect 26200 11296 26206 11308
rect 28994 11296 29000 11308
rect 29052 11296 29058 11348
rect 29546 11296 29552 11348
rect 29604 11336 29610 11348
rect 30374 11336 30380 11348
rect 29604 11308 30380 11336
rect 29604 11296 29610 11308
rect 30374 11296 30380 11308
rect 30432 11296 30438 11348
rect 26748 11203 26806 11209
rect 26748 11200 26760 11203
rect 23891 11172 24256 11200
rect 25332 11172 26760 11200
rect 23891 11169 23903 11172
rect 23845 11163 23903 11169
rect 17313 11104 18920 11132
rect 18969 11135 19027 11141
rect 17313 11101 17325 11104
rect 17267 11095 17325 11101
rect 18969 11101 18981 11135
rect 19015 11101 19027 11135
rect 18969 11095 19027 11101
rect 11790 11024 11796 11076
rect 11848 11024 11854 11076
rect 12250 11024 12256 11076
rect 12308 11024 12314 11076
rect 11563 10968 11744 10996
rect 12452 10996 12480 11092
rect 14642 11024 14648 11076
rect 14700 11024 14706 11076
rect 14918 11024 14924 11076
rect 14976 11024 14982 11076
rect 15470 11024 15476 11076
rect 15528 11064 15534 11076
rect 16206 11064 16212 11076
rect 15528 11036 16212 11064
rect 15528 11024 15534 11036
rect 16206 11024 16212 11036
rect 16264 11024 16270 11076
rect 18690 11024 18696 11076
rect 18748 11064 18754 11076
rect 18984 11064 19012 11095
rect 19150 11092 19156 11144
rect 19208 11132 19214 11144
rect 19432 11135 19490 11141
rect 19432 11132 19444 11135
rect 19208 11104 19444 11132
rect 19208 11092 19214 11104
rect 19432 11101 19444 11104
rect 19478 11101 19490 11135
rect 19432 11095 19490 11101
rect 21542 11092 21548 11144
rect 21600 11132 21606 11144
rect 21729 11135 21787 11141
rect 21729 11132 21741 11135
rect 21600 11104 21741 11132
rect 21600 11092 21606 11104
rect 21729 11101 21741 11104
rect 21775 11132 21787 11135
rect 22002 11132 22008 11144
rect 21775 11104 22008 11132
rect 21775 11101 21787 11104
rect 21729 11095 21787 11101
rect 22002 11092 22008 11104
rect 22060 11092 22066 11144
rect 22094 11092 22100 11144
rect 22152 11092 22158 11144
rect 22235 11135 22293 11141
rect 22235 11101 22247 11135
rect 22281 11132 22293 11135
rect 22370 11132 22376 11144
rect 22281 11104 22376 11132
rect 22281 11101 22293 11104
rect 22235 11095 22293 11101
rect 22370 11092 22376 11104
rect 22428 11092 22434 11144
rect 22465 11135 22523 11141
rect 22465 11101 22477 11135
rect 22511 11132 22523 11135
rect 23566 11132 23572 11144
rect 22511 11104 23572 11132
rect 22511 11101 22523 11104
rect 22465 11095 22523 11101
rect 23566 11092 23572 11104
rect 23624 11092 23630 11144
rect 23937 11135 23995 11141
rect 23937 11132 23949 11135
rect 23768 11104 23949 11132
rect 18748 11036 19012 11064
rect 18748 11024 18754 11036
rect 13538 10996 13544 11008
rect 12452 10968 13544 10996
rect 11563 10965 11575 10968
rect 11517 10959 11575 10965
rect 13538 10956 13544 10968
rect 13596 10956 13602 11008
rect 14182 10956 14188 11008
rect 14240 10996 14246 11008
rect 14277 10999 14335 11005
rect 14277 10996 14289 10999
rect 14240 10968 14289 10996
rect 14240 10956 14246 10968
rect 14277 10965 14289 10968
rect 14323 10965 14335 10999
rect 14277 10959 14335 10965
rect 18966 10956 18972 11008
rect 19024 10996 19030 11008
rect 21174 10996 21180 11008
rect 19024 10968 21180 10996
rect 19024 10956 19030 10968
rect 21174 10956 21180 10968
rect 21232 10956 21238 11008
rect 21266 10956 21272 11008
rect 21324 10956 21330 11008
rect 21634 10956 21640 11008
rect 21692 10996 21698 11008
rect 22094 10996 22100 11008
rect 21692 10968 22100 10996
rect 21692 10956 21698 10968
rect 22094 10956 22100 10968
rect 22152 10956 22158 11008
rect 22646 10956 22652 11008
rect 22704 10996 22710 11008
rect 23768 10996 23796 11104
rect 23937 11101 23949 11104
rect 23983 11132 23995 11135
rect 24118 11132 24124 11144
rect 23983 11104 24124 11132
rect 23983 11101 23995 11104
rect 23937 11095 23995 11101
rect 24118 11092 24124 11104
rect 24176 11092 24182 11144
rect 24228 11132 24256 11172
rect 26620 11144 26648 11172
rect 26748 11169 26760 11172
rect 26794 11169 26806 11203
rect 26748 11163 26806 11169
rect 28166 11160 28172 11212
rect 28224 11200 28230 11212
rect 28629 11203 28687 11209
rect 28629 11200 28641 11203
rect 28224 11172 28641 11200
rect 28224 11160 28230 11172
rect 28629 11169 28641 11172
rect 28675 11169 28687 11203
rect 28629 11163 28687 11169
rect 28905 11203 28963 11209
rect 28905 11169 28917 11203
rect 28951 11200 28963 11203
rect 30190 11200 30196 11212
rect 28951 11172 30196 11200
rect 28951 11169 28963 11172
rect 28905 11163 28963 11169
rect 30190 11160 30196 11172
rect 30248 11160 30254 11212
rect 30392 11200 30420 11296
rect 30561 11203 30619 11209
rect 30561 11200 30573 11203
rect 30392 11172 30573 11200
rect 30561 11169 30573 11172
rect 30607 11169 30619 11203
rect 30561 11163 30619 11169
rect 24400 11135 24458 11141
rect 24400 11132 24412 11135
rect 24228 11104 24412 11132
rect 24400 11101 24412 11104
rect 24446 11101 24458 11135
rect 24400 11095 24458 11101
rect 24670 11092 24676 11144
rect 24728 11092 24734 11144
rect 26418 11092 26424 11144
rect 26476 11092 26482 11144
rect 26602 11092 26608 11144
rect 26660 11092 26666 11144
rect 26878 11092 26884 11144
rect 26936 11092 26942 11144
rect 27157 11135 27215 11141
rect 27157 11101 27169 11135
rect 27203 11132 27215 11135
rect 27522 11132 27528 11144
rect 27203 11104 27528 11132
rect 27203 11101 27215 11104
rect 27157 11095 27215 11101
rect 27522 11092 27528 11104
rect 27580 11092 27586 11144
rect 28442 11092 28448 11144
rect 28500 11132 28506 11144
rect 28500 11104 30420 11132
rect 28500 11092 28506 11104
rect 28074 11024 28080 11076
rect 28132 11064 28138 11076
rect 28261 11067 28319 11073
rect 28261 11064 28273 11067
rect 28132 11036 28273 11064
rect 28132 11024 28138 11036
rect 28261 11033 28273 11036
rect 28307 11033 28319 11067
rect 28261 11027 28319 11033
rect 30006 11024 30012 11076
rect 30064 11024 30070 11076
rect 30392 11073 30420 11104
rect 30377 11067 30435 11073
rect 30377 11033 30389 11067
rect 30423 11033 30435 11067
rect 30377 11027 30435 11033
rect 22704 10968 23796 10996
rect 22704 10956 22710 10968
rect 23842 10956 23848 11008
rect 23900 10996 23906 11008
rect 30098 10996 30104 11008
rect 23900 10968 30104 10996
rect 23900 10956 23906 10968
rect 30098 10956 30104 10968
rect 30156 10956 30162 11008
rect 552 10906 30912 10928
rect 552 10854 4193 10906
rect 4245 10854 4257 10906
rect 4309 10854 4321 10906
rect 4373 10854 4385 10906
rect 4437 10854 4449 10906
rect 4501 10854 11783 10906
rect 11835 10854 11847 10906
rect 11899 10854 11911 10906
rect 11963 10854 11975 10906
rect 12027 10854 12039 10906
rect 12091 10854 19373 10906
rect 19425 10854 19437 10906
rect 19489 10854 19501 10906
rect 19553 10854 19565 10906
rect 19617 10854 19629 10906
rect 19681 10854 26963 10906
rect 27015 10854 27027 10906
rect 27079 10854 27091 10906
rect 27143 10854 27155 10906
rect 27207 10854 27219 10906
rect 27271 10854 30912 10906
rect 552 10832 30912 10854
rect 5074 10792 5080 10804
rect 2976 10764 5080 10792
rect 937 10659 995 10665
rect 937 10625 949 10659
rect 983 10656 995 10659
rect 1302 10656 1308 10668
rect 983 10628 1308 10656
rect 983 10625 995 10628
rect 937 10619 995 10625
rect 1302 10616 1308 10628
rect 1360 10616 1366 10668
rect 1443 10657 1501 10663
rect 1443 10623 1455 10657
rect 1489 10656 1501 10657
rect 2976 10656 3004 10764
rect 5074 10752 5080 10764
rect 5132 10752 5138 10804
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10792 5319 10795
rect 6086 10792 6092 10804
rect 5307 10764 6092 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 6086 10752 6092 10764
rect 6144 10752 6150 10804
rect 7742 10752 7748 10804
rect 7800 10792 7806 10804
rect 8113 10795 8171 10801
rect 8113 10792 8125 10795
rect 7800 10764 8125 10792
rect 7800 10752 7806 10764
rect 8113 10761 8125 10764
rect 8159 10792 8171 10795
rect 8846 10792 8852 10804
rect 8159 10764 8852 10792
rect 8159 10761 8171 10764
rect 8113 10755 8171 10761
rect 8846 10752 8852 10764
rect 8904 10752 8910 10804
rect 9232 10764 11100 10792
rect 9232 10724 9260 10764
rect 8870 10696 9260 10724
rect 11072 10724 11100 10764
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 16025 10795 16083 10801
rect 11204 10764 15976 10792
rect 11204 10752 11210 10764
rect 13354 10724 13360 10736
rect 11072 10696 13360 10724
rect 1489 10628 3004 10656
rect 3053 10659 3111 10665
rect 1489 10623 1501 10628
rect 1443 10617 1501 10623
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3700 10659 3758 10665
rect 3700 10656 3712 10659
rect 3099 10628 3712 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3700 10625 3712 10628
rect 3746 10625 3758 10659
rect 4430 10656 4436 10668
rect 3700 10619 3758 10625
rect 3804 10628 4436 10656
rect 842 10548 848 10600
rect 900 10588 906 10600
rect 1673 10591 1731 10597
rect 1673 10588 1685 10591
rect 900 10560 1685 10588
rect 900 10548 906 10560
rect 1673 10557 1685 10560
rect 1719 10557 1731 10591
rect 1673 10551 1731 10557
rect 3234 10548 3240 10600
rect 3292 10548 3298 10600
rect 3804 10588 3832 10628
rect 4430 10616 4436 10628
rect 4488 10616 4494 10668
rect 6000 10659 6058 10665
rect 6000 10656 6012 10659
rect 5828 10628 6012 10656
rect 5828 10600 5856 10628
rect 6000 10625 6012 10628
rect 6046 10625 6058 10659
rect 6000 10619 6058 10625
rect 6196 10628 7972 10656
rect 3344 10560 3832 10588
rect 3973 10591 4031 10597
rect 1403 10455 1461 10461
rect 1403 10421 1415 10455
rect 1449 10452 1461 10455
rect 1762 10452 1768 10464
rect 1449 10424 1768 10452
rect 1449 10421 1461 10424
rect 1403 10415 1461 10421
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 2038 10412 2044 10464
rect 2096 10452 2102 10464
rect 3344 10452 3372 10560
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 4614 10588 4620 10600
rect 4019 10560 4620 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 5534 10548 5540 10600
rect 5592 10548 5598 10600
rect 5810 10548 5816 10600
rect 5868 10548 5874 10600
rect 5902 10548 5908 10600
rect 5960 10588 5966 10600
rect 6196 10588 6224 10628
rect 5960 10560 6224 10588
rect 5960 10548 5966 10560
rect 6270 10548 6276 10600
rect 6328 10548 6334 10600
rect 7944 10597 7972 10628
rect 7929 10591 7987 10597
rect 7929 10557 7941 10591
rect 7975 10557 7987 10591
rect 7929 10551 7987 10557
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8662 10588 8668 10600
rect 8435 10560 8668 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 8870 10597 8898 10696
rect 13354 10684 13360 10696
rect 13412 10684 13418 10736
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 9677 10659 9735 10665
rect 9677 10656 9689 10659
rect 9456 10628 9689 10656
rect 9456 10616 9462 10628
rect 9677 10625 9689 10628
rect 9723 10625 9735 10659
rect 9677 10619 9735 10625
rect 9858 10616 9864 10668
rect 9916 10616 9922 10668
rect 10042 10665 10048 10668
rect 10004 10659 10048 10665
rect 10004 10625 10016 10659
rect 10004 10619 10048 10625
rect 10042 10616 10048 10619
rect 10100 10616 10106 10668
rect 10140 10659 10198 10665
rect 10140 10625 10152 10659
rect 10186 10625 10198 10659
rect 10140 10619 10198 10625
rect 10413 10659 10471 10665
rect 10413 10625 10425 10659
rect 10459 10656 10471 10659
rect 11054 10656 11060 10668
rect 10459 10628 11060 10656
rect 10459 10625 10471 10628
rect 10413 10619 10471 10625
rect 8849 10591 8907 10597
rect 8849 10557 8861 10591
rect 8895 10557 8907 10591
rect 8849 10551 8907 10557
rect 9306 10548 9312 10600
rect 9364 10548 9370 10600
rect 9876 10588 9904 10616
rect 10155 10588 10183 10619
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 11793 10659 11851 10665
rect 11793 10625 11805 10659
rect 11839 10656 11851 10659
rect 13814 10656 13820 10668
rect 11839 10628 13820 10656
rect 11839 10625 11851 10628
rect 11793 10619 11851 10625
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 14047 10659 14105 10665
rect 14047 10625 14059 10659
rect 14093 10656 14105 10659
rect 14182 10656 14188 10668
rect 14093 10628 14188 10656
rect 14093 10625 14105 10628
rect 14047 10619 14105 10625
rect 14182 10616 14188 10628
rect 14240 10616 14246 10668
rect 15948 10656 15976 10764
rect 16025 10761 16037 10795
rect 16071 10792 16083 10795
rect 16758 10792 16764 10804
rect 16071 10764 16764 10792
rect 16071 10761 16083 10764
rect 16025 10755 16083 10761
rect 16758 10752 16764 10764
rect 16816 10752 16822 10804
rect 16942 10752 16948 10804
rect 17000 10792 17006 10804
rect 17000 10764 19104 10792
rect 17000 10752 17006 10764
rect 19076 10733 19104 10764
rect 19242 10752 19248 10804
rect 19300 10752 19306 10804
rect 21542 10792 21548 10804
rect 19536 10764 21548 10792
rect 19061 10727 19119 10733
rect 19061 10693 19073 10727
rect 19107 10724 19119 10727
rect 19536 10724 19564 10764
rect 21542 10752 21548 10764
rect 21600 10752 21606 10804
rect 21729 10795 21787 10801
rect 21729 10761 21741 10795
rect 21775 10792 21787 10795
rect 22278 10792 22284 10804
rect 21775 10764 22284 10792
rect 21775 10761 21787 10764
rect 21729 10755 21787 10761
rect 22278 10752 22284 10764
rect 22336 10752 22342 10804
rect 26605 10795 26663 10801
rect 26605 10761 26617 10795
rect 26651 10792 26663 10795
rect 26786 10792 26792 10804
rect 26651 10764 26792 10792
rect 26651 10761 26663 10764
rect 26605 10755 26663 10761
rect 26786 10752 26792 10764
rect 26844 10752 26850 10804
rect 28629 10795 28687 10801
rect 28629 10761 28641 10795
rect 28675 10792 28687 10795
rect 30558 10792 30564 10804
rect 28675 10764 30564 10792
rect 28675 10761 28687 10764
rect 28629 10755 28687 10761
rect 30558 10752 30564 10764
rect 30616 10752 30622 10804
rect 19107 10696 19564 10724
rect 19107 10693 19119 10696
rect 19061 10687 19119 10693
rect 16758 10656 16764 10668
rect 15948 10628 16764 10656
rect 16758 10616 16764 10628
rect 16816 10616 16822 10668
rect 17494 10656 17500 10668
rect 16874 10641 17500 10656
rect 16874 10610 16901 10641
rect 16889 10607 16901 10610
rect 16935 10628 17500 10641
rect 16935 10607 16947 10628
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 19536 10665 19564 10696
rect 21266 10684 21272 10736
rect 21324 10724 21330 10736
rect 21910 10724 21916 10736
rect 21324 10696 21916 10724
rect 21324 10684 21330 10696
rect 21910 10684 21916 10696
rect 21968 10684 21974 10736
rect 19521 10659 19579 10665
rect 19521 10625 19533 10659
rect 19567 10625 19579 10659
rect 19521 10619 19579 10625
rect 19886 10616 19892 10668
rect 19944 10616 19950 10668
rect 20027 10657 20085 10663
rect 20027 10623 20039 10657
rect 20073 10656 20085 10657
rect 20714 10656 20720 10668
rect 20073 10628 20720 10656
rect 20073 10623 20085 10628
rect 20027 10617 20085 10623
rect 20714 10616 20720 10628
rect 20772 10616 20778 10668
rect 21450 10616 21456 10668
rect 21508 10656 21514 10668
rect 21637 10659 21695 10665
rect 21637 10656 21649 10659
rect 21508 10628 21649 10656
rect 21508 10616 21514 10628
rect 21637 10625 21649 10628
rect 21683 10625 21695 10659
rect 21637 10619 21695 10625
rect 21726 10616 21732 10668
rect 21784 10656 21790 10668
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 21784 10628 22017 10656
rect 21784 10616 21790 10628
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 22922 10656 22928 10668
rect 22005 10619 22063 10625
rect 22210 10628 22928 10656
rect 16889 10601 16947 10607
rect 9585 10567 9643 10573
rect 7650 10480 7656 10532
rect 7708 10480 7714 10532
rect 7834 10480 7840 10532
rect 7892 10520 7898 10532
rect 9125 10523 9183 10529
rect 9125 10520 9137 10523
rect 7892 10492 9137 10520
rect 7892 10480 7898 10492
rect 9125 10489 9137 10492
rect 9171 10520 9183 10523
rect 9324 10520 9352 10548
rect 9585 10533 9597 10567
rect 9631 10533 9643 10567
rect 9876 10560 10183 10588
rect 10318 10548 10324 10600
rect 10376 10588 10382 10600
rect 12158 10588 12164 10600
rect 10376 10560 12164 10588
rect 10376 10548 10382 10560
rect 12158 10548 12164 10560
rect 12216 10548 12222 10600
rect 12342 10548 12348 10600
rect 12400 10588 12406 10600
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 12400 10560 12449 10588
rect 12400 10548 12406 10560
rect 12437 10557 12449 10560
rect 12483 10557 12495 10591
rect 12437 10551 12495 10557
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 12894 10588 12900 10600
rect 12676 10560 12900 10588
rect 12676 10548 12682 10560
rect 12894 10548 12900 10560
rect 12952 10548 12958 10600
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10588 13415 10591
rect 13446 10588 13452 10600
rect 13403 10560 13452 10588
rect 13403 10557 13415 10560
rect 13357 10551 13415 10557
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 13538 10548 13544 10600
rect 13596 10548 13602 10600
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 13648 10560 14289 10588
rect 9585 10527 9643 10533
rect 9171 10492 9352 10520
rect 9171 10489 9183 10492
rect 9125 10483 9183 10489
rect 2096 10424 3372 10452
rect 3703 10455 3761 10461
rect 2096 10412 2102 10424
rect 3703 10421 3715 10455
rect 3749 10452 3761 10455
rect 3970 10452 3976 10464
rect 3749 10424 3976 10452
rect 3749 10421 3761 10424
rect 3703 10415 3761 10421
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 4430 10412 4436 10464
rect 4488 10452 4494 10464
rect 4706 10452 4712 10464
rect 4488 10424 4712 10452
rect 4488 10412 4494 10424
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 6003 10455 6061 10461
rect 6003 10421 6015 10455
rect 6049 10452 6061 10455
rect 6178 10452 6184 10464
rect 6049 10424 6184 10452
rect 6049 10421 6061 10424
rect 6003 10415 6061 10421
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 8573 10455 8631 10461
rect 8573 10421 8585 10455
rect 8619 10452 8631 10455
rect 8754 10452 8760 10464
rect 8619 10424 8760 10452
rect 8619 10421 8631 10424
rect 8573 10415 8631 10421
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 9398 10412 9404 10464
rect 9456 10412 9462 10464
rect 9600 10452 9628 10527
rect 11977 10523 12035 10529
rect 11977 10489 11989 10523
rect 12023 10520 12035 10523
rect 13556 10520 13584 10548
rect 12023 10492 13584 10520
rect 12023 10489 12035 10492
rect 11977 10483 12035 10489
rect 10410 10452 10416 10464
rect 9600 10424 10416 10452
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 12066 10412 12072 10464
rect 12124 10452 12130 10464
rect 12434 10452 12440 10464
rect 12124 10424 12440 10452
rect 12124 10412 12130 10424
rect 12434 10412 12440 10424
rect 12492 10412 12498 10464
rect 12618 10412 12624 10464
rect 12676 10412 12682 10464
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 13078 10452 13084 10464
rect 12943 10424 13084 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 13078 10412 13084 10424
rect 13136 10412 13142 10464
rect 13173 10455 13231 10461
rect 13173 10421 13185 10455
rect 13219 10452 13231 10455
rect 13648 10452 13676 10560
rect 14277 10557 14289 10560
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 16393 10591 16451 10597
rect 16393 10557 16405 10591
rect 16439 10588 16451 10591
rect 16482 10588 16488 10600
rect 16439 10560 16488 10588
rect 16439 10557 16451 10560
rect 16393 10551 16451 10557
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 17129 10591 17187 10597
rect 17129 10557 17141 10591
rect 17175 10588 17187 10591
rect 19150 10588 19156 10600
rect 17175 10560 19156 10588
rect 17175 10557 17187 10560
rect 17129 10551 17187 10557
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 19429 10591 19487 10597
rect 19429 10588 19441 10591
rect 19306 10560 19441 10588
rect 18509 10523 18567 10529
rect 18509 10489 18521 10523
rect 18555 10520 18567 10523
rect 18690 10520 18696 10532
rect 18555 10492 18696 10520
rect 18555 10489 18567 10492
rect 18509 10483 18567 10489
rect 18690 10480 18696 10492
rect 18748 10480 18754 10532
rect 18782 10480 18788 10532
rect 18840 10480 18846 10532
rect 13219 10424 13676 10452
rect 13219 10421 13231 10424
rect 13173 10415 13231 10421
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 14007 10455 14065 10461
rect 14007 10452 14019 10455
rect 13964 10424 14019 10452
rect 13964 10412 13970 10424
rect 14007 10421 14019 10424
rect 14053 10421 14065 10455
rect 14007 10415 14065 10421
rect 15286 10412 15292 10464
rect 15344 10452 15350 10464
rect 15381 10455 15439 10461
rect 15381 10452 15393 10455
rect 15344 10424 15393 10452
rect 15344 10412 15350 10424
rect 15381 10421 15393 10424
rect 15427 10421 15439 10455
rect 15381 10415 15439 10421
rect 16666 10412 16672 10464
rect 16724 10452 16730 10464
rect 16850 10452 16856 10464
rect 16908 10461 16914 10464
rect 16724 10424 16856 10452
rect 16724 10412 16730 10424
rect 16850 10412 16856 10424
rect 16908 10415 16917 10461
rect 16908 10412 16914 10415
rect 17034 10412 17040 10464
rect 17092 10452 17098 10464
rect 19306 10452 19334 10560
rect 19429 10557 19441 10560
rect 19475 10588 19487 10591
rect 19904 10588 19932 10616
rect 19475 10560 19932 10588
rect 19475 10557 19487 10560
rect 19429 10551 19487 10557
rect 20254 10548 20260 10600
rect 20312 10548 20318 10600
rect 21818 10548 21824 10600
rect 21876 10588 21882 10600
rect 21913 10591 21971 10597
rect 21913 10588 21925 10591
rect 21876 10560 21925 10588
rect 21876 10548 21882 10560
rect 21913 10557 21925 10560
rect 21959 10557 21971 10591
rect 22210 10588 22238 10628
rect 22922 10616 22928 10628
rect 22980 10616 22986 10668
rect 23474 10616 23480 10668
rect 23532 10616 23538 10668
rect 24946 10665 24952 10668
rect 24908 10659 24952 10665
rect 23584 10628 24716 10656
rect 21913 10551 21971 10557
rect 22020 10560 22238 10588
rect 22281 10591 22339 10597
rect 20990 10480 20996 10532
rect 21048 10520 21054 10532
rect 21542 10520 21548 10532
rect 21048 10492 21548 10520
rect 21048 10480 21054 10492
rect 21542 10480 21548 10492
rect 21600 10480 21606 10532
rect 17092 10424 19334 10452
rect 17092 10412 17098 10424
rect 19610 10412 19616 10464
rect 19668 10452 19674 10464
rect 19987 10455 20045 10461
rect 19987 10452 19999 10455
rect 19668 10424 19999 10452
rect 19668 10412 19674 10424
rect 19987 10421 19999 10424
rect 20033 10452 20045 10455
rect 22020 10452 22048 10560
rect 22281 10557 22293 10591
rect 22327 10588 22339 10591
rect 22327 10560 22968 10588
rect 22327 10557 22339 10560
rect 22281 10551 22339 10557
rect 22940 10520 22968 10560
rect 23014 10548 23020 10600
rect 23072 10588 23078 10600
rect 23584 10588 23612 10628
rect 23072 10560 23612 10588
rect 23937 10591 23995 10597
rect 23072 10548 23078 10560
rect 23937 10557 23949 10591
rect 23983 10588 23995 10591
rect 24302 10588 24308 10600
rect 23983 10560 24308 10588
rect 23983 10557 23995 10560
rect 23937 10551 23995 10557
rect 23842 10520 23848 10532
rect 22940 10492 23848 10520
rect 23842 10480 23848 10492
rect 23900 10480 23906 10532
rect 20033 10424 22048 10452
rect 20033 10421 20045 10424
rect 19987 10415 20045 10421
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 23952 10452 23980 10551
rect 24302 10548 24308 10560
rect 24360 10588 24366 10600
rect 24581 10591 24639 10597
rect 24581 10588 24593 10591
rect 24360 10560 24593 10588
rect 24360 10548 24366 10560
rect 24581 10557 24593 10560
rect 24627 10557 24639 10591
rect 24688 10588 24716 10628
rect 24908 10625 24920 10659
rect 24908 10619 24952 10625
rect 24946 10616 24952 10619
rect 25004 10616 25010 10668
rect 25087 10659 25145 10665
rect 25087 10625 25099 10659
rect 25133 10656 25145 10659
rect 26789 10659 26847 10665
rect 25133 10628 25728 10656
rect 25133 10625 25145 10628
rect 25087 10619 25145 10625
rect 25700 10600 25728 10628
rect 26789 10625 26801 10659
rect 26835 10656 26847 10659
rect 27798 10656 27804 10668
rect 26835 10628 27804 10656
rect 26835 10625 26847 10628
rect 26789 10619 26847 10625
rect 27798 10616 27804 10628
rect 27856 10616 27862 10668
rect 29178 10616 29184 10668
rect 29236 10656 29242 10668
rect 29730 10656 29736 10668
rect 29236 10628 29736 10656
rect 29236 10616 29242 10628
rect 29730 10616 29736 10628
rect 29788 10656 29794 10668
rect 29788 10628 30144 10656
rect 29788 10616 29794 10628
rect 25317 10591 25375 10597
rect 25317 10588 25329 10591
rect 24688 10560 25329 10588
rect 24581 10551 24639 10557
rect 25317 10557 25329 10560
rect 25363 10557 25375 10591
rect 25317 10551 25375 10557
rect 25682 10548 25688 10600
rect 25740 10548 25746 10600
rect 25774 10548 25780 10600
rect 25832 10588 25838 10600
rect 27065 10591 27123 10597
rect 27065 10588 27077 10591
rect 25832 10560 27077 10588
rect 25832 10548 25838 10560
rect 27065 10557 27077 10560
rect 27111 10557 27123 10591
rect 27065 10551 27123 10557
rect 28813 10591 28871 10597
rect 28813 10557 28825 10591
rect 28859 10588 28871 10591
rect 29454 10588 29460 10600
rect 28859 10560 29460 10588
rect 28859 10557 28871 10560
rect 28813 10551 28871 10557
rect 29454 10548 29460 10560
rect 29512 10548 29518 10600
rect 29546 10548 29552 10600
rect 29604 10548 29610 10600
rect 30116 10597 30144 10628
rect 30101 10591 30159 10597
rect 30101 10557 30113 10591
rect 30147 10557 30159 10591
rect 30101 10551 30159 10557
rect 24118 10480 24124 10532
rect 24176 10480 24182 10532
rect 29089 10523 29147 10529
rect 29089 10489 29101 10523
rect 29135 10520 29147 10523
rect 29564 10520 29592 10548
rect 29135 10492 29592 10520
rect 29641 10523 29699 10529
rect 29135 10489 29147 10492
rect 29089 10483 29147 10489
rect 29641 10489 29653 10523
rect 29687 10520 29699 10523
rect 29687 10492 30144 10520
rect 29687 10489 29699 10492
rect 29641 10483 29699 10489
rect 22152 10424 23980 10452
rect 22152 10412 22158 10424
rect 24026 10412 24032 10464
rect 24084 10412 24090 10464
rect 24136 10452 24164 10480
rect 30116 10464 30144 10492
rect 25130 10452 25136 10464
rect 24136 10424 25136 10452
rect 25130 10412 25136 10424
rect 25188 10412 25194 10464
rect 25406 10412 25412 10464
rect 25464 10452 25470 10464
rect 28169 10455 28227 10461
rect 28169 10452 28181 10455
rect 25464 10424 28181 10452
rect 25464 10412 25470 10424
rect 28169 10421 28181 10424
rect 28215 10421 28227 10455
rect 28169 10415 28227 10421
rect 28994 10412 29000 10464
rect 29052 10452 29058 10464
rect 29181 10455 29239 10461
rect 29181 10452 29193 10455
rect 29052 10424 29193 10452
rect 29052 10412 29058 10424
rect 29181 10421 29193 10424
rect 29227 10421 29239 10455
rect 29181 10415 29239 10421
rect 29362 10412 29368 10464
rect 29420 10452 29426 10464
rect 29733 10455 29791 10461
rect 29733 10452 29745 10455
rect 29420 10424 29745 10452
rect 29420 10412 29426 10424
rect 29733 10421 29745 10424
rect 29779 10421 29791 10455
rect 29733 10415 29791 10421
rect 30098 10412 30104 10464
rect 30156 10412 30162 10464
rect 30282 10412 30288 10464
rect 30340 10412 30346 10464
rect 552 10362 31072 10384
rect 552 10310 7988 10362
rect 8040 10310 8052 10362
rect 8104 10310 8116 10362
rect 8168 10310 8180 10362
rect 8232 10310 8244 10362
rect 8296 10310 15578 10362
rect 15630 10310 15642 10362
rect 15694 10310 15706 10362
rect 15758 10310 15770 10362
rect 15822 10310 15834 10362
rect 15886 10310 23168 10362
rect 23220 10310 23232 10362
rect 23284 10310 23296 10362
rect 23348 10310 23360 10362
rect 23412 10310 23424 10362
rect 23476 10310 30758 10362
rect 30810 10310 30822 10362
rect 30874 10310 30886 10362
rect 30938 10310 30950 10362
rect 31002 10310 31014 10362
rect 31066 10310 31072 10362
rect 552 10288 31072 10310
rect 1587 10251 1645 10257
rect 1587 10217 1599 10251
rect 1633 10248 1645 10251
rect 1762 10248 1768 10260
rect 1633 10220 1768 10248
rect 1633 10217 1645 10220
rect 1587 10211 1645 10217
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 3795 10251 3853 10257
rect 3795 10217 3807 10251
rect 3841 10248 3853 10251
rect 3970 10248 3976 10260
rect 3841 10220 3976 10248
rect 3841 10217 3853 10220
rect 3795 10211 3853 10217
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 6454 10248 6460 10260
rect 5592 10220 6460 10248
rect 5592 10208 5598 10220
rect 6454 10208 6460 10220
rect 6512 10208 6518 10260
rect 6822 10248 6828 10260
rect 6564 10220 6828 10248
rect 5445 10183 5503 10189
rect 5445 10149 5457 10183
rect 5491 10180 5503 10183
rect 5810 10180 5816 10192
rect 5491 10152 5816 10180
rect 5491 10149 5503 10152
rect 5445 10143 5503 10149
rect 5810 10140 5816 10152
rect 5868 10140 5874 10192
rect 6178 10140 6184 10192
rect 6236 10180 6242 10192
rect 6564 10180 6592 10220
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 6923 10251 6981 10257
rect 6923 10217 6935 10251
rect 6969 10248 6981 10251
rect 7834 10248 7840 10260
rect 6969 10220 7840 10248
rect 6969 10217 6981 10220
rect 6923 10211 6981 10217
rect 7834 10208 7840 10220
rect 7892 10208 7898 10260
rect 9490 10248 9496 10260
rect 8496 10220 9496 10248
rect 6236 10152 6592 10180
rect 6236 10140 6242 10152
rect 1029 10115 1087 10121
rect 1029 10081 1041 10115
rect 1075 10112 1087 10115
rect 3237 10115 3295 10121
rect 1075 10084 1440 10112
rect 1075 10081 1087 10084
rect 1029 10075 1087 10081
rect 1412 10056 1440 10084
rect 1786 10084 2774 10112
rect 1121 10047 1179 10053
rect 1121 10013 1133 10047
rect 1167 10044 1179 10047
rect 1302 10044 1308 10056
rect 1167 10016 1308 10044
rect 1167 10013 1179 10016
rect 1121 10007 1179 10013
rect 1302 10004 1308 10016
rect 1360 10004 1366 10056
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 1627 10047 1685 10053
rect 1627 10013 1639 10047
rect 1673 10044 1685 10047
rect 1786 10044 1814 10084
rect 1673 10016 1814 10044
rect 1857 10047 1915 10053
rect 1673 10013 1685 10016
rect 1627 10007 1685 10013
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 1903 10016 2544 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 845 9911 903 9917
rect 845 9877 857 9911
rect 891 9908 903 9911
rect 2516 9908 2544 10016
rect 891 9880 2544 9908
rect 2746 9908 2774 10084
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 4065 10115 4123 10121
rect 3283 10084 3832 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 3326 10004 3332 10056
rect 3384 10004 3390 10056
rect 3804 10053 3832 10084
rect 4065 10081 4077 10115
rect 4111 10112 4123 10115
rect 4522 10112 4528 10124
rect 4111 10084 4528 10112
rect 4111 10081 4123 10084
rect 4065 10075 4123 10081
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 5626 10072 5632 10124
rect 5684 10112 5690 10124
rect 5905 10115 5963 10121
rect 5905 10112 5917 10115
rect 5684 10084 5917 10112
rect 5684 10072 5690 10084
rect 5905 10081 5917 10084
rect 5951 10081 5963 10115
rect 5905 10075 5963 10081
rect 6457 10115 6515 10121
rect 6457 10081 6469 10115
rect 6503 10112 6515 10115
rect 6730 10112 6736 10124
rect 6503 10084 6736 10112
rect 6503 10081 6515 10084
rect 6457 10075 6515 10081
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 6840 10084 7328 10112
rect 3792 10047 3850 10053
rect 3792 10013 3804 10047
rect 3838 10013 3850 10047
rect 6840 10044 6868 10084
rect 7300 10056 7328 10084
rect 8496 10056 8524 10220
rect 9490 10208 9496 10220
rect 9548 10248 9554 10260
rect 12066 10248 12072 10260
rect 9548 10220 12072 10248
rect 9548 10208 9554 10220
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 13354 10208 13360 10260
rect 13412 10208 13418 10260
rect 13446 10208 13452 10260
rect 13504 10248 13510 10260
rect 15470 10248 15476 10260
rect 13504 10220 15476 10248
rect 13504 10208 13510 10220
rect 15470 10208 15476 10220
rect 15528 10248 15534 10260
rect 16206 10248 16212 10260
rect 15528 10220 16212 10248
rect 15528 10208 15534 10220
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 16853 10251 16911 10257
rect 16853 10217 16865 10251
rect 16899 10217 16911 10251
rect 16853 10211 16911 10217
rect 16868 10180 16896 10211
rect 17126 10208 17132 10260
rect 17184 10248 17190 10260
rect 17595 10251 17653 10257
rect 17595 10248 17607 10251
rect 17184 10220 17607 10248
rect 17184 10208 17190 10220
rect 17595 10217 17607 10220
rect 17641 10248 17653 10251
rect 17641 10220 18834 10248
rect 17641 10217 17653 10220
rect 17595 10211 17653 10217
rect 16040 10152 16436 10180
rect 16868 10152 17264 10180
rect 8573 10115 8631 10121
rect 8573 10081 8585 10115
rect 8619 10112 8631 10115
rect 8619 10084 9168 10112
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 3792 10007 3850 10013
rect 6196 10016 6868 10044
rect 6963 10047 7021 10053
rect 5718 9936 5724 9988
rect 5776 9976 5782 9988
rect 6196 9976 6224 10016
rect 6963 10013 6975 10047
rect 7009 10044 7021 10047
rect 7098 10044 7104 10056
rect 7009 10016 7104 10044
rect 7009 10013 7021 10016
rect 6963 10007 7021 10013
rect 7098 10004 7104 10016
rect 7156 10004 7162 10056
rect 7190 10004 7196 10056
rect 7248 10004 7254 10056
rect 7282 10004 7288 10056
rect 7340 10004 7346 10056
rect 8478 10004 8484 10056
rect 8536 10044 8542 10056
rect 9030 10053 9036 10056
rect 8665 10047 8723 10053
rect 8665 10044 8677 10047
rect 8536 10016 8677 10044
rect 8536 10004 8542 10016
rect 8665 10013 8677 10016
rect 8711 10013 8723 10047
rect 8665 10007 8723 10013
rect 8992 10047 9036 10053
rect 8992 10013 9004 10047
rect 8992 10007 9036 10013
rect 9030 10004 9036 10007
rect 9088 10004 9094 10056
rect 9140 10053 9168 10084
rect 9398 10072 9404 10124
rect 9456 10072 9462 10124
rect 9674 10072 9680 10124
rect 9732 10112 9738 10124
rect 10226 10112 10232 10124
rect 9732 10084 10232 10112
rect 9732 10072 9738 10084
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 10594 10072 10600 10124
rect 10652 10112 10658 10124
rect 11701 10115 11759 10121
rect 11701 10112 11713 10115
rect 10652 10084 11713 10112
rect 10652 10072 10658 10084
rect 11701 10081 11713 10084
rect 11747 10081 11759 10115
rect 11701 10075 11759 10081
rect 12894 10072 12900 10124
rect 12952 10112 12958 10124
rect 13265 10115 13323 10121
rect 13265 10112 13277 10115
rect 12952 10084 13277 10112
rect 12952 10072 12958 10084
rect 13265 10081 13277 10084
rect 13311 10081 13323 10115
rect 13265 10075 13323 10081
rect 13538 10072 13544 10124
rect 13596 10072 13602 10124
rect 15470 10072 15476 10124
rect 15528 10112 15534 10124
rect 15528 10084 15884 10112
rect 15528 10072 15534 10084
rect 9128 10047 9186 10053
rect 9128 10013 9140 10047
rect 9174 10013 9186 10047
rect 9128 10007 9186 10013
rect 10778 10004 10784 10056
rect 10836 10044 10842 10056
rect 11330 10053 11336 10056
rect 10965 10047 11023 10053
rect 10965 10044 10977 10047
rect 10836 10016 10977 10044
rect 10836 10004 10842 10016
rect 10965 10013 10977 10016
rect 11011 10013 11023 10047
rect 10965 10007 11023 10013
rect 11292 10047 11336 10053
rect 11292 10013 11304 10047
rect 11292 10007 11336 10013
rect 11330 10004 11336 10007
rect 11388 10004 11394 10056
rect 11422 10004 11428 10056
rect 11480 10004 11486 10056
rect 13906 10053 13912 10056
rect 13868 10047 13912 10053
rect 13868 10013 13880 10047
rect 13868 10007 13912 10013
rect 13906 10004 13912 10007
rect 13964 10004 13970 10056
rect 13998 10004 14004 10056
rect 14056 10055 14062 10056
rect 14056 10049 14078 10055
rect 14066 10015 14078 10049
rect 14056 10009 14078 10015
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10044 14335 10047
rect 15856 10044 15884 10084
rect 15930 10072 15936 10124
rect 15988 10121 15994 10124
rect 15988 10112 15999 10121
rect 16040 10112 16068 10152
rect 15988 10084 16068 10112
rect 16301 10115 16359 10121
rect 15988 10075 15999 10084
rect 16301 10081 16313 10115
rect 16347 10081 16359 10115
rect 16301 10075 16359 10081
rect 15988 10072 15994 10075
rect 16316 10044 16344 10075
rect 16408 10056 16436 10152
rect 16761 10115 16819 10121
rect 16761 10081 16773 10115
rect 16807 10081 16819 10115
rect 16761 10075 16819 10081
rect 14323 10016 15792 10044
rect 15856 10016 16344 10044
rect 14323 10013 14335 10016
rect 14056 10004 14062 10009
rect 14277 10007 14335 10013
rect 5776 9948 6224 9976
rect 5776 9936 5782 9948
rect 8570 9936 8576 9988
rect 8628 9936 8634 9988
rect 15764 9985 15792 10016
rect 16390 10004 16396 10056
rect 16448 10004 16454 10056
rect 15749 9979 15807 9985
rect 15749 9945 15761 9979
rect 15795 9945 15807 9979
rect 16776 9976 16804 10075
rect 16942 10072 16948 10124
rect 17000 10072 17006 10124
rect 17034 10072 17040 10124
rect 17092 10072 17098 10124
rect 17236 10112 17264 10152
rect 18690 10140 18696 10192
rect 18748 10140 18754 10192
rect 18806 10180 18834 10220
rect 19058 10208 19064 10260
rect 19116 10248 19122 10260
rect 19153 10251 19211 10257
rect 19153 10248 19165 10251
rect 19116 10220 19165 10248
rect 19116 10208 19122 10220
rect 19153 10217 19165 10220
rect 19199 10217 19211 10251
rect 19153 10211 19211 10217
rect 19981 10251 20039 10257
rect 19981 10217 19993 10251
rect 20027 10248 20039 10251
rect 20254 10248 20260 10260
rect 20027 10220 20260 10248
rect 20027 10217 20039 10220
rect 19981 10211 20039 10217
rect 20254 10208 20260 10220
rect 20312 10208 20318 10260
rect 20990 10208 20996 10260
rect 21048 10208 21054 10260
rect 22646 10248 22652 10260
rect 21284 10220 22652 10248
rect 19610 10180 19616 10192
rect 18806 10152 19616 10180
rect 19610 10140 19616 10152
rect 19668 10140 19674 10192
rect 20622 10180 20628 10192
rect 20180 10152 20628 10180
rect 17865 10115 17923 10121
rect 17865 10112 17877 10115
rect 17236 10084 17877 10112
rect 17865 10081 17877 10084
rect 17911 10081 17923 10115
rect 17865 10075 17923 10081
rect 16960 10044 16988 10072
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 16960 10016 17141 10044
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 17635 10047 17693 10053
rect 17635 10013 17647 10047
rect 17681 10044 17693 10047
rect 17770 10044 17776 10056
rect 17681 10016 17776 10044
rect 17681 10013 17693 10016
rect 17635 10007 17693 10013
rect 17770 10004 17776 10016
rect 17828 10004 17834 10056
rect 18708 9976 18736 10140
rect 19337 10115 19395 10121
rect 19337 10081 19349 10115
rect 19383 10112 19395 10115
rect 19518 10112 19524 10124
rect 19383 10084 19524 10112
rect 19383 10081 19395 10084
rect 19337 10075 19395 10081
rect 19518 10072 19524 10084
rect 19576 10072 19582 10124
rect 19702 10072 19708 10124
rect 19760 10112 19766 10124
rect 20180 10121 20208 10152
rect 20622 10140 20628 10152
rect 20680 10140 20686 10192
rect 20165 10115 20223 10121
rect 20165 10112 20177 10115
rect 19760 10084 20177 10112
rect 19760 10072 19766 10084
rect 20165 10081 20177 10084
rect 20211 10081 20223 10115
rect 20165 10075 20223 10081
rect 20254 10072 20260 10124
rect 20312 10112 20318 10124
rect 20441 10115 20499 10121
rect 20441 10112 20453 10115
rect 20312 10084 20453 10112
rect 20312 10072 20318 10084
rect 20441 10081 20453 10084
rect 20487 10081 20499 10115
rect 20441 10075 20499 10081
rect 18782 10004 18788 10056
rect 18840 10044 18846 10056
rect 21284 10053 21312 10220
rect 22646 10208 22652 10220
rect 22704 10208 22710 10260
rect 22830 10208 22836 10260
rect 22888 10248 22894 10260
rect 23109 10251 23167 10257
rect 23109 10248 23121 10251
rect 22888 10220 23121 10248
rect 22888 10208 22894 10220
rect 23109 10217 23121 10220
rect 23155 10217 23167 10251
rect 23109 10211 23167 10217
rect 23477 10251 23535 10257
rect 23477 10217 23489 10251
rect 23523 10248 23535 10251
rect 23566 10248 23572 10260
rect 23523 10220 23572 10248
rect 23523 10217 23535 10220
rect 23477 10211 23535 10217
rect 23566 10208 23572 10220
rect 23624 10208 23630 10260
rect 23845 10251 23903 10257
rect 23845 10217 23857 10251
rect 23891 10248 23903 10251
rect 24670 10248 24676 10260
rect 23891 10220 24676 10248
rect 23891 10217 23903 10220
rect 23845 10211 23903 10217
rect 24670 10208 24676 10220
rect 24728 10208 24734 10260
rect 24946 10208 24952 10260
rect 25004 10248 25010 10260
rect 25004 10220 25544 10248
rect 25004 10208 25010 10220
rect 22922 10140 22928 10192
rect 22980 10180 22986 10192
rect 25516 10180 25544 10220
rect 26326 10208 26332 10260
rect 26384 10248 26390 10260
rect 30009 10251 30067 10257
rect 30009 10248 30021 10251
rect 26384 10220 30021 10248
rect 26384 10208 26390 10220
rect 30009 10217 30021 10220
rect 30055 10217 30067 10251
rect 30009 10211 30067 10217
rect 26510 10180 26516 10192
rect 22980 10152 24164 10180
rect 25516 10152 26516 10180
rect 22980 10140 22986 10152
rect 21634 10121 21640 10124
rect 21596 10115 21640 10121
rect 21596 10081 21608 10115
rect 21596 10075 21640 10081
rect 21634 10072 21640 10075
rect 21692 10072 21698 10124
rect 22002 10072 22008 10124
rect 22060 10072 22066 10124
rect 23661 10115 23719 10121
rect 23661 10112 23673 10115
rect 23584 10084 23673 10112
rect 21269 10047 21327 10053
rect 21269 10044 21281 10047
rect 18840 10016 21281 10044
rect 18840 10004 18846 10016
rect 21269 10013 21281 10016
rect 21315 10013 21327 10047
rect 21269 10007 21327 10013
rect 21450 10004 21456 10056
rect 21508 10044 21514 10056
rect 21732 10047 21790 10053
rect 21732 10044 21744 10047
rect 21508 10016 21744 10044
rect 21508 10004 21514 10016
rect 21732 10013 21744 10016
rect 21778 10013 21790 10047
rect 21732 10007 21790 10013
rect 21910 10004 21916 10056
rect 21968 10044 21974 10056
rect 23474 10044 23480 10056
rect 21968 10016 23480 10044
rect 21968 10004 21974 10016
rect 23474 10004 23480 10016
rect 23532 10004 23538 10056
rect 23584 9988 23612 10084
rect 23661 10081 23673 10084
rect 23707 10112 23719 10115
rect 24029 10115 24087 10121
rect 24029 10112 24041 10115
rect 23707 10084 24041 10112
rect 23707 10081 23719 10084
rect 23661 10075 23719 10081
rect 24029 10081 24041 10084
rect 24075 10081 24087 10115
rect 24136 10112 24164 10152
rect 26510 10140 26516 10152
rect 26568 10140 26574 10192
rect 30282 10140 30288 10192
rect 30340 10180 30346 10192
rect 30340 10152 30604 10180
rect 30340 10140 30346 10152
rect 24486 10121 24492 10124
rect 24448 10115 24492 10121
rect 24448 10112 24460 10115
rect 24136 10084 24460 10112
rect 24029 10075 24087 10081
rect 24448 10081 24460 10084
rect 24448 10075 24492 10081
rect 24486 10072 24492 10075
rect 24544 10072 24550 10124
rect 24599 10084 24992 10112
rect 24599 10053 24627 10084
rect 24964 10056 24992 10084
rect 25130 10072 25136 10124
rect 25188 10072 25194 10124
rect 26237 10115 26295 10121
rect 26237 10081 26249 10115
rect 26283 10112 26295 10115
rect 26283 10084 26924 10112
rect 26283 10081 26295 10084
rect 26237 10075 26295 10081
rect 24121 10047 24179 10053
rect 24121 10013 24133 10047
rect 24167 10013 24179 10047
rect 24599 10047 24658 10053
rect 24599 10016 24612 10047
rect 24121 10007 24179 10013
rect 24600 10013 24612 10016
rect 24646 10013 24658 10047
rect 24600 10007 24658 10013
rect 16776 9948 17172 9976
rect 18708 9948 20392 9976
rect 15749 9939 15807 9945
rect 8588 9908 8616 9936
rect 2746 9880 8616 9908
rect 10689 9911 10747 9917
rect 891 9877 903 9880
rect 845 9871 903 9877
rect 10689 9877 10701 9911
rect 10735 9908 10747 9911
rect 11146 9908 11152 9920
rect 10735 9880 11152 9908
rect 10735 9877 10747 9880
rect 10689 9871 10747 9877
rect 11146 9868 11152 9880
rect 11204 9868 11210 9920
rect 12158 9868 12164 9920
rect 12216 9908 12222 9920
rect 12805 9911 12863 9917
rect 12805 9908 12817 9911
rect 12216 9880 12817 9908
rect 12216 9868 12222 9880
rect 12805 9877 12817 9880
rect 12851 9877 12863 9911
rect 12805 9871 12863 9877
rect 15378 9868 15384 9920
rect 15436 9868 15442 9920
rect 16114 9868 16120 9920
rect 16172 9868 16178 9920
rect 16577 9911 16635 9917
rect 16577 9877 16589 9911
rect 16623 9908 16635 9911
rect 16942 9908 16948 9920
rect 16623 9880 16948 9908
rect 16623 9877 16635 9880
rect 16577 9871 16635 9877
rect 16942 9868 16948 9880
rect 17000 9868 17006 9920
rect 17144 9908 17172 9948
rect 18046 9908 18052 9920
rect 17144 9880 18052 9908
rect 18046 9868 18052 9880
rect 18104 9868 18110 9920
rect 19518 9868 19524 9920
rect 19576 9908 19582 9920
rect 19978 9908 19984 9920
rect 19576 9880 19984 9908
rect 19576 9868 19582 9880
rect 19978 9868 19984 9880
rect 20036 9868 20042 9920
rect 20364 9908 20392 9948
rect 23566 9936 23572 9988
rect 23624 9936 23630 9988
rect 23658 9908 23664 9920
rect 20364 9880 23664 9908
rect 23658 9868 23664 9880
rect 23716 9868 23722 9920
rect 24136 9908 24164 10007
rect 24854 10004 24860 10056
rect 24912 10004 24918 10056
rect 24946 10004 24952 10056
rect 25004 10004 25010 10056
rect 25148 10044 25176 10072
rect 26418 10044 26424 10056
rect 25148 10016 26424 10044
rect 26418 10004 26424 10016
rect 26476 10004 26482 10056
rect 26602 10004 26608 10056
rect 26660 10044 26666 10056
rect 26896 10053 26924 10084
rect 28166 10072 28172 10124
rect 28224 10112 28230 10124
rect 28629 10115 28687 10121
rect 28629 10112 28641 10115
rect 28224 10084 28641 10112
rect 28224 10072 28230 10084
rect 28629 10081 28641 10084
rect 28675 10081 28687 10115
rect 28629 10075 28687 10081
rect 28902 10072 28908 10124
rect 28960 10072 28966 10124
rect 30576 10121 30604 10152
rect 30561 10115 30619 10121
rect 30561 10081 30573 10115
rect 30607 10081 30619 10115
rect 30561 10075 30619 10081
rect 26748 10047 26806 10053
rect 26748 10044 26760 10047
rect 26660 10016 26760 10044
rect 26660 10004 26666 10016
rect 26748 10013 26760 10016
rect 26794 10013 26806 10047
rect 26748 10007 26806 10013
rect 26884 10047 26942 10053
rect 26884 10013 26896 10047
rect 26930 10013 26942 10047
rect 26884 10007 26942 10013
rect 27157 10047 27215 10053
rect 27157 10013 27169 10047
rect 27203 10044 27215 10047
rect 28258 10044 28264 10056
rect 27203 10016 28264 10044
rect 27203 10013 27215 10016
rect 27157 10007 27215 10013
rect 28258 10004 28264 10016
rect 28316 10004 28322 10056
rect 24302 9908 24308 9920
rect 24136 9880 24308 9908
rect 24302 9868 24308 9880
rect 24360 9908 24366 9920
rect 26050 9908 26056 9920
rect 24360 9880 26056 9908
rect 24360 9868 24366 9880
rect 26050 9868 26056 9880
rect 26108 9868 26114 9920
rect 28166 9868 28172 9920
rect 28224 9908 28230 9920
rect 28261 9911 28319 9917
rect 28261 9908 28273 9911
rect 28224 9880 28273 9908
rect 28224 9868 28230 9880
rect 28261 9877 28273 9880
rect 28307 9877 28319 9911
rect 28261 9871 28319 9877
rect 30374 9868 30380 9920
rect 30432 9868 30438 9920
rect 552 9818 30912 9840
rect 552 9766 4193 9818
rect 4245 9766 4257 9818
rect 4309 9766 4321 9818
rect 4373 9766 4385 9818
rect 4437 9766 4449 9818
rect 4501 9766 11783 9818
rect 11835 9766 11847 9818
rect 11899 9766 11911 9818
rect 11963 9766 11975 9818
rect 12027 9766 12039 9818
rect 12091 9766 19373 9818
rect 19425 9766 19437 9818
rect 19489 9766 19501 9818
rect 19553 9766 19565 9818
rect 19617 9766 19629 9818
rect 19681 9766 26963 9818
rect 27015 9766 27027 9818
rect 27079 9766 27091 9818
rect 27143 9766 27155 9818
rect 27207 9766 27219 9818
rect 27271 9766 30912 9818
rect 552 9744 30912 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 2038 9704 2044 9716
rect 1452 9676 2044 9704
rect 1452 9664 1458 9676
rect 2038 9664 2044 9676
rect 2096 9664 2102 9716
rect 2590 9664 2596 9716
rect 2648 9704 2654 9716
rect 5718 9704 5724 9716
rect 2648 9676 5724 9704
rect 2648 9664 2654 9676
rect 5718 9664 5724 9676
rect 5776 9664 5782 9716
rect 5813 9707 5871 9713
rect 5813 9673 5825 9707
rect 5859 9704 5871 9707
rect 6270 9704 6276 9716
rect 5859 9676 6276 9704
rect 5859 9673 5871 9676
rect 5813 9667 5871 9673
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 6454 9664 6460 9716
rect 6512 9704 6518 9716
rect 8754 9704 8760 9716
rect 6512 9676 7512 9704
rect 6512 9664 6518 9676
rect 7484 9636 7512 9676
rect 8312 9676 8760 9704
rect 8312 9636 8340 9676
rect 8754 9664 8760 9676
rect 8812 9664 8818 9716
rect 8846 9664 8852 9716
rect 8904 9704 8910 9716
rect 10318 9704 10324 9716
rect 8904 9676 10324 9704
rect 8904 9664 8910 9676
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 12802 9704 12808 9716
rect 10612 9676 12808 9704
rect 7484 9608 8340 9636
rect 937 9571 995 9577
rect 937 9537 949 9571
rect 983 9568 995 9571
rect 1302 9568 1308 9580
rect 983 9540 1308 9568
rect 983 9537 995 9540
rect 937 9531 995 9537
rect 1302 9528 1308 9540
rect 1360 9528 1366 9580
rect 1443 9571 1501 9577
rect 1443 9537 1455 9571
rect 1489 9568 1501 9571
rect 3053 9571 3111 9577
rect 1489 9540 2774 9568
rect 1489 9537 1501 9540
rect 1443 9531 1501 9537
rect 1026 9460 1032 9512
rect 1084 9500 1090 9512
rect 1673 9503 1731 9509
rect 1673 9500 1685 9503
rect 1084 9472 1685 9500
rect 1084 9460 1090 9472
rect 1673 9469 1685 9472
rect 1719 9469 1731 9503
rect 1673 9463 1731 9469
rect 2746 9432 2774 9540
rect 3053 9537 3065 9571
rect 3099 9568 3111 9571
rect 4068 9571 4126 9577
rect 4068 9568 4080 9571
rect 3099 9540 4080 9568
rect 3099 9537 3111 9540
rect 3053 9531 3111 9537
rect 4068 9537 4080 9540
rect 4114 9537 4126 9571
rect 4068 9531 4126 9537
rect 4706 9528 4712 9580
rect 4764 9568 4770 9580
rect 6454 9568 6460 9580
rect 4764 9540 6460 9568
rect 4764 9528 4770 9540
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 3970 9509 3976 9512
rect 3605 9503 3663 9509
rect 3605 9500 3617 9503
rect 3476 9472 3617 9500
rect 3476 9460 3482 9472
rect 3605 9469 3617 9472
rect 3651 9469 3663 9503
rect 3605 9463 3663 9469
rect 3932 9503 3976 9509
rect 3932 9469 3944 9503
rect 3932 9463 3976 9469
rect 3970 9460 3976 9463
rect 4028 9460 4034 9512
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9500 4399 9503
rect 5166 9500 5172 9512
rect 4387 9472 5172 9500
rect 4387 9469 4399 9472
rect 4341 9463 4399 9469
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 6012 9509 6040 9540
rect 6454 9528 6460 9540
rect 6512 9528 6518 9580
rect 6595 9571 6653 9577
rect 6595 9537 6607 9571
rect 6641 9568 6653 9571
rect 7006 9568 7012 9580
rect 6641 9540 7012 9568
rect 6641 9537 6653 9540
rect 6595 9531 6653 9537
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 8573 9571 8631 9577
rect 8573 9568 8585 9571
rect 8536 9540 8585 9568
rect 8536 9528 8542 9540
rect 8573 9537 8585 9540
rect 8619 9537 8631 9571
rect 8573 9531 8631 9537
rect 9079 9571 9137 9577
rect 9079 9537 9091 9571
rect 9125 9568 9137 9571
rect 9125 9540 9260 9568
rect 9125 9537 9137 9540
rect 9079 9531 9137 9537
rect 9232 9512 9260 9540
rect 10502 9528 10508 9580
rect 10560 9528 10566 9580
rect 5997 9503 6055 9509
rect 5997 9469 6009 9503
rect 6043 9469 6055 9503
rect 5997 9463 6055 9469
rect 6089 9503 6147 9509
rect 6089 9469 6101 9503
rect 6135 9500 6147 9503
rect 6730 9500 6736 9512
rect 6135 9472 6736 9500
rect 6135 9469 6147 9472
rect 6089 9463 6147 9469
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 8386 9500 8392 9512
rect 6871 9472 8392 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 9214 9460 9220 9512
rect 9272 9460 9278 9512
rect 9309 9503 9367 9509
rect 9309 9469 9321 9503
rect 9355 9500 9367 9503
rect 10520 9500 10548 9528
rect 9355 9472 10548 9500
rect 9355 9469 9367 9472
rect 9309 9463 9367 9469
rect 2746 9404 3556 9432
rect 1403 9367 1461 9373
rect 1403 9333 1415 9367
rect 1449 9364 1461 9367
rect 1762 9364 1768 9376
rect 1449 9336 1768 9364
rect 1449 9333 1461 9336
rect 1403 9327 1461 9333
rect 1762 9324 1768 9336
rect 1820 9324 1826 9376
rect 1946 9324 1952 9376
rect 2004 9364 2010 9376
rect 3418 9364 3424 9376
rect 2004 9336 3424 9364
rect 2004 9324 2010 9336
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 3528 9373 3556 9404
rect 5074 9392 5080 9444
rect 5132 9392 5138 9444
rect 5721 9435 5779 9441
rect 5721 9401 5733 9435
rect 5767 9432 5779 9435
rect 5902 9432 5908 9444
rect 5767 9404 5908 9432
rect 5767 9401 5779 9404
rect 5721 9395 5779 9401
rect 5902 9392 5908 9404
rect 5960 9392 5966 9444
rect 7834 9392 7840 9444
rect 7892 9392 7898 9444
rect 8205 9435 8263 9441
rect 8205 9401 8217 9435
rect 8251 9401 8263 9435
rect 8205 9395 8263 9401
rect 3513 9367 3571 9373
rect 3513 9333 3525 9367
rect 3559 9364 3571 9367
rect 5092 9364 5120 9392
rect 3559 9336 5120 9364
rect 3559 9333 3571 9336
rect 3513 9327 3571 9333
rect 5350 9324 5356 9376
rect 5408 9364 5414 9376
rect 6362 9364 6368 9376
rect 5408 9336 6368 9364
rect 5408 9324 5414 9336
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 6555 9367 6613 9373
rect 6555 9333 6567 9367
rect 6601 9364 6613 9367
rect 7852 9364 7880 9392
rect 6601 9336 7880 9364
rect 8220 9364 8248 9395
rect 8938 9364 8944 9376
rect 8220 9336 8944 9364
rect 6601 9333 6613 9336
rect 6555 9327 6613 9333
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9030 9324 9036 9376
rect 9088 9373 9094 9376
rect 9088 9364 9097 9373
rect 9582 9364 9588 9376
rect 9088 9336 9588 9364
rect 9088 9327 9097 9336
rect 9088 9324 9094 9327
rect 9582 9324 9588 9336
rect 9640 9364 9646 9376
rect 10612 9364 10640 9676
rect 12802 9664 12808 9676
rect 12860 9664 12866 9716
rect 12986 9664 12992 9716
rect 13044 9704 13050 9716
rect 13446 9704 13452 9716
rect 13044 9676 13452 9704
rect 13044 9664 13050 9676
rect 13446 9664 13452 9676
rect 13504 9704 13510 9716
rect 15470 9704 15476 9716
rect 13504 9676 15476 9704
rect 13504 9664 13510 9676
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 17770 9664 17776 9716
rect 17828 9664 17834 9716
rect 19150 9664 19156 9716
rect 19208 9704 19214 9716
rect 23750 9704 23756 9716
rect 19208 9676 23756 9704
rect 19208 9664 19214 9676
rect 23750 9664 23756 9676
rect 23808 9664 23814 9716
rect 25222 9704 25228 9716
rect 23860 9676 25228 9704
rect 17788 9636 17816 9664
rect 18233 9639 18291 9645
rect 18233 9636 18245 9639
rect 17788 9608 18245 9636
rect 18233 9605 18245 9608
rect 18279 9605 18291 9639
rect 18233 9599 18291 9605
rect 20530 9596 20536 9648
rect 20588 9596 20594 9648
rect 22370 9596 22376 9648
rect 22428 9636 22434 9648
rect 22741 9639 22799 9645
rect 22741 9636 22753 9639
rect 22428 9608 22753 9636
rect 22428 9596 22434 9608
rect 22741 9605 22753 9608
rect 22787 9605 22799 9639
rect 22741 9599 22799 9605
rect 23106 9596 23112 9648
rect 23164 9636 23170 9648
rect 23201 9639 23259 9645
rect 23201 9636 23213 9639
rect 23164 9608 23213 9636
rect 23164 9596 23170 9608
rect 23201 9605 23213 9608
rect 23247 9605 23259 9639
rect 23201 9599 23259 9605
rect 23477 9639 23535 9645
rect 23477 9605 23489 9639
rect 23523 9636 23535 9639
rect 23860 9636 23888 9676
rect 25222 9664 25228 9676
rect 25280 9664 25286 9716
rect 25682 9664 25688 9716
rect 25740 9664 25746 9716
rect 28258 9664 28264 9716
rect 28316 9664 28322 9716
rect 29454 9704 29460 9716
rect 29012 9676 29460 9704
rect 23523 9608 23888 9636
rect 23523 9605 23535 9608
rect 23477 9599 23535 9605
rect 27522 9596 27528 9648
rect 27580 9636 27586 9648
rect 28537 9639 28595 9645
rect 28537 9636 28549 9639
rect 27580 9608 28549 9636
rect 27580 9596 27586 9608
rect 28537 9605 28549 9608
rect 28583 9605 28595 9639
rect 28537 9599 28595 9605
rect 10689 9571 10747 9577
rect 10689 9537 10701 9571
rect 10735 9568 10747 9571
rect 10735 9540 11008 9568
rect 10735 9537 10747 9540
rect 10689 9531 10747 9537
rect 10778 9460 10784 9512
rect 10836 9460 10842 9512
rect 10980 9500 11008 9540
rect 11054 9528 11060 9580
rect 11112 9577 11118 9580
rect 11112 9571 11166 9577
rect 11112 9537 11120 9571
rect 11154 9537 11166 9571
rect 11112 9531 11166 9537
rect 11112 9528 11118 9531
rect 11238 9528 11244 9580
rect 11296 9528 11302 9580
rect 11422 9528 11428 9580
rect 11480 9528 11486 9580
rect 13170 9568 13176 9580
rect 13096 9540 13176 9568
rect 11440 9500 11468 9528
rect 10980 9472 11468 9500
rect 11514 9460 11520 9512
rect 11572 9460 11578 9512
rect 13096 9509 13124 9540
rect 13170 9528 13176 9540
rect 13228 9528 13234 9580
rect 13262 9528 13268 9580
rect 13320 9528 13326 9580
rect 13538 9528 13544 9580
rect 13596 9528 13602 9580
rect 14004 9569 14062 9575
rect 14004 9535 14016 9569
rect 14050 9568 14062 9569
rect 14090 9568 14096 9580
rect 14050 9540 14096 9568
rect 14050 9535 14062 9540
rect 14004 9529 14062 9535
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 14277 9571 14335 9577
rect 14277 9537 14289 9571
rect 14323 9568 14335 9571
rect 14642 9568 14648 9580
rect 14323 9540 14648 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 16856 9571 16914 9577
rect 16856 9537 16868 9571
rect 16902 9568 16914 9571
rect 19199 9571 19257 9577
rect 16902 9540 18644 9568
rect 16902 9537 16914 9540
rect 16856 9531 16914 9537
rect 13081 9503 13139 9509
rect 13081 9469 13093 9503
rect 13127 9469 13139 9503
rect 13280 9500 13308 9528
rect 15749 9503 15807 9509
rect 15749 9500 15761 9503
rect 13280 9472 15761 9500
rect 13081 9463 13139 9469
rect 15749 9469 15761 9472
rect 15795 9469 15807 9503
rect 15749 9463 15807 9469
rect 16393 9503 16451 9509
rect 16393 9469 16405 9503
rect 16439 9500 16451 9503
rect 16758 9500 16764 9512
rect 16439 9472 16764 9500
rect 16439 9469 16451 9472
rect 16393 9463 16451 9469
rect 16758 9460 16764 9472
rect 16816 9460 16822 9512
rect 17126 9460 17132 9512
rect 17184 9460 17190 9512
rect 9640 9336 10640 9364
rect 10796 9364 10824 9460
rect 18616 9444 18644 9540
rect 19199 9537 19211 9571
rect 19245 9568 19257 9571
rect 19245 9540 19932 9568
rect 19245 9537 19257 9540
rect 19199 9531 19257 9537
rect 19904 9512 19932 9540
rect 21174 9528 21180 9580
rect 21232 9568 21238 9580
rect 21364 9569 21422 9575
rect 21232 9566 21312 9568
rect 21364 9566 21376 9569
rect 21232 9540 21376 9566
rect 21232 9528 21238 9540
rect 21284 9538 21376 9540
rect 21364 9535 21376 9538
rect 21410 9535 21422 9569
rect 21364 9529 21422 9535
rect 21634 9528 21640 9580
rect 21692 9528 21698 9580
rect 23842 9568 23848 9580
rect 22572 9540 23848 9568
rect 22572 9512 22600 9540
rect 23842 9528 23848 9540
rect 23900 9568 23906 9580
rect 24026 9568 24032 9580
rect 23900 9540 24032 9568
rect 23900 9528 23906 9540
rect 24026 9528 24032 9540
rect 24084 9528 24090 9580
rect 24351 9571 24409 9577
rect 24351 9537 24363 9571
rect 24397 9568 24409 9571
rect 25314 9568 25320 9580
rect 24397 9540 25320 9568
rect 24397 9537 24409 9540
rect 24351 9531 24409 9537
rect 25314 9528 25320 9540
rect 25372 9528 25378 9580
rect 26516 9571 26574 9577
rect 26516 9568 26528 9571
rect 25884 9540 26528 9568
rect 18690 9460 18696 9512
rect 18748 9500 18754 9512
rect 19334 9500 19340 9512
rect 18748 9472 19340 9500
rect 18748 9460 18754 9472
rect 19334 9460 19340 9472
rect 19392 9460 19398 9512
rect 19426 9460 19432 9512
rect 19484 9460 19490 9512
rect 19886 9460 19892 9512
rect 19944 9460 19950 9512
rect 20901 9503 20959 9509
rect 20901 9469 20913 9503
rect 20947 9500 20959 9503
rect 22554 9500 22560 9512
rect 20947 9472 22560 9500
rect 20947 9469 20959 9472
rect 20901 9463 20959 9469
rect 12176 9404 12756 9432
rect 11146 9364 11152 9376
rect 10796 9336 11152 9364
rect 9640 9324 9646 9336
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 12176 9364 12204 9404
rect 11388 9336 12204 9364
rect 11388 9324 11394 9336
rect 12618 9324 12624 9376
rect 12676 9324 12682 9376
rect 12728 9364 12756 9404
rect 13170 9392 13176 9444
rect 13228 9432 13234 9444
rect 13265 9435 13323 9441
rect 13265 9432 13277 9435
rect 13228 9404 13277 9432
rect 13228 9392 13234 9404
rect 13265 9401 13277 9404
rect 13311 9432 13323 9435
rect 13354 9432 13360 9444
rect 13311 9404 13360 9432
rect 13311 9401 13323 9404
rect 13265 9395 13323 9401
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 15657 9435 15715 9441
rect 15657 9401 15669 9435
rect 15703 9432 15715 9435
rect 15930 9432 15936 9444
rect 15703 9404 15936 9432
rect 15703 9401 15715 9404
rect 15657 9395 15715 9401
rect 15930 9392 15936 9404
rect 15988 9392 15994 9444
rect 16025 9435 16083 9441
rect 16025 9401 16037 9435
rect 16071 9401 16083 9435
rect 16025 9395 16083 9401
rect 13906 9364 13912 9376
rect 12728 9336 13912 9364
rect 13906 9324 13912 9336
rect 13964 9364 13970 9376
rect 14007 9367 14065 9373
rect 14007 9364 14019 9367
rect 13964 9336 14019 9364
rect 13964 9324 13970 9336
rect 14007 9333 14019 9336
rect 14053 9364 14065 9367
rect 16040 9364 16068 9395
rect 18598 9392 18604 9444
rect 18656 9392 18662 9444
rect 14053 9336 16068 9364
rect 16859 9367 16917 9373
rect 14053 9333 14065 9336
rect 14007 9327 14065 9333
rect 16859 9333 16871 9367
rect 16905 9364 16917 9367
rect 17218 9364 17224 9376
rect 16905 9336 17224 9364
rect 16905 9333 16917 9336
rect 16859 9327 16917 9333
rect 17218 9324 17224 9336
rect 17276 9364 17282 9376
rect 19058 9364 19064 9376
rect 17276 9336 19064 9364
rect 17276 9324 17282 9336
rect 19058 9324 19064 9336
rect 19116 9364 19122 9376
rect 19159 9367 19217 9373
rect 19159 9364 19171 9367
rect 19116 9336 19171 9364
rect 19116 9324 19122 9336
rect 19159 9333 19171 9336
rect 19205 9333 19217 9367
rect 19159 9327 19217 9333
rect 19334 9324 19340 9376
rect 19392 9364 19398 9376
rect 20916 9364 20944 9463
rect 22554 9460 22560 9472
rect 22612 9460 22618 9512
rect 23385 9503 23443 9509
rect 23385 9469 23397 9503
rect 23431 9469 23443 9503
rect 23385 9463 23443 9469
rect 22370 9392 22376 9444
rect 22428 9432 22434 9444
rect 23400 9432 23428 9463
rect 23474 9460 23480 9512
rect 23532 9500 23538 9512
rect 23661 9503 23719 9509
rect 23661 9500 23673 9503
rect 23532 9472 23673 9500
rect 23532 9460 23538 9472
rect 23661 9469 23673 9472
rect 23707 9469 23719 9503
rect 24486 9500 24492 9512
rect 23661 9463 23719 9469
rect 23768 9472 24492 9500
rect 23768 9432 23796 9472
rect 24486 9460 24492 9472
rect 24544 9460 24550 9512
rect 24581 9503 24639 9509
rect 24581 9469 24593 9503
rect 24627 9500 24639 9503
rect 25682 9500 25688 9512
rect 24627 9472 25688 9500
rect 24627 9469 24639 9472
rect 24581 9463 24639 9469
rect 25682 9460 25688 9472
rect 25740 9460 25746 9512
rect 22428 9404 23796 9432
rect 22428 9392 22434 9404
rect 25884 9376 25912 9540
rect 26516 9537 26528 9540
rect 26562 9537 26574 9571
rect 26516 9531 26574 9537
rect 26970 9528 26976 9580
rect 27028 9568 27034 9580
rect 28902 9568 28908 9580
rect 27028 9540 28908 9568
rect 27028 9528 27034 9540
rect 26050 9460 26056 9512
rect 26108 9460 26114 9512
rect 26418 9460 26424 9512
rect 26476 9500 26482 9512
rect 28460 9509 28488 9540
rect 28902 9528 28908 9540
rect 28960 9528 28966 9580
rect 26789 9503 26847 9509
rect 26789 9500 26801 9503
rect 26476 9472 26801 9500
rect 26476 9460 26482 9472
rect 26789 9469 26801 9472
rect 26835 9469 26847 9503
rect 26789 9463 26847 9469
rect 28445 9503 28503 9509
rect 28445 9469 28457 9503
rect 28491 9469 28503 9503
rect 28445 9463 28503 9469
rect 28721 9503 28779 9509
rect 28721 9469 28733 9503
rect 28767 9500 28779 9503
rect 29012 9500 29040 9676
rect 29454 9664 29460 9676
rect 29512 9704 29518 9716
rect 30282 9704 30288 9716
rect 29512 9676 30288 9704
rect 29512 9664 29518 9676
rect 30282 9664 30288 9676
rect 30340 9664 30346 9716
rect 30009 9639 30067 9645
rect 30009 9605 30021 9639
rect 30055 9636 30067 9639
rect 30650 9636 30656 9648
rect 30055 9608 30656 9636
rect 30055 9605 30067 9608
rect 30009 9599 30067 9605
rect 30650 9596 30656 9608
rect 30708 9596 30714 9648
rect 29086 9528 29092 9580
rect 29144 9568 29150 9580
rect 29144 9540 30236 9568
rect 29144 9528 29150 9540
rect 30208 9509 30236 9540
rect 28767 9472 29040 9500
rect 29181 9503 29239 9509
rect 28767 9469 28779 9472
rect 28721 9463 28779 9469
rect 29181 9469 29193 9503
rect 29227 9500 29239 9503
rect 30193 9503 30251 9509
rect 29227 9472 29408 9500
rect 29227 9469 29239 9472
rect 29181 9463 29239 9469
rect 27522 9392 27528 9444
rect 27580 9432 27586 9444
rect 28736 9432 28764 9463
rect 27580 9404 28764 9432
rect 27580 9392 27586 9404
rect 29380 9376 29408 9472
rect 30193 9469 30205 9503
rect 30239 9469 30251 9503
rect 30193 9463 30251 9469
rect 30469 9503 30527 9509
rect 30469 9469 30481 9503
rect 30515 9469 30527 9503
rect 30469 9463 30527 9469
rect 30484 9432 30512 9463
rect 30116 9404 30512 9432
rect 30116 9376 30144 9404
rect 19392 9336 20944 9364
rect 19392 9324 19398 9336
rect 21358 9324 21364 9376
rect 21416 9373 21422 9376
rect 21416 9364 21425 9373
rect 21416 9336 21461 9364
rect 21416 9327 21425 9336
rect 21416 9324 21422 9327
rect 23750 9324 23756 9376
rect 23808 9364 23814 9376
rect 24311 9367 24369 9373
rect 24311 9364 24323 9367
rect 23808 9336 24323 9364
rect 23808 9324 23814 9336
rect 24311 9333 24323 9336
rect 24357 9333 24369 9367
rect 24311 9327 24369 9333
rect 24486 9324 24492 9376
rect 24544 9364 24550 9376
rect 25774 9364 25780 9376
rect 24544 9336 25780 9364
rect 24544 9324 24550 9336
rect 25774 9324 25780 9336
rect 25832 9324 25838 9376
rect 25866 9324 25872 9376
rect 25924 9324 25930 9376
rect 26510 9324 26516 9376
rect 26568 9373 26574 9376
rect 26568 9327 26577 9373
rect 26568 9324 26574 9327
rect 27890 9324 27896 9376
rect 27948 9324 27954 9376
rect 28994 9324 29000 9376
rect 29052 9324 29058 9376
rect 29362 9324 29368 9376
rect 29420 9324 29426 9376
rect 30098 9324 30104 9376
rect 30156 9324 30162 9376
rect 30282 9324 30288 9376
rect 30340 9324 30346 9376
rect 552 9274 31072 9296
rect 552 9222 7988 9274
rect 8040 9222 8052 9274
rect 8104 9222 8116 9274
rect 8168 9222 8180 9274
rect 8232 9222 8244 9274
rect 8296 9222 15578 9274
rect 15630 9222 15642 9274
rect 15694 9222 15706 9274
rect 15758 9222 15770 9274
rect 15822 9222 15834 9274
rect 15886 9222 23168 9274
rect 23220 9222 23232 9274
rect 23284 9222 23296 9274
rect 23348 9222 23360 9274
rect 23412 9222 23424 9274
rect 23476 9222 30758 9274
rect 30810 9222 30822 9274
rect 30874 9222 30886 9274
rect 30938 9222 30950 9274
rect 31002 9222 31014 9274
rect 31066 9222 31072 9274
rect 552 9200 31072 9222
rect 1302 9120 1308 9172
rect 1360 9120 1366 9172
rect 2866 9120 2872 9172
rect 2924 9169 2930 9172
rect 2924 9160 2933 9169
rect 2924 9132 2969 9160
rect 2924 9123 2933 9132
rect 2924 9120 2930 9123
rect 4614 9120 4620 9172
rect 4672 9120 4678 9172
rect 4724 9132 7144 9160
rect 1029 9095 1087 9101
rect 1029 9092 1041 9095
rect 860 9064 1041 9092
rect 860 8956 888 9064
rect 1029 9061 1041 9064
rect 1075 9061 1087 9095
rect 1946 9092 1952 9104
rect 1029 9055 1087 9061
rect 1596 9064 1952 9092
rect 1596 8956 1624 9064
rect 1946 9052 1952 9064
rect 2004 9052 2010 9104
rect 4525 9095 4583 9101
rect 4525 9061 4537 9095
rect 4571 9092 4583 9095
rect 4724 9092 4752 9132
rect 7116 9092 7144 9132
rect 7190 9120 7196 9172
rect 7248 9160 7254 9172
rect 7285 9163 7343 9169
rect 7285 9160 7297 9163
rect 7248 9132 7297 9160
rect 7248 9120 7254 9132
rect 7285 9129 7297 9132
rect 7331 9129 7343 9163
rect 7285 9123 7343 9129
rect 7558 9120 7564 9172
rect 7616 9120 7622 9172
rect 7650 9120 7656 9172
rect 7708 9120 7714 9172
rect 7834 9120 7840 9172
rect 7892 9160 7898 9172
rect 8027 9163 8085 9169
rect 8027 9160 8039 9163
rect 7892 9132 8039 9160
rect 7892 9120 7898 9132
rect 8027 9129 8039 9132
rect 8073 9129 8085 9163
rect 8027 9123 8085 9129
rect 9214 9120 9220 9172
rect 9272 9160 9278 9172
rect 9401 9163 9459 9169
rect 9401 9160 9413 9163
rect 9272 9132 9413 9160
rect 9272 9120 9278 9132
rect 9401 9129 9413 9132
rect 9447 9129 9459 9163
rect 9401 9123 9459 9129
rect 10321 9163 10379 9169
rect 10321 9129 10333 9163
rect 10367 9160 10379 9163
rect 11514 9160 11520 9172
rect 10367 9132 11520 9160
rect 10367 9129 10379 9132
rect 10321 9123 10379 9129
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 13357 9163 13415 9169
rect 13357 9160 13369 9163
rect 12406 9132 13369 9160
rect 7576 9092 7604 9120
rect 4571 9064 4752 9092
rect 4816 9064 6224 9092
rect 7116 9064 7604 9092
rect 4571 9061 4583 9064
rect 4525 9055 4583 9061
rect 1673 9027 1731 9033
rect 1673 8993 1685 9027
rect 1719 8993 1731 9027
rect 1673 8987 1731 8993
rect 860 8928 1624 8956
rect 1688 8888 1716 8987
rect 1762 8984 1768 9036
rect 1820 8984 1826 9036
rect 2406 8984 2412 9036
rect 2464 8984 2470 9036
rect 4816 9033 4844 9064
rect 5644 9033 5672 9064
rect 4801 9027 4859 9033
rect 4801 9024 4813 9027
rect 2792 8996 4813 9024
rect 1780 8956 1808 8984
rect 1857 8959 1915 8965
rect 1857 8956 1869 8959
rect 1780 8928 1869 8956
rect 1857 8925 1869 8928
rect 1903 8925 1915 8959
rect 2792 8956 2820 8996
rect 4801 8993 4813 8996
rect 4847 8993 4859 9027
rect 4801 8987 4859 8993
rect 5077 9027 5135 9033
rect 5077 8993 5089 9027
rect 5123 8993 5135 9027
rect 5077 8987 5135 8993
rect 5361 9027 5419 9033
rect 5361 8993 5373 9027
rect 5407 8993 5419 9027
rect 5361 8987 5419 8993
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 8993 5687 9027
rect 5997 9027 6055 9033
rect 5997 9024 6009 9027
rect 5629 8987 5687 8993
rect 5736 8996 6009 9024
rect 2958 8967 2964 8968
rect 1857 8919 1915 8925
rect 1964 8928 2820 8956
rect 2915 8961 2964 8967
rect 1964 8900 1992 8928
rect 2915 8927 2927 8961
rect 2961 8927 2964 8961
rect 2915 8921 2964 8927
rect 2958 8916 2964 8921
rect 3016 8916 3022 8968
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8956 3203 8959
rect 3326 8956 3332 8968
rect 3191 8928 3332 8956
rect 3191 8925 3203 8928
rect 3145 8919 3203 8925
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 5092 8900 5120 8987
rect 5368 8900 5396 8987
rect 1762 8888 1768 8900
rect 1688 8860 1768 8888
rect 1762 8848 1768 8860
rect 1820 8848 1826 8900
rect 1946 8848 1952 8900
rect 2004 8848 2010 8900
rect 3804 8860 4844 8888
rect 1670 8780 1676 8832
rect 1728 8820 1734 8832
rect 3804 8820 3832 8860
rect 4816 8832 4844 8860
rect 5074 8848 5080 8900
rect 5132 8888 5138 8900
rect 5132 8860 5304 8888
rect 5132 8848 5138 8860
rect 1728 8792 3832 8820
rect 1728 8780 1734 8792
rect 4798 8780 4804 8832
rect 4856 8780 4862 8832
rect 4890 8780 4896 8832
rect 4948 8780 4954 8832
rect 4982 8780 4988 8832
rect 5040 8820 5046 8832
rect 5169 8823 5227 8829
rect 5169 8820 5181 8823
rect 5040 8792 5181 8820
rect 5040 8780 5046 8792
rect 5169 8789 5181 8792
rect 5215 8789 5227 8823
rect 5276 8820 5304 8860
rect 5350 8848 5356 8900
rect 5408 8848 5414 8900
rect 5442 8848 5448 8900
rect 5500 8848 5506 8900
rect 5736 8820 5764 8996
rect 5997 8993 6009 8996
rect 6043 9024 6055 9027
rect 6086 9024 6092 9036
rect 6043 8996 6092 9024
rect 6043 8993 6055 8996
rect 5997 8987 6055 8993
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 6196 8956 6224 9064
rect 6362 8984 6368 9036
rect 6420 8984 6426 9036
rect 6638 8984 6644 9036
rect 6696 8984 6702 9036
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 8993 6975 9027
rect 6917 8987 6975 8993
rect 6932 8956 6960 8987
rect 7190 8984 7196 9036
rect 7248 8984 7254 9036
rect 7466 8984 7472 9036
rect 7524 8984 7530 9036
rect 6196 8928 6960 8956
rect 6181 8891 6239 8897
rect 6181 8857 6193 8891
rect 6227 8888 6239 8891
rect 6270 8888 6276 8900
rect 6227 8860 6276 8888
rect 6227 8857 6239 8860
rect 6181 8851 6239 8857
rect 6270 8848 6276 8860
rect 6328 8848 6334 8900
rect 6733 8891 6791 8897
rect 6733 8888 6745 8891
rect 6380 8860 6745 8888
rect 6380 8832 6408 8860
rect 6733 8857 6745 8860
rect 6779 8857 6791 8891
rect 6932 8888 6960 8928
rect 7006 8916 7012 8968
rect 7064 8956 7070 8968
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 7064 8928 7573 8956
rect 7064 8916 7070 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7668 8956 7696 9120
rect 12406 9036 12434 9132
rect 13357 9129 13369 9132
rect 13403 9129 13415 9163
rect 13357 9123 13415 9129
rect 13906 9120 13912 9172
rect 13964 9160 13970 9172
rect 14007 9163 14065 9169
rect 14007 9160 14019 9163
rect 13964 9132 14019 9160
rect 13964 9120 13970 9132
rect 14007 9129 14019 9132
rect 14053 9129 14065 9163
rect 14007 9123 14065 9129
rect 15654 9120 15660 9172
rect 15712 9160 15718 9172
rect 16114 9160 16120 9172
rect 15712 9132 16120 9160
rect 15712 9120 15718 9132
rect 16114 9120 16120 9132
rect 16172 9120 16178 9172
rect 16577 9163 16635 9169
rect 16577 9129 16589 9163
rect 16623 9160 16635 9163
rect 17126 9160 17132 9172
rect 16623 9132 17132 9160
rect 16623 9129 16635 9132
rect 16577 9123 16635 9129
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 17218 9120 17224 9172
rect 17276 9160 17282 9172
rect 17319 9163 17377 9169
rect 17319 9160 17331 9163
rect 17276 9132 17331 9160
rect 17276 9120 17282 9132
rect 17319 9129 17331 9132
rect 17365 9129 17377 9163
rect 17319 9123 17377 9129
rect 17862 9120 17868 9172
rect 17920 9160 17926 9172
rect 18693 9163 18751 9169
rect 18693 9160 18705 9163
rect 17920 9132 18705 9160
rect 17920 9120 17926 9132
rect 18693 9129 18705 9132
rect 18739 9129 18751 9163
rect 18693 9123 18751 9129
rect 19061 9163 19119 9169
rect 19061 9129 19073 9163
rect 19107 9160 19119 9163
rect 19426 9160 19432 9172
rect 19107 9132 19432 9160
rect 19107 9129 19119 9132
rect 19061 9123 19119 9129
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 20257 9163 20315 9169
rect 20257 9129 20269 9163
rect 20303 9160 20315 9163
rect 20438 9160 20444 9172
rect 20303 9132 20444 9160
rect 20303 9129 20315 9132
rect 20257 9123 20315 9129
rect 20438 9120 20444 9132
rect 20496 9120 20502 9172
rect 21269 9163 21327 9169
rect 21269 9129 21281 9163
rect 21315 9160 21327 9163
rect 21634 9160 21640 9172
rect 21315 9132 21640 9160
rect 21315 9129 21327 9132
rect 21269 9123 21327 9129
rect 21634 9120 21640 9132
rect 21692 9120 21698 9172
rect 22002 9120 22008 9172
rect 22060 9160 22066 9172
rect 23566 9160 23572 9172
rect 22060 9132 23572 9160
rect 22060 9120 22066 9132
rect 23566 9120 23572 9132
rect 23624 9120 23630 9172
rect 23658 9120 23664 9172
rect 23716 9160 23722 9172
rect 23716 9132 24348 9160
rect 23716 9120 23722 9132
rect 19150 9052 19156 9104
rect 19208 9092 19214 9104
rect 20625 9095 20683 9101
rect 20625 9092 20637 9095
rect 19208 9064 20637 9092
rect 19208 9052 19214 9064
rect 20625 9061 20637 9064
rect 20671 9092 20683 9095
rect 21358 9092 21364 9104
rect 20671 9064 21364 9092
rect 20671 9061 20683 9064
rect 20625 9055 20683 9061
rect 21358 9052 21364 9064
rect 21416 9092 21422 9104
rect 21416 9064 23060 9092
rect 21416 9052 21422 9064
rect 8202 8984 8208 9036
rect 8260 9024 8266 9036
rect 9861 9027 9919 9033
rect 9861 9024 9873 9027
rect 8260 8996 9873 9024
rect 8260 8984 8266 8996
rect 9861 8993 9873 8996
rect 9907 8993 9919 9027
rect 9861 8987 9919 8993
rect 10502 8984 10508 9036
rect 10560 8984 10566 9036
rect 11330 9033 11336 9036
rect 10781 9027 10839 9033
rect 10781 8993 10793 9027
rect 10827 9024 10839 9027
rect 11292 9027 11336 9033
rect 10827 8996 10916 9024
rect 10827 8993 10839 8996
rect 10781 8987 10839 8993
rect 8024 8977 8082 8983
rect 8024 8956 8036 8977
rect 7668 8943 8036 8956
rect 8070 8943 8082 8977
rect 10888 8968 10916 8996
rect 11292 8993 11304 9027
rect 11292 8987 11336 8993
rect 11330 8984 11336 8987
rect 11388 8984 11394 9036
rect 11606 8984 11612 9036
rect 11664 9024 11670 9036
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 11664 8996 11713 9024
rect 11664 8984 11670 8996
rect 11701 8993 11713 8996
rect 11747 8993 11759 9027
rect 11701 8987 11759 8993
rect 12342 8984 12348 9036
rect 12400 8996 12434 9036
rect 12400 8984 12406 8996
rect 12710 8984 12716 9036
rect 12768 9024 12774 9036
rect 13173 9027 13231 9033
rect 13173 9024 13185 9027
rect 12768 8996 13185 9024
rect 12768 8984 12774 8996
rect 13173 8993 13185 8996
rect 13219 8993 13231 9027
rect 13173 8987 13231 8993
rect 13538 8984 13544 9036
rect 13596 8984 13602 9036
rect 14277 9027 14335 9033
rect 14277 8993 14289 9027
rect 14323 9024 14335 9027
rect 14918 9024 14924 9036
rect 14323 8996 14924 9024
rect 14323 8993 14335 8996
rect 14277 8987 14335 8993
rect 14918 8984 14924 8996
rect 14976 8984 14982 9036
rect 15470 8984 15476 9036
rect 15528 9024 15534 9036
rect 15933 9027 15991 9033
rect 15933 9024 15945 9027
rect 15528 8996 15945 9024
rect 15528 8984 15534 8996
rect 15933 8993 15945 8996
rect 15979 8993 15991 9027
rect 15933 8987 15991 8993
rect 16114 8984 16120 9036
rect 16172 9024 16178 9036
rect 16482 9024 16488 9036
rect 16172 8996 16488 9024
rect 16172 8984 16178 8996
rect 16482 8984 16488 8996
rect 16540 8984 16546 9036
rect 16666 8984 16672 9036
rect 16724 9024 16730 9036
rect 16761 9027 16819 9033
rect 16761 9024 16773 9027
rect 16724 8996 16773 9024
rect 16724 8984 16730 8996
rect 16761 8993 16773 8996
rect 16807 8993 16819 9027
rect 16761 8987 16819 8993
rect 16942 8984 16948 9036
rect 17000 9024 17006 9036
rect 17589 9027 17647 9033
rect 17589 9024 17601 9027
rect 17000 8996 17601 9024
rect 17000 8984 17006 8996
rect 17589 8993 17601 8996
rect 17635 8993 17647 9027
rect 17589 8987 17647 8993
rect 18782 8984 18788 9036
rect 18840 9024 18846 9036
rect 19245 9027 19303 9033
rect 19245 9024 19257 9027
rect 18840 8996 19257 9024
rect 18840 8984 18846 8996
rect 19245 8993 19257 8996
rect 19291 8993 19303 9027
rect 19245 8987 19303 8993
rect 19521 9027 19579 9033
rect 19521 8993 19533 9027
rect 19567 9024 19579 9027
rect 19567 8996 19748 9024
rect 19567 8993 19579 8996
rect 19521 8987 19579 8993
rect 7668 8937 8082 8943
rect 7668 8928 8067 8937
rect 7561 8919 7619 8925
rect 8294 8916 8300 8968
rect 8352 8916 8358 8968
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 10870 8956 10876 8968
rect 8536 8928 9168 8956
rect 8536 8916 8542 8928
rect 9140 8888 9168 8928
rect 9508 8928 10876 8956
rect 9398 8888 9404 8900
rect 6932 8860 7144 8888
rect 9140 8860 9404 8888
rect 6733 8851 6791 8857
rect 5276 8792 5764 8820
rect 5169 8783 5227 8789
rect 5810 8780 5816 8832
rect 5868 8780 5874 8832
rect 6362 8780 6368 8832
rect 6420 8780 6426 8832
rect 6454 8780 6460 8832
rect 6512 8780 6518 8832
rect 7006 8780 7012 8832
rect 7064 8780 7070 8832
rect 7116 8820 7144 8860
rect 9398 8848 9404 8860
rect 9456 8848 9462 8900
rect 8478 8820 8484 8832
rect 7116 8792 8484 8820
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 8662 8780 8668 8832
rect 8720 8820 8726 8832
rect 9508 8820 9536 8928
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8956 11023 8959
rect 11146 8956 11152 8968
rect 11011 8928 11152 8956
rect 11011 8925 11023 8928
rect 10965 8919 11023 8925
rect 11146 8916 11152 8928
rect 11204 8916 11210 8968
rect 11428 8961 11486 8967
rect 11428 8927 11440 8961
rect 11474 8956 11486 8961
rect 11514 8956 11520 8968
rect 11474 8928 11520 8956
rect 11474 8927 11486 8928
rect 11428 8921 11486 8927
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 12802 8916 12808 8968
rect 12860 8956 12866 8968
rect 13078 8956 13084 8968
rect 12860 8928 13084 8956
rect 12860 8916 12866 8928
rect 13078 8916 13084 8928
rect 13136 8916 13142 8968
rect 14047 8959 14105 8965
rect 14047 8925 14059 8959
rect 14093 8956 14105 8959
rect 15194 8956 15200 8968
rect 14093 8928 15200 8956
rect 14093 8925 14105 8928
rect 14047 8919 14105 8925
rect 15194 8916 15200 8928
rect 15252 8916 15258 8968
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8956 16911 8959
rect 17126 8956 17132 8968
rect 16899 8928 17132 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 17359 8959 17417 8965
rect 17359 8925 17371 8959
rect 17405 8956 17417 8959
rect 17405 8928 19472 8956
rect 17405 8925 17417 8928
rect 17359 8919 17417 8925
rect 10594 8848 10600 8900
rect 10652 8848 10658 8900
rect 15470 8848 15476 8900
rect 15528 8888 15534 8900
rect 15749 8891 15807 8897
rect 15749 8888 15761 8891
rect 15528 8860 15761 8888
rect 15528 8848 15534 8860
rect 15749 8857 15761 8860
rect 15795 8857 15807 8891
rect 15749 8851 15807 8857
rect 8720 8792 9536 8820
rect 10137 8823 10195 8829
rect 8720 8780 8726 8792
rect 10137 8789 10149 8823
rect 10183 8820 10195 8823
rect 11330 8820 11336 8832
rect 10183 8792 11336 8820
rect 10183 8789 10195 8792
rect 10137 8783 10195 8789
rect 11330 8780 11336 8792
rect 11388 8780 11394 8832
rect 12342 8780 12348 8832
rect 12400 8820 12406 8832
rect 12805 8823 12863 8829
rect 12805 8820 12817 8823
rect 12400 8792 12817 8820
rect 12400 8780 12406 8792
rect 12805 8789 12817 8792
rect 12851 8789 12863 8823
rect 12805 8783 12863 8789
rect 15562 8780 15568 8832
rect 15620 8780 15626 8832
rect 16393 8823 16451 8829
rect 16393 8789 16405 8823
rect 16439 8820 16451 8823
rect 16482 8820 16488 8832
rect 16439 8792 16488 8820
rect 16439 8789 16451 8792
rect 16393 8783 16451 8789
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 19242 8780 19248 8832
rect 19300 8820 19306 8832
rect 19337 8823 19395 8829
rect 19337 8820 19349 8823
rect 19300 8792 19349 8820
rect 19300 8780 19306 8792
rect 19337 8789 19349 8792
rect 19383 8789 19395 8823
rect 19444 8820 19472 8928
rect 19720 8900 19748 8996
rect 19978 8984 19984 9036
rect 20036 9024 20042 9036
rect 20349 9027 20407 9033
rect 20349 9024 20361 9027
rect 20036 8996 20361 9024
rect 20036 8984 20042 8996
rect 20349 8993 20361 8996
rect 20395 8993 20407 9027
rect 20349 8987 20407 8993
rect 20364 8956 20392 8987
rect 20530 8984 20536 9036
rect 20588 9024 20594 9036
rect 21453 9027 21511 9033
rect 21453 9024 21465 9027
rect 20588 8996 21465 9024
rect 20588 8984 20594 8996
rect 21453 8993 21465 8996
rect 21499 9024 21511 9027
rect 22002 9024 22008 9036
rect 21499 8996 22008 9024
rect 21499 8993 21511 8996
rect 21453 8987 21511 8993
rect 22002 8984 22008 8996
rect 22060 8984 22066 9036
rect 22189 9027 22247 9033
rect 22189 8993 22201 9027
rect 22235 9024 22247 9027
rect 22278 9024 22284 9036
rect 22235 8996 22284 9024
rect 22235 8993 22247 8996
rect 22189 8987 22247 8993
rect 22278 8984 22284 8996
rect 22336 8984 22342 9036
rect 22465 9027 22523 9033
rect 22465 8993 22477 9027
rect 22511 8993 22523 9027
rect 22465 8987 22523 8993
rect 20622 8956 20628 8968
rect 20364 8928 20628 8956
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 19702 8848 19708 8900
rect 19760 8848 19766 8900
rect 19889 8891 19947 8897
rect 19889 8857 19901 8891
rect 19935 8888 19947 8891
rect 20346 8888 20352 8900
rect 19935 8860 20352 8888
rect 19935 8857 19947 8860
rect 19889 8851 19947 8857
rect 20346 8848 20352 8860
rect 20404 8848 20410 8900
rect 21910 8848 21916 8900
rect 21968 8888 21974 8900
rect 22480 8888 22508 8987
rect 22554 8984 22560 9036
rect 22612 9024 22618 9036
rect 22925 9027 22983 9033
rect 22925 9024 22937 9027
rect 22612 8996 22937 9024
rect 22612 8984 22618 8996
rect 22925 8993 22937 8996
rect 22971 8993 22983 9027
rect 23032 9024 23060 9064
rect 23252 9027 23310 9033
rect 23252 9024 23264 9027
rect 23032 8996 23264 9024
rect 22925 8987 22983 8993
rect 23252 8993 23264 8996
rect 23298 9024 23310 9027
rect 23750 9024 23756 9036
rect 23298 8996 23756 9024
rect 23298 8993 23310 8996
rect 23252 8987 23310 8993
rect 23750 8984 23756 8996
rect 23808 8984 23814 9036
rect 24320 9024 24348 9132
rect 24854 9120 24860 9172
rect 24912 9120 24918 9172
rect 24946 9120 24952 9172
rect 25004 9120 25010 9172
rect 25682 9120 25688 9172
rect 25740 9120 25746 9172
rect 25961 9163 26019 9169
rect 25961 9129 25973 9163
rect 26007 9129 26019 9163
rect 27522 9160 27528 9172
rect 25961 9123 26019 9129
rect 26068 9132 27528 9160
rect 24872 9092 24900 9120
rect 25976 9092 26004 9123
rect 24872 9064 26004 9092
rect 25317 9027 25375 9033
rect 24320 8996 25268 9024
rect 23431 8959 23489 8965
rect 23431 8925 23443 8959
rect 23477 8956 23489 8959
rect 23566 8956 23572 8968
rect 23477 8928 23572 8956
rect 23477 8925 23489 8928
rect 23431 8919 23489 8925
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 23661 8959 23719 8965
rect 23661 8925 23673 8959
rect 23707 8956 23719 8959
rect 23707 8928 25176 8956
rect 23707 8925 23719 8928
rect 23661 8919 23719 8925
rect 21968 8860 22508 8888
rect 21968 8848 21974 8860
rect 22646 8848 22652 8900
rect 22704 8848 22710 8900
rect 25148 8897 25176 8928
rect 25133 8891 25191 8897
rect 25133 8857 25145 8891
rect 25179 8857 25191 8891
rect 25240 8888 25268 8996
rect 25317 8993 25329 9027
rect 25363 9024 25375 9027
rect 25363 8996 25544 9024
rect 25363 8993 25375 8996
rect 25317 8987 25375 8993
rect 25516 8968 25544 8996
rect 25590 8984 25596 9036
rect 25648 8984 25654 9036
rect 25774 8984 25780 9036
rect 25832 9024 25838 9036
rect 25869 9027 25927 9033
rect 25869 9024 25881 9027
rect 25832 8996 25881 9024
rect 25832 8984 25838 8996
rect 25869 8993 25881 8996
rect 25915 9024 25927 9027
rect 26068 9024 26096 9132
rect 27522 9120 27528 9132
rect 27580 9120 27586 9172
rect 27890 9120 27896 9172
rect 27948 9120 27954 9172
rect 28994 9160 29000 9172
rect 28092 9132 29000 9160
rect 25915 8996 26096 9024
rect 25915 8993 25927 8996
rect 25869 8987 25927 8993
rect 26142 8984 26148 9036
rect 26200 8984 26206 9036
rect 26326 8984 26332 9036
rect 26384 9024 26390 9036
rect 26421 9027 26479 9033
rect 26421 9024 26433 9027
rect 26384 8996 26433 9024
rect 26384 8984 26390 8996
rect 26421 8993 26433 8996
rect 26467 8993 26479 9027
rect 27908 9024 27936 9120
rect 26421 8987 26479 8993
rect 27080 8996 27936 9024
rect 25498 8916 25504 8968
rect 25556 8956 25562 8968
rect 26160 8956 26188 8984
rect 25556 8928 26188 8956
rect 25556 8916 25562 8928
rect 26602 8916 26608 8968
rect 26660 8956 26666 8968
rect 26748 8959 26806 8965
rect 26748 8956 26760 8959
rect 26660 8928 26760 8956
rect 26660 8916 26666 8928
rect 26748 8925 26760 8928
rect 26794 8925 26806 8959
rect 26748 8919 26806 8925
rect 26927 8959 26985 8965
rect 26927 8925 26939 8959
rect 26973 8956 26985 8959
rect 27080 8956 27108 8996
rect 26973 8928 27108 8956
rect 27157 8959 27215 8965
rect 26973 8925 26985 8928
rect 26927 8919 26985 8925
rect 27157 8925 27169 8959
rect 27203 8956 27215 8959
rect 28092 8956 28120 9132
rect 28994 9120 29000 9132
rect 29052 9120 29058 9172
rect 29270 9120 29276 9172
rect 29328 9160 29334 9172
rect 30009 9163 30067 9169
rect 30009 9160 30021 9163
rect 29328 9132 30021 9160
rect 29328 9120 29334 9132
rect 30009 9129 30021 9132
rect 30055 9129 30067 9163
rect 30009 9123 30067 9129
rect 30377 9163 30435 9169
rect 30377 9129 30389 9163
rect 30423 9160 30435 9163
rect 30466 9160 30472 9172
rect 30423 9132 30472 9160
rect 30423 9129 30435 9132
rect 30377 9123 30435 9129
rect 30466 9120 30472 9132
rect 30524 9120 30530 9172
rect 29822 9052 29828 9104
rect 29880 9092 29886 9104
rect 30190 9092 30196 9104
rect 29880 9064 30196 9092
rect 29880 9052 29886 9064
rect 30190 9052 30196 9064
rect 30248 9092 30254 9104
rect 30248 9064 30604 9092
rect 30248 9052 30254 9064
rect 28626 8984 28632 9036
rect 28684 8984 28690 9036
rect 28905 9027 28963 9033
rect 28905 8993 28917 9027
rect 28951 9024 28963 9027
rect 30006 9024 30012 9036
rect 28951 8996 30012 9024
rect 28951 8993 28963 8996
rect 28905 8987 28963 8993
rect 30006 8984 30012 8996
rect 30064 8984 30070 9036
rect 30576 9033 30604 9064
rect 30561 9027 30619 9033
rect 30561 8993 30573 9027
rect 30607 8993 30619 9027
rect 30561 8987 30619 8993
rect 27203 8928 28120 8956
rect 27203 8925 27215 8928
rect 27157 8919 27215 8925
rect 29362 8916 29368 8968
rect 29420 8956 29426 8968
rect 29546 8956 29552 8968
rect 29420 8928 29552 8956
rect 29420 8916 29426 8928
rect 29546 8916 29552 8928
rect 29604 8916 29610 8968
rect 25240 8860 25544 8888
rect 25133 8851 25191 8857
rect 20806 8820 20812 8832
rect 19444 8792 20812 8820
rect 19337 8783 19395 8789
rect 20806 8780 20812 8792
rect 20864 8780 20870 8832
rect 22005 8823 22063 8829
rect 22005 8789 22017 8823
rect 22051 8820 22063 8823
rect 22186 8820 22192 8832
rect 22051 8792 22192 8820
rect 22051 8789 22063 8792
rect 22005 8783 22063 8789
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 25406 8780 25412 8832
rect 25464 8780 25470 8832
rect 25516 8820 25544 8860
rect 26878 8820 26884 8832
rect 25516 8792 26884 8820
rect 26878 8780 26884 8792
rect 26936 8780 26942 8832
rect 28258 8780 28264 8832
rect 28316 8780 28322 8832
rect 28902 8780 28908 8832
rect 28960 8820 28966 8832
rect 29362 8820 29368 8832
rect 28960 8792 29368 8820
rect 28960 8780 28966 8792
rect 29362 8780 29368 8792
rect 29420 8780 29426 8832
rect 30006 8780 30012 8832
rect 30064 8820 30070 8832
rect 30466 8820 30472 8832
rect 30064 8792 30472 8820
rect 30064 8780 30070 8792
rect 30466 8780 30472 8792
rect 30524 8780 30530 8832
rect 552 8730 30912 8752
rect 552 8678 4193 8730
rect 4245 8678 4257 8730
rect 4309 8678 4321 8730
rect 4373 8678 4385 8730
rect 4437 8678 4449 8730
rect 4501 8678 11783 8730
rect 11835 8678 11847 8730
rect 11899 8678 11911 8730
rect 11963 8678 11975 8730
rect 12027 8678 12039 8730
rect 12091 8678 19373 8730
rect 19425 8678 19437 8730
rect 19489 8678 19501 8730
rect 19553 8678 19565 8730
rect 19617 8678 19629 8730
rect 19681 8678 26963 8730
rect 27015 8678 27027 8730
rect 27079 8678 27091 8730
rect 27143 8678 27155 8730
rect 27207 8678 27219 8730
rect 27271 8678 30912 8730
rect 552 8656 30912 8678
rect 934 8576 940 8628
rect 992 8616 998 8628
rect 992 8588 2452 8616
rect 992 8576 998 8588
rect 2424 8560 2452 8588
rect 2774 8576 2780 8628
rect 2832 8576 2838 8628
rect 5460 8588 7052 8616
rect 2406 8508 2412 8560
rect 2464 8548 2470 8560
rect 3234 8548 3240 8560
rect 2464 8520 3240 8548
rect 2464 8508 2470 8520
rect 3234 8508 3240 8520
rect 3292 8508 3298 8560
rect 4706 8508 4712 8560
rect 4764 8548 4770 8560
rect 5077 8551 5135 8557
rect 5077 8548 5089 8551
rect 4764 8520 5089 8548
rect 4764 8508 4770 8520
rect 5077 8517 5089 8520
rect 5123 8517 5135 8551
rect 5077 8511 5135 8517
rect 1443 8483 1501 8489
rect 1443 8449 1455 8483
rect 1489 8480 1501 8483
rect 1489 8452 2728 8480
rect 1489 8449 1501 8452
rect 1443 8443 1501 8449
rect 750 8372 756 8424
rect 808 8412 814 8424
rect 937 8415 995 8421
rect 937 8412 949 8415
rect 808 8384 949 8412
rect 808 8372 814 8384
rect 937 8381 949 8384
rect 983 8381 995 8415
rect 937 8375 995 8381
rect 1264 8415 1322 8421
rect 1264 8381 1276 8415
rect 1310 8412 1322 8415
rect 1578 8412 1584 8424
rect 1310 8384 1584 8412
rect 1310 8381 1322 8384
rect 1264 8375 1322 8381
rect 1578 8372 1584 8384
rect 1636 8372 1642 8424
rect 1670 8372 1676 8424
rect 1728 8372 1734 8424
rect 2700 8356 2728 8452
rect 2958 8440 2964 8492
rect 3016 8440 3022 8492
rect 3050 8440 3056 8492
rect 3108 8480 3114 8492
rect 3700 8483 3758 8489
rect 3700 8480 3712 8483
rect 3108 8452 3712 8480
rect 3108 8440 3114 8452
rect 3700 8449 3712 8452
rect 3746 8449 3758 8483
rect 3700 8443 3758 8449
rect 2682 8304 2688 8356
rect 2740 8304 2746 8356
rect 2976 8344 3004 8440
rect 3234 8372 3240 8424
rect 3292 8372 3298 8424
rect 3602 8421 3608 8424
rect 3564 8415 3608 8421
rect 3564 8412 3576 8415
rect 3344 8384 3576 8412
rect 3344 8344 3372 8384
rect 3564 8381 3576 8384
rect 3564 8375 3608 8381
rect 3602 8372 3608 8375
rect 3660 8372 3666 8424
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 5460 8412 5488 8588
rect 7024 8548 7052 8588
rect 7098 8576 7104 8628
rect 7156 8616 7162 8628
rect 7377 8619 7435 8625
rect 7377 8616 7389 8619
rect 7156 8588 7389 8616
rect 7156 8576 7162 8588
rect 7377 8585 7389 8588
rect 7423 8585 7435 8619
rect 8021 8619 8079 8625
rect 7377 8579 7435 8585
rect 7668 8588 7972 8616
rect 7668 8548 7696 8588
rect 7024 8520 7696 8548
rect 7745 8551 7803 8557
rect 7745 8517 7757 8551
rect 7791 8517 7803 8551
rect 7745 8511 7803 8517
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 5902 8440 5908 8492
rect 5960 8480 5966 8492
rect 6000 8483 6058 8489
rect 6000 8480 6012 8483
rect 5960 8452 6012 8480
rect 5960 8440 5966 8452
rect 6000 8449 6012 8452
rect 6046 8449 6058 8483
rect 6000 8443 6058 8449
rect 6730 8440 6736 8492
rect 6788 8480 6794 8492
rect 7760 8480 7788 8511
rect 6788 8452 7788 8480
rect 7944 8480 7972 8588
rect 8021 8585 8033 8619
rect 8067 8616 8079 8619
rect 8294 8616 8300 8628
rect 8067 8588 8300 8616
rect 8067 8585 8079 8588
rect 8021 8579 8079 8585
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 8386 8576 8392 8628
rect 8444 8576 8450 8628
rect 8478 8576 8484 8628
rect 8536 8616 8542 8628
rect 9122 8616 9128 8628
rect 8536 8588 9128 8616
rect 8536 8576 8542 8588
rect 9122 8576 9128 8588
rect 9180 8616 9186 8628
rect 9180 8588 11106 8616
rect 9180 8576 9186 8588
rect 8754 8548 8760 8560
rect 8220 8520 8760 8548
rect 7944 8452 8156 8480
rect 6788 8440 6794 8452
rect 4019 8384 5488 8412
rect 5828 8412 5856 8440
rect 6273 8415 6331 8421
rect 6273 8412 6285 8415
rect 5828 8384 6285 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 6273 8381 6285 8384
rect 6319 8381 6331 8415
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 6273 8375 6331 8381
rect 7852 8384 7941 8412
rect 2976 8316 3372 8344
rect 7852 8288 7880 8384
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 7929 8375 7987 8381
rect 5994 8236 6000 8288
rect 6052 8285 6058 8288
rect 6052 8239 6061 8285
rect 6052 8236 6058 8239
rect 7834 8236 7840 8288
rect 7892 8236 7898 8288
rect 8128 8276 8156 8452
rect 8220 8421 8248 8520
rect 8754 8508 8760 8520
rect 8812 8548 8818 8560
rect 9306 8548 9312 8560
rect 8812 8520 9312 8548
rect 8812 8508 8818 8520
rect 9306 8508 9312 8520
rect 9364 8508 9370 8560
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 8536 8452 8616 8480
rect 8536 8440 8542 8452
rect 8588 8421 8616 8452
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 8720 8452 9076 8480
rect 8720 8440 8726 8452
rect 9048 8421 9076 8452
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9956 8483 10014 8489
rect 9956 8480 9968 8483
rect 9180 8452 9968 8480
rect 9180 8440 9186 8452
rect 9956 8449 9968 8452
rect 10002 8449 10014 8483
rect 9956 8443 10014 8449
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10962 8480 10968 8492
rect 10275 8452 10968 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10962 8440 10968 8452
rect 11020 8440 11026 8492
rect 11078 8480 11106 8588
rect 11514 8576 11520 8628
rect 11572 8576 11578 8628
rect 12069 8619 12127 8625
rect 12069 8585 12081 8619
rect 12115 8616 12127 8619
rect 13357 8619 13415 8625
rect 12115 8588 13216 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 11146 8508 11152 8560
rect 11204 8548 11210 8560
rect 12084 8548 12112 8579
rect 11204 8520 12112 8548
rect 11204 8508 11210 8520
rect 12526 8508 12532 8560
rect 12584 8548 12590 8560
rect 12805 8551 12863 8557
rect 12805 8548 12817 8551
rect 12584 8520 12817 8548
rect 12584 8508 12590 8520
rect 12805 8517 12817 8520
rect 12851 8517 12863 8551
rect 12805 8511 12863 8517
rect 13078 8508 13084 8560
rect 13136 8508 13142 8560
rect 13188 8548 13216 8588
rect 13357 8585 13369 8619
rect 13403 8616 13415 8619
rect 16022 8616 16028 8628
rect 13403 8588 15148 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 15120 8560 15148 8588
rect 15488 8588 16028 8616
rect 13188 8520 13584 8548
rect 13556 8492 13584 8520
rect 15102 8508 15108 8560
rect 15160 8508 15166 8560
rect 15194 8508 15200 8560
rect 15252 8548 15258 8560
rect 15381 8551 15439 8557
rect 15381 8548 15393 8551
rect 15252 8520 15393 8548
rect 15252 8508 15258 8520
rect 15381 8517 15393 8520
rect 15427 8517 15439 8551
rect 15381 8511 15439 8517
rect 11078 8452 13216 8480
rect 8205 8415 8263 8421
rect 8205 8381 8217 8415
rect 8251 8381 8263 8415
rect 8205 8375 8263 8381
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 9033 8415 9091 8421
rect 9033 8381 9045 8415
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 9214 8372 9220 8424
rect 9272 8412 9278 8424
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 9272 8384 9321 8412
rect 9272 8372 9278 8384
rect 9309 8381 9321 8384
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 9490 8372 9496 8424
rect 9548 8372 9554 8424
rect 9582 8372 9588 8424
rect 9640 8412 9646 8424
rect 9820 8415 9878 8421
rect 9820 8412 9832 8415
rect 9640 8384 9832 8412
rect 9640 8372 9646 8384
rect 9820 8381 9832 8384
rect 9866 8381 9878 8415
rect 9820 8375 9878 8381
rect 11330 8372 11336 8424
rect 11388 8372 11394 8424
rect 11698 8372 11704 8424
rect 11756 8412 11762 8424
rect 12636 8421 12664 8452
rect 13188 8421 13216 8452
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 13906 8489 13912 8492
rect 13868 8483 13912 8489
rect 13868 8449 13880 8483
rect 13868 8443 13912 8449
rect 13906 8440 13912 8443
rect 13964 8440 13970 8492
rect 14047 8483 14105 8489
rect 14047 8449 14059 8483
rect 14093 8480 14105 8483
rect 15488 8480 15516 8588
rect 16022 8576 16028 8588
rect 16080 8576 16086 8628
rect 16666 8576 16672 8628
rect 16724 8616 16730 8628
rect 16724 8588 17540 8616
rect 16724 8576 16730 8588
rect 15562 8508 15568 8560
rect 15620 8508 15626 8560
rect 17512 8548 17540 8588
rect 17586 8576 17592 8628
rect 17644 8576 17650 8628
rect 18598 8576 18604 8628
rect 18656 8616 18662 8628
rect 18656 8588 20116 8616
rect 18656 8576 18662 8588
rect 17954 8548 17960 8560
rect 17512 8520 17960 8548
rect 17954 8508 17960 8520
rect 18012 8508 18018 8560
rect 14093 8452 15516 8480
rect 15580 8480 15608 8508
rect 16212 8483 16270 8489
rect 16212 8480 16224 8483
rect 15580 8452 16224 8480
rect 14093 8449 14105 8452
rect 14047 8443 14105 8449
rect 16212 8449 16224 8452
rect 16258 8449 16270 8483
rect 16212 8443 16270 8449
rect 17126 8440 17132 8492
rect 17184 8480 17190 8492
rect 18690 8480 18696 8492
rect 17184 8452 18696 8480
rect 17184 8440 17190 8452
rect 12345 8415 12403 8421
rect 12345 8412 12357 8415
rect 11756 8384 12357 8412
rect 11756 8372 11762 8384
rect 12345 8381 12357 8384
rect 12391 8381 12403 8415
rect 12345 8375 12403 8381
rect 12621 8415 12679 8421
rect 12621 8381 12633 8415
rect 12667 8381 12679 8415
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12621 8375 12679 8381
rect 12820 8384 12909 8412
rect 11348 8344 11376 8372
rect 11793 8347 11851 8353
rect 11793 8344 11805 8347
rect 8772 8316 9260 8344
rect 11348 8316 11805 8344
rect 8772 8276 8800 8316
rect 8128 8248 8800 8276
rect 8849 8279 8907 8285
rect 8849 8245 8861 8279
rect 8895 8276 8907 8279
rect 9030 8276 9036 8288
rect 8895 8248 9036 8276
rect 8895 8245 8907 8248
rect 8849 8239 8907 8245
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 9122 8236 9128 8288
rect 9180 8236 9186 8288
rect 9232 8276 9260 8316
rect 11793 8313 11805 8316
rect 11839 8313 11851 8347
rect 11793 8307 11851 8313
rect 11606 8276 11612 8288
rect 9232 8248 11612 8276
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 12066 8236 12072 8288
rect 12124 8276 12130 8288
rect 12437 8279 12495 8285
rect 12437 8276 12449 8279
rect 12124 8248 12449 8276
rect 12124 8236 12130 8248
rect 12437 8245 12449 8248
rect 12483 8245 12495 8279
rect 12820 8276 12848 8384
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 13173 8415 13231 8421
rect 13173 8381 13185 8415
rect 13219 8412 13231 8415
rect 14182 8412 14188 8424
rect 13219 8384 14188 8412
rect 13219 8381 13231 8384
rect 13173 8375 13231 8381
rect 14182 8372 14188 8384
rect 14240 8372 14246 8424
rect 14277 8415 14335 8421
rect 14277 8381 14289 8415
rect 14323 8412 14335 8415
rect 15654 8412 15660 8424
rect 14323 8384 15660 8412
rect 14323 8381 14335 8384
rect 14277 8375 14335 8381
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 15749 8415 15807 8421
rect 15749 8381 15761 8415
rect 15795 8381 15807 8415
rect 15749 8375 15807 8381
rect 16485 8415 16543 8421
rect 16485 8381 16497 8415
rect 16531 8412 16543 8415
rect 17586 8412 17592 8424
rect 16531 8384 17592 8412
rect 16531 8381 16543 8384
rect 16485 8375 16543 8381
rect 15764 8344 15792 8375
rect 17586 8372 17592 8384
rect 17644 8372 17650 8424
rect 18064 8421 18092 8452
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 19058 8489 19064 8492
rect 19020 8483 19064 8489
rect 19020 8449 19032 8483
rect 19020 8443 19064 8449
rect 19058 8440 19064 8443
rect 19116 8440 19122 8492
rect 19150 8440 19156 8492
rect 19208 8480 19214 8492
rect 19208 8452 19253 8480
rect 19208 8440 19214 8452
rect 19334 8440 19340 8492
rect 19392 8480 19398 8492
rect 19429 8483 19487 8489
rect 19429 8480 19441 8483
rect 19392 8452 19441 8480
rect 19392 8440 19398 8452
rect 19429 8449 19441 8452
rect 19475 8449 19487 8483
rect 20088 8480 20116 8588
rect 20714 8576 20720 8628
rect 20772 8576 20778 8628
rect 22278 8576 22284 8628
rect 22336 8616 22342 8628
rect 25590 8616 25596 8628
rect 22336 8588 25596 8616
rect 22336 8576 22342 8588
rect 25590 8576 25596 8588
rect 25648 8576 25654 8628
rect 25866 8576 25872 8628
rect 25924 8576 25930 8628
rect 26053 8619 26111 8625
rect 26053 8585 26065 8619
rect 26099 8616 26111 8619
rect 26418 8616 26424 8628
rect 26099 8588 26424 8616
rect 26099 8585 26111 8588
rect 26053 8579 26111 8585
rect 26418 8576 26424 8588
rect 26476 8576 26482 8628
rect 27798 8616 27804 8628
rect 26712 8588 27804 8616
rect 25406 8508 25412 8560
rect 25464 8508 25470 8560
rect 20714 8480 20720 8492
rect 20088 8452 20720 8480
rect 19429 8443 19487 8449
rect 20714 8440 20720 8452
rect 20772 8440 20778 8492
rect 22002 8440 22008 8492
rect 22060 8489 22066 8492
rect 22060 8483 22109 8489
rect 22060 8449 22063 8483
rect 22097 8480 22109 8483
rect 22097 8452 22153 8480
rect 22097 8449 22109 8452
rect 22060 8443 22109 8449
rect 22060 8440 22066 8443
rect 22186 8440 22192 8492
rect 22244 8480 22250 8492
rect 22281 8483 22339 8489
rect 22281 8480 22293 8483
rect 22244 8452 22293 8480
rect 22244 8440 22250 8452
rect 22281 8449 22293 8452
rect 22327 8449 22339 8483
rect 22281 8443 22339 8449
rect 23661 8483 23719 8489
rect 23661 8449 23673 8483
rect 23707 8480 23719 8483
rect 24308 8483 24366 8489
rect 24308 8480 24320 8483
rect 23707 8452 24320 8480
rect 23707 8449 23719 8452
rect 23661 8443 23719 8449
rect 24308 8449 24320 8452
rect 24354 8449 24366 8483
rect 24308 8443 24366 8449
rect 24581 8483 24639 8489
rect 24581 8449 24593 8483
rect 24627 8480 24639 8483
rect 25424 8480 25452 8508
rect 24627 8452 25452 8480
rect 24627 8449 24639 8452
rect 24581 8443 24639 8449
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 18414 8372 18420 8424
rect 18472 8412 18478 8424
rect 21450 8412 21456 8424
rect 18472 8384 21456 8412
rect 18472 8372 18478 8384
rect 21450 8372 21456 8384
rect 21508 8412 21514 8424
rect 21545 8415 21603 8421
rect 21545 8412 21557 8415
rect 21508 8384 21557 8412
rect 21508 8372 21514 8384
rect 21545 8381 21557 8384
rect 21591 8412 21603 8415
rect 21910 8412 21916 8424
rect 21591 8384 21916 8412
rect 21591 8381 21603 8384
rect 21545 8375 21603 8381
rect 21910 8372 21916 8384
rect 21968 8412 21974 8424
rect 22922 8412 22928 8424
rect 21968 8384 22928 8412
rect 21968 8372 21974 8384
rect 22922 8372 22928 8384
rect 22980 8372 22986 8424
rect 23750 8372 23756 8424
rect 23808 8372 23814 8424
rect 23842 8372 23848 8424
rect 23900 8372 23906 8424
rect 24172 8415 24230 8421
rect 24172 8412 24184 8415
rect 23952 8384 24184 8412
rect 14936 8316 15792 8344
rect 23768 8344 23796 8372
rect 23952 8344 23980 8384
rect 24172 8381 24184 8384
rect 24218 8381 24230 8415
rect 25608 8412 25636 8576
rect 26712 8480 26740 8588
rect 27798 8576 27804 8588
rect 27856 8576 27862 8628
rect 28534 8576 28540 8628
rect 28592 8576 28598 8628
rect 29178 8576 29184 8628
rect 29236 8616 29242 8628
rect 30285 8619 30343 8625
rect 30285 8616 30297 8619
rect 29236 8588 30297 8616
rect 29236 8576 29242 8588
rect 30285 8585 30297 8588
rect 30331 8585 30343 8619
rect 30285 8579 30343 8585
rect 28626 8508 28632 8560
rect 28684 8548 28690 8560
rect 29825 8551 29883 8557
rect 29825 8548 29837 8551
rect 28684 8520 29837 8548
rect 28684 8508 28690 8520
rect 29825 8517 29837 8520
rect 29871 8517 29883 8551
rect 29825 8511 29883 8517
rect 27024 8483 27082 8489
rect 27024 8480 27036 8483
rect 26620 8452 27036 8480
rect 26237 8415 26295 8421
rect 26237 8412 26249 8415
rect 25608 8384 26249 8412
rect 24172 8375 24230 8381
rect 26237 8381 26249 8384
rect 26283 8412 26295 8415
rect 26510 8412 26516 8424
rect 26283 8384 26516 8412
rect 26283 8381 26295 8384
rect 26237 8375 26295 8381
rect 26510 8372 26516 8384
rect 26568 8372 26574 8424
rect 23768 8316 23980 8344
rect 26620 8344 26648 8452
rect 27024 8449 27036 8452
rect 27070 8449 27082 8483
rect 27024 8443 27082 8449
rect 27203 8483 27261 8489
rect 27203 8449 27215 8483
rect 27249 8480 27261 8483
rect 28074 8480 28080 8492
rect 27249 8452 28080 8480
rect 27249 8449 27261 8452
rect 27203 8443 27261 8449
rect 28074 8440 28080 8452
rect 28132 8440 28138 8492
rect 30374 8480 30380 8492
rect 28920 8452 30380 8480
rect 26697 8415 26755 8421
rect 26697 8381 26709 8415
rect 26743 8412 26755 8415
rect 27338 8412 27344 8424
rect 26743 8384 27344 8412
rect 26743 8381 26755 8384
rect 26697 8375 26755 8381
rect 27338 8372 27344 8384
rect 27396 8372 27402 8424
rect 27433 8415 27491 8421
rect 27433 8381 27445 8415
rect 27479 8412 27491 8415
rect 28920 8412 28948 8452
rect 30374 8440 30380 8452
rect 30432 8440 30438 8492
rect 27479 8384 28948 8412
rect 29089 8415 29147 8421
rect 27479 8381 27491 8384
rect 27433 8375 27491 8381
rect 29089 8381 29101 8415
rect 29135 8381 29147 8415
rect 29089 8375 29147 8381
rect 29641 8415 29699 8421
rect 29641 8381 29653 8415
rect 29687 8381 29699 8415
rect 29641 8375 29699 8381
rect 30101 8415 30159 8421
rect 30101 8381 30113 8415
rect 30147 8412 30159 8415
rect 30190 8412 30196 8424
rect 30147 8384 30196 8412
rect 30147 8381 30159 8384
rect 30101 8375 30159 8381
rect 26786 8344 26792 8356
rect 26620 8316 26792 8344
rect 13630 8276 13636 8288
rect 12820 8248 13636 8276
rect 12437 8239 12495 8245
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 14550 8236 14556 8288
rect 14608 8276 14614 8288
rect 14936 8276 14964 8316
rect 26786 8304 26792 8316
rect 26844 8304 26850 8356
rect 28810 8304 28816 8356
rect 28868 8344 28874 8356
rect 29104 8344 29132 8375
rect 28868 8316 29132 8344
rect 29656 8344 29684 8375
rect 30190 8372 30196 8384
rect 30248 8372 30254 8424
rect 31202 8344 31208 8356
rect 29656 8316 31208 8344
rect 28868 8304 28874 8316
rect 31202 8304 31208 8316
rect 31260 8304 31266 8356
rect 14608 8248 14964 8276
rect 14608 8236 14614 8248
rect 16022 8236 16028 8288
rect 16080 8276 16086 8288
rect 16215 8279 16273 8285
rect 16215 8276 16227 8279
rect 16080 8248 16227 8276
rect 16080 8236 16086 8248
rect 16215 8245 16227 8248
rect 16261 8245 16273 8279
rect 16215 8239 16273 8245
rect 19058 8236 19064 8288
rect 19116 8276 19122 8288
rect 21634 8276 21640 8288
rect 19116 8248 21640 8276
rect 19116 8236 19122 8248
rect 21634 8236 21640 8248
rect 21692 8276 21698 8288
rect 21910 8276 21916 8288
rect 21692 8248 21916 8276
rect 21692 8236 21698 8248
rect 21910 8236 21916 8248
rect 21968 8276 21974 8288
rect 22011 8279 22069 8285
rect 22011 8276 22023 8279
rect 21968 8248 22023 8276
rect 21968 8236 21974 8248
rect 22011 8245 22023 8248
rect 22057 8245 22069 8279
rect 22011 8239 22069 8245
rect 22554 8236 22560 8288
rect 22612 8276 22618 8288
rect 25038 8276 25044 8288
rect 22612 8248 25044 8276
rect 22612 8236 22618 8248
rect 25038 8236 25044 8248
rect 25096 8236 25102 8288
rect 28074 8236 28080 8288
rect 28132 8276 28138 8288
rect 29178 8276 29184 8288
rect 28132 8248 29184 8276
rect 28132 8236 28138 8248
rect 29178 8236 29184 8248
rect 29236 8236 29242 8288
rect 552 8186 31072 8208
rect 552 8134 7988 8186
rect 8040 8134 8052 8186
rect 8104 8134 8116 8186
rect 8168 8134 8180 8186
rect 8232 8134 8244 8186
rect 8296 8134 15578 8186
rect 15630 8134 15642 8186
rect 15694 8134 15706 8186
rect 15758 8134 15770 8186
rect 15822 8134 15834 8186
rect 15886 8134 23168 8186
rect 23220 8134 23232 8186
rect 23284 8134 23296 8186
rect 23348 8134 23360 8186
rect 23412 8134 23424 8186
rect 23476 8134 30758 8186
rect 30810 8134 30822 8186
rect 30874 8134 30886 8186
rect 30938 8134 30950 8186
rect 31002 8134 31014 8186
rect 31066 8134 31072 8186
rect 552 8112 31072 8134
rect 1397 8075 1455 8081
rect 1397 8041 1409 8075
rect 1443 8072 1455 8075
rect 2222 8072 2228 8084
rect 1443 8044 2228 8072
rect 1443 8041 1455 8044
rect 1397 8035 1455 8041
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 2875 8075 2933 8081
rect 2875 8072 2887 8075
rect 2424 8044 2887 8072
rect 2038 8004 2044 8016
rect 1872 7976 2044 8004
rect 1029 7939 1087 7945
rect 1029 7905 1041 7939
rect 1075 7936 1087 7939
rect 1578 7936 1584 7948
rect 1075 7908 1584 7936
rect 1075 7905 1087 7908
rect 1029 7899 1087 7905
rect 1578 7896 1584 7908
rect 1636 7896 1642 7948
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 1762 7936 1768 7948
rect 1719 7908 1768 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 1762 7896 1768 7908
rect 1820 7896 1826 7948
rect 1486 7828 1492 7880
rect 1544 7868 1550 7880
rect 1872 7877 1900 7976
rect 2038 7964 2044 7976
rect 2096 8004 2102 8016
rect 2424 8004 2452 8044
rect 2875 8041 2887 8044
rect 2921 8041 2933 8075
rect 2875 8035 2933 8041
rect 5166 8032 5172 8084
rect 5224 8032 5230 8084
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 6638 8072 6644 8084
rect 5776 8044 6644 8072
rect 5776 8032 5782 8044
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 7650 8032 7656 8084
rect 7708 8032 7714 8084
rect 9674 8072 9680 8084
rect 8128 8044 9680 8072
rect 5810 8004 5816 8016
rect 2096 7976 2452 8004
rect 5644 7976 5816 8004
rect 2096 7964 2102 7976
rect 3145 7939 3203 7945
rect 3145 7936 3157 7939
rect 1964 7908 3157 7936
rect 1857 7871 1915 7877
rect 1857 7868 1869 7871
rect 1544 7840 1869 7868
rect 1544 7828 1550 7840
rect 1857 7837 1869 7840
rect 1903 7837 1915 7871
rect 1857 7831 1915 7837
rect 1302 7760 1308 7812
rect 1360 7800 1366 7812
rect 1964 7800 1992 7908
rect 3145 7905 3157 7908
rect 3191 7905 3203 7939
rect 3145 7899 3203 7905
rect 3234 7896 3240 7948
rect 3292 7936 3298 7948
rect 4709 7939 4767 7945
rect 4709 7936 4721 7939
rect 3292 7908 4721 7936
rect 3292 7896 3298 7908
rect 4709 7905 4721 7908
rect 4755 7905 4767 7939
rect 4709 7899 4767 7905
rect 5166 7896 5172 7948
rect 5224 7936 5230 7948
rect 5644 7945 5672 7976
rect 5810 7964 5816 7976
rect 5868 7964 5874 8016
rect 5353 7939 5411 7945
rect 5353 7936 5365 7939
rect 5224 7908 5365 7936
rect 5224 7896 5230 7908
rect 5353 7905 5365 7908
rect 5399 7905 5411 7939
rect 5353 7899 5411 7905
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7905 5687 7939
rect 6549 7939 6607 7945
rect 6549 7936 6561 7939
rect 5629 7899 5687 7905
rect 5736 7908 6561 7936
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 2915 7871 2973 7877
rect 2915 7837 2927 7871
rect 2961 7868 2973 7871
rect 5534 7868 5540 7880
rect 2961 7840 5540 7868
rect 2961 7837 2973 7840
rect 2915 7831 2973 7837
rect 1360 7772 1992 7800
rect 1360 7760 1366 7772
rect 845 7735 903 7741
rect 845 7701 857 7735
rect 891 7732 903 7735
rect 1118 7732 1124 7744
rect 891 7704 1124 7732
rect 891 7701 903 7704
rect 845 7695 903 7701
rect 1118 7692 1124 7704
rect 1176 7692 1182 7744
rect 2424 7732 2452 7831
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 4985 7803 5043 7809
rect 4985 7769 4997 7803
rect 5031 7800 5043 7803
rect 5258 7800 5264 7812
rect 5031 7772 5264 7800
rect 5031 7769 5043 7772
rect 4985 7763 5043 7769
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 5445 7803 5503 7809
rect 5445 7769 5457 7803
rect 5491 7800 5503 7803
rect 5736 7800 5764 7908
rect 6549 7905 6561 7908
rect 6595 7905 6607 7939
rect 6549 7899 6607 7905
rect 5810 7828 5816 7880
rect 5868 7828 5874 7880
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 6140 7871 6198 7877
rect 6140 7868 6152 7871
rect 6052 7840 6152 7868
rect 6052 7828 6058 7840
rect 6140 7837 6152 7840
rect 6186 7837 6198 7871
rect 6140 7831 6198 7837
rect 6319 7871 6377 7877
rect 6319 7837 6331 7871
rect 6365 7868 6377 7871
rect 8128 7868 8156 8044
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 11330 8032 11336 8084
rect 11388 8072 11394 8084
rect 13541 8075 13599 8081
rect 11388 8044 13492 8072
rect 11388 8032 11394 8044
rect 10318 7964 10324 8016
rect 10376 8004 10382 8016
rect 10376 7976 11008 8004
rect 10376 7964 10382 7976
rect 8205 7939 8263 7945
rect 8205 7905 8217 7939
rect 8251 7905 8263 7939
rect 8205 7899 8263 7905
rect 8297 7939 8355 7945
rect 8297 7905 8309 7939
rect 8343 7936 8355 7939
rect 8386 7936 8392 7948
rect 8343 7908 8392 7936
rect 8343 7905 8355 7908
rect 8297 7899 8355 7905
rect 6365 7840 8156 7868
rect 6365 7837 6377 7840
rect 6319 7831 6377 7837
rect 5491 7772 5764 7800
rect 5491 7769 5503 7772
rect 5445 7763 5503 7769
rect 7834 7760 7840 7812
rect 7892 7800 7898 7812
rect 8220 7800 8248 7899
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 9033 7939 9091 7945
rect 9033 7905 9045 7939
rect 9079 7936 9091 7939
rect 9122 7936 9128 7948
rect 9079 7908 9128 7936
rect 9079 7905 9091 7908
rect 9033 7899 9091 7905
rect 9122 7896 9128 7908
rect 9180 7896 9186 7948
rect 9306 7896 9312 7948
rect 9364 7936 9370 7948
rect 10980 7945 11008 7976
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 9364 7908 10517 7936
rect 9364 7896 9370 7908
rect 10505 7905 10517 7908
rect 10551 7905 10563 7939
rect 10505 7899 10563 7905
rect 10965 7939 11023 7945
rect 10965 7905 10977 7939
rect 11011 7905 11023 7939
rect 10965 7899 11023 7905
rect 8570 7828 8576 7880
rect 8628 7877 8634 7880
rect 8628 7871 8682 7877
rect 8628 7837 8636 7871
rect 8670 7837 8682 7871
rect 8628 7831 8682 7837
rect 8803 7871 8861 7877
rect 8803 7837 8815 7871
rect 8849 7868 8861 7871
rect 10594 7868 10600 7880
rect 8849 7840 10600 7868
rect 8849 7837 8861 7840
rect 8803 7831 8861 7837
rect 8628 7828 8634 7831
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 10980 7868 11008 7899
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 11296 7908 12081 7936
rect 11296 7896 11302 7908
rect 12069 7905 12081 7908
rect 12115 7905 12127 7939
rect 13464 7936 13492 8044
rect 13541 8041 13553 8075
rect 13587 8041 13599 8075
rect 13541 8035 13599 8041
rect 14283 8075 14341 8081
rect 14283 8041 14295 8075
rect 14329 8072 14341 8075
rect 14826 8072 14832 8084
rect 14329 8044 14832 8072
rect 14329 8041 14341 8044
rect 14283 8035 14341 8041
rect 13556 8004 13584 8035
rect 14826 8032 14832 8044
rect 14884 8072 14890 8084
rect 16022 8072 16028 8084
rect 14884 8044 16028 8072
rect 14884 8032 14890 8044
rect 16022 8032 16028 8044
rect 16080 8032 16086 8084
rect 16666 8032 16672 8084
rect 16724 8072 16730 8084
rect 17037 8075 17095 8081
rect 17037 8072 17049 8075
rect 16724 8044 17049 8072
rect 16724 8032 16730 8044
rect 17037 8041 17049 8044
rect 17083 8072 17095 8075
rect 17083 8044 17356 8072
rect 17083 8041 17095 8044
rect 17037 8035 17095 8041
rect 13556 7976 13952 8004
rect 13464 7908 13676 7936
rect 12069 7899 12127 7905
rect 11146 7868 11152 7880
rect 10980 7840 11152 7868
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 11330 7828 11336 7880
rect 11388 7828 11394 7880
rect 11698 7877 11704 7880
rect 11660 7871 11704 7877
rect 11660 7837 11672 7871
rect 11660 7831 11704 7837
rect 11698 7828 11704 7831
rect 11756 7828 11762 7880
rect 11790 7828 11796 7880
rect 11848 7877 11854 7880
rect 11848 7871 11887 7877
rect 11875 7837 11887 7871
rect 13648 7868 13676 7908
rect 13722 7896 13728 7948
rect 13780 7896 13786 7948
rect 13924 7936 13952 7976
rect 16206 7964 16212 8016
rect 16264 7964 16270 8016
rect 16298 7964 16304 8016
rect 16356 8004 16362 8016
rect 17328 8004 17356 8044
rect 17586 8032 17592 8084
rect 17644 8032 17650 8084
rect 18515 8075 18573 8081
rect 18515 8041 18527 8075
rect 18561 8072 18573 8075
rect 19058 8072 19064 8084
rect 18561 8044 19064 8072
rect 18561 8041 18573 8044
rect 18515 8035 18573 8041
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 19886 8032 19892 8084
rect 19944 8032 19950 8084
rect 21910 8032 21916 8084
rect 21968 8072 21974 8084
rect 21968 8044 22968 8072
rect 21968 8032 21974 8044
rect 21266 8004 21272 8016
rect 16356 7976 17264 8004
rect 17328 7976 18184 8004
rect 16356 7964 16362 7976
rect 14553 7939 14611 7945
rect 14553 7936 14565 7939
rect 13924 7908 14565 7936
rect 14553 7905 14565 7908
rect 14599 7905 14611 7939
rect 14553 7899 14611 7905
rect 16390 7896 16396 7948
rect 16448 7936 16454 7948
rect 17236 7945 17264 7976
rect 18156 7948 18184 7976
rect 20462 7976 20668 8004
rect 16761 7939 16819 7945
rect 16761 7936 16773 7939
rect 16448 7908 16773 7936
rect 16448 7896 16454 7908
rect 16761 7905 16773 7908
rect 16807 7905 16819 7939
rect 16761 7899 16819 7905
rect 17221 7939 17279 7945
rect 17221 7905 17233 7939
rect 17267 7905 17279 7939
rect 17221 7899 17279 7905
rect 17773 7939 17831 7945
rect 17773 7905 17785 7939
rect 17819 7905 17831 7939
rect 17773 7899 17831 7905
rect 13817 7871 13875 7877
rect 13817 7868 13829 7871
rect 13648 7840 13829 7868
rect 11848 7831 11887 7837
rect 13817 7837 13829 7840
rect 13863 7837 13875 7871
rect 13817 7831 13875 7837
rect 14323 7871 14381 7877
rect 14323 7837 14335 7871
rect 14369 7868 14381 7871
rect 15378 7868 15384 7880
rect 14369 7840 15384 7868
rect 14369 7837 14381 7840
rect 14323 7831 14381 7837
rect 11848 7828 11854 7831
rect 8294 7800 8300 7812
rect 7892 7772 8300 7800
rect 7892 7760 7898 7772
rect 8294 7760 8300 7772
rect 8352 7760 8358 7812
rect 13832 7744 13860 7831
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 17405 7803 17463 7809
rect 17405 7800 17417 7803
rect 15212 7772 17417 7800
rect 3234 7732 3240 7744
rect 2424 7704 3240 7732
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 4249 7735 4307 7741
rect 4249 7732 4261 7735
rect 4120 7704 4261 7732
rect 4120 7692 4126 7704
rect 4249 7701 4261 7704
rect 4295 7701 4307 7735
rect 4249 7695 4307 7701
rect 5994 7692 6000 7744
rect 6052 7732 6058 7744
rect 7558 7732 7564 7744
rect 6052 7704 7564 7732
rect 6052 7692 6058 7704
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 8938 7732 8944 7744
rect 8067 7704 8944 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 8938 7692 8944 7704
rect 8996 7692 9002 7744
rect 10318 7692 10324 7744
rect 10376 7692 10382 7744
rect 10686 7692 10692 7744
rect 10744 7692 10750 7744
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 11149 7735 11207 7741
rect 11149 7732 11161 7735
rect 10836 7704 11161 7732
rect 10836 7692 10842 7704
rect 11149 7701 11161 7704
rect 11195 7701 11207 7735
rect 11149 7695 11207 7701
rect 13170 7692 13176 7744
rect 13228 7692 13234 7744
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 14550 7732 14556 7744
rect 13872 7704 14556 7732
rect 13872 7692 13878 7704
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 15212 7732 15240 7772
rect 17405 7769 17417 7772
rect 17451 7800 17463 7803
rect 17788 7800 17816 7899
rect 18138 7896 18144 7948
rect 18196 7896 18202 7948
rect 20462 7936 20490 7976
rect 20640 7948 20668 7976
rect 21100 7976 21272 8004
rect 18708 7920 20490 7936
rect 18570 7908 20490 7920
rect 18570 7895 18736 7908
rect 20530 7896 20536 7948
rect 20588 7896 20594 7948
rect 20622 7896 20628 7948
rect 20680 7896 20686 7948
rect 21100 7945 21128 7976
rect 21266 7964 21272 7976
rect 21324 7964 21330 8016
rect 21085 7939 21143 7945
rect 21085 7905 21097 7939
rect 21131 7905 21143 7939
rect 22005 7939 22063 7945
rect 22005 7936 22017 7939
rect 21085 7899 21143 7905
rect 21192 7908 22017 7936
rect 18545 7892 18736 7895
rect 18545 7889 18603 7892
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7868 18107 7871
rect 18414 7868 18420 7880
rect 18095 7840 18420 7868
rect 18095 7837 18107 7840
rect 18049 7831 18107 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 18545 7855 18557 7889
rect 18591 7855 18603 7889
rect 18545 7849 18603 7855
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7868 18843 7871
rect 18874 7868 18880 7880
rect 18831 7840 18880 7868
rect 18831 7837 18843 7840
rect 18785 7831 18843 7837
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 17451 7772 17816 7800
rect 20349 7803 20407 7809
rect 17451 7769 17463 7772
rect 17405 7763 17463 7769
rect 20349 7769 20361 7803
rect 20395 7800 20407 7803
rect 21192 7800 21220 7908
rect 22005 7905 22017 7908
rect 22051 7905 22063 7939
rect 22940 7936 22968 8044
rect 23014 8032 23020 8084
rect 23072 8072 23078 8084
rect 23109 8075 23167 8081
rect 23109 8072 23121 8075
rect 23072 8044 23121 8072
rect 23072 8032 23078 8044
rect 23109 8041 23121 8044
rect 23155 8041 23167 8075
rect 23109 8035 23167 8041
rect 25314 8032 25320 8084
rect 25372 8032 25378 8084
rect 27798 8032 27804 8084
rect 27856 8072 27862 8084
rect 28175 8075 28233 8081
rect 28175 8072 28187 8075
rect 27856 8044 28187 8072
rect 27856 8032 27862 8044
rect 28175 8041 28187 8044
rect 28221 8041 28233 8075
rect 28175 8035 28233 8041
rect 28350 8032 28356 8084
rect 28408 8072 28414 8084
rect 29549 8075 29607 8081
rect 29549 8072 29561 8075
rect 28408 8044 29561 8072
rect 28408 8032 28414 8044
rect 29549 8041 29561 8044
rect 29595 8041 29607 8075
rect 29549 8035 29607 8041
rect 25038 7964 25044 8016
rect 25096 7964 25102 8016
rect 29362 7964 29368 8016
rect 29420 8004 29426 8016
rect 29420 7976 30604 8004
rect 29420 7964 29426 7976
rect 23804 7939 23862 7945
rect 23804 7936 23816 7939
rect 22940 7908 23816 7936
rect 22005 7899 22063 7905
rect 23804 7905 23816 7908
rect 23850 7905 23862 7939
rect 23804 7899 23862 7905
rect 24486 7896 24492 7948
rect 24544 7896 24550 7948
rect 25056 7936 25084 7964
rect 25685 7939 25743 7945
rect 25685 7936 25697 7939
rect 25056 7908 25697 7936
rect 25685 7905 25697 7908
rect 25731 7936 25743 7939
rect 26418 7936 26424 7948
rect 25731 7908 26424 7936
rect 25731 7905 25743 7908
rect 25685 7899 25743 7905
rect 26418 7896 26424 7908
rect 26476 7936 26482 7948
rect 27522 7936 27528 7948
rect 26476 7908 27528 7936
rect 26476 7896 26482 7908
rect 27522 7896 27528 7908
rect 27580 7896 27586 7948
rect 27617 7939 27675 7945
rect 27617 7905 27629 7939
rect 27663 7936 27675 7939
rect 28074 7936 28080 7948
rect 27663 7908 28080 7936
rect 27663 7905 27675 7908
rect 27617 7899 27675 7905
rect 28074 7896 28080 7908
rect 28132 7896 28138 7948
rect 28442 7896 28448 7948
rect 28500 7896 28506 7948
rect 29546 7896 29552 7948
rect 29604 7936 29610 7948
rect 29914 7936 29920 7948
rect 29604 7908 29920 7936
rect 29604 7896 29610 7908
rect 29914 7896 29920 7908
rect 29972 7936 29978 7948
rect 30576 7945 30604 7976
rect 30285 7939 30343 7945
rect 30285 7936 30297 7939
rect 29972 7908 30297 7936
rect 29972 7896 29978 7908
rect 30285 7905 30297 7908
rect 30331 7905 30343 7939
rect 30285 7899 30343 7905
rect 30561 7939 30619 7945
rect 30561 7905 30573 7939
rect 30607 7905 30619 7939
rect 30561 7899 30619 7905
rect 21269 7871 21327 7877
rect 21269 7837 21281 7871
rect 21315 7868 21327 7871
rect 21450 7868 21456 7880
rect 21315 7840 21456 7868
rect 21315 7837 21327 7840
rect 21269 7831 21327 7837
rect 21450 7828 21456 7840
rect 21508 7828 21514 7880
rect 21634 7877 21640 7880
rect 21596 7871 21640 7877
rect 21596 7837 21608 7871
rect 21596 7831 21640 7837
rect 21634 7828 21640 7831
rect 21692 7828 21698 7880
rect 21775 7871 21833 7877
rect 21775 7837 21787 7871
rect 21821 7868 21833 7871
rect 21821 7840 22876 7868
rect 21821 7837 21833 7840
rect 21775 7831 21833 7837
rect 20395 7772 21220 7800
rect 20395 7769 20407 7772
rect 20349 7763 20407 7769
rect 14792 7704 15240 7732
rect 14792 7692 14798 7704
rect 15654 7692 15660 7744
rect 15712 7692 15718 7744
rect 15746 7692 15752 7744
rect 15804 7732 15810 7744
rect 16301 7735 16359 7741
rect 16301 7732 16313 7735
rect 15804 7704 16313 7732
rect 15804 7692 15810 7704
rect 16301 7701 16313 7704
rect 16347 7732 16359 7735
rect 16758 7732 16764 7744
rect 16347 7704 16764 7732
rect 16347 7701 16359 7704
rect 16301 7695 16359 7701
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 17494 7692 17500 7744
rect 17552 7732 17558 7744
rect 20438 7732 20444 7744
rect 17552 7704 20444 7732
rect 17552 7692 17558 7704
rect 20438 7692 20444 7704
rect 20496 7692 20502 7744
rect 20901 7735 20959 7741
rect 20901 7701 20913 7735
rect 20947 7732 20959 7735
rect 22186 7732 22192 7744
rect 20947 7704 22192 7732
rect 20947 7701 20959 7704
rect 20901 7695 20959 7701
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 22848 7732 22876 7840
rect 22922 7828 22928 7880
rect 22980 7868 22986 7880
rect 23477 7871 23535 7877
rect 23477 7868 23489 7871
rect 22980 7840 23489 7868
rect 22980 7828 22986 7840
rect 23477 7837 23489 7840
rect 23523 7837 23535 7871
rect 23477 7831 23535 7837
rect 23658 7828 23664 7880
rect 23716 7868 23722 7880
rect 23983 7871 24041 7877
rect 23983 7868 23995 7871
rect 23716 7840 23995 7868
rect 23716 7828 23722 7840
rect 23983 7837 23995 7840
rect 24029 7837 24041 7871
rect 23983 7831 24041 7837
rect 24118 7828 24124 7880
rect 24176 7868 24182 7880
rect 24213 7871 24271 7877
rect 24213 7868 24225 7871
rect 24176 7840 24225 7868
rect 24176 7828 24182 7840
rect 24213 7837 24225 7840
rect 24259 7837 24271 7871
rect 24504 7868 24532 7896
rect 25869 7871 25927 7877
rect 25869 7868 25881 7871
rect 24504 7840 25881 7868
rect 24213 7831 24271 7837
rect 25869 7837 25881 7840
rect 25915 7868 25927 7871
rect 26602 7868 26608 7880
rect 25915 7840 26608 7868
rect 25915 7837 25927 7840
rect 25869 7831 25927 7837
rect 26602 7828 26608 7840
rect 26660 7828 26666 7880
rect 27246 7828 27252 7880
rect 27304 7868 27310 7880
rect 27706 7868 27712 7880
rect 27304 7840 27712 7868
rect 27304 7828 27310 7840
rect 27706 7828 27712 7840
rect 27764 7828 27770 7880
rect 28166 7828 28172 7880
rect 28224 7868 28230 7880
rect 28224 7840 28269 7868
rect 28224 7828 28230 7840
rect 30101 7803 30159 7809
rect 30101 7800 30113 7803
rect 29104 7772 30113 7800
rect 25222 7732 25228 7744
rect 22848 7704 25228 7732
rect 25222 7692 25228 7704
rect 25280 7692 25286 7744
rect 27430 7692 27436 7744
rect 27488 7692 27494 7744
rect 28810 7692 28816 7744
rect 28868 7732 28874 7744
rect 29104 7732 29132 7772
rect 30101 7769 30113 7772
rect 30147 7769 30159 7803
rect 30101 7763 30159 7769
rect 28868 7704 29132 7732
rect 28868 7692 28874 7704
rect 30374 7692 30380 7744
rect 30432 7692 30438 7744
rect 552 7642 30912 7664
rect 552 7590 4193 7642
rect 4245 7590 4257 7642
rect 4309 7590 4321 7642
rect 4373 7590 4385 7642
rect 4437 7590 4449 7642
rect 4501 7590 11783 7642
rect 11835 7590 11847 7642
rect 11899 7590 11911 7642
rect 11963 7590 11975 7642
rect 12027 7590 12039 7642
rect 12091 7590 19373 7642
rect 19425 7590 19437 7642
rect 19489 7590 19501 7642
rect 19553 7590 19565 7642
rect 19617 7590 19629 7642
rect 19681 7590 26963 7642
rect 27015 7590 27027 7642
rect 27079 7590 27091 7642
rect 27143 7590 27155 7642
rect 27207 7590 27219 7642
rect 27271 7590 30912 7642
rect 552 7568 30912 7590
rect 2746 7500 7420 7528
rect 1118 7352 1124 7404
rect 1176 7392 1182 7404
rect 1443 7395 1501 7401
rect 1176 7364 1384 7392
rect 1176 7352 1182 7364
rect 750 7284 756 7336
rect 808 7324 814 7336
rect 937 7327 995 7333
rect 937 7324 949 7327
rect 808 7296 949 7324
rect 808 7284 814 7296
rect 937 7293 949 7296
rect 983 7293 995 7327
rect 1264 7327 1322 7333
rect 1264 7324 1276 7327
rect 937 7287 995 7293
rect 1044 7296 1276 7324
rect 1044 7188 1072 7296
rect 1264 7293 1276 7296
rect 1310 7293 1322 7327
rect 1356 7324 1384 7364
rect 1443 7361 1455 7395
rect 1489 7392 1501 7395
rect 2746 7392 2774 7500
rect 7392 7469 7420 7500
rect 7650 7488 7656 7540
rect 7708 7528 7714 7540
rect 10229 7531 10287 7537
rect 10229 7528 10241 7531
rect 7708 7500 10241 7528
rect 7708 7488 7714 7500
rect 10229 7497 10241 7500
rect 10275 7497 10287 7531
rect 13170 7528 13176 7540
rect 10229 7491 10287 7497
rect 10336 7500 13176 7528
rect 7377 7463 7435 7469
rect 7377 7429 7389 7463
rect 7423 7429 7435 7463
rect 7377 7423 7435 7429
rect 7558 7420 7564 7472
rect 7616 7420 7622 7472
rect 3564 7395 3622 7401
rect 3564 7392 3576 7395
rect 1489 7364 2774 7392
rect 2884 7364 3576 7392
rect 1489 7361 1501 7364
rect 1443 7355 1501 7361
rect 1673 7327 1731 7333
rect 1673 7324 1685 7327
rect 1356 7296 1685 7324
rect 1264 7287 1322 7293
rect 1673 7293 1685 7296
rect 1719 7293 1731 7327
rect 1673 7287 1731 7293
rect 2038 7284 2044 7336
rect 2096 7324 2102 7336
rect 2884 7324 2912 7364
rect 3564 7361 3576 7364
rect 3610 7361 3622 7395
rect 3564 7355 3622 7361
rect 3743 7395 3801 7401
rect 3743 7361 3755 7395
rect 3789 7392 3801 7395
rect 3789 7364 5028 7392
rect 3789 7361 3801 7364
rect 3743 7355 3801 7361
rect 2096 7296 2912 7324
rect 2096 7284 2102 7296
rect 3234 7284 3240 7336
rect 3292 7284 3298 7336
rect 3326 7284 3332 7336
rect 3384 7324 3390 7336
rect 3973 7327 4031 7333
rect 3973 7324 3985 7327
rect 3384 7296 3985 7324
rect 3384 7284 3390 7296
rect 3973 7293 3985 7296
rect 4019 7293 4031 7327
rect 3973 7287 4031 7293
rect 3050 7216 3056 7268
rect 3108 7216 3114 7268
rect 5000 7256 5028 7364
rect 5258 7352 5264 7404
rect 5316 7392 5322 7404
rect 5442 7392 5448 7404
rect 5316 7364 5448 7392
rect 5316 7352 5322 7364
rect 5442 7352 5448 7364
rect 5500 7392 5506 7404
rect 5902 7401 5908 7404
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 5500 7364 5549 7392
rect 5500 7352 5506 7364
rect 5537 7361 5549 7364
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 5864 7395 5908 7401
rect 5864 7361 5876 7395
rect 5864 7355 5908 7361
rect 5902 7352 5908 7355
rect 5960 7352 5966 7404
rect 6043 7395 6101 7401
rect 6043 7361 6055 7395
rect 6089 7392 6101 7395
rect 6730 7392 6736 7404
rect 6089 7364 6736 7392
rect 6089 7361 6101 7364
rect 6043 7355 6101 7361
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 7576 7392 7604 7420
rect 7929 7395 7987 7401
rect 7929 7392 7941 7395
rect 7576 7364 7941 7392
rect 7929 7361 7941 7364
rect 7975 7392 7987 7395
rect 8570 7392 8576 7404
rect 7975 7364 8576 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 8570 7352 8576 7364
rect 8628 7392 8634 7404
rect 8716 7395 8774 7401
rect 8716 7392 8728 7395
rect 8628 7364 8728 7392
rect 8628 7352 8634 7364
rect 8716 7361 8728 7364
rect 8762 7361 8774 7395
rect 8716 7355 8774 7361
rect 8895 7393 8953 7399
rect 8895 7359 8907 7393
rect 8941 7390 8953 7393
rect 8941 7362 9035 7390
rect 8941 7359 8953 7362
rect 8895 7353 8953 7359
rect 5074 7284 5080 7336
rect 5132 7324 5138 7336
rect 6273 7327 6331 7333
rect 6273 7324 6285 7327
rect 5132 7296 6285 7324
rect 5132 7284 5138 7296
rect 6273 7293 6285 7296
rect 6319 7293 6331 7327
rect 6273 7287 6331 7293
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7324 7803 7327
rect 7834 7324 7840 7336
rect 7791 7296 7840 7324
rect 7791 7293 7803 7296
rect 7745 7287 7803 7293
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 8386 7284 8392 7336
rect 8444 7284 8450 7336
rect 9007 7324 9035 7362
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 10336 7324 10364 7500
rect 13170 7488 13176 7500
rect 13228 7488 13234 7540
rect 15746 7528 15752 7540
rect 14022 7500 15752 7528
rect 10965 7463 11023 7469
rect 10965 7429 10977 7463
rect 11011 7460 11023 7463
rect 11238 7460 11244 7472
rect 11011 7432 11244 7460
rect 11011 7429 11023 7432
rect 10965 7423 11023 7429
rect 11238 7420 11244 7432
rect 11296 7420 11302 7472
rect 11747 7395 11805 7401
rect 11747 7361 11759 7395
rect 11793 7392 11805 7395
rect 12618 7392 12624 7404
rect 11793 7364 12624 7392
rect 11793 7361 11805 7364
rect 11747 7355 11805 7361
rect 12618 7352 12624 7364
rect 12676 7352 12682 7404
rect 13170 7392 13176 7404
rect 12912 7364 13176 7392
rect 10873 7327 10931 7333
rect 10873 7324 10885 7327
rect 9007 7296 10364 7324
rect 10520 7296 10885 7324
rect 5000 7228 5672 7256
rect 1486 7188 1492 7200
rect 1044 7160 1492 7188
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 1762 7148 1768 7200
rect 1820 7188 1826 7200
rect 4430 7188 4436 7200
rect 1820 7160 4436 7188
rect 1820 7148 1826 7160
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 4614 7148 4620 7200
rect 4672 7188 4678 7200
rect 5077 7191 5135 7197
rect 5077 7188 5089 7191
rect 4672 7160 5089 7188
rect 4672 7148 4678 7160
rect 5077 7157 5089 7160
rect 5123 7157 5135 7191
rect 5644 7188 5672 7228
rect 10520 7200 10548 7296
rect 10873 7293 10885 7296
rect 10919 7293 10931 7327
rect 10873 7287 10931 7293
rect 10962 7284 10968 7336
rect 11020 7324 11026 7336
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 11020 7296 11161 7324
rect 11020 7284 11026 7296
rect 11149 7293 11161 7296
rect 11195 7293 11207 7327
rect 11149 7287 11207 7293
rect 11238 7284 11244 7336
rect 11296 7284 11302 7336
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11348 7296 11989 7324
rect 11348 7256 11376 7296
rect 11977 7293 11989 7296
rect 12023 7293 12035 7327
rect 11977 7287 12035 7293
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 12912 7324 12940 7364
rect 13170 7352 13176 7364
rect 13228 7392 13234 7404
rect 14022 7392 14050 7500
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 16206 7488 16212 7540
rect 16264 7488 16270 7540
rect 17770 7488 17776 7540
rect 17828 7488 17834 7540
rect 18874 7528 18880 7540
rect 18708 7500 18880 7528
rect 14093 7463 14151 7469
rect 14093 7429 14105 7463
rect 14139 7429 14151 7463
rect 18708 7460 18736 7500
rect 18874 7488 18880 7500
rect 18932 7528 18938 7540
rect 19886 7528 19892 7540
rect 18932 7500 19892 7528
rect 18932 7488 18938 7500
rect 19886 7488 19892 7500
rect 19944 7488 19950 7540
rect 20717 7531 20775 7537
rect 20717 7497 20729 7531
rect 20763 7528 20775 7531
rect 20806 7528 20812 7540
rect 20763 7500 20812 7528
rect 20763 7497 20775 7500
rect 20717 7491 20775 7497
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 21269 7531 21327 7537
rect 21269 7497 21281 7531
rect 21315 7528 21327 7531
rect 21315 7500 23152 7528
rect 21315 7497 21327 7500
rect 21269 7491 21327 7497
rect 14093 7423 14151 7429
rect 18064 7432 18736 7460
rect 23124 7460 23152 7500
rect 23566 7488 23572 7540
rect 23624 7488 23630 7540
rect 24118 7488 24124 7540
rect 24176 7488 24182 7540
rect 27522 7488 27528 7540
rect 27580 7528 27586 7540
rect 28997 7531 29055 7537
rect 28997 7528 29009 7531
rect 27580 7500 29009 7528
rect 27580 7488 27586 7500
rect 28997 7497 29009 7500
rect 29043 7497 29055 7531
rect 28997 7491 29055 7497
rect 24136 7460 24164 7488
rect 23124 7432 24164 7460
rect 25961 7463 26019 7469
rect 13228 7364 14050 7392
rect 14108 7392 14136 7423
rect 14875 7395 14933 7401
rect 14108 7364 14688 7392
rect 13228 7352 13234 7364
rect 12492 7296 12940 7324
rect 12492 7284 12498 7296
rect 12986 7284 12992 7336
rect 13044 7324 13050 7336
rect 13262 7324 13268 7336
rect 13044 7296 13268 7324
rect 13044 7284 13050 7296
rect 13262 7284 13268 7296
rect 13320 7324 13326 7336
rect 13541 7327 13599 7333
rect 13541 7324 13553 7327
rect 13320 7296 13553 7324
rect 13320 7284 13326 7296
rect 13541 7293 13553 7296
rect 13587 7293 13599 7327
rect 14022 7324 14050 7364
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 14022 7296 14289 7324
rect 13541 7287 13599 7293
rect 14277 7293 14289 7296
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 14369 7327 14427 7333
rect 14369 7293 14381 7327
rect 14415 7324 14427 7327
rect 14458 7324 14464 7336
rect 14415 7296 14464 7324
rect 14415 7293 14427 7296
rect 14369 7287 14427 7293
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 14660 7324 14688 7364
rect 14875 7361 14887 7395
rect 14921 7392 14933 7395
rect 15286 7392 15292 7404
rect 14921 7364 15292 7392
rect 14921 7361 14933 7364
rect 14875 7355 14933 7361
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 15620 7364 17448 7392
rect 15620 7352 15626 7364
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 14660 7296 15117 7324
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 16574 7284 16580 7336
rect 16632 7324 16638 7336
rect 16669 7327 16727 7333
rect 16669 7324 16681 7327
rect 16632 7296 16681 7324
rect 16632 7284 16638 7296
rect 16669 7293 16681 7296
rect 16715 7293 16727 7327
rect 16669 7287 16727 7293
rect 16758 7284 16764 7336
rect 16816 7324 16822 7336
rect 17126 7324 17132 7336
rect 16816 7296 17132 7324
rect 16816 7284 16822 7296
rect 17126 7284 17132 7296
rect 17184 7284 17190 7336
rect 17420 7333 17448 7364
rect 17405 7327 17463 7333
rect 17405 7293 17417 7327
rect 17451 7324 17463 7327
rect 17494 7324 17500 7336
rect 17451 7296 17500 7324
rect 17451 7293 17463 7296
rect 17405 7287 17463 7293
rect 17494 7284 17500 7296
rect 17552 7284 17558 7336
rect 18064 7333 18092 7432
rect 25961 7429 25973 7463
rect 26007 7429 26019 7463
rect 25961 7423 26019 7429
rect 18325 7395 18383 7401
rect 18325 7361 18337 7395
rect 18371 7392 18383 7395
rect 18506 7392 18512 7404
rect 18371 7364 18512 7392
rect 18371 7361 18383 7364
rect 18325 7355 18383 7361
rect 18506 7352 18512 7364
rect 18564 7392 18570 7404
rect 19058 7401 19064 7404
rect 19020 7395 19064 7401
rect 19020 7392 19032 7395
rect 18564 7364 19032 7392
rect 18564 7352 18570 7364
rect 19020 7361 19032 7364
rect 19020 7355 19064 7361
rect 19058 7352 19064 7355
rect 19116 7352 19122 7404
rect 19189 7395 19247 7401
rect 19189 7361 19201 7395
rect 19235 7392 19247 7395
rect 21726 7392 21732 7404
rect 19235 7364 21732 7392
rect 19235 7361 19247 7364
rect 19189 7355 19247 7361
rect 21726 7352 21732 7364
rect 21784 7352 21790 7404
rect 21910 7401 21916 7404
rect 21872 7395 21916 7401
rect 21872 7361 21884 7395
rect 21872 7355 21916 7361
rect 21910 7352 21916 7355
rect 21968 7352 21974 7404
rect 22002 7352 22008 7404
rect 22060 7352 22066 7404
rect 22186 7352 22192 7404
rect 22244 7392 22250 7404
rect 22281 7395 22339 7401
rect 22281 7392 22293 7395
rect 22244 7364 22293 7392
rect 22244 7352 22250 7364
rect 22281 7361 22293 7364
rect 22327 7361 22339 7395
rect 22281 7355 22339 7361
rect 22646 7352 22652 7404
rect 22704 7392 22710 7404
rect 24118 7392 24124 7404
rect 22704 7364 24124 7392
rect 22704 7352 22710 7364
rect 24118 7352 24124 7364
rect 24176 7352 24182 7404
rect 24394 7352 24400 7404
rect 24452 7392 24458 7404
rect 24584 7395 24642 7401
rect 24584 7392 24596 7395
rect 24452 7364 24596 7392
rect 24452 7352 24458 7364
rect 24584 7361 24596 7364
rect 24630 7361 24642 7395
rect 25976 7392 26004 7423
rect 26792 7395 26850 7401
rect 26792 7392 26804 7395
rect 24584 7355 24642 7361
rect 24780 7364 26004 7392
rect 26068 7364 26804 7392
rect 22008 7343 22020 7352
rect 22054 7343 22066 7352
rect 22008 7337 22066 7343
rect 17957 7327 18015 7333
rect 17957 7293 17969 7327
rect 18003 7293 18015 7327
rect 17957 7287 18015 7293
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 13817 7259 13875 7265
rect 13817 7256 13829 7259
rect 10704 7228 11376 7256
rect 13004 7228 13829 7256
rect 7650 7188 7656 7200
rect 5644 7160 7656 7188
rect 5077 7151 5135 7157
rect 7650 7148 7656 7160
rect 7708 7148 7714 7200
rect 10502 7148 10508 7200
rect 10560 7148 10566 7200
rect 10704 7197 10732 7228
rect 10689 7191 10747 7197
rect 10689 7157 10701 7191
rect 10735 7157 10747 7191
rect 10689 7151 10747 7157
rect 11698 7148 11704 7200
rect 11756 7197 11762 7200
rect 11756 7188 11765 7197
rect 13004 7188 13032 7228
rect 13817 7225 13829 7228
rect 13863 7225 13875 7259
rect 17972 7256 18000 7287
rect 18414 7284 18420 7336
rect 18472 7324 18478 7336
rect 18693 7327 18751 7333
rect 18693 7324 18705 7327
rect 18472 7296 18705 7324
rect 18472 7284 18478 7296
rect 18693 7293 18705 7296
rect 18739 7293 18751 7327
rect 19429 7327 19487 7333
rect 19429 7324 19441 7327
rect 18693 7287 18751 7293
rect 18800 7320 19104 7324
rect 19168 7320 19441 7324
rect 18800 7296 19441 7320
rect 18598 7256 18604 7268
rect 13817 7219 13875 7225
rect 15764 7228 17356 7256
rect 17972 7228 18604 7256
rect 11756 7160 13032 7188
rect 11756 7151 11765 7160
rect 11756 7148 11762 7151
rect 13078 7148 13084 7200
rect 13136 7148 13142 7200
rect 13832 7188 13860 7219
rect 14182 7188 14188 7200
rect 13832 7160 14188 7188
rect 14182 7148 14188 7160
rect 14240 7188 14246 7200
rect 14826 7188 14832 7200
rect 14884 7197 14890 7200
rect 14240 7160 14832 7188
rect 14240 7148 14246 7160
rect 14826 7148 14832 7160
rect 14884 7188 14893 7197
rect 14884 7160 14929 7188
rect 14884 7151 14893 7160
rect 14884 7148 14890 7151
rect 15010 7148 15016 7200
rect 15068 7188 15074 7200
rect 15764 7188 15792 7228
rect 15068 7160 15792 7188
rect 15068 7148 15074 7160
rect 16758 7148 16764 7200
rect 16816 7148 16822 7200
rect 17328 7197 17356 7228
rect 18598 7216 18604 7228
rect 18656 7216 18662 7268
rect 17313 7191 17371 7197
rect 17313 7157 17325 7191
rect 17359 7157 17371 7191
rect 17313 7151 17371 7157
rect 17586 7148 17592 7200
rect 17644 7148 17650 7200
rect 17770 7148 17776 7200
rect 17828 7188 17834 7200
rect 18800 7188 18828 7296
rect 19076 7292 19196 7296
rect 19429 7293 19441 7296
rect 19475 7293 19487 7327
rect 19429 7287 19487 7293
rect 20438 7284 20444 7336
rect 20496 7324 20502 7336
rect 20898 7324 20904 7336
rect 20496 7296 20904 7324
rect 20496 7284 20502 7296
rect 20898 7284 20904 7296
rect 20956 7284 20962 7336
rect 21453 7327 21511 7333
rect 21453 7293 21465 7327
rect 21499 7293 21511 7327
rect 21453 7287 21511 7293
rect 17828 7160 18828 7188
rect 21468 7188 21496 7287
rect 21542 7284 21548 7336
rect 21600 7284 21606 7336
rect 24780 7324 24808 7364
rect 24228 7296 24808 7324
rect 22370 7188 22376 7200
rect 21468 7160 22376 7188
rect 17828 7148 17834 7160
rect 22370 7148 22376 7160
rect 22428 7148 22434 7200
rect 22554 7148 22560 7200
rect 22612 7188 22618 7200
rect 24228 7188 24256 7296
rect 24854 7284 24860 7336
rect 24912 7284 24918 7336
rect 26068 7324 26096 7364
rect 26792 7361 26804 7364
rect 26838 7361 26850 7395
rect 26792 7355 26850 7361
rect 25608 7296 26096 7324
rect 22612 7160 24256 7188
rect 22612 7148 22618 7160
rect 24486 7148 24492 7200
rect 24544 7188 24550 7200
rect 24587 7191 24645 7197
rect 24587 7188 24599 7191
rect 24544 7160 24599 7188
rect 24544 7148 24550 7160
rect 24587 7157 24599 7160
rect 24633 7157 24645 7191
rect 24587 7151 24645 7157
rect 24762 7148 24768 7200
rect 24820 7188 24826 7200
rect 25608 7188 25636 7296
rect 26142 7284 26148 7336
rect 26200 7324 26206 7336
rect 26329 7327 26387 7333
rect 26329 7324 26341 7327
rect 26200 7296 26341 7324
rect 26200 7284 26206 7296
rect 26329 7293 26341 7296
rect 26375 7293 26387 7327
rect 27065 7327 27123 7333
rect 27065 7324 27077 7327
rect 26329 7287 26387 7293
rect 26436 7296 27077 7324
rect 25682 7216 25688 7268
rect 25740 7256 25746 7268
rect 26436 7256 26464 7296
rect 27065 7293 27077 7296
rect 27111 7293 27123 7327
rect 28721 7327 28779 7333
rect 28721 7324 28733 7327
rect 27065 7287 27123 7293
rect 28644 7296 28733 7324
rect 25740 7228 26464 7256
rect 25740 7216 25746 7228
rect 28644 7200 28672 7296
rect 28721 7293 28733 7296
rect 28767 7293 28779 7327
rect 28721 7287 28779 7293
rect 29181 7327 29239 7333
rect 29181 7293 29193 7327
rect 29227 7324 29239 7327
rect 29270 7324 29276 7336
rect 29227 7296 29276 7324
rect 29227 7293 29239 7296
rect 29181 7287 29239 7293
rect 29270 7284 29276 7296
rect 29328 7284 29334 7336
rect 29454 7284 29460 7336
rect 29512 7284 29518 7336
rect 24820 7160 25636 7188
rect 24820 7148 24826 7160
rect 26602 7148 26608 7200
rect 26660 7188 26666 7200
rect 26795 7191 26853 7197
rect 26795 7188 26807 7191
rect 26660 7160 26807 7188
rect 26660 7148 26666 7160
rect 26795 7157 26807 7160
rect 26841 7157 26853 7191
rect 26795 7151 26853 7157
rect 26970 7148 26976 7200
rect 27028 7188 27034 7200
rect 28169 7191 28227 7197
rect 28169 7188 28181 7191
rect 27028 7160 28181 7188
rect 27028 7148 27034 7160
rect 28169 7157 28181 7160
rect 28215 7157 28227 7191
rect 28169 7151 28227 7157
rect 28534 7148 28540 7200
rect 28592 7148 28598 7200
rect 28626 7148 28632 7200
rect 28684 7148 28690 7200
rect 29273 7191 29331 7197
rect 29273 7157 29285 7191
rect 29319 7188 29331 7191
rect 29730 7188 29736 7200
rect 29319 7160 29736 7188
rect 29319 7157 29331 7160
rect 29273 7151 29331 7157
rect 29730 7148 29736 7160
rect 29788 7148 29794 7200
rect 552 7098 31072 7120
rect 552 7046 7988 7098
rect 8040 7046 8052 7098
rect 8104 7046 8116 7098
rect 8168 7046 8180 7098
rect 8232 7046 8244 7098
rect 8296 7046 15578 7098
rect 15630 7046 15642 7098
rect 15694 7046 15706 7098
rect 15758 7046 15770 7098
rect 15822 7046 15834 7098
rect 15886 7046 23168 7098
rect 23220 7046 23232 7098
rect 23284 7046 23296 7098
rect 23348 7046 23360 7098
rect 23412 7046 23424 7098
rect 23476 7046 30758 7098
rect 30810 7046 30822 7098
rect 30874 7046 30886 7098
rect 30938 7046 30950 7098
rect 31002 7046 31014 7098
rect 31066 7046 31072 7098
rect 552 7024 31072 7046
rect 3234 6984 3240 6996
rect 768 6956 3240 6984
rect 768 6928 796 6956
rect 750 6876 756 6928
rect 808 6876 814 6928
rect 1121 6851 1179 6857
rect 1121 6817 1133 6851
rect 1167 6848 1179 6851
rect 1167 6820 1354 6848
rect 1167 6817 1179 6820
rect 1121 6811 1179 6817
rect 934 6604 940 6656
rect 992 6604 998 6656
rect 1210 6604 1216 6656
rect 1268 6604 1274 6656
rect 1326 6644 1354 6820
rect 1394 6808 1400 6860
rect 1452 6808 1458 6860
rect 1489 6851 1547 6857
rect 1489 6817 1501 6851
rect 1535 6817 1547 6851
rect 1596 6848 1624 6956
rect 3234 6944 3240 6956
rect 3292 6984 3298 6996
rect 3418 6984 3424 6996
rect 3292 6956 3424 6984
rect 3292 6944 3298 6956
rect 3418 6944 3424 6956
rect 3476 6944 3482 6996
rect 5074 6944 5080 6996
rect 5132 6984 5138 6996
rect 5169 6987 5227 6993
rect 5169 6984 5181 6987
rect 5132 6956 5181 6984
rect 5132 6944 5138 6956
rect 5169 6953 5181 6956
rect 5215 6953 5227 6987
rect 5169 6947 5227 6953
rect 5442 6944 5448 6996
rect 5500 6984 5506 6996
rect 5810 6984 5816 6996
rect 5500 6956 5816 6984
rect 5500 6944 5506 6956
rect 5810 6944 5816 6956
rect 5868 6984 5874 6996
rect 5868 6956 8248 6984
rect 5868 6944 5874 6956
rect 1762 6876 1768 6928
rect 1820 6876 1826 6928
rect 2038 6876 2044 6928
rect 2096 6916 2102 6928
rect 2096 6888 2176 6916
rect 2096 6876 2102 6888
rect 2148 6848 2176 6888
rect 3602 6876 3608 6928
rect 3660 6916 3666 6928
rect 3970 6916 3976 6928
rect 3660 6888 3976 6916
rect 3660 6876 3666 6888
rect 3970 6876 3976 6888
rect 4028 6916 4034 6928
rect 4525 6919 4583 6925
rect 4525 6916 4537 6919
rect 4028 6888 4537 6916
rect 4028 6876 4034 6888
rect 4525 6885 4537 6888
rect 4571 6885 4583 6919
rect 4525 6879 4583 6885
rect 4614 6876 4620 6928
rect 4672 6916 4678 6928
rect 4672 6888 5212 6916
rect 4672 6876 4678 6888
rect 2368 6851 2426 6857
rect 2368 6848 2380 6851
rect 1596 6820 1900 6848
rect 2148 6820 2380 6848
rect 1489 6811 1547 6817
rect 1412 6712 1440 6808
rect 1504 6780 1532 6811
rect 1670 6780 1676 6792
rect 1504 6752 1676 6780
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 1872 6780 1900 6820
rect 2368 6817 2380 6820
rect 2414 6817 2426 6851
rect 4249 6851 4307 6857
rect 2368 6811 2426 6817
rect 2700 6820 3372 6848
rect 2537 6801 2595 6807
rect 2537 6798 2549 6801
rect 2041 6783 2099 6789
rect 2041 6780 2053 6783
rect 1872 6752 2053 6780
rect 2041 6749 2053 6752
rect 2087 6749 2099 6783
rect 2516 6767 2549 6798
rect 2583 6780 2595 6801
rect 2700 6780 2728 6820
rect 2583 6767 2728 6780
rect 2516 6752 2728 6767
rect 2777 6783 2835 6789
rect 2041 6743 2099 6749
rect 2777 6749 2789 6783
rect 2823 6780 2835 6783
rect 3234 6780 3240 6792
rect 2823 6752 3240 6780
rect 2823 6749 2835 6752
rect 2777 6743 2835 6749
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3344 6780 3372 6820
rect 4249 6817 4261 6851
rect 4295 6848 4307 6851
rect 4338 6848 4344 6860
rect 4295 6820 4344 6848
rect 4295 6817 4307 6820
rect 4249 6811 4307 6817
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 5074 6848 5080 6860
rect 5000 6820 5080 6848
rect 3878 6780 3884 6792
rect 3344 6752 3884 6780
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 5000 6780 5028 6820
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 5184 6852 5212 6888
rect 5184 6848 5304 6852
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 5184 6824 5365 6848
rect 5276 6820 5365 6824
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 5626 6808 5632 6860
rect 5684 6808 5690 6860
rect 5828 6857 5856 6944
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6817 5871 6851
rect 5813 6811 5871 6817
rect 5902 6808 5908 6860
rect 5960 6848 5966 6860
rect 8220 6857 8248 6956
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 8671 6987 8729 6993
rect 8671 6984 8683 6987
rect 8628 6956 8683 6984
rect 8628 6944 8634 6956
rect 8671 6953 8683 6956
rect 8717 6953 8729 6987
rect 8671 6947 8729 6953
rect 11149 6987 11207 6993
rect 11149 6953 11161 6987
rect 11195 6953 11207 6987
rect 11149 6947 11207 6953
rect 11164 6916 11192 6947
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 11891 6987 11949 6993
rect 11891 6984 11903 6987
rect 11756 6956 11903 6984
rect 11756 6944 11762 6956
rect 11891 6953 11903 6956
rect 11937 6953 11949 6987
rect 11891 6947 11949 6953
rect 17770 6944 17776 6996
rect 17828 6944 17834 6996
rect 18506 6944 18512 6996
rect 18564 6993 18570 6996
rect 18564 6984 18573 6993
rect 18564 6956 18609 6984
rect 18564 6947 18573 6956
rect 18564 6944 18570 6947
rect 18690 6944 18696 6996
rect 18748 6984 18754 6996
rect 20070 6984 20076 6996
rect 18748 6956 20076 6984
rect 18748 6944 18754 6956
rect 20070 6944 20076 6956
rect 20128 6944 20134 6996
rect 21008 6956 23520 6984
rect 17126 6916 17132 6928
rect 11164 6888 11468 6916
rect 6140 6851 6198 6857
rect 6140 6848 6152 6851
rect 5960 6820 6152 6848
rect 5960 6808 5966 6820
rect 6140 6817 6152 6820
rect 6186 6817 6198 6851
rect 6140 6811 6198 6817
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6848 8263 6851
rect 8478 6848 8484 6860
rect 8251 6820 8484 6848
rect 8251 6817 8263 6820
rect 8205 6811 8263 6817
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 10597 6851 10655 6857
rect 8864 6820 10548 6848
rect 6276 6801 6334 6807
rect 5442 6780 5448 6792
rect 5000 6752 5448 6780
rect 1854 6712 1860 6724
rect 1412 6684 1860 6712
rect 1854 6672 1860 6684
rect 1912 6672 1918 6724
rect 5000 6712 5028 6752
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 6276 6767 6288 6801
rect 6322 6780 6334 6801
rect 6362 6780 6368 6792
rect 6322 6767 6368 6780
rect 6276 6761 6368 6767
rect 6291 6752 6368 6761
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 6546 6740 6552 6792
rect 6604 6740 6610 6792
rect 8711 6783 8769 6789
rect 8711 6749 8723 6783
rect 8757 6780 8769 6783
rect 8864 6780 8892 6820
rect 8757 6752 8892 6780
rect 8757 6749 8769 6752
rect 8711 6743 8769 6749
rect 8938 6740 8944 6792
rect 8996 6740 9002 6792
rect 3436 6684 5028 6712
rect 3436 6644 3464 6684
rect 1326 6616 3464 6644
rect 3878 6604 3884 6656
rect 3936 6604 3942 6656
rect 4893 6647 4951 6653
rect 4893 6613 4905 6647
rect 4939 6644 4951 6647
rect 5350 6644 5356 6656
rect 4939 6616 5356 6644
rect 4939 6613 4951 6616
rect 4893 6607 4951 6613
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 5442 6604 5448 6656
rect 5500 6604 5506 6656
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 7653 6647 7711 6653
rect 7653 6644 7665 6647
rect 5868 6616 7665 6644
rect 5868 6604 5874 6616
rect 7653 6613 7665 6616
rect 7699 6613 7711 6647
rect 7653 6607 7711 6613
rect 7742 6604 7748 6656
rect 7800 6644 7806 6656
rect 10045 6647 10103 6653
rect 10045 6644 10057 6647
rect 7800 6616 10057 6644
rect 7800 6604 7806 6616
rect 10045 6613 10057 6616
rect 10091 6613 10103 6647
rect 10045 6607 10103 6613
rect 10410 6604 10416 6656
rect 10468 6604 10474 6656
rect 10520 6644 10548 6820
rect 10597 6817 10609 6851
rect 10643 6848 10655 6851
rect 11146 6848 11152 6860
rect 10643 6820 11152 6848
rect 10643 6817 10655 6820
rect 10597 6811 10655 6817
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 11238 6808 11244 6860
rect 11296 6808 11302 6860
rect 11330 6808 11336 6860
rect 11388 6808 11394 6860
rect 11440 6848 11468 6888
rect 16316 6888 16626 6916
rect 12161 6851 12219 6857
rect 12161 6848 12173 6851
rect 11440 6820 12173 6848
rect 12161 6817 12173 6820
rect 12207 6817 12219 6851
rect 12161 6811 12219 6817
rect 13814 6808 13820 6860
rect 13872 6808 13878 6860
rect 13906 6808 13912 6860
rect 13964 6808 13970 6860
rect 14182 6857 14188 6860
rect 14144 6851 14188 6857
rect 14144 6817 14156 6851
rect 14144 6811 14188 6817
rect 14182 6808 14188 6811
rect 14240 6808 14246 6860
rect 15930 6848 15936 6860
rect 14476 6820 15936 6848
rect 11054 6644 11060 6656
rect 10520 6616 11060 6644
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11164 6644 11192 6808
rect 11256 6780 11284 6808
rect 11425 6783 11483 6789
rect 11425 6780 11437 6783
rect 11256 6752 11437 6780
rect 11425 6749 11437 6752
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 11931 6785 11989 6791
rect 11931 6751 11943 6785
rect 11977 6780 11989 6785
rect 12342 6780 12348 6792
rect 11977 6752 12348 6780
rect 11977 6751 11989 6752
rect 11931 6745 11989 6751
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 13924 6780 13952 6808
rect 12820 6752 13952 6780
rect 14323 6783 14381 6789
rect 12820 6644 12848 6752
rect 14323 6749 14335 6783
rect 14369 6780 14381 6783
rect 14476 6780 14504 6820
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 16022 6808 16028 6860
rect 16080 6848 16086 6860
rect 16316 6857 16344 6888
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 16080 6820 16313 6848
rect 16080 6808 16086 6820
rect 16301 6817 16313 6820
rect 16347 6817 16359 6851
rect 16301 6811 16359 6817
rect 16390 6808 16396 6860
rect 16448 6808 16454 6860
rect 14369 6752 14504 6780
rect 14553 6783 14611 6789
rect 14369 6749 14381 6752
rect 14323 6743 14381 6749
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 16598 6780 16626 6888
rect 16684 6888 17132 6916
rect 16684 6857 16712 6888
rect 17126 6876 17132 6888
rect 17184 6916 17190 6928
rect 21008 6916 21036 6956
rect 22094 6916 22100 6928
rect 17184 6888 17264 6916
rect 17184 6876 17190 6888
rect 17236 6857 17264 6888
rect 17880 6888 18092 6916
rect 16661 6851 16719 6857
rect 16661 6817 16673 6851
rect 16707 6817 16719 6851
rect 16661 6811 16719 6817
rect 16945 6851 17003 6857
rect 16945 6817 16957 6851
rect 16991 6817 17003 6851
rect 16945 6811 17003 6817
rect 17221 6851 17279 6857
rect 17221 6817 17233 6851
rect 17267 6817 17279 6851
rect 17586 6848 17592 6860
rect 17221 6811 17279 6817
rect 17420 6820 17592 6848
rect 16758 6780 16764 6792
rect 14599 6752 16160 6780
rect 16598 6752 16764 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 15654 6672 15660 6724
rect 15712 6672 15718 6724
rect 16132 6721 16160 6752
rect 16758 6740 16764 6752
rect 16816 6780 16822 6792
rect 16960 6780 16988 6811
rect 17310 6780 17316 6792
rect 16816 6752 17316 6780
rect 16816 6740 16822 6752
rect 17310 6740 17316 6752
rect 17368 6740 17374 6792
rect 16117 6715 16175 6721
rect 16117 6681 16129 6715
rect 16163 6681 16175 6715
rect 16117 6675 16175 6681
rect 16390 6672 16396 6724
rect 16448 6712 16454 6724
rect 17129 6715 17187 6721
rect 16448 6684 16896 6712
rect 16448 6672 16454 6684
rect 11164 6616 12848 6644
rect 13262 6604 13268 6656
rect 13320 6604 13326 6656
rect 13722 6604 13728 6656
rect 13780 6644 13786 6656
rect 16206 6644 16212 6656
rect 13780 6616 16212 6644
rect 13780 6604 13786 6616
rect 16206 6604 16212 6616
rect 16264 6604 16270 6656
rect 16577 6647 16635 6653
rect 16577 6613 16589 6647
rect 16623 6644 16635 6647
rect 16666 6644 16672 6656
rect 16623 6616 16672 6644
rect 16623 6613 16635 6616
rect 16577 6607 16635 6613
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 16868 6653 16896 6684
rect 17129 6681 17141 6715
rect 17175 6712 17187 6715
rect 17420 6712 17448 6820
rect 17586 6808 17592 6820
rect 17644 6808 17650 6860
rect 17681 6851 17739 6857
rect 17681 6817 17693 6851
rect 17727 6848 17739 6851
rect 17770 6848 17776 6860
rect 17727 6820 17776 6848
rect 17727 6817 17739 6820
rect 17681 6811 17739 6817
rect 17770 6808 17776 6820
rect 17828 6808 17834 6860
rect 17880 6780 17908 6888
rect 17957 6851 18015 6857
rect 17957 6817 17969 6851
rect 18003 6817 18015 6851
rect 18064 6848 18092 6888
rect 20364 6888 21036 6916
rect 18785 6851 18843 6857
rect 18785 6848 18797 6851
rect 18064 6820 18797 6848
rect 17957 6811 18015 6817
rect 18785 6817 18797 6820
rect 18831 6817 18843 6851
rect 19702 6848 19708 6860
rect 18785 6811 18843 6817
rect 18892 6820 19708 6848
rect 17512 6752 17908 6780
rect 17512 6721 17540 6752
rect 17175 6684 17448 6712
rect 17497 6715 17555 6721
rect 17175 6681 17187 6684
rect 17129 6675 17187 6681
rect 17497 6681 17509 6715
rect 17543 6681 17555 6715
rect 17972 6712 18000 6811
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6780 18107 6783
rect 18414 6780 18420 6792
rect 18095 6752 18420 6780
rect 18095 6749 18107 6752
rect 18049 6743 18107 6749
rect 18414 6740 18420 6752
rect 18472 6740 18478 6792
rect 18598 6791 18604 6792
rect 18555 6785 18604 6791
rect 18555 6751 18567 6785
rect 18601 6751 18604 6785
rect 18555 6745 18604 6751
rect 18598 6740 18604 6745
rect 18656 6740 18662 6792
rect 18690 6740 18696 6792
rect 18748 6780 18754 6792
rect 18892 6780 18920 6820
rect 19702 6808 19708 6820
rect 19760 6848 19766 6860
rect 20364 6848 20392 6888
rect 19760 6820 20392 6848
rect 20441 6851 20499 6857
rect 19760 6808 19766 6820
rect 20441 6817 20453 6851
rect 20487 6817 20499 6851
rect 20441 6811 20499 6817
rect 18748 6752 18920 6780
rect 18748 6740 18754 6752
rect 18966 6740 18972 6792
rect 19024 6780 19030 6792
rect 20456 6780 20484 6811
rect 20530 6808 20536 6860
rect 20588 6848 20594 6860
rect 21008 6857 21036 6888
rect 21092 6888 22100 6916
rect 20717 6851 20775 6857
rect 20717 6848 20729 6851
rect 20588 6820 20729 6848
rect 20588 6808 20594 6820
rect 20717 6817 20729 6820
rect 20763 6817 20775 6851
rect 20717 6811 20775 6817
rect 20993 6851 21051 6857
rect 20993 6817 21005 6851
rect 21039 6817 21051 6851
rect 20993 6811 21051 6817
rect 21092 6792 21120 6888
rect 22094 6876 22100 6888
rect 22152 6876 22158 6928
rect 23492 6916 23520 6956
rect 23658 6944 23664 6996
rect 23716 6984 23722 6996
rect 30006 6984 30012 6996
rect 23716 6956 30012 6984
rect 23716 6944 23722 6956
rect 30006 6944 30012 6956
rect 30064 6944 30070 6996
rect 23492 6888 23704 6916
rect 23676 6860 23704 6888
rect 24504 6888 24716 6916
rect 22922 6808 22928 6860
rect 22980 6848 22986 6860
rect 22980 6820 23152 6848
rect 22980 6808 22986 6820
rect 21082 6780 21088 6792
rect 19024 6752 21088 6780
rect 19024 6740 19030 6752
rect 21082 6740 21088 6752
rect 21140 6740 21146 6792
rect 22094 6740 22100 6792
rect 22152 6740 22158 6792
rect 22462 6789 22468 6792
rect 22424 6783 22468 6789
rect 22424 6749 22436 6783
rect 22424 6743 22468 6749
rect 22462 6740 22468 6743
rect 22520 6740 22526 6792
rect 22603 6783 22661 6789
rect 22603 6749 22615 6783
rect 22649 6780 22661 6783
rect 22738 6780 22744 6792
rect 22649 6752 22744 6780
rect 22649 6749 22661 6752
rect 22603 6743 22661 6749
rect 22738 6740 22744 6752
rect 22796 6740 22802 6792
rect 22833 6783 22891 6789
rect 22833 6749 22845 6783
rect 22879 6780 22891 6783
rect 23014 6780 23020 6792
rect 22879 6752 23020 6780
rect 22879 6749 22891 6752
rect 22833 6743 22891 6749
rect 23014 6740 23020 6752
rect 23072 6740 23078 6792
rect 23124 6780 23152 6820
rect 23658 6808 23664 6860
rect 23716 6808 23722 6860
rect 24504 6857 24532 6888
rect 24489 6851 24547 6857
rect 24489 6817 24501 6851
rect 24535 6817 24547 6851
rect 24489 6811 24547 6817
rect 24578 6808 24584 6860
rect 24636 6808 24642 6860
rect 24688 6848 24716 6888
rect 26142 6876 26148 6928
rect 26200 6916 26206 6928
rect 27249 6919 27307 6925
rect 27249 6916 27261 6919
rect 26200 6888 27261 6916
rect 26200 6876 26206 6888
rect 27249 6885 27261 6888
rect 27295 6885 27307 6919
rect 27249 6879 27307 6885
rect 27338 6876 27344 6928
rect 27396 6916 27402 6928
rect 27614 6916 27620 6928
rect 27396 6888 27620 6916
rect 27396 6876 27402 6888
rect 27614 6876 27620 6888
rect 27672 6876 27678 6928
rect 27798 6876 27804 6928
rect 27856 6876 27862 6928
rect 24688 6820 26096 6848
rect 24857 6783 24915 6789
rect 24857 6780 24869 6783
rect 23124 6752 24869 6780
rect 24857 6749 24869 6752
rect 24903 6749 24915 6783
rect 24857 6743 24915 6749
rect 24946 6740 24952 6792
rect 25004 6780 25010 6792
rect 25004 6752 26004 6780
rect 25004 6740 25010 6752
rect 17972 6684 18092 6712
rect 17497 6675 17555 6681
rect 18064 6656 18092 6684
rect 16853 6647 16911 6653
rect 16853 6613 16865 6647
rect 16899 6613 16911 6647
rect 16853 6607 16911 6613
rect 17402 6604 17408 6656
rect 17460 6604 17466 6656
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 18414 6644 18420 6656
rect 18104 6616 18420 6644
rect 18104 6604 18110 6616
rect 18414 6604 18420 6616
rect 18472 6604 18478 6656
rect 19150 6604 19156 6656
rect 19208 6644 19214 6656
rect 19889 6647 19947 6653
rect 19889 6644 19901 6647
rect 19208 6616 19901 6644
rect 19208 6604 19214 6616
rect 19889 6613 19901 6616
rect 19935 6613 19947 6647
rect 19889 6607 19947 6613
rect 20254 6604 20260 6656
rect 20312 6604 20318 6656
rect 20346 6604 20352 6656
rect 20404 6644 20410 6656
rect 20533 6647 20591 6653
rect 20533 6644 20545 6647
rect 20404 6616 20545 6644
rect 20404 6604 20410 6616
rect 20533 6613 20545 6616
rect 20579 6613 20591 6647
rect 20533 6607 20591 6613
rect 20809 6647 20867 6653
rect 20809 6613 20821 6647
rect 20855 6644 20867 6647
rect 21542 6644 21548 6656
rect 20855 6616 21548 6644
rect 20855 6613 20867 6616
rect 20809 6607 20867 6613
rect 21542 6604 21548 6616
rect 21600 6604 21606 6656
rect 22370 6604 22376 6656
rect 22428 6644 22434 6656
rect 23290 6644 23296 6656
rect 22428 6616 23296 6644
rect 22428 6604 22434 6616
rect 23290 6604 23296 6616
rect 23348 6604 23354 6656
rect 24118 6604 24124 6656
rect 24176 6604 24182 6656
rect 24305 6647 24363 6653
rect 24305 6613 24317 6647
rect 24351 6644 24363 6647
rect 24854 6644 24860 6656
rect 24351 6616 24860 6644
rect 24351 6613 24363 6616
rect 24305 6607 24363 6613
rect 24854 6604 24860 6616
rect 24912 6604 24918 6656
rect 25976 6644 26004 6752
rect 26068 6712 26096 6820
rect 26234 6808 26240 6860
rect 26292 6848 26298 6860
rect 26513 6851 26571 6857
rect 26513 6848 26525 6851
rect 26292 6820 26525 6848
rect 26292 6808 26298 6820
rect 26513 6817 26525 6820
rect 26559 6817 26571 6851
rect 26513 6811 26571 6817
rect 26694 6808 26700 6860
rect 26752 6808 26758 6860
rect 27706 6808 27712 6860
rect 27764 6808 27770 6860
rect 27816 6848 27844 6876
rect 28036 6851 28094 6857
rect 28036 6848 28048 6851
rect 27816 6820 28048 6848
rect 28036 6817 28048 6820
rect 28082 6817 28094 6851
rect 28036 6811 28094 6817
rect 28445 6851 28503 6857
rect 28445 6817 28457 6851
rect 28491 6848 28503 6851
rect 30282 6848 30288 6860
rect 28491 6820 30288 6848
rect 28491 6817 28503 6820
rect 28445 6811 28503 6817
rect 30282 6808 30288 6820
rect 30340 6808 30346 6860
rect 26145 6783 26203 6789
rect 26145 6749 26157 6783
rect 26191 6780 26203 6783
rect 26712 6780 26740 6808
rect 26191 6752 26740 6780
rect 28205 6801 28263 6807
rect 28205 6767 28217 6801
rect 28251 6792 28263 6801
rect 28251 6767 28264 6792
rect 28205 6761 28264 6767
rect 28230 6752 28264 6761
rect 26191 6749 26203 6752
rect 26145 6743 26203 6749
rect 28258 6740 28264 6752
rect 28316 6740 28322 6792
rect 26789 6715 26847 6721
rect 26789 6712 26801 6715
rect 26068 6684 26801 6712
rect 26789 6681 26801 6684
rect 26835 6712 26847 6715
rect 27338 6712 27344 6724
rect 26835 6684 27344 6712
rect 26835 6681 26847 6684
rect 26789 6675 26847 6681
rect 27338 6672 27344 6684
rect 27396 6672 27402 6724
rect 29546 6672 29552 6724
rect 29604 6672 29610 6724
rect 28902 6644 28908 6656
rect 25976 6616 28908 6644
rect 28902 6604 28908 6616
rect 28960 6604 28966 6656
rect 552 6554 30912 6576
rect 552 6502 4193 6554
rect 4245 6502 4257 6554
rect 4309 6502 4321 6554
rect 4373 6502 4385 6554
rect 4437 6502 4449 6554
rect 4501 6502 11783 6554
rect 11835 6502 11847 6554
rect 11899 6502 11911 6554
rect 11963 6502 11975 6554
rect 12027 6502 12039 6554
rect 12091 6502 19373 6554
rect 19425 6502 19437 6554
rect 19489 6502 19501 6554
rect 19553 6502 19565 6554
rect 19617 6502 19629 6554
rect 19681 6502 26963 6554
rect 27015 6502 27027 6554
rect 27079 6502 27091 6554
rect 27143 6502 27155 6554
rect 27207 6502 27219 6554
rect 27271 6502 30912 6554
rect 552 6480 30912 6502
rect 1210 6400 1216 6452
rect 1268 6440 1274 6452
rect 1268 6412 2360 6440
rect 1268 6400 1274 6412
rect 2332 6372 2360 6412
rect 2774 6400 2780 6452
rect 2832 6400 2838 6452
rect 9858 6440 9864 6452
rect 3252 6412 5304 6440
rect 3252 6372 3280 6412
rect 2332 6344 3280 6372
rect 1443 6307 1501 6313
rect 1443 6273 1455 6307
rect 1489 6304 1501 6307
rect 2130 6304 2136 6316
rect 1489 6276 2136 6304
rect 1489 6273 1501 6276
rect 1443 6267 1501 6273
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 3743 6307 3801 6313
rect 3743 6273 3755 6307
rect 3789 6304 3801 6307
rect 4062 6304 4068 6316
rect 3789 6276 4068 6304
rect 3789 6273 3801 6276
rect 3743 6267 3801 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 5276 6304 5304 6412
rect 7944 6412 9864 6440
rect 5718 6304 5724 6316
rect 5276 6276 5724 6304
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 5902 6313 5908 6316
rect 5864 6307 5908 6313
rect 5864 6273 5876 6307
rect 5864 6267 5908 6273
rect 5902 6264 5908 6267
rect 5960 6264 5966 6316
rect 6086 6313 6092 6316
rect 6043 6307 6092 6313
rect 6043 6273 6055 6307
rect 6089 6273 6092 6307
rect 6043 6267 6092 6273
rect 6086 6264 6092 6267
rect 6144 6264 6150 6316
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6304 6331 6307
rect 6454 6304 6460 6316
rect 6319 6276 6460 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 6454 6264 6460 6276
rect 6512 6264 6518 6316
rect 750 6196 756 6248
rect 808 6236 814 6248
rect 937 6239 995 6245
rect 937 6236 949 6239
rect 808 6208 949 6236
rect 808 6196 814 6208
rect 937 6205 949 6208
rect 983 6205 995 6239
rect 937 6199 995 6205
rect 1264 6239 1322 6245
rect 1264 6205 1276 6239
rect 1310 6236 1322 6239
rect 1578 6236 1584 6248
rect 1310 6208 1584 6236
rect 1310 6205 1322 6208
rect 1264 6199 1322 6205
rect 1578 6196 1584 6208
rect 1636 6196 1642 6248
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 2590 6236 2596 6248
rect 1719 6208 2596 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 2866 6196 2872 6248
rect 2924 6236 2930 6248
rect 3237 6239 3295 6245
rect 3237 6236 3249 6239
rect 2924 6208 3249 6236
rect 2924 6196 2930 6208
rect 3237 6205 3249 6208
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 3973 6239 4031 6245
rect 3973 6236 3985 6239
rect 3660 6208 3985 6236
rect 3660 6196 3666 6208
rect 3973 6205 3985 6208
rect 4019 6205 4031 6239
rect 3973 6199 4031 6205
rect 5258 6196 5264 6248
rect 5316 6236 5322 6248
rect 5537 6239 5595 6245
rect 5537 6236 5549 6239
rect 5316 6208 5549 6236
rect 5316 6196 5322 6208
rect 5537 6205 5549 6208
rect 5583 6205 5595 6239
rect 5537 6199 5595 6205
rect 7742 6128 7748 6180
rect 7800 6168 7806 6180
rect 7837 6171 7895 6177
rect 7837 6168 7849 6171
rect 7800 6140 7849 6168
rect 7800 6128 7806 6140
rect 7837 6137 7849 6140
rect 7883 6137 7895 6171
rect 7837 6131 7895 6137
rect 2130 6060 2136 6112
rect 2188 6100 2194 6112
rect 3703 6103 3761 6109
rect 3703 6100 3715 6103
rect 2188 6072 3715 6100
rect 2188 6060 2194 6072
rect 3703 6069 3715 6072
rect 3749 6100 3761 6103
rect 4246 6100 4252 6112
rect 3749 6072 4252 6100
rect 3749 6069 3761 6072
rect 3703 6063 3761 6069
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 5074 6060 5080 6112
rect 5132 6060 5138 6112
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 7377 6103 7435 6109
rect 7377 6100 7389 6103
rect 5592 6072 7389 6100
rect 5592 6060 5598 6072
rect 7377 6069 7389 6072
rect 7423 6069 7435 6103
rect 7377 6063 7435 6069
rect 7650 6060 7656 6112
rect 7708 6100 7714 6112
rect 7944 6109 7972 6412
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 10594 6400 10600 6452
rect 10652 6440 10658 6452
rect 13262 6440 13268 6452
rect 10652 6412 13268 6440
rect 10652 6400 10658 6412
rect 13262 6400 13268 6412
rect 13320 6400 13326 6452
rect 13446 6400 13452 6452
rect 13504 6400 13510 6452
rect 13817 6443 13875 6449
rect 13817 6409 13829 6443
rect 13863 6440 13875 6443
rect 14550 6440 14556 6452
rect 13863 6412 14556 6440
rect 13863 6409 13875 6412
rect 13817 6403 13875 6409
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 14642 6400 14648 6452
rect 14700 6440 14706 6452
rect 16022 6440 16028 6452
rect 14700 6412 16028 6440
rect 14700 6400 14706 6412
rect 16022 6400 16028 6412
rect 16080 6400 16086 6452
rect 16206 6400 16212 6452
rect 16264 6400 16270 6452
rect 20622 6440 20628 6452
rect 16868 6412 20628 6440
rect 13464 6372 13492 6400
rect 13188 6344 14320 6372
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 8716 6307 8774 6313
rect 8716 6304 8728 6307
rect 8628 6276 8728 6304
rect 8628 6264 8634 6276
rect 8716 6273 8728 6276
rect 8762 6273 8774 6307
rect 8716 6267 8774 6273
rect 8895 6307 8953 6313
rect 8895 6273 8907 6307
rect 8941 6304 8953 6307
rect 8941 6276 10916 6304
rect 8941 6273 8953 6276
rect 8895 6267 8953 6273
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 8478 6236 8484 6248
rect 8435 6208 8484 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 8478 6196 8484 6208
rect 8536 6196 8542 6248
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 10410 6236 10416 6248
rect 9171 6208 10416 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 10597 6239 10655 6245
rect 10597 6236 10609 6239
rect 10560 6208 10609 6236
rect 10560 6196 10566 6208
rect 10597 6205 10609 6208
rect 10643 6205 10655 6239
rect 10888 6236 10916 6276
rect 11054 6264 11060 6316
rect 11112 6304 11118 6316
rect 13078 6304 13084 6316
rect 11112 6276 11157 6304
rect 11256 6276 13084 6304
rect 11112 6264 11118 6276
rect 11256 6236 11284 6276
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 10888 6208 11284 6236
rect 10597 6199 10655 6205
rect 11330 6196 11336 6248
rect 11388 6196 11394 6248
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 12989 6239 13047 6245
rect 12989 6236 13001 6239
rect 12768 6208 13001 6236
rect 12768 6196 12774 6208
rect 12989 6205 13001 6208
rect 13035 6236 13047 6239
rect 13188 6236 13216 6344
rect 13354 6264 13360 6316
rect 13412 6304 13418 6316
rect 13412 6276 13860 6304
rect 13412 6264 13418 6276
rect 13035 6208 13216 6236
rect 13265 6239 13323 6245
rect 13035 6205 13047 6208
rect 12989 6199 13047 6205
rect 13265 6205 13277 6239
rect 13311 6236 13323 6239
rect 13372 6236 13400 6264
rect 13311 6208 13400 6236
rect 13725 6239 13783 6245
rect 13311 6205 13323 6208
rect 13265 6199 13323 6205
rect 13725 6205 13737 6239
rect 13771 6205 13783 6239
rect 13832 6236 13860 6276
rect 14292 6245 14320 6344
rect 14366 6264 14372 6316
rect 14424 6264 14430 6316
rect 14734 6264 14740 6316
rect 14792 6264 14798 6316
rect 14875 6307 14933 6313
rect 14875 6273 14887 6307
rect 14921 6304 14933 6307
rect 15194 6304 15200 6316
rect 14921 6276 15200 6304
rect 14921 6273 14933 6276
rect 14875 6267 14933 6273
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 15470 6264 15476 6316
rect 15528 6264 15534 6316
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13832 6208 14013 6236
rect 13725 6199 13783 6205
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 14277 6239 14335 6245
rect 14277 6205 14289 6239
rect 14323 6205 14335 6239
rect 14752 6236 14780 6264
rect 14277 6199 14335 6205
rect 14384 6208 14780 6236
rect 15105 6239 15163 6245
rect 13740 6168 13768 6199
rect 13906 6168 13912 6180
rect 11992 6140 13912 6168
rect 7929 6103 7987 6109
rect 7929 6100 7941 6103
rect 7708 6072 7941 6100
rect 7708 6060 7714 6072
rect 7929 6069 7941 6072
rect 7975 6069 7987 6103
rect 7929 6063 7987 6069
rect 8938 6060 8944 6112
rect 8996 6100 9002 6112
rect 10229 6103 10287 6109
rect 10229 6100 10241 6103
rect 8996 6072 10241 6100
rect 8996 6060 9002 6072
rect 10229 6069 10241 6072
rect 10275 6069 10287 6103
rect 10229 6063 10287 6069
rect 11063 6103 11121 6109
rect 11063 6069 11075 6103
rect 11109 6100 11121 6103
rect 11238 6100 11244 6112
rect 11109 6072 11244 6100
rect 11109 6069 11121 6072
rect 11063 6063 11121 6069
rect 11238 6060 11244 6072
rect 11296 6060 11302 6112
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 11992 6100 12020 6140
rect 13906 6128 13912 6140
rect 13964 6168 13970 6180
rect 14384 6168 14412 6208
rect 15105 6205 15117 6239
rect 15151 6236 15163 6239
rect 15488 6236 15516 6264
rect 16868 6245 16896 6412
rect 20622 6400 20628 6412
rect 20680 6400 20686 6452
rect 20714 6400 20720 6452
rect 20772 6400 20778 6452
rect 22738 6400 22744 6452
rect 22796 6400 22802 6452
rect 23216 6412 28580 6440
rect 17034 6332 17040 6384
rect 17092 6372 17098 6384
rect 17681 6375 17739 6381
rect 17681 6372 17693 6375
rect 17092 6344 17693 6372
rect 17092 6332 17098 6344
rect 17681 6341 17693 6344
rect 17727 6341 17739 6375
rect 17681 6335 17739 6341
rect 17770 6332 17776 6384
rect 17828 6372 17834 6384
rect 18690 6372 18696 6384
rect 17828 6344 18696 6372
rect 17828 6332 17834 6344
rect 17788 6304 17816 6332
rect 17374 6276 17816 6304
rect 15151 6208 15516 6236
rect 16853 6239 16911 6245
rect 15151 6205 15163 6208
rect 15105 6199 15163 6205
rect 16853 6205 16865 6239
rect 16899 6205 16911 6239
rect 16853 6199 16911 6205
rect 17126 6196 17132 6248
rect 17184 6196 17190 6248
rect 17374 6241 17402 6276
rect 17374 6235 17439 6241
rect 17374 6204 17393 6235
rect 17381 6201 17393 6204
rect 17427 6201 17439 6235
rect 17381 6195 17439 6201
rect 17494 6196 17500 6248
rect 17552 6196 17558 6248
rect 17954 6196 17960 6248
rect 18012 6196 18018 6248
rect 18049 6239 18107 6245
rect 18049 6205 18061 6239
rect 18095 6236 18107 6239
rect 18138 6236 18144 6248
rect 18095 6208 18144 6236
rect 18095 6205 18107 6208
rect 18049 6199 18107 6205
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 18524 6245 18552 6344
rect 18690 6332 18696 6344
rect 18748 6332 18754 6384
rect 19242 6313 19248 6316
rect 19199 6307 19248 6313
rect 19199 6273 19211 6307
rect 19245 6273 19248 6307
rect 19199 6267 19248 6273
rect 19242 6264 19248 6267
rect 19300 6264 19306 6316
rect 21364 6307 21422 6313
rect 21364 6304 21376 6307
rect 20548 6276 21376 6304
rect 20548 6248 20576 6276
rect 21364 6273 21376 6276
rect 21410 6273 21422 6307
rect 21364 6267 21422 6273
rect 18509 6239 18567 6245
rect 18509 6205 18521 6239
rect 18555 6205 18567 6239
rect 18509 6199 18567 6205
rect 18598 6196 18604 6248
rect 18656 6236 18662 6248
rect 18693 6239 18751 6245
rect 18693 6236 18705 6239
rect 18656 6208 18705 6236
rect 18656 6196 18662 6208
rect 18693 6205 18705 6208
rect 18739 6205 18751 6239
rect 19429 6239 19487 6245
rect 19429 6236 19441 6239
rect 18693 6199 18751 6205
rect 18800 6208 19441 6236
rect 18800 6168 18828 6208
rect 19429 6205 19441 6208
rect 19475 6205 19487 6239
rect 19429 6199 19487 6205
rect 20530 6196 20536 6248
rect 20588 6196 20594 6248
rect 20901 6239 20959 6245
rect 20901 6205 20913 6239
rect 20947 6236 20959 6239
rect 21174 6236 21180 6248
rect 20947 6208 21180 6236
rect 20947 6205 20959 6208
rect 20901 6199 20959 6205
rect 21174 6196 21180 6208
rect 21232 6196 21238 6248
rect 21542 6196 21548 6248
rect 21600 6236 21606 6248
rect 21637 6239 21695 6245
rect 21637 6236 21649 6239
rect 21600 6208 21649 6236
rect 21600 6196 21606 6208
rect 21637 6205 21649 6208
rect 21683 6205 21695 6239
rect 21637 6199 21695 6205
rect 21726 6196 21732 6248
rect 21784 6236 21790 6248
rect 23216 6236 23244 6412
rect 23290 6332 23296 6384
rect 23348 6332 23354 6384
rect 28552 6381 28580 6412
rect 28537 6375 28595 6381
rect 28537 6341 28549 6375
rect 28583 6341 28595 6375
rect 28537 6335 28595 6341
rect 23308 6245 23336 6332
rect 24302 6264 24308 6316
rect 24360 6304 24366 6316
rect 24492 6307 24550 6313
rect 24492 6304 24504 6307
rect 24360 6276 24504 6304
rect 24360 6264 24366 6276
rect 24492 6273 24504 6276
rect 24538 6273 24550 6307
rect 24492 6267 24550 6273
rect 24688 6276 26096 6304
rect 21784 6208 23244 6236
rect 23293 6239 23351 6245
rect 21784 6196 21790 6208
rect 23293 6205 23305 6239
rect 23339 6205 23351 6239
rect 23293 6199 23351 6205
rect 23842 6196 23848 6248
rect 23900 6236 23906 6248
rect 24029 6239 24087 6245
rect 24029 6236 24041 6239
rect 23900 6208 24041 6236
rect 23900 6196 23906 6208
rect 24029 6205 24041 6208
rect 24075 6236 24087 6239
rect 24688 6236 24716 6276
rect 24075 6208 24716 6236
rect 24765 6239 24823 6245
rect 24075 6205 24087 6208
rect 24029 6199 24087 6205
rect 24765 6205 24777 6239
rect 24811 6236 24823 6239
rect 25498 6236 25504 6248
rect 24811 6208 25504 6236
rect 24811 6205 24823 6208
rect 24765 6199 24823 6205
rect 25498 6196 25504 6208
rect 25556 6196 25562 6248
rect 13964 6140 14412 6168
rect 17788 6140 18828 6168
rect 13964 6128 13970 6140
rect 11848 6072 12020 6100
rect 11848 6060 11854 6072
rect 12434 6060 12440 6112
rect 12492 6060 12498 6112
rect 12802 6060 12808 6112
rect 12860 6060 12866 6112
rect 13078 6060 13084 6112
rect 13136 6060 13142 6112
rect 13538 6060 13544 6112
rect 13596 6060 13602 6112
rect 14093 6103 14151 6109
rect 14093 6069 14105 6103
rect 14139 6100 14151 6103
rect 14458 6100 14464 6112
rect 14139 6072 14464 6100
rect 14139 6069 14151 6072
rect 14093 6063 14151 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 14826 6060 14832 6112
rect 14884 6109 14890 6112
rect 14884 6100 14893 6109
rect 16669 6103 16727 6109
rect 14884 6072 14929 6100
rect 14884 6063 14893 6072
rect 16669 6069 16681 6103
rect 16715 6100 16727 6103
rect 16850 6100 16856 6112
rect 16715 6072 16856 6100
rect 16715 6069 16727 6072
rect 16669 6063 16727 6069
rect 14884 6060 14890 6063
rect 16850 6060 16856 6072
rect 16908 6060 16914 6112
rect 16942 6060 16948 6112
rect 17000 6060 17006 6112
rect 17218 6060 17224 6112
rect 17276 6060 17282 6112
rect 17788 6109 17816 6140
rect 17773 6103 17831 6109
rect 17773 6069 17785 6103
rect 17819 6069 17831 6103
rect 17773 6063 17831 6069
rect 18046 6060 18052 6112
rect 18104 6100 18110 6112
rect 18233 6103 18291 6109
rect 18233 6100 18245 6103
rect 18104 6072 18245 6100
rect 18104 6060 18110 6072
rect 18233 6069 18245 6072
rect 18279 6069 18291 6103
rect 18233 6063 18291 6069
rect 18325 6103 18383 6109
rect 18325 6069 18337 6103
rect 18371 6100 18383 6103
rect 18966 6100 18972 6112
rect 18371 6072 18972 6100
rect 18371 6069 18383 6072
rect 18325 6063 18383 6069
rect 18966 6060 18972 6072
rect 19024 6060 19030 6112
rect 19058 6060 19064 6112
rect 19116 6100 19122 6112
rect 19159 6103 19217 6109
rect 19159 6100 19171 6103
rect 19116 6072 19171 6100
rect 19116 6060 19122 6072
rect 19159 6069 19171 6072
rect 19205 6069 19217 6103
rect 19159 6063 19217 6069
rect 21367 6103 21425 6109
rect 21367 6069 21379 6103
rect 21413 6100 21425 6103
rect 21542 6100 21548 6112
rect 21413 6072 21548 6100
rect 21413 6069 21425 6072
rect 21367 6063 21425 6069
rect 21542 6060 21548 6072
rect 21600 6060 21606 6112
rect 22830 6060 22836 6112
rect 22888 6100 22894 6112
rect 23109 6103 23167 6109
rect 23109 6100 23121 6103
rect 22888 6072 23121 6100
rect 22888 6060 22894 6072
rect 23109 6069 23121 6072
rect 23155 6069 23167 6103
rect 23109 6063 23167 6069
rect 24394 6060 24400 6112
rect 24452 6100 24458 6112
rect 24495 6103 24553 6109
rect 24495 6100 24507 6103
rect 24452 6072 24507 6100
rect 24452 6060 24458 6072
rect 24495 6069 24507 6072
rect 24541 6100 24553 6103
rect 25774 6100 25780 6112
rect 24541 6072 25780 6100
rect 24541 6069 24553 6072
rect 24495 6063 24553 6069
rect 25774 6060 25780 6072
rect 25832 6060 25838 6112
rect 25866 6060 25872 6112
rect 25924 6060 25930 6112
rect 26068 6100 26096 6276
rect 26142 6264 26148 6316
rect 26200 6304 26206 6316
rect 26694 6304 26700 6316
rect 26200 6276 26700 6304
rect 26200 6264 26206 6276
rect 26694 6264 26700 6276
rect 26752 6264 26758 6316
rect 26878 6264 26884 6316
rect 26936 6304 26942 6316
rect 27160 6307 27218 6313
rect 27160 6304 27172 6307
rect 26936 6276 27172 6304
rect 26936 6264 26942 6276
rect 27160 6273 27172 6276
rect 27206 6273 27218 6307
rect 27160 6267 27218 6273
rect 27430 6264 27436 6316
rect 27488 6264 27494 6316
rect 26510 6196 26516 6248
rect 26568 6236 26574 6248
rect 26605 6239 26663 6245
rect 26605 6236 26617 6239
rect 26568 6208 26617 6236
rect 26568 6196 26574 6208
rect 26605 6205 26617 6208
rect 26651 6236 26663 6239
rect 26651 6208 26740 6236
rect 26651 6205 26663 6208
rect 26605 6199 26663 6205
rect 26712 6168 26740 6208
rect 27890 6196 27896 6248
rect 27948 6236 27954 6248
rect 27948 6208 29684 6236
rect 27948 6196 27954 6208
rect 26786 6168 26792 6180
rect 26712 6140 26792 6168
rect 26786 6128 26792 6140
rect 26844 6128 26850 6180
rect 29656 6112 29684 6208
rect 26326 6100 26332 6112
rect 26068 6072 26332 6100
rect 26326 6060 26332 6072
rect 26384 6060 26390 6112
rect 26418 6060 26424 6112
rect 26476 6060 26482 6112
rect 26602 6060 26608 6112
rect 26660 6100 26666 6112
rect 27163 6103 27221 6109
rect 27163 6100 27175 6103
rect 26660 6072 27175 6100
rect 26660 6060 26666 6072
rect 27163 6069 27175 6072
rect 27209 6069 27221 6103
rect 27163 6063 27221 6069
rect 29638 6060 29644 6112
rect 29696 6060 29702 6112
rect 552 6010 31072 6032
rect 552 5958 7988 6010
rect 8040 5958 8052 6010
rect 8104 5958 8116 6010
rect 8168 5958 8180 6010
rect 8232 5958 8244 6010
rect 8296 5958 15578 6010
rect 15630 5958 15642 6010
rect 15694 5958 15706 6010
rect 15758 5958 15770 6010
rect 15822 5958 15834 6010
rect 15886 5958 23168 6010
rect 23220 5958 23232 6010
rect 23284 5958 23296 6010
rect 23348 5958 23360 6010
rect 23412 5958 23424 6010
rect 23476 5958 30758 6010
rect 30810 5958 30822 6010
rect 30874 5958 30886 6010
rect 30938 5958 30950 6010
rect 31002 5958 31014 6010
rect 31066 5958 31072 6010
rect 552 5936 31072 5958
rect 937 5899 995 5905
rect 937 5865 949 5899
rect 983 5896 995 5899
rect 1026 5896 1032 5908
rect 983 5868 1032 5896
rect 983 5865 995 5868
rect 937 5859 995 5865
rect 1026 5856 1032 5868
rect 1084 5856 1090 5908
rect 1762 5856 1768 5908
rect 1820 5905 1826 5908
rect 1820 5896 1829 5905
rect 2130 5896 2136 5908
rect 1820 5868 2136 5896
rect 1820 5859 1829 5868
rect 1820 5856 1826 5859
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 3878 5896 3884 5908
rect 2746 5868 3884 5896
rect 658 5720 664 5772
rect 716 5720 722 5772
rect 1121 5763 1179 5769
rect 1121 5729 1133 5763
rect 1167 5760 1179 5763
rect 1394 5760 1400 5772
rect 1167 5732 1400 5760
rect 1167 5729 1179 5732
rect 1121 5723 1179 5729
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 2746 5760 2774 5868
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 3970 5856 3976 5908
rect 4028 5905 4034 5908
rect 4028 5896 4037 5905
rect 4028 5868 4073 5896
rect 4028 5859 4037 5868
rect 4028 5856 4034 5859
rect 5442 5856 5448 5908
rect 5500 5856 5506 5908
rect 6086 5856 6092 5908
rect 6144 5896 6150 5908
rect 6279 5899 6337 5905
rect 6279 5896 6291 5899
rect 6144 5868 6291 5896
rect 6144 5856 6150 5868
rect 6279 5865 6291 5868
rect 6325 5896 6337 5899
rect 7558 5896 7564 5908
rect 6325 5868 7564 5896
rect 6325 5865 6337 5868
rect 6279 5859 6337 5865
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 8487 5899 8545 5905
rect 8487 5865 8499 5899
rect 8533 5896 8545 5899
rect 8662 5896 8668 5908
rect 8533 5868 8668 5896
rect 8533 5865 8545 5868
rect 8487 5859 8545 5865
rect 8662 5856 8668 5868
rect 8720 5856 8726 5908
rect 10594 5856 10600 5908
rect 10652 5896 10658 5908
rect 10965 5899 11023 5905
rect 10965 5896 10977 5899
rect 10652 5868 10977 5896
rect 10652 5856 10658 5868
rect 10965 5865 10977 5868
rect 11011 5865 11023 5899
rect 12710 5896 12716 5908
rect 10965 5859 11023 5865
rect 11164 5868 12716 5896
rect 5460 5760 5488 5856
rect 11164 5769 11192 5868
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 13538 5856 13544 5908
rect 13596 5856 13602 5908
rect 20346 5856 20352 5908
rect 20404 5856 20410 5908
rect 21082 5856 21088 5908
rect 21140 5856 21146 5908
rect 21542 5856 21548 5908
rect 21600 5896 21606 5908
rect 21735 5899 21793 5905
rect 21735 5896 21747 5899
rect 21600 5868 21747 5896
rect 21600 5856 21606 5868
rect 21735 5865 21747 5868
rect 21781 5865 21793 5899
rect 21735 5859 21793 5865
rect 22462 5856 22468 5908
rect 22520 5896 22526 5908
rect 23943 5899 24001 5905
rect 23943 5896 23955 5899
rect 22520 5868 23955 5896
rect 22520 5856 22526 5868
rect 23943 5865 23955 5868
rect 23989 5865 24001 5899
rect 23943 5859 24001 5865
rect 25682 5856 25688 5908
rect 25740 5856 25746 5908
rect 25774 5856 25780 5908
rect 25832 5896 25838 5908
rect 26887 5899 26945 5905
rect 26887 5896 26899 5899
rect 25832 5868 26899 5896
rect 25832 5856 25838 5868
rect 26887 5865 26899 5868
rect 26933 5865 26945 5899
rect 26887 5859 26945 5865
rect 29270 5856 29276 5908
rect 29328 5856 29334 5908
rect 29454 5856 29460 5908
rect 29512 5856 29518 5908
rect 6196 5760 6408 5764
rect 6549 5763 6607 5769
rect 6549 5760 6561 5763
rect 1964 5732 2774 5760
rect 3436 5732 5028 5760
rect 5460 5736 6561 5760
rect 5460 5732 6224 5736
rect 6380 5732 6561 5736
rect 676 5692 704 5720
rect 1801 5713 1859 5719
rect 1305 5695 1363 5701
rect 1305 5692 1317 5695
rect 676 5664 1317 5692
rect 1305 5661 1317 5664
rect 1351 5661 1363 5695
rect 1801 5679 1813 5713
rect 1847 5692 1859 5713
rect 1964 5692 1992 5732
rect 1847 5679 1992 5692
rect 1801 5673 1992 5679
rect 1826 5664 1992 5673
rect 2041 5695 2099 5701
rect 1305 5655 1363 5661
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 3436 5692 3464 5732
rect 5000 5704 5028 5732
rect 6549 5729 6561 5732
rect 6595 5729 6607 5763
rect 10413 5763 10471 5769
rect 10413 5760 10425 5763
rect 6549 5723 6607 5729
rect 6748 5732 10425 5760
rect 6748 5704 6776 5732
rect 10413 5729 10425 5732
rect 10459 5760 10471 5763
rect 10781 5763 10839 5769
rect 10781 5760 10793 5763
rect 10459 5732 10793 5760
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 10781 5729 10793 5732
rect 10827 5729 10839 5763
rect 10781 5723 10839 5729
rect 11149 5763 11207 5769
rect 11149 5729 11161 5763
rect 11195 5729 11207 5763
rect 11149 5723 11207 5729
rect 2087 5664 3464 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 3510 5652 3516 5704
rect 3568 5652 3574 5704
rect 4062 5701 4068 5704
rect 4019 5695 4068 5701
rect 4019 5661 4031 5695
rect 4065 5661 4068 5695
rect 4019 5655 4068 5661
rect 4062 5652 4068 5655
rect 4120 5652 4126 5704
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 4614 5692 4620 5704
rect 4295 5664 4620 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 4982 5652 4988 5704
rect 5040 5652 5046 5704
rect 5810 5652 5816 5704
rect 5868 5652 5874 5704
rect 6270 5652 6276 5704
rect 6328 5652 6334 5704
rect 6730 5652 6736 5704
rect 6788 5652 6794 5704
rect 7742 5652 7748 5704
rect 7800 5692 7806 5704
rect 8021 5695 8079 5701
rect 8021 5692 8033 5695
rect 7800 5664 8033 5692
rect 7800 5652 7806 5664
rect 8021 5661 8033 5664
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 8478 5652 8484 5704
rect 8536 5652 8542 5704
rect 8754 5652 8760 5704
rect 8812 5652 8818 5704
rect 10796 5692 10824 5723
rect 11422 5720 11428 5772
rect 11480 5720 11486 5772
rect 11514 5720 11520 5772
rect 11572 5760 11578 5772
rect 11936 5763 11994 5769
rect 11936 5760 11948 5763
rect 11572 5732 11948 5760
rect 11572 5720 11578 5732
rect 11936 5729 11948 5732
rect 11982 5729 11994 5763
rect 12434 5760 12440 5772
rect 11936 5723 11994 5729
rect 12268 5732 12440 5760
rect 10796 5664 11560 5692
rect 10597 5627 10655 5633
rect 10597 5593 10609 5627
rect 10643 5624 10655 5627
rect 11330 5624 11336 5636
rect 10643 5596 11336 5624
rect 10643 5593 10655 5596
rect 10597 5587 10655 5593
rect 11330 5584 11336 5596
rect 11388 5584 11394 5636
rect 3329 5559 3387 5565
rect 3329 5525 3341 5559
rect 3375 5556 3387 5559
rect 3970 5556 3976 5568
rect 3375 5528 3976 5556
rect 3375 5525 3387 5528
rect 3329 5519 3387 5525
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 4246 5516 4252 5568
rect 4304 5556 4310 5568
rect 4982 5556 4988 5568
rect 4304 5528 4988 5556
rect 4304 5516 4310 5528
rect 4982 5516 4988 5528
rect 5040 5516 5046 5568
rect 5537 5559 5595 5565
rect 5537 5525 5549 5559
rect 5583 5556 5595 5559
rect 6454 5556 6460 5568
rect 5583 5528 6460 5556
rect 5583 5525 5595 5528
rect 5537 5519 5595 5525
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 7006 5516 7012 5568
rect 7064 5556 7070 5568
rect 7653 5559 7711 5565
rect 7653 5556 7665 5559
rect 7064 5528 7665 5556
rect 7064 5516 7070 5528
rect 7653 5525 7665 5528
rect 7699 5525 7711 5559
rect 7653 5519 7711 5525
rect 9582 5516 9588 5568
rect 9640 5556 9646 5568
rect 9861 5559 9919 5565
rect 9861 5556 9873 5559
rect 9640 5528 9873 5556
rect 9640 5516 9646 5528
rect 9861 5525 9873 5528
rect 9907 5525 9919 5559
rect 9861 5519 9919 5525
rect 10226 5516 10232 5568
rect 10284 5516 10290 5568
rect 10318 5516 10324 5568
rect 10376 5556 10382 5568
rect 11241 5559 11299 5565
rect 11241 5556 11253 5559
rect 10376 5528 11253 5556
rect 10376 5516 10382 5528
rect 11241 5525 11253 5528
rect 11287 5525 11299 5559
rect 11532 5556 11560 5664
rect 11606 5652 11612 5704
rect 11664 5652 11670 5704
rect 12115 5695 12173 5701
rect 12115 5661 12127 5695
rect 12161 5692 12173 5695
rect 12268 5692 12296 5732
rect 12434 5720 12440 5732
rect 12492 5720 12498 5772
rect 12161 5664 12296 5692
rect 12345 5695 12403 5701
rect 12161 5661 12173 5664
rect 12115 5655 12173 5661
rect 12345 5661 12357 5695
rect 12391 5692 12403 5695
rect 13556 5692 13584 5856
rect 13722 5720 13728 5772
rect 13780 5760 13786 5772
rect 13780 5732 14320 5760
rect 13780 5720 13786 5732
rect 14292 5719 14320 5732
rect 14458 5720 14464 5772
rect 14516 5760 14522 5772
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 14516 5732 14565 5760
rect 14516 5720 14522 5732
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 15933 5763 15991 5769
rect 15933 5729 15945 5763
rect 15979 5760 15991 5763
rect 15979 5732 16712 5760
rect 15979 5729 15991 5732
rect 15933 5723 15991 5729
rect 14292 5713 14354 5719
rect 12391 5664 13584 5692
rect 12391 5661 12403 5664
rect 12345 5655 12403 5661
rect 13814 5652 13820 5704
rect 13872 5652 13878 5704
rect 13998 5652 14004 5704
rect 14056 5692 14062 5704
rect 14144 5695 14202 5701
rect 14144 5692 14156 5695
rect 14056 5664 14156 5692
rect 14056 5652 14062 5664
rect 14144 5661 14156 5664
rect 14190 5661 14202 5695
rect 14292 5682 14308 5713
rect 14296 5679 14308 5682
rect 14342 5679 14354 5713
rect 14296 5673 14354 5679
rect 14144 5655 14202 5661
rect 16206 5652 16212 5704
rect 16264 5652 16270 5704
rect 16574 5701 16580 5704
rect 16536 5695 16580 5701
rect 16536 5661 16548 5695
rect 16536 5655 16580 5661
rect 16574 5652 16580 5655
rect 16632 5652 16638 5704
rect 16684 5701 16712 5732
rect 16850 5720 16856 5772
rect 16908 5760 16914 5772
rect 16945 5763 17003 5769
rect 16945 5760 16957 5763
rect 16908 5732 16957 5760
rect 16908 5720 16914 5732
rect 16945 5729 16957 5732
rect 16991 5729 17003 5763
rect 16945 5723 17003 5729
rect 18325 5763 18383 5769
rect 18325 5729 18337 5763
rect 18371 5760 18383 5763
rect 19153 5763 19211 5769
rect 18371 5732 18920 5760
rect 18371 5729 18383 5732
rect 18325 5723 18383 5729
rect 18782 5701 18788 5704
rect 16672 5695 16730 5701
rect 16672 5661 16684 5695
rect 16718 5661 16730 5695
rect 18417 5695 18475 5701
rect 18417 5692 18429 5695
rect 16672 5655 16730 5661
rect 18340 5664 18429 5692
rect 18340 5568 18368 5664
rect 18417 5661 18429 5664
rect 18463 5661 18475 5695
rect 18417 5655 18475 5661
rect 18744 5695 18788 5701
rect 18744 5661 18756 5695
rect 18744 5655 18788 5661
rect 18782 5652 18788 5655
rect 18840 5652 18846 5704
rect 18892 5701 18920 5732
rect 19153 5729 19165 5763
rect 19199 5760 19211 5763
rect 20364 5760 20392 5856
rect 20622 5788 20628 5840
rect 20680 5788 20686 5840
rect 19199 5732 20392 5760
rect 20640 5760 20668 5788
rect 21100 5769 21128 5856
rect 20809 5763 20867 5769
rect 20809 5760 20821 5763
rect 20640 5732 20821 5760
rect 19199 5729 19211 5732
rect 19153 5723 19211 5729
rect 20809 5729 20821 5732
rect 20855 5729 20867 5763
rect 20809 5723 20867 5729
rect 21077 5763 21135 5769
rect 21077 5729 21089 5763
rect 21123 5729 21135 5763
rect 21077 5723 21135 5729
rect 21174 5720 21180 5772
rect 21232 5760 21238 5772
rect 21269 5763 21327 5769
rect 21269 5760 21281 5763
rect 21232 5732 21281 5760
rect 21232 5720 21238 5732
rect 21269 5729 21281 5732
rect 21315 5729 21327 5763
rect 21269 5723 21327 5729
rect 21818 5720 21824 5772
rect 21876 5760 21882 5772
rect 22005 5763 22063 5769
rect 22005 5760 22017 5763
rect 21876 5732 22017 5760
rect 21876 5720 21882 5732
rect 22005 5729 22017 5732
rect 22051 5729 22063 5763
rect 22005 5723 22063 5729
rect 23385 5763 23443 5769
rect 23385 5729 23397 5763
rect 23431 5760 23443 5763
rect 25869 5763 25927 5769
rect 23431 5732 23980 5760
rect 23431 5729 23443 5732
rect 23385 5723 23443 5729
rect 18880 5695 18938 5701
rect 18880 5661 18892 5695
rect 18926 5661 18938 5695
rect 18880 5655 18938 5661
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5692 20591 5695
rect 21732 5695 21790 5701
rect 21732 5692 21744 5695
rect 20579 5664 21744 5692
rect 20579 5661 20591 5664
rect 20533 5655 20591 5661
rect 21732 5661 21744 5664
rect 21778 5661 21790 5695
rect 21732 5655 21790 5661
rect 22186 5652 22192 5704
rect 22244 5692 22250 5704
rect 23952 5701 23980 5732
rect 25869 5729 25881 5763
rect 25915 5729 25927 5763
rect 25869 5723 25927 5729
rect 23477 5695 23535 5701
rect 23477 5692 23489 5695
rect 22244 5664 23489 5692
rect 22244 5652 22250 5664
rect 23477 5661 23489 5664
rect 23523 5661 23535 5695
rect 23477 5655 23535 5661
rect 23940 5695 23998 5701
rect 23940 5661 23952 5695
rect 23986 5661 23998 5695
rect 23940 5655 23998 5661
rect 24210 5652 24216 5704
rect 24268 5652 24274 5704
rect 25884 5692 25912 5723
rect 26050 5720 26056 5772
rect 26108 5760 26114 5772
rect 26145 5763 26203 5769
rect 26145 5760 26157 5763
rect 26108 5732 26157 5760
rect 26108 5720 26114 5732
rect 26145 5729 26157 5732
rect 26191 5729 26203 5763
rect 26145 5723 26203 5729
rect 26326 5720 26332 5772
rect 26384 5760 26390 5772
rect 26421 5763 26479 5769
rect 26421 5760 26433 5763
rect 26384 5732 26433 5760
rect 26384 5720 26390 5732
rect 26421 5729 26433 5732
rect 26467 5729 26479 5763
rect 28629 5763 28687 5769
rect 28629 5760 28641 5763
rect 26421 5723 26479 5729
rect 26712 5732 28641 5760
rect 26712 5692 26740 5732
rect 28629 5729 28641 5732
rect 28675 5760 28687 5763
rect 29086 5760 29092 5772
rect 28675 5732 29092 5760
rect 28675 5729 28687 5732
rect 28629 5723 28687 5729
rect 29086 5720 29092 5732
rect 29144 5720 29150 5772
rect 29181 5763 29239 5769
rect 29181 5729 29193 5763
rect 29227 5760 29239 5763
rect 29288 5760 29316 5856
rect 29472 5769 29500 5856
rect 29227 5732 29316 5760
rect 29457 5763 29515 5769
rect 29227 5729 29239 5732
rect 29181 5723 29239 5729
rect 29457 5729 29469 5763
rect 29503 5729 29515 5763
rect 29457 5723 29515 5729
rect 25884 5664 26740 5692
rect 26786 5652 26792 5704
rect 26844 5692 26850 5704
rect 26884 5695 26942 5701
rect 26884 5692 26896 5695
rect 26844 5664 26896 5692
rect 26844 5652 26850 5664
rect 26884 5661 26896 5664
rect 26930 5661 26942 5695
rect 26884 5655 26942 5661
rect 27154 5652 27160 5704
rect 27212 5652 27218 5704
rect 27246 5652 27252 5704
rect 27304 5692 27310 5704
rect 29472 5692 29500 5723
rect 27304 5664 29500 5692
rect 27304 5652 27310 5664
rect 20622 5584 20628 5636
rect 20680 5584 20686 5636
rect 28350 5584 28356 5636
rect 28408 5624 28414 5636
rect 28408 5596 29040 5624
rect 28408 5584 28414 5596
rect 11790 5556 11796 5568
rect 11532 5528 11796 5556
rect 11241 5519 11299 5525
rect 11790 5516 11796 5528
rect 11848 5516 11854 5568
rect 13633 5559 13691 5565
rect 13633 5525 13645 5559
rect 13679 5556 13691 5559
rect 14274 5556 14280 5568
rect 13679 5528 14280 5556
rect 13679 5525 13691 5528
rect 13633 5519 13691 5525
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 15470 5516 15476 5568
rect 15528 5556 15534 5568
rect 16390 5556 16396 5568
rect 15528 5528 16396 5556
rect 15528 5516 15534 5528
rect 16390 5516 16396 5528
rect 16448 5516 16454 5568
rect 18322 5516 18328 5568
rect 18380 5516 18386 5568
rect 18598 5516 18604 5568
rect 18656 5556 18662 5568
rect 20806 5556 20812 5568
rect 18656 5528 20812 5556
rect 18656 5516 18662 5528
rect 20806 5516 20812 5528
rect 20864 5516 20870 5568
rect 20901 5559 20959 5565
rect 20901 5525 20913 5559
rect 20947 5556 20959 5559
rect 21450 5556 21456 5568
rect 20947 5528 21456 5556
rect 20947 5525 20959 5528
rect 20901 5519 20959 5525
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 23106 5516 23112 5568
rect 23164 5556 23170 5568
rect 24210 5556 24216 5568
rect 23164 5528 24216 5556
rect 23164 5516 23170 5528
rect 24210 5516 24216 5528
rect 24268 5516 24274 5568
rect 24946 5516 24952 5568
rect 25004 5556 25010 5568
rect 25317 5559 25375 5565
rect 25317 5556 25329 5559
rect 25004 5528 25329 5556
rect 25004 5516 25010 5528
rect 25317 5525 25329 5528
rect 25363 5525 25375 5559
rect 25317 5519 25375 5525
rect 25958 5516 25964 5568
rect 26016 5516 26022 5568
rect 26050 5516 26056 5568
rect 26108 5556 26114 5568
rect 27154 5556 27160 5568
rect 26108 5528 27160 5556
rect 26108 5516 26114 5528
rect 27154 5516 27160 5528
rect 27212 5516 27218 5568
rect 28258 5516 28264 5568
rect 28316 5516 28322 5568
rect 28442 5516 28448 5568
rect 28500 5556 28506 5568
rect 29012 5565 29040 5596
rect 28813 5559 28871 5565
rect 28813 5556 28825 5559
rect 28500 5528 28825 5556
rect 28500 5516 28506 5528
rect 28813 5525 28825 5528
rect 28859 5525 28871 5559
rect 28813 5519 28871 5525
rect 28997 5559 29055 5565
rect 28997 5525 29009 5559
rect 29043 5525 29055 5559
rect 28997 5519 29055 5525
rect 29270 5516 29276 5568
rect 29328 5516 29334 5568
rect 552 5466 30912 5488
rect 552 5414 4193 5466
rect 4245 5414 4257 5466
rect 4309 5414 4321 5466
rect 4373 5414 4385 5466
rect 4437 5414 4449 5466
rect 4501 5414 11783 5466
rect 11835 5414 11847 5466
rect 11899 5414 11911 5466
rect 11963 5414 11975 5466
rect 12027 5414 12039 5466
rect 12091 5414 19373 5466
rect 19425 5414 19437 5466
rect 19489 5414 19501 5466
rect 19553 5414 19565 5466
rect 19617 5414 19629 5466
rect 19681 5414 26963 5466
rect 27015 5414 27027 5466
rect 27079 5414 27091 5466
rect 27143 5414 27155 5466
rect 27207 5414 27219 5466
rect 27271 5414 30912 5466
rect 552 5392 30912 5414
rect 2866 5352 2872 5364
rect 952 5324 2872 5352
rect 658 5176 664 5228
rect 716 5216 722 5228
rect 952 5225 980 5324
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 2961 5355 3019 5361
rect 2961 5321 2973 5355
rect 3007 5352 3019 5355
rect 4062 5352 4068 5364
rect 3007 5324 4068 5352
rect 3007 5321 3019 5324
rect 2961 5315 3019 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 6270 5352 6276 5364
rect 5951 5324 6276 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 10226 5352 10232 5364
rect 7484 5324 10232 5352
rect 3418 5244 3424 5296
rect 3476 5284 3482 5296
rect 3513 5287 3571 5293
rect 3513 5284 3525 5287
rect 3476 5256 3525 5284
rect 3476 5244 3482 5256
rect 3513 5253 3525 5256
rect 3559 5253 3571 5287
rect 3513 5247 3571 5253
rect 6086 5244 6092 5296
rect 6144 5244 6150 5296
rect 937 5219 995 5225
rect 937 5216 949 5219
rect 716 5188 949 5216
rect 716 5176 722 5188
rect 937 5185 949 5188
rect 983 5185 995 5219
rect 4246 5216 4252 5228
rect 1448 5207 4252 5216
rect 937 5179 995 5185
rect 1433 5201 4252 5207
rect 1433 5167 1445 5201
rect 1479 5188 4252 5201
rect 1479 5167 1491 5188
rect 4246 5176 4252 5188
rect 4304 5176 4310 5228
rect 4387 5219 4445 5225
rect 4387 5185 4399 5219
rect 4433 5216 4445 5219
rect 5074 5216 5080 5228
rect 4433 5188 5080 5216
rect 4433 5185 4445 5188
rect 4387 5179 4445 5185
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 6104 5216 6132 5244
rect 6270 5216 6276 5228
rect 6104 5188 6276 5216
rect 6270 5176 6276 5188
rect 6328 5176 6334 5228
rect 6595 5219 6653 5225
rect 6595 5185 6607 5219
rect 6641 5216 6653 5219
rect 7006 5216 7012 5228
rect 6641 5188 7012 5216
rect 6641 5185 6653 5188
rect 6595 5179 6653 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 1433 5161 1491 5167
rect 1670 5108 1676 5160
rect 1728 5108 1734 5160
rect 3510 5108 3516 5160
rect 3568 5148 3574 5160
rect 3881 5151 3939 5157
rect 3881 5148 3893 5151
rect 3568 5120 3893 5148
rect 3568 5108 3574 5120
rect 3881 5117 3893 5120
rect 3927 5117 3939 5151
rect 4617 5151 4675 5157
rect 4617 5148 4629 5151
rect 3881 5111 3939 5117
rect 3988 5120 4629 5148
rect 2866 5040 2872 5092
rect 2924 5080 2930 5092
rect 3329 5083 3387 5089
rect 3329 5080 3341 5083
rect 2924 5052 3341 5080
rect 2924 5040 2930 5052
rect 3329 5049 3341 5052
rect 3375 5080 3387 5083
rect 3694 5080 3700 5092
rect 3375 5052 3700 5080
rect 3375 5049 3387 5052
rect 3329 5043 3387 5049
rect 3694 5040 3700 5052
rect 3752 5040 3758 5092
rect 3786 5040 3792 5092
rect 3844 5080 3850 5092
rect 3988 5080 4016 5120
rect 4617 5117 4629 5120
rect 4663 5117 4675 5151
rect 4617 5111 4675 5117
rect 5350 5108 5356 5160
rect 5408 5108 5414 5160
rect 6089 5151 6147 5157
rect 6089 5117 6101 5151
rect 6135 5148 6147 5151
rect 6730 5148 6736 5160
rect 6135 5120 6736 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 6730 5108 6736 5120
rect 6788 5108 6794 5160
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 7484 5148 7512 5324
rect 10226 5312 10232 5324
rect 10284 5312 10290 5364
rect 13265 5355 13323 5361
rect 11164 5324 13216 5352
rect 7558 5176 7564 5228
rect 7616 5216 7622 5228
rect 8573 5219 8631 5225
rect 8573 5216 8585 5219
rect 7616 5188 8585 5216
rect 7616 5176 7622 5188
rect 8573 5185 8585 5188
rect 8619 5216 8631 5219
rect 8846 5216 8852 5228
rect 8619 5188 8852 5216
rect 8619 5185 8631 5188
rect 8573 5179 8631 5185
rect 8846 5176 8852 5188
rect 8904 5176 8910 5228
rect 9398 5225 9404 5228
rect 9360 5219 9404 5225
rect 9360 5185 9372 5219
rect 9360 5179 9404 5185
rect 9398 5176 9404 5179
rect 9456 5176 9462 5228
rect 9496 5217 9554 5223
rect 9496 5183 9508 5217
rect 9542 5216 9554 5217
rect 9582 5216 9588 5228
rect 9542 5188 9588 5216
rect 9542 5183 9554 5188
rect 9496 5177 9554 5183
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 11054 5216 11060 5228
rect 9692 5188 11060 5216
rect 6871 5120 7512 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 7834 5108 7840 5160
rect 7892 5148 7898 5160
rect 8389 5151 8447 5157
rect 8389 5148 8401 5151
rect 7892 5120 8401 5148
rect 7892 5108 7898 5120
rect 8389 5117 8401 5120
rect 8435 5148 8447 5151
rect 8938 5148 8944 5160
rect 8435 5120 8944 5148
rect 8435 5117 8447 5120
rect 8389 5111 8447 5117
rect 8938 5108 8944 5120
rect 8996 5108 9002 5160
rect 9030 5108 9036 5160
rect 9088 5108 9094 5160
rect 9692 5148 9720 5188
rect 11054 5176 11060 5188
rect 11112 5176 11118 5228
rect 9140 5120 9720 5148
rect 3844 5052 4016 5080
rect 3844 5040 3850 5052
rect 1403 5015 1461 5021
rect 1403 4981 1415 5015
rect 1449 5012 1461 5015
rect 1762 5012 1768 5024
rect 1449 4984 1768 5012
rect 1449 4981 1461 4984
rect 1403 4975 1461 4981
rect 1762 4972 1768 4984
rect 1820 5012 1826 5024
rect 2130 5012 2136 5024
rect 1820 4984 2136 5012
rect 1820 4972 1826 4984
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 3878 4972 3884 5024
rect 3936 5012 3942 5024
rect 4347 5015 4405 5021
rect 4347 5012 4359 5015
rect 3936 4984 4359 5012
rect 3936 4972 3942 4984
rect 4347 4981 4359 4984
rect 4393 4981 4405 5015
rect 5368 5012 5396 5108
rect 6362 5012 6368 5024
rect 5368 4984 6368 5012
rect 4347 4975 4405 4981
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 6546 4972 6552 5024
rect 6604 5021 6610 5024
rect 6604 5012 6613 5021
rect 8113 5015 8171 5021
rect 6604 4984 6649 5012
rect 6604 4975 6613 4984
rect 8113 4981 8125 5015
rect 8159 5012 8171 5015
rect 9140 5012 9168 5120
rect 9766 5108 9772 5160
rect 9824 5108 9830 5160
rect 11164 5148 11192 5324
rect 13188 5284 13216 5324
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13722 5352 13728 5364
rect 13311 5324 13728 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 21726 5352 21732 5364
rect 14022 5324 21732 5352
rect 14022 5284 14050 5324
rect 21726 5312 21732 5324
rect 21784 5312 21790 5364
rect 23014 5312 23020 5364
rect 23072 5352 23078 5364
rect 23385 5355 23443 5361
rect 23385 5352 23397 5355
rect 23072 5324 23397 5352
rect 23072 5312 23078 5324
rect 23385 5321 23397 5324
rect 23431 5321 23443 5355
rect 29181 5355 29239 5361
rect 29181 5352 29193 5355
rect 23385 5315 23443 5321
rect 23492 5324 29193 5352
rect 13188 5256 14050 5284
rect 23106 5244 23112 5296
rect 23164 5244 23170 5296
rect 11241 5219 11299 5225
rect 11241 5185 11253 5219
rect 11287 5216 11299 5219
rect 11422 5216 11428 5228
rect 11287 5188 11428 5216
rect 11287 5185 11299 5188
rect 11241 5179 11299 5185
rect 11422 5176 11428 5188
rect 11480 5216 11486 5228
rect 11606 5216 11612 5228
rect 11480 5188 11612 5216
rect 11480 5176 11486 5188
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 11698 5176 11704 5228
rect 11756 5216 11762 5228
rect 11977 5219 12035 5225
rect 11756 5188 11801 5216
rect 11756 5176 11762 5188
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 12802 5216 12808 5228
rect 12023 5188 12808 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 12802 5176 12808 5188
rect 12860 5176 12866 5228
rect 13630 5176 13636 5228
rect 13688 5176 13694 5228
rect 14001 5219 14059 5225
rect 14001 5216 14013 5219
rect 13832 5188 14013 5216
rect 10980 5120 11192 5148
rect 8159 4984 9168 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 6604 4972 6610 4975
rect 9490 4972 9496 5024
rect 9548 5012 9554 5024
rect 10980 5012 11008 5120
rect 11882 5108 11888 5160
rect 11940 5148 11946 5160
rect 13648 5148 13676 5176
rect 13832 5160 13860 5188
rect 14001 5185 14013 5188
rect 14047 5185 14059 5219
rect 14464 5219 14522 5225
rect 14464 5216 14476 5219
rect 14001 5179 14059 5185
rect 14108 5188 14476 5216
rect 11940 5120 13676 5148
rect 11940 5108 11946 5120
rect 13814 5108 13820 5160
rect 13872 5108 13878 5160
rect 13906 5108 13912 5160
rect 13964 5108 13970 5160
rect 11146 5040 11152 5092
rect 11204 5040 11210 5092
rect 14108 5080 14136 5188
rect 14464 5185 14476 5188
rect 14510 5185 14522 5219
rect 14464 5179 14522 5185
rect 14550 5176 14556 5228
rect 14608 5216 14614 5228
rect 14737 5219 14795 5225
rect 14737 5216 14749 5219
rect 14608 5188 14749 5216
rect 14608 5176 14614 5188
rect 14737 5185 14749 5188
rect 14783 5185 14795 5219
rect 14737 5179 14795 5185
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 16672 5219 16730 5225
rect 16672 5216 16684 5219
rect 16163 5188 16684 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 16672 5185 16684 5188
rect 16718 5185 16730 5219
rect 16672 5179 16730 5185
rect 16942 5176 16948 5228
rect 17000 5176 17006 5228
rect 18325 5219 18383 5225
rect 18325 5185 18337 5219
rect 18371 5216 18383 5219
rect 19156 5219 19214 5225
rect 19156 5216 19168 5219
rect 18371 5188 19168 5216
rect 18371 5185 18383 5188
rect 18325 5179 18383 5185
rect 19156 5185 19168 5188
rect 19202 5185 19214 5219
rect 19156 5179 19214 5185
rect 19429 5219 19487 5225
rect 19429 5185 19441 5219
rect 19475 5216 19487 5219
rect 20254 5216 20260 5228
rect 19475 5188 20260 5216
rect 19475 5185 19487 5188
rect 19429 5179 19487 5185
rect 20254 5176 20260 5188
rect 20312 5176 20318 5228
rect 20809 5219 20867 5225
rect 20809 5185 20821 5219
rect 20855 5216 20867 5219
rect 21364 5219 21422 5225
rect 21364 5216 21376 5219
rect 20855 5188 21376 5216
rect 20855 5185 20867 5188
rect 20809 5179 20867 5185
rect 21364 5185 21376 5188
rect 21410 5185 21422 5219
rect 21364 5179 21422 5185
rect 21450 5176 21456 5228
rect 21508 5216 21514 5228
rect 21637 5219 21695 5225
rect 21637 5216 21649 5219
rect 21508 5188 21649 5216
rect 21508 5176 21514 5188
rect 21637 5185 21649 5188
rect 21683 5185 21695 5219
rect 21637 5179 21695 5185
rect 16209 5151 16267 5157
rect 16209 5117 16221 5151
rect 16255 5148 16267 5151
rect 16298 5148 16304 5160
rect 16255 5120 16304 5148
rect 16255 5117 16267 5120
rect 16209 5111 16267 5117
rect 16298 5108 16304 5120
rect 16356 5108 16362 5160
rect 18693 5151 18751 5157
rect 18693 5148 18705 5151
rect 18340 5120 18705 5148
rect 18340 5092 18368 5120
rect 18693 5117 18705 5120
rect 18739 5117 18751 5151
rect 18693 5111 18751 5117
rect 18806 5120 20668 5148
rect 13648 5052 14136 5080
rect 13648 5024 13676 5052
rect 18322 5040 18328 5092
rect 18380 5040 18386 5092
rect 18806 5080 18834 5120
rect 18708 5052 18834 5080
rect 9548 4984 11008 5012
rect 9548 4972 9554 4984
rect 11514 4972 11520 5024
rect 11572 5012 11578 5024
rect 11707 5015 11765 5021
rect 11707 5012 11719 5015
rect 11572 4984 11719 5012
rect 11572 4972 11578 4984
rect 11707 4981 11719 4984
rect 11753 4981 11765 5015
rect 11707 4975 11765 4981
rect 13630 4972 13636 5024
rect 13688 4972 13694 5024
rect 13722 4972 13728 5024
rect 13780 4972 13786 5024
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 14467 5015 14525 5021
rect 14467 5012 14479 5015
rect 14056 4984 14479 5012
rect 14056 4972 14062 4984
rect 14467 4981 14479 4984
rect 14513 4981 14525 5015
rect 14467 4975 14525 4981
rect 16574 4972 16580 5024
rect 16632 5012 16638 5024
rect 16675 5015 16733 5021
rect 16675 5012 16687 5015
rect 16632 4984 16687 5012
rect 16632 4972 16638 4984
rect 16675 4981 16687 4984
rect 16721 5012 16733 5015
rect 16850 5012 16856 5024
rect 16721 4984 16856 5012
rect 16721 4981 16733 4984
rect 16675 4975 16733 4981
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 17310 4972 17316 5024
rect 17368 5012 17374 5024
rect 18708 5012 18736 5052
rect 17368 4984 18736 5012
rect 17368 4972 17374 4984
rect 18782 4972 18788 5024
rect 18840 5012 18846 5024
rect 19159 5015 19217 5021
rect 19159 5012 19171 5015
rect 18840 4984 19171 5012
rect 18840 4972 18846 4984
rect 19159 4981 19171 4984
rect 19205 4981 19217 5015
rect 20640 5012 20668 5120
rect 20714 5108 20720 5160
rect 20772 5148 20778 5160
rect 20901 5151 20959 5157
rect 20901 5148 20913 5151
rect 20772 5120 20913 5148
rect 20772 5108 20778 5120
rect 20901 5117 20913 5120
rect 20947 5148 20959 5151
rect 21174 5148 21180 5160
rect 20947 5120 21180 5148
rect 20947 5117 20959 5120
rect 20901 5111 20959 5117
rect 21174 5108 21180 5120
rect 21232 5108 21238 5160
rect 22738 5108 22744 5160
rect 22796 5148 22802 5160
rect 23293 5151 23351 5157
rect 23293 5148 23305 5151
rect 22796 5120 23305 5148
rect 22796 5108 22802 5120
rect 23293 5117 23305 5120
rect 23339 5117 23351 5151
rect 23293 5111 23351 5117
rect 23492 5080 23520 5324
rect 29181 5321 29193 5324
rect 29227 5321 29239 5355
rect 29181 5315 29239 5321
rect 29362 5312 29368 5364
rect 29420 5312 29426 5364
rect 25498 5244 25504 5296
rect 25556 5284 25562 5296
rect 26237 5287 26295 5293
rect 26237 5284 26249 5287
rect 25556 5256 26249 5284
rect 25556 5244 25562 5256
rect 26237 5253 26249 5256
rect 26283 5253 26295 5287
rect 29380 5284 29408 5312
rect 26237 5247 26295 5253
rect 28966 5256 29408 5284
rect 24535 5219 24593 5225
rect 24535 5185 24547 5219
rect 24581 5216 24593 5219
rect 24946 5216 24952 5228
rect 24581 5188 24952 5216
rect 24581 5185 24593 5188
rect 24535 5179 24593 5185
rect 24946 5176 24952 5188
rect 25004 5176 25010 5228
rect 25958 5176 25964 5228
rect 26016 5176 26022 5228
rect 26602 5176 26608 5228
rect 26660 5216 26666 5228
rect 27024 5219 27082 5225
rect 27024 5216 27036 5219
rect 26660 5188 27036 5216
rect 26660 5176 26666 5188
rect 27024 5185 27036 5188
rect 27070 5185 27082 5219
rect 27433 5219 27491 5225
rect 27208 5207 27384 5216
rect 27024 5179 27082 5185
rect 27193 5201 27384 5207
rect 23569 5151 23627 5157
rect 23569 5117 23581 5151
rect 23615 5117 23627 5151
rect 23569 5111 23627 5117
rect 22664 5052 23520 5080
rect 23584 5080 23612 5111
rect 23842 5108 23848 5160
rect 23900 5148 23906 5160
rect 24029 5151 24087 5157
rect 24029 5148 24041 5151
rect 23900 5120 24041 5148
rect 23900 5108 23906 5120
rect 24029 5117 24041 5120
rect 24075 5117 24087 5151
rect 24029 5111 24087 5117
rect 24765 5151 24823 5157
rect 24765 5117 24777 5151
rect 24811 5148 24823 5151
rect 25976 5148 26004 5176
rect 27193 5167 27205 5201
rect 27239 5188 27384 5201
rect 27239 5167 27251 5188
rect 27193 5161 27251 5167
rect 24811 5120 26004 5148
rect 26421 5151 26479 5157
rect 24811 5117 24823 5120
rect 24765 5111 24823 5117
rect 26421 5117 26433 5151
rect 26467 5117 26479 5151
rect 26421 5111 26479 5117
rect 23658 5080 23664 5092
rect 23584 5052 23664 5080
rect 21266 5012 21272 5024
rect 20640 4984 21272 5012
rect 19159 4975 19217 4981
rect 21266 4972 21272 4984
rect 21324 4972 21330 5024
rect 21367 5015 21425 5021
rect 21367 4981 21379 5015
rect 21413 5012 21425 5015
rect 21542 5012 21548 5024
rect 21413 4984 21548 5012
rect 21413 4981 21425 4984
rect 21367 4975 21425 4981
rect 21542 4972 21548 4984
rect 21600 4972 21606 5024
rect 21634 4972 21640 5024
rect 21692 5012 21698 5024
rect 22664 5012 22692 5052
rect 23658 5040 23664 5052
rect 23716 5040 23722 5092
rect 26145 5083 26203 5089
rect 26145 5049 26157 5083
rect 26191 5080 26203 5083
rect 26326 5080 26332 5092
rect 26191 5052 26332 5080
rect 26191 5049 26203 5052
rect 26145 5043 26203 5049
rect 26326 5040 26332 5052
rect 26384 5040 26390 5092
rect 26436 5080 26464 5111
rect 26694 5108 26700 5160
rect 26752 5108 26758 5160
rect 27356 5148 27384 5188
rect 27433 5185 27445 5219
rect 27479 5216 27491 5219
rect 27522 5216 27528 5228
rect 27479 5188 27528 5216
rect 27479 5185 27491 5188
rect 27433 5179 27491 5185
rect 27522 5176 27528 5188
rect 27580 5176 27586 5228
rect 27798 5176 27804 5228
rect 27856 5216 27862 5228
rect 28966 5216 28994 5256
rect 27856 5188 28994 5216
rect 27856 5176 27862 5188
rect 29086 5176 29092 5228
rect 29144 5176 29150 5228
rect 28989 5151 29047 5157
rect 27356 5120 28672 5148
rect 26510 5080 26516 5092
rect 26436 5052 26516 5080
rect 26510 5040 26516 5052
rect 26568 5040 26574 5092
rect 21692 4984 22692 5012
rect 21692 4972 21698 4984
rect 22738 4972 22744 5024
rect 22796 4972 22802 5024
rect 24394 4972 24400 5024
rect 24452 5012 24458 5024
rect 24495 5015 24553 5021
rect 24495 5012 24507 5015
rect 24452 4984 24507 5012
rect 24452 4972 24458 4984
rect 24495 4981 24507 4984
rect 24541 4981 24553 5015
rect 24495 4975 24553 4981
rect 25222 4972 25228 5024
rect 25280 5012 25286 5024
rect 28537 5015 28595 5021
rect 28537 5012 28549 5015
rect 25280 4984 28549 5012
rect 25280 4972 25286 4984
rect 28537 4981 28549 4984
rect 28583 4981 28595 5015
rect 28644 5012 28672 5120
rect 28989 5117 29001 5151
rect 29035 5148 29047 5151
rect 29104 5148 29132 5176
rect 29035 5120 29132 5148
rect 29273 5151 29331 5157
rect 29035 5117 29047 5120
rect 28989 5111 29047 5117
rect 29273 5117 29285 5151
rect 29319 5148 29331 5151
rect 29380 5148 29408 5256
rect 29319 5120 29408 5148
rect 29319 5117 29331 5120
rect 29273 5111 29331 5117
rect 28994 5012 29000 5024
rect 28644 4984 29000 5012
rect 28537 4975 28595 4981
rect 28994 4972 29000 4984
rect 29052 4972 29058 5024
rect 29454 4972 29460 5024
rect 29512 4972 29518 5024
rect 552 4922 31072 4944
rect 552 4870 7988 4922
rect 8040 4870 8052 4922
rect 8104 4870 8116 4922
rect 8168 4870 8180 4922
rect 8232 4870 8244 4922
rect 8296 4870 15578 4922
rect 15630 4870 15642 4922
rect 15694 4870 15706 4922
rect 15758 4870 15770 4922
rect 15822 4870 15834 4922
rect 15886 4870 23168 4922
rect 23220 4870 23232 4922
rect 23284 4870 23296 4922
rect 23348 4870 23360 4922
rect 23412 4870 23424 4922
rect 23476 4870 30758 4922
rect 30810 4870 30822 4922
rect 30874 4870 30886 4922
rect 30938 4870 30950 4922
rect 31002 4870 31014 4922
rect 31066 4870 31072 4922
rect 552 4848 31072 4870
rect 842 4768 848 4820
rect 900 4808 906 4820
rect 1029 4811 1087 4817
rect 1029 4808 1041 4811
rect 900 4780 1041 4808
rect 900 4768 906 4780
rect 1029 4777 1041 4780
rect 1075 4777 1087 4811
rect 1946 4808 1952 4820
rect 1029 4771 1087 4777
rect 1228 4780 1952 4808
rect 1228 4681 1256 4780
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 3878 4768 3884 4820
rect 3936 4808 3942 4820
rect 3979 4811 4037 4817
rect 3979 4808 3991 4811
rect 3936 4780 3991 4808
rect 3936 4768 3942 4780
rect 3979 4777 3991 4780
rect 4025 4777 4037 4811
rect 3979 4771 4037 4777
rect 6270 4768 6276 4820
rect 6328 4817 6334 4820
rect 6328 4808 6337 4817
rect 8487 4811 8545 4817
rect 6328 4780 6373 4808
rect 6328 4771 6337 4780
rect 8487 4777 8499 4811
rect 8533 4808 8545 4811
rect 8662 4808 8668 4820
rect 8533 4780 8668 4808
rect 8533 4777 8545 4780
rect 8487 4771 8545 4777
rect 6328 4768 6334 4771
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 8846 4768 8852 4820
rect 8904 4808 8910 4820
rect 8904 4780 9674 4808
rect 8904 4768 8910 4780
rect 9646 4740 9674 4780
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 10597 4811 10655 4817
rect 10597 4808 10609 4811
rect 9824 4780 10609 4808
rect 9824 4768 9830 4780
rect 10597 4777 10609 4780
rect 10643 4777 10655 4811
rect 10597 4771 10655 4777
rect 10870 4768 10876 4820
rect 10928 4768 10934 4820
rect 10962 4768 10968 4820
rect 11020 4768 11026 4820
rect 11330 4808 11336 4820
rect 11256 4780 11336 4808
rect 10888 4740 10916 4768
rect 9646 4712 10916 4740
rect 1213 4675 1271 4681
rect 1213 4641 1225 4675
rect 1259 4641 1271 4675
rect 2774 4672 2780 4684
rect 1213 4635 1271 4641
rect 1964 4644 2780 4672
rect 1801 4625 1859 4631
rect 842 4564 848 4616
rect 900 4604 906 4616
rect 1305 4607 1363 4613
rect 1305 4604 1317 4607
rect 900 4576 1317 4604
rect 900 4564 906 4576
rect 1305 4573 1317 4576
rect 1351 4573 1363 4607
rect 1305 4567 1363 4573
rect 1486 4564 1492 4616
rect 1544 4604 1550 4616
rect 1632 4607 1690 4613
rect 1632 4604 1644 4607
rect 1544 4576 1644 4604
rect 1544 4564 1550 4576
rect 1632 4573 1644 4576
rect 1678 4573 1690 4607
rect 1801 4591 1813 4625
rect 1847 4604 1859 4625
rect 1964 4604 1992 4644
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 5629 4675 5687 4681
rect 2976 4644 4292 4672
rect 1847 4591 1992 4604
rect 1801 4585 1992 4591
rect 1816 4576 1992 4585
rect 1632 4567 1690 4573
rect 2038 4564 2044 4616
rect 2096 4564 2102 4616
rect 952 4508 1348 4536
rect 952 4480 980 4508
rect 934 4428 940 4480
rect 992 4428 998 4480
rect 1320 4468 1348 4508
rect 2976 4468 3004 4644
rect 3142 4564 3148 4616
rect 3200 4604 3206 4616
rect 3418 4604 3424 4616
rect 3200 4576 3424 4604
rect 3200 4564 3206 4576
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 3528 4480 3556 4567
rect 3970 4564 3976 4616
rect 4028 4604 4034 4616
rect 4264 4613 4292 4644
rect 5629 4641 5641 4675
rect 5675 4672 5687 4675
rect 5675 4656 6086 4672
rect 6196 4656 6319 4676
rect 5675 4648 6319 4656
rect 5675 4644 6224 4648
rect 5675 4641 5687 4644
rect 5629 4635 5687 4641
rect 6058 4628 6224 4644
rect 4249 4607 4307 4613
rect 4028 4576 4073 4604
rect 4028 4564 4034 4576
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 5810 4604 5816 4616
rect 5316 4576 5816 4604
rect 5316 4564 5322 4576
rect 5810 4564 5816 4576
rect 5868 4564 5874 4616
rect 6291 4615 6319 4648
rect 7929 4675 7987 4681
rect 7929 4641 7941 4675
rect 7975 4672 7987 4675
rect 7975 4644 8156 4672
rect 7975 4641 7987 4644
rect 7929 4635 7987 4641
rect 6276 4609 6334 4615
rect 6276 4575 6288 4609
rect 6322 4575 6334 4609
rect 6276 4569 6334 4575
rect 6362 4564 6368 4616
rect 6420 4604 6426 4616
rect 6549 4607 6607 4613
rect 6549 4604 6561 4607
rect 6420 4576 6561 4604
rect 6420 4564 6426 4576
rect 6549 4573 6561 4576
rect 6595 4573 6607 4607
rect 6549 4567 6607 4573
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 7742 4604 7748 4616
rect 6788 4576 7748 4604
rect 6788 4564 6794 4576
rect 7742 4564 7748 4576
rect 7800 4604 7806 4616
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 7800 4576 8033 4604
rect 7800 4564 7806 4576
rect 8021 4573 8033 4576
rect 8067 4573 8079 4607
rect 8128 4604 8156 4644
rect 8570 4632 8576 4684
rect 8628 4672 8634 4684
rect 8628 4644 8800 4672
rect 8628 4632 8634 4644
rect 8772 4613 8800 4644
rect 8846 4632 8852 4684
rect 8904 4672 8910 4684
rect 10413 4675 10471 4681
rect 10413 4672 10425 4675
rect 8904 4644 10425 4672
rect 8904 4632 8910 4644
rect 10413 4641 10425 4644
rect 10459 4641 10471 4675
rect 10413 4635 10471 4641
rect 10781 4675 10839 4681
rect 10781 4641 10793 4675
rect 10827 4672 10839 4675
rect 10980 4672 11008 4768
rect 10827 4644 11008 4672
rect 10827 4641 10839 4644
rect 10781 4635 10839 4641
rect 8484 4607 8542 4613
rect 8484 4604 8496 4607
rect 8128 4576 8496 4604
rect 8021 4567 8079 4573
rect 8484 4573 8496 4576
rect 8530 4573 8542 4607
rect 8484 4567 8542 4573
rect 8757 4607 8815 4613
rect 8757 4573 8769 4607
rect 8803 4573 8815 4607
rect 10428 4604 10456 4635
rect 11054 4632 11060 4684
rect 11112 4672 11118 4684
rect 11256 4681 11284 4780
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 11514 4768 11520 4820
rect 11572 4808 11578 4820
rect 12075 4811 12133 4817
rect 12075 4808 12087 4811
rect 11572 4780 12087 4808
rect 11572 4768 11578 4780
rect 12075 4777 12087 4780
rect 12121 4777 12133 4811
rect 12075 4771 12133 4777
rect 13630 4768 13636 4820
rect 13688 4768 13694 4820
rect 13722 4768 13728 4820
rect 13780 4768 13786 4820
rect 16675 4811 16733 4817
rect 16675 4777 16687 4811
rect 16721 4808 16733 4811
rect 16850 4808 16856 4820
rect 16721 4780 16856 4808
rect 16721 4777 16733 4780
rect 16675 4771 16733 4777
rect 16850 4768 16856 4780
rect 16908 4768 16914 4820
rect 17770 4768 17776 4820
rect 17828 4808 17834 4820
rect 21634 4808 21640 4820
rect 17828 4780 21640 4808
rect 17828 4768 17834 4780
rect 21634 4768 21640 4780
rect 21692 4768 21698 4820
rect 21726 4768 21732 4820
rect 21784 4768 21790 4820
rect 21818 4768 21824 4820
rect 21876 4808 21882 4820
rect 22005 4811 22063 4817
rect 22005 4808 22017 4811
rect 21876 4780 22017 4808
rect 21876 4768 21882 4780
rect 22005 4777 22017 4780
rect 22051 4777 22063 4811
rect 22005 4771 22063 4777
rect 22462 4768 22468 4820
rect 22520 4808 22526 4820
rect 22563 4811 22621 4817
rect 22563 4808 22575 4811
rect 22520 4780 22575 4808
rect 22520 4768 22526 4780
rect 22563 4777 22575 4780
rect 22609 4777 22621 4811
rect 22563 4771 22621 4777
rect 24489 4811 24547 4817
rect 24489 4777 24501 4811
rect 24535 4808 24547 4811
rect 26050 4808 26056 4820
rect 24535 4780 26056 4808
rect 24535 4777 24547 4780
rect 24489 4771 24547 4777
rect 26050 4768 26056 4780
rect 26108 4768 26114 4820
rect 28442 4808 28448 4820
rect 26896 4780 28448 4808
rect 11241 4675 11299 4681
rect 11241 4672 11253 4675
rect 11112 4644 11253 4672
rect 11112 4632 11118 4644
rect 11241 4641 11253 4644
rect 11287 4641 11299 4675
rect 11517 4675 11575 4681
rect 11517 4672 11529 4675
rect 11241 4635 11299 4641
rect 11348 4644 11529 4672
rect 11348 4604 11376 4644
rect 11517 4641 11529 4644
rect 11563 4672 11575 4675
rect 11882 4672 11888 4684
rect 11563 4644 11888 4672
rect 11563 4641 11575 4644
rect 11517 4635 11575 4641
rect 11882 4632 11888 4644
rect 11940 4632 11946 4684
rect 12345 4675 12403 4681
rect 12345 4641 12357 4675
rect 12391 4672 12403 4675
rect 13078 4672 13084 4684
rect 12391 4644 13084 4672
rect 12391 4641 12403 4644
rect 12345 4635 12403 4641
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13740 4672 13768 4768
rect 20530 4700 20536 4752
rect 20588 4700 20594 4752
rect 21266 4700 21272 4752
rect 21324 4740 21330 4752
rect 24213 4743 24271 4749
rect 21324 4712 21588 4740
rect 21324 4700 21330 4712
rect 14553 4675 14611 4681
rect 14553 4672 14565 4675
rect 13740 4644 14565 4672
rect 14553 4641 14565 4644
rect 14599 4641 14611 4675
rect 14553 4635 14611 4641
rect 15933 4675 15991 4681
rect 15933 4641 15945 4675
rect 15979 4672 15991 4675
rect 16945 4675 17003 4681
rect 15979 4644 16712 4672
rect 15979 4641 15991 4644
rect 15933 4635 15991 4641
rect 10428 4576 11376 4604
rect 8757 4567 8815 4573
rect 11422 4564 11428 4616
rect 11480 4604 11486 4616
rect 11609 4607 11667 4613
rect 11609 4604 11621 4607
rect 11480 4576 11621 4604
rect 11480 4564 11486 4576
rect 11609 4573 11621 4576
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 12066 4564 12072 4616
rect 12124 4606 12130 4616
rect 12124 4578 12167 4606
rect 12124 4564 12130 4578
rect 13814 4564 13820 4616
rect 13872 4564 13878 4616
rect 13998 4564 14004 4616
rect 14056 4604 14062 4616
rect 14144 4607 14202 4613
rect 14144 4604 14156 4607
rect 14056 4576 14156 4604
rect 14056 4564 14062 4576
rect 14144 4573 14156 4576
rect 14190 4573 14202 4607
rect 14144 4567 14202 4573
rect 14274 4564 14280 4616
rect 14332 4604 14338 4616
rect 16209 4607 16267 4613
rect 14332 4576 14377 4604
rect 14332 4564 14338 4576
rect 16209 4573 16221 4607
rect 16255 4604 16267 4607
rect 16390 4604 16396 4616
rect 16255 4576 16396 4604
rect 16255 4573 16267 4576
rect 16209 4567 16267 4573
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 16684 4613 16712 4644
rect 16945 4641 16957 4675
rect 16991 4672 17003 4675
rect 17218 4672 17224 4684
rect 16991 4644 17224 4672
rect 16991 4641 17003 4644
rect 16945 4635 17003 4641
rect 17218 4632 17224 4644
rect 17276 4632 17282 4684
rect 18325 4675 18383 4681
rect 18325 4641 18337 4675
rect 18371 4672 18383 4675
rect 18371 4644 18920 4672
rect 18371 4641 18383 4644
rect 18325 4635 18383 4641
rect 18782 4613 18788 4616
rect 16672 4607 16730 4613
rect 16672 4573 16684 4607
rect 16718 4573 16730 4607
rect 18417 4607 18475 4613
rect 18417 4604 18429 4607
rect 16672 4567 16730 4573
rect 18340 4576 18429 4604
rect 9490 4496 9496 4548
rect 9548 4536 9554 4548
rect 10229 4539 10287 4545
rect 10229 4536 10241 4539
rect 9548 4508 10241 4536
rect 9548 4496 9554 4508
rect 10229 4505 10241 4508
rect 10275 4505 10287 4539
rect 10229 4499 10287 4505
rect 11057 4539 11115 4545
rect 11057 4505 11069 4539
rect 11103 4536 11115 4539
rect 11514 4536 11520 4548
rect 11103 4508 11520 4536
rect 11103 4505 11115 4508
rect 11057 4499 11115 4505
rect 11514 4496 11520 4508
rect 11572 4496 11578 4548
rect 18340 4480 18368 4576
rect 18417 4573 18429 4576
rect 18463 4573 18475 4607
rect 18417 4567 18475 4573
rect 18744 4607 18788 4613
rect 18744 4573 18756 4607
rect 18744 4567 18788 4573
rect 18782 4564 18788 4567
rect 18840 4564 18846 4616
rect 18892 4613 18920 4644
rect 18966 4632 18972 4684
rect 19024 4672 19030 4684
rect 19153 4675 19211 4681
rect 19153 4672 19165 4675
rect 19024 4644 19165 4672
rect 19024 4632 19030 4644
rect 19153 4641 19165 4644
rect 19199 4641 19211 4675
rect 19153 4635 19211 4641
rect 20806 4632 20812 4684
rect 20864 4672 20870 4684
rect 21085 4675 21143 4681
rect 21085 4672 21097 4675
rect 20864 4644 21097 4672
rect 20864 4632 20870 4644
rect 21085 4641 21097 4644
rect 21131 4672 21143 4675
rect 21174 4672 21180 4684
rect 21131 4644 21180 4672
rect 21131 4641 21143 4644
rect 21085 4635 21143 4641
rect 21174 4632 21180 4644
rect 21232 4632 21238 4684
rect 21358 4632 21364 4684
rect 21416 4672 21422 4684
rect 21560 4681 21588 4712
rect 24213 4709 24225 4743
rect 24259 4740 24271 4743
rect 24302 4740 24308 4752
rect 24259 4712 24308 4740
rect 24259 4709 24271 4712
rect 24213 4703 24271 4709
rect 24302 4700 24308 4712
rect 24360 4700 24366 4752
rect 26896 4740 26924 4780
rect 28442 4768 28448 4780
rect 28500 4768 28506 4820
rect 29638 4768 29644 4820
rect 29696 4808 29702 4820
rect 29733 4811 29791 4817
rect 29733 4808 29745 4811
rect 29696 4780 29745 4808
rect 29696 4768 29702 4780
rect 29733 4777 29745 4780
rect 29779 4777 29791 4811
rect 29733 4771 29791 4777
rect 24780 4712 26924 4740
rect 21453 4675 21511 4681
rect 21453 4672 21465 4675
rect 21416 4644 21465 4672
rect 21416 4632 21422 4644
rect 21453 4641 21465 4644
rect 21499 4641 21511 4675
rect 21453 4635 21511 4641
rect 21545 4675 21603 4681
rect 21545 4641 21557 4675
rect 21591 4672 21603 4675
rect 21821 4675 21879 4681
rect 21821 4672 21833 4675
rect 21591 4644 21833 4672
rect 21591 4641 21603 4644
rect 21545 4635 21603 4641
rect 21821 4641 21833 4644
rect 21867 4641 21879 4675
rect 21821 4635 21879 4641
rect 22097 4675 22155 4681
rect 22097 4641 22109 4675
rect 22143 4672 22155 4675
rect 22186 4672 22192 4684
rect 22143 4644 22192 4672
rect 22143 4641 22155 4644
rect 22097 4635 22155 4641
rect 22186 4632 22192 4644
rect 22244 4632 22250 4684
rect 22738 4632 22744 4684
rect 22796 4632 22802 4684
rect 22830 4632 22836 4684
rect 22888 4632 22894 4684
rect 23658 4632 23664 4684
rect 23716 4672 23722 4684
rect 24673 4675 24731 4681
rect 24673 4672 24685 4675
rect 23716 4644 24685 4672
rect 23716 4632 23722 4644
rect 24673 4641 24685 4644
rect 24719 4672 24731 4675
rect 24780 4672 24808 4712
rect 24719 4644 24808 4672
rect 24719 4641 24731 4644
rect 24673 4635 24731 4641
rect 26142 4632 26148 4684
rect 26200 4672 26206 4684
rect 26896 4681 26924 4712
rect 27154 4700 27160 4752
rect 27212 4740 27218 4752
rect 27212 4712 28028 4740
rect 27212 4700 27218 4712
rect 26605 4675 26663 4681
rect 26605 4672 26617 4675
rect 26200 4644 26617 4672
rect 26200 4632 26206 4644
rect 26605 4641 26617 4644
rect 26651 4641 26663 4675
rect 26605 4635 26663 4641
rect 26881 4675 26939 4681
rect 26881 4641 26893 4675
rect 26927 4641 26939 4675
rect 26881 4635 26939 4641
rect 27065 4675 27123 4681
rect 27065 4641 27077 4675
rect 27111 4672 27123 4675
rect 27798 4672 27804 4684
rect 27111 4644 27804 4672
rect 27111 4641 27123 4644
rect 27065 4635 27123 4641
rect 27798 4632 27804 4644
rect 27856 4632 27862 4684
rect 27890 4632 27896 4684
rect 27948 4632 27954 4684
rect 28000 4672 28028 4712
rect 28000 4644 28399 4672
rect 18880 4607 18938 4613
rect 18880 4573 18892 4607
rect 18926 4573 18938 4607
rect 18880 4567 18938 4573
rect 19242 4564 19248 4616
rect 19300 4604 19306 4616
rect 22603 4607 22661 4613
rect 19300 4576 22094 4604
rect 19300 4564 19306 4576
rect 20625 4539 20683 4545
rect 20625 4536 20637 4539
rect 19812 4508 20637 4536
rect 1320 4440 3004 4468
rect 3142 4428 3148 4480
rect 3200 4428 3206 4480
rect 3510 4428 3516 4480
rect 3568 4468 3574 4480
rect 8846 4468 8852 4480
rect 3568 4440 8852 4468
rect 3568 4428 3574 4440
rect 8846 4428 8852 4440
rect 8904 4428 8910 4480
rect 10042 4428 10048 4480
rect 10100 4428 10106 4480
rect 11333 4471 11391 4477
rect 11333 4437 11345 4471
rect 11379 4468 11391 4471
rect 12158 4468 12164 4480
rect 11379 4440 12164 4468
rect 11379 4437 11391 4440
rect 11333 4431 11391 4437
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 12250 4428 12256 4480
rect 12308 4468 12314 4480
rect 16666 4468 16672 4480
rect 12308 4440 16672 4468
rect 12308 4428 12314 4440
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 18322 4428 18328 4480
rect 18380 4428 18386 4480
rect 19058 4428 19064 4480
rect 19116 4468 19122 4480
rect 19812 4468 19840 4508
rect 20625 4505 20637 4508
rect 20671 4505 20683 4539
rect 20625 4499 20683 4505
rect 19116 4440 19840 4468
rect 20901 4471 20959 4477
rect 19116 4428 19122 4440
rect 20901 4437 20913 4471
rect 20947 4468 20959 4471
rect 20990 4468 20996 4480
rect 20947 4440 20996 4468
rect 20947 4437 20959 4440
rect 20901 4431 20959 4437
rect 20990 4428 20996 4440
rect 21048 4428 21054 4480
rect 21269 4471 21327 4477
rect 21269 4437 21281 4471
rect 21315 4468 21327 4471
rect 21450 4468 21456 4480
rect 21315 4440 21456 4468
rect 21315 4437 21327 4440
rect 21269 4431 21327 4437
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 22066 4468 22094 4576
rect 22603 4573 22615 4607
rect 22649 4604 22661 4607
rect 22756 4604 22784 4632
rect 22649 4576 22784 4604
rect 22649 4573 22661 4576
rect 22603 4567 22661 4573
rect 26510 4564 26516 4616
rect 26568 4604 26574 4616
rect 28166 4604 28172 4616
rect 26568 4576 28172 4604
rect 26568 4564 26574 4576
rect 28166 4564 28172 4576
rect 28224 4613 28230 4616
rect 28371 4615 28399 4644
rect 28534 4632 28540 4684
rect 28592 4672 28598 4684
rect 28629 4675 28687 4681
rect 28629 4672 28641 4675
rect 28592 4644 28641 4672
rect 28592 4632 28598 4644
rect 28629 4641 28641 4644
rect 28675 4641 28687 4675
rect 28629 4635 28687 4641
rect 28224 4607 28278 4613
rect 28224 4573 28232 4607
rect 28266 4573 28278 4607
rect 28371 4609 28430 4615
rect 28371 4578 28384 4609
rect 28224 4567 28278 4573
rect 28372 4575 28384 4578
rect 28418 4575 28430 4609
rect 28372 4569 28430 4575
rect 28224 4564 28230 4567
rect 26786 4496 26792 4548
rect 26844 4536 26850 4548
rect 27890 4536 27896 4548
rect 26844 4508 27896 4536
rect 26844 4496 26850 4508
rect 27890 4496 27896 4508
rect 27948 4496 27954 4548
rect 24762 4468 24768 4480
rect 22066 4440 24768 4468
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 26421 4471 26479 4477
rect 26421 4437 26433 4471
rect 26467 4468 26479 4471
rect 26602 4468 26608 4480
rect 26467 4440 26608 4468
rect 26467 4437 26479 4440
rect 26421 4431 26479 4437
rect 26602 4428 26608 4440
rect 26660 4428 26666 4480
rect 26694 4428 26700 4480
rect 26752 4428 26758 4480
rect 26878 4428 26884 4480
rect 26936 4468 26942 4480
rect 27249 4471 27307 4477
rect 27249 4468 27261 4471
rect 26936 4440 27261 4468
rect 26936 4428 26942 4440
rect 27249 4437 27261 4440
rect 27295 4437 27307 4471
rect 27249 4431 27307 4437
rect 552 4378 30912 4400
rect 552 4326 4193 4378
rect 4245 4326 4257 4378
rect 4309 4326 4321 4378
rect 4373 4326 4385 4378
rect 4437 4326 4449 4378
rect 4501 4326 11783 4378
rect 11835 4326 11847 4378
rect 11899 4326 11911 4378
rect 11963 4326 11975 4378
rect 12027 4326 12039 4378
rect 12091 4326 19373 4378
rect 19425 4326 19437 4378
rect 19489 4326 19501 4378
rect 19553 4326 19565 4378
rect 19617 4326 19629 4378
rect 19681 4326 26963 4378
rect 27015 4326 27027 4378
rect 27079 4326 27091 4378
rect 27143 4326 27155 4378
rect 27207 4326 27219 4378
rect 27271 4326 30912 4378
rect 552 4304 30912 4326
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3108 4236 6040 4264
rect 3108 4224 3114 4236
rect 842 4088 848 4140
rect 900 4088 906 4140
rect 1302 4088 1308 4140
rect 1360 4119 1366 4140
rect 1360 4113 1399 4119
rect 1320 4082 1353 4088
rect 1341 4079 1353 4082
rect 1387 4079 1399 4113
rect 1578 4088 1584 4140
rect 1636 4088 1642 4140
rect 1670 4088 1676 4140
rect 1728 4128 1734 4140
rect 3970 4128 3976 4140
rect 1728 4100 3976 4128
rect 1728 4088 1734 4100
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 4252 4129 4310 4135
rect 4252 4095 4264 4129
rect 4298 4128 4310 4129
rect 4338 4128 4344 4140
rect 4298 4100 4344 4128
rect 4298 4095 4310 4100
rect 4252 4089 4310 4095
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 4522 4088 4528 4140
rect 4580 4088 4586 4140
rect 5902 4088 5908 4140
rect 5960 4088 5966 4140
rect 6012 4128 6040 4236
rect 7558 4224 7564 4276
rect 7616 4264 7622 4276
rect 7616 4236 11560 4264
rect 7616 4224 7622 4236
rect 9030 4156 9036 4208
rect 9088 4196 9094 4208
rect 11532 4196 11560 4236
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 11977 4267 12035 4273
rect 11977 4264 11989 4267
rect 11756 4236 11989 4264
rect 11756 4224 11762 4236
rect 11977 4233 11989 4236
rect 12023 4233 12035 4267
rect 26878 4264 26884 4276
rect 11977 4227 12035 4233
rect 15580 4236 26884 4264
rect 12250 4196 12256 4208
rect 9088 4168 9812 4196
rect 11532 4168 12256 4196
rect 9088 4156 9094 4168
rect 6012 4100 6132 4128
rect 1341 4073 1399 4079
rect 2958 4020 2964 4072
rect 3016 4020 3022 4072
rect 3789 4063 3847 4069
rect 3789 4029 3801 4063
rect 3835 4060 3847 4063
rect 5442 4060 5448 4072
rect 3835 4032 5448 4060
rect 3835 4029 3847 4032
rect 3789 4023 3847 4029
rect 3804 3992 3832 4023
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5626 4020 5632 4072
rect 5684 4060 5690 4072
rect 5997 4063 6055 4069
rect 5997 4060 6009 4063
rect 5684 4032 6009 4060
rect 5684 4020 5690 4032
rect 5997 4029 6009 4032
rect 6043 4029 6055 4063
rect 6104 4060 6132 4100
rect 6178 4088 6184 4140
rect 6236 4128 6242 4140
rect 6324 4131 6382 4137
rect 6324 4128 6336 4131
rect 6236 4100 6336 4128
rect 6236 4088 6242 4100
rect 6324 4097 6336 4100
rect 6370 4097 6382 4131
rect 6324 4091 6382 4097
rect 6460 4129 6518 4135
rect 6460 4095 6472 4129
rect 6506 4095 6518 4129
rect 9674 4128 9680 4140
rect 6460 4089 6518 4095
rect 6748 4100 9680 4128
rect 6475 4060 6503 4089
rect 6748 4069 6776 4100
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 6104 4032 6503 4060
rect 6733 4063 6791 4069
rect 5997 4023 6055 4029
rect 6733 4029 6745 4063
rect 6779 4029 6791 4063
rect 6733 4023 6791 4029
rect 8389 4063 8447 4069
rect 8389 4029 8401 4063
rect 8435 4060 8447 4063
rect 8938 4060 8944 4072
rect 8435 4032 8944 4060
rect 8435 4029 8447 4032
rect 8389 4023 8447 4029
rect 2240 3964 3832 3992
rect 1311 3927 1369 3933
rect 1311 3893 1323 3927
rect 1357 3924 1369 3927
rect 1486 3924 1492 3936
rect 1357 3896 1492 3924
rect 1357 3893 1369 3896
rect 1311 3887 1369 3893
rect 1486 3884 1492 3896
rect 1544 3884 1550 3936
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 2240 3924 2268 3964
rect 1636 3896 2268 3924
rect 1636 3884 1642 3896
rect 3050 3884 3056 3936
rect 3108 3924 3114 3936
rect 3421 3927 3479 3933
rect 3421 3924 3433 3927
rect 3108 3896 3433 3924
rect 3108 3884 3114 3896
rect 3421 3893 3433 3896
rect 3467 3893 3479 3927
rect 3421 3887 3479 3893
rect 3694 3884 3700 3936
rect 3752 3924 3758 3936
rect 4255 3927 4313 3933
rect 4255 3924 4267 3927
rect 3752 3896 4267 3924
rect 3752 3884 3758 3896
rect 4255 3893 4267 3896
rect 4301 3924 4313 3927
rect 5626 3924 5632 3936
rect 4301 3896 5632 3924
rect 4301 3893 4313 3896
rect 4255 3887 4313 3893
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 6012 3924 6040 4023
rect 8938 4020 8944 4032
rect 8996 4020 9002 4072
rect 9585 4063 9643 4069
rect 9585 4060 9597 4063
rect 9324 4032 9597 4060
rect 7484 3964 8340 3992
rect 7484 3924 7512 3964
rect 6012 3896 7512 3924
rect 7834 3884 7840 3936
rect 7892 3884 7898 3936
rect 8312 3924 8340 3964
rect 8662 3952 8668 4004
rect 8720 3952 8726 4004
rect 8846 3952 8852 4004
rect 8904 3992 8910 4004
rect 9033 3995 9091 4001
rect 9033 3992 9045 3995
rect 8904 3964 9045 3992
rect 8904 3952 8910 3964
rect 9033 3961 9045 3964
rect 9079 3961 9091 3995
rect 9033 3955 9091 3961
rect 9125 3927 9183 3933
rect 9125 3924 9137 3927
rect 8312 3896 9137 3924
rect 9125 3893 9137 3896
rect 9171 3893 9183 3927
rect 9324 3924 9352 4032
rect 9585 4029 9597 4032
rect 9631 4029 9643 4063
rect 9784 4060 9812 4168
rect 12250 4156 12256 4168
rect 12308 4156 12314 4208
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10600 4131 10658 4137
rect 10600 4128 10612 4131
rect 10100 4100 10612 4128
rect 10100 4088 10106 4100
rect 10600 4097 10612 4100
rect 10646 4097 10658 4131
rect 10600 4091 10658 4097
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 10873 4131 10931 4137
rect 10873 4128 10885 4131
rect 10744 4100 10885 4128
rect 10744 4088 10750 4100
rect 10873 4097 10885 4100
rect 10919 4097 10931 4131
rect 10873 4091 10931 4097
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4128 13323 4131
rect 13814 4128 13820 4140
rect 13311 4100 13820 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 13909 4131 13967 4137
rect 13909 4097 13921 4131
rect 13955 4128 13967 4131
rect 14642 4128 14648 4140
rect 13955 4100 14648 4128
rect 13955 4097 13967 4100
rect 13909 4091 13967 4097
rect 14642 4088 14648 4100
rect 14700 4137 14706 4140
rect 14700 4131 14749 4137
rect 14700 4097 14703 4131
rect 14737 4128 14749 4131
rect 15580 4128 15608 4236
rect 26878 4224 26884 4236
rect 26936 4224 26942 4276
rect 19242 4196 19248 4208
rect 18524 4168 19248 4196
rect 17862 4128 17868 4140
rect 14737 4100 14793 4128
rect 15028 4100 15608 4128
rect 15672 4100 16528 4128
rect 14737 4097 14749 4100
rect 14700 4091 14749 4097
rect 14700 4088 14706 4091
rect 10137 4063 10195 4069
rect 10137 4060 10149 4063
rect 9784 4032 10149 4060
rect 9585 4023 9643 4029
rect 10137 4029 10149 4032
rect 10183 4060 10195 4063
rect 10502 4060 10508 4072
rect 10183 4032 10508 4060
rect 10183 4029 10195 4032
rect 10137 4023 10195 4029
rect 10502 4020 10508 4032
rect 10560 4020 10566 4072
rect 12802 4020 12808 4072
rect 12860 4060 12866 4072
rect 14185 4063 14243 4069
rect 14185 4060 14197 4063
rect 12860 4032 14197 4060
rect 12860 4020 12866 4032
rect 14185 4029 14197 4032
rect 14231 4029 14243 4063
rect 14185 4023 14243 4029
rect 14512 4063 14570 4069
rect 14512 4029 14524 4063
rect 14558 4060 14570 4063
rect 14826 4060 14832 4072
rect 14558 4032 14832 4060
rect 14558 4029 14570 4032
rect 14512 4023 14570 4029
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 14921 4063 14979 4069
rect 14921 4029 14933 4063
rect 14967 4060 14979 4063
rect 15028 4060 15056 4100
rect 14967 4032 15056 4060
rect 14967 4029 14979 4032
rect 14921 4023 14979 4029
rect 15194 4020 15200 4072
rect 15252 4060 15258 4072
rect 15672 4060 15700 4100
rect 16500 4072 16528 4100
rect 16874 4113 17868 4128
rect 16874 4082 16901 4113
rect 16889 4079 16901 4082
rect 16935 4100 17868 4113
rect 16935 4079 16947 4100
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 18524 4137 18552 4168
rect 19242 4156 19248 4168
rect 19300 4156 19306 4208
rect 18509 4131 18567 4137
rect 18509 4097 18521 4131
rect 18555 4097 18567 4131
rect 18509 4091 18567 4097
rect 18782 4088 18788 4140
rect 18840 4128 18846 4140
rect 19981 4131 20039 4137
rect 19981 4128 19993 4131
rect 18840 4100 19993 4128
rect 18840 4088 18846 4100
rect 19981 4097 19993 4100
rect 20027 4097 20039 4131
rect 19981 4091 20039 4097
rect 20349 4131 20407 4137
rect 20349 4097 20361 4131
rect 20395 4128 20407 4131
rect 20714 4128 20720 4140
rect 20395 4100 20720 4128
rect 20395 4097 20407 4100
rect 20349 4091 20407 4097
rect 20714 4088 20720 4100
rect 20772 4088 20778 4140
rect 20806 4088 20812 4140
rect 20864 4128 20870 4140
rect 20864 4100 20909 4128
rect 20864 4088 20870 4100
rect 20990 4088 20996 4140
rect 21048 4128 21054 4140
rect 21085 4131 21143 4137
rect 21085 4128 21097 4131
rect 21048 4100 21097 4128
rect 21048 4088 21054 4100
rect 21085 4097 21097 4100
rect 21131 4097 21143 4131
rect 21085 4091 21143 4097
rect 22462 4088 22468 4140
rect 22520 4128 22526 4140
rect 22833 4131 22891 4137
rect 22833 4128 22845 4131
rect 22520 4100 22845 4128
rect 22520 4088 22526 4100
rect 22833 4097 22845 4100
rect 22879 4097 22891 4131
rect 23750 4128 23756 4140
rect 22833 4091 22891 4097
rect 23308 4100 23756 4128
rect 16889 4073 16947 4079
rect 15252 4032 15700 4060
rect 15252 4020 15258 4032
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 16393 4063 16451 4069
rect 16393 4060 16405 4063
rect 16264 4032 16405 4060
rect 16264 4020 16270 4032
rect 16393 4029 16405 4032
rect 16439 4029 16451 4063
rect 16393 4023 16451 4029
rect 16482 4020 16488 4072
rect 16540 4020 16546 4072
rect 17129 4063 17187 4069
rect 17129 4029 17141 4063
rect 17175 4060 17187 4063
rect 17770 4060 17776 4072
rect 17175 4032 17776 4060
rect 17175 4029 17187 4032
rect 17129 4023 17187 4029
rect 17770 4020 17776 4032
rect 17828 4020 17834 4072
rect 18690 4020 18696 4072
rect 18748 4060 18754 4072
rect 19797 4063 19855 4069
rect 19797 4060 19809 4063
rect 18748 4032 19104 4060
rect 18748 4020 18754 4032
rect 9398 3952 9404 4004
rect 9456 3992 9462 4004
rect 9861 3995 9919 4001
rect 9861 3992 9873 3995
rect 9456 3964 9873 3992
rect 9456 3952 9462 3964
rect 9861 3961 9873 3964
rect 9907 3961 9919 3995
rect 9861 3955 9919 3961
rect 12437 3995 12495 4001
rect 12437 3961 12449 3995
rect 12483 3992 12495 3995
rect 12894 3992 12900 4004
rect 12483 3964 12900 3992
rect 12483 3961 12495 3964
rect 12437 3955 12495 3961
rect 9766 3924 9772 3936
rect 9324 3896 9772 3924
rect 9125 3887 9183 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 9876 3924 9904 3955
rect 12894 3952 12900 3964
rect 12952 3952 12958 4004
rect 12989 3995 13047 4001
rect 12989 3961 13001 3995
rect 13035 3992 13047 3995
rect 13035 3964 14326 3992
rect 13035 3961 13047 3964
rect 12989 3955 13047 3961
rect 10603 3927 10661 3933
rect 10603 3924 10615 3927
rect 9876 3896 10615 3924
rect 10603 3893 10615 3896
rect 10649 3924 10661 3927
rect 11238 3924 11244 3936
rect 10649 3896 11244 3924
rect 10649 3893 10661 3896
rect 10603 3887 10661 3893
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 12529 3927 12587 3933
rect 12529 3924 12541 3927
rect 11388 3896 12541 3924
rect 11388 3884 11394 3896
rect 12529 3893 12541 3896
rect 12575 3893 12587 3927
rect 14298 3924 14326 3964
rect 16298 3952 16304 4004
rect 16356 3952 16362 4004
rect 16390 3924 16396 3936
rect 14298 3896 16396 3924
rect 12529 3887 12587 3893
rect 16390 3884 16396 3896
rect 16448 3884 16454 3936
rect 16500 3924 16528 4020
rect 18874 3952 18880 4004
rect 18932 3992 18938 4004
rect 18969 3995 19027 4001
rect 18969 3992 18981 3995
rect 18932 3964 18981 3992
rect 18932 3952 18938 3964
rect 18969 3961 18981 3964
rect 19015 3961 19027 3995
rect 18969 3955 19027 3961
rect 16666 3924 16672 3936
rect 16500 3896 16672 3924
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 16859 3927 16917 3933
rect 16859 3924 16871 3927
rect 16816 3896 16871 3924
rect 16816 3884 16822 3896
rect 16859 3893 16871 3896
rect 16905 3893 16917 3927
rect 19076 3924 19104 4032
rect 19536 4032 19809 4060
rect 19242 3952 19248 4004
rect 19300 3992 19306 4004
rect 19337 3995 19395 4001
rect 19337 3992 19349 3995
rect 19300 3964 19349 3992
rect 19300 3952 19306 3964
rect 19337 3961 19349 3964
rect 19383 3961 19395 3995
rect 19337 3955 19395 3961
rect 19536 3924 19564 4032
rect 19797 4029 19809 4032
rect 19843 4060 19855 4063
rect 19886 4060 19892 4072
rect 19843 4032 19892 4060
rect 19843 4029 19855 4032
rect 19797 4023 19855 4029
rect 19886 4020 19892 4032
rect 19944 4020 19950 4072
rect 21174 4020 21180 4072
rect 21232 4060 21238 4072
rect 22649 4063 22707 4069
rect 21232 4032 21791 4060
rect 21232 4020 21238 4032
rect 21763 3992 21791 4032
rect 22649 4029 22661 4063
rect 22695 4060 22707 4063
rect 23308 4060 23336 4100
rect 23750 4088 23756 4100
rect 23808 4088 23814 4140
rect 24995 4131 25053 4137
rect 24412 4100 24900 4128
rect 22695 4032 23336 4060
rect 23385 4063 23443 4069
rect 22695 4029 22707 4032
rect 22649 4023 22707 4029
rect 23385 4029 23397 4063
rect 23431 4060 23443 4063
rect 23566 4060 23572 4072
rect 23431 4032 23572 4060
rect 23431 4029 23443 4032
rect 23385 4023 23443 4029
rect 23400 3992 23428 4023
rect 23566 4020 23572 4032
rect 23624 4020 23630 4072
rect 23661 4063 23719 4069
rect 23661 4029 23673 4063
rect 23707 4060 23719 4063
rect 24412 4060 24440 4100
rect 23707 4032 24440 4060
rect 24489 4063 24547 4069
rect 23707 4029 23719 4032
rect 23661 4023 23719 4029
rect 24489 4029 24501 4063
rect 24535 4060 24547 4063
rect 24762 4060 24768 4072
rect 24535 4032 24768 4060
rect 24535 4029 24547 4032
rect 24489 4023 24547 4029
rect 24762 4020 24768 4032
rect 24820 4020 24826 4072
rect 24872 4060 24900 4100
rect 24995 4097 25007 4131
rect 25041 4128 25053 4131
rect 25866 4128 25872 4140
rect 25041 4100 25872 4128
rect 25041 4097 25053 4100
rect 24995 4091 25053 4097
rect 25866 4088 25872 4100
rect 25924 4088 25930 4140
rect 26418 4088 26424 4140
rect 26476 4088 26482 4140
rect 26510 4088 26516 4140
rect 26568 4128 26574 4140
rect 27024 4131 27082 4137
rect 27246 4135 27252 4140
rect 27024 4128 27036 4131
rect 26568 4100 27036 4128
rect 26568 4088 26574 4100
rect 27024 4097 27036 4100
rect 27070 4097 27082 4131
rect 27024 4091 27082 4097
rect 27193 4129 27252 4135
rect 27193 4095 27205 4129
rect 27239 4095 27252 4129
rect 27193 4089 27252 4095
rect 27246 4088 27252 4089
rect 27304 4088 27310 4140
rect 27433 4131 27491 4137
rect 27433 4097 27445 4131
rect 27479 4128 27491 4131
rect 30374 4128 30380 4140
rect 27479 4100 30380 4128
rect 27479 4097 27491 4100
rect 27433 4091 27491 4097
rect 30374 4088 30380 4100
rect 30432 4088 30438 4140
rect 25130 4060 25136 4072
rect 24872 4032 25136 4060
rect 25130 4020 25136 4032
rect 25188 4020 25194 4072
rect 25225 4063 25283 4069
rect 25225 4029 25237 4063
rect 25271 4060 25283 4063
rect 26436 4060 26464 4088
rect 25271 4032 26464 4060
rect 26697 4063 26755 4069
rect 25271 4029 25283 4032
rect 25225 4023 25283 4029
rect 26697 4029 26709 4063
rect 26743 4060 26755 4063
rect 26786 4060 26792 4072
rect 26743 4032 26792 4060
rect 26743 4029 26755 4032
rect 26697 4023 26755 4029
rect 26786 4020 26792 4032
rect 26844 4020 26850 4072
rect 28997 4063 29055 4069
rect 28997 4029 29009 4063
rect 29043 4060 29055 4063
rect 29178 4060 29184 4072
rect 29043 4032 29184 4060
rect 29043 4029 29055 4032
rect 28997 4023 29055 4029
rect 29178 4020 29184 4032
rect 29236 4020 29242 4072
rect 24394 3992 24400 4004
rect 21763 3964 23428 3992
rect 23492 3964 24400 3992
rect 19076 3896 19564 3924
rect 19613 3927 19671 3933
rect 16859 3887 16917 3893
rect 19613 3893 19625 3927
rect 19659 3924 19671 3927
rect 19794 3924 19800 3936
rect 19659 3896 19800 3924
rect 19659 3893 19671 3896
rect 19613 3887 19671 3893
rect 19794 3884 19800 3896
rect 19852 3884 19858 3936
rect 20815 3927 20873 3933
rect 20815 3893 20827 3927
rect 20861 3924 20873 3927
rect 21542 3924 21548 3936
rect 20861 3896 21548 3924
rect 20861 3893 20873 3896
rect 20815 3887 20873 3893
rect 21542 3884 21548 3896
rect 21600 3884 21606 3936
rect 22373 3927 22431 3933
rect 22373 3893 22385 3927
rect 22419 3924 22431 3927
rect 22462 3924 22468 3936
rect 22419 3896 22468 3924
rect 22419 3893 22431 3896
rect 22373 3887 22431 3893
rect 22462 3884 22468 3896
rect 22520 3884 22526 3936
rect 23014 3884 23020 3936
rect 23072 3924 23078 3936
rect 23492 3933 23520 3964
rect 24394 3952 24400 3964
rect 24452 3952 24458 4004
rect 29086 3952 29092 4004
rect 29144 3992 29150 4004
rect 29144 3964 29224 3992
rect 29144 3952 29150 3964
rect 23201 3927 23259 3933
rect 23201 3924 23213 3927
rect 23072 3896 23213 3924
rect 23072 3884 23078 3896
rect 23201 3893 23213 3896
rect 23247 3893 23259 3927
rect 23201 3887 23259 3893
rect 23477 3927 23535 3933
rect 23477 3893 23489 3927
rect 23523 3893 23535 3927
rect 23477 3887 23535 3893
rect 23658 3884 23664 3936
rect 23716 3924 23722 3936
rect 24029 3927 24087 3933
rect 24029 3924 24041 3927
rect 23716 3896 24041 3924
rect 23716 3884 23722 3896
rect 24029 3893 24041 3896
rect 24075 3893 24087 3927
rect 24029 3887 24087 3893
rect 24955 3927 25013 3933
rect 24955 3893 24967 3927
rect 25001 3924 25013 3927
rect 26050 3924 26056 3936
rect 25001 3896 26056 3924
rect 25001 3893 25013 3896
rect 24955 3887 25013 3893
rect 26050 3884 26056 3896
rect 26108 3884 26114 3936
rect 26510 3884 26516 3936
rect 26568 3884 26574 3936
rect 28074 3884 28080 3936
rect 28132 3924 28138 3936
rect 29196 3933 29224 3964
rect 28537 3927 28595 3933
rect 28537 3924 28549 3927
rect 28132 3896 28549 3924
rect 28132 3884 28138 3896
rect 28537 3893 28549 3896
rect 28583 3893 28595 3927
rect 28537 3887 28595 3893
rect 29181 3927 29239 3933
rect 29181 3893 29193 3927
rect 29227 3893 29239 3927
rect 29181 3887 29239 3893
rect 29454 3884 29460 3936
rect 29512 3924 29518 3936
rect 30193 3927 30251 3933
rect 30193 3924 30205 3927
rect 29512 3896 30205 3924
rect 29512 3884 29518 3896
rect 30193 3893 30205 3896
rect 30239 3893 30251 3927
rect 30193 3887 30251 3893
rect 552 3834 31072 3856
rect 552 3782 7988 3834
rect 8040 3782 8052 3834
rect 8104 3782 8116 3834
rect 8168 3782 8180 3834
rect 8232 3782 8244 3834
rect 8296 3782 15578 3834
rect 15630 3782 15642 3834
rect 15694 3782 15706 3834
rect 15758 3782 15770 3834
rect 15822 3782 15834 3834
rect 15886 3782 23168 3834
rect 23220 3782 23232 3834
rect 23284 3782 23296 3834
rect 23348 3782 23360 3834
rect 23412 3782 23424 3834
rect 23476 3782 30758 3834
rect 30810 3782 30822 3834
rect 30874 3782 30886 3834
rect 30938 3782 30950 3834
rect 31002 3782 31014 3834
rect 31066 3782 31072 3834
rect 552 3760 31072 3782
rect 1029 3723 1087 3729
rect 1029 3689 1041 3723
rect 1075 3720 1087 3723
rect 3786 3720 3792 3732
rect 1075 3692 3792 3720
rect 1075 3689 1087 3692
rect 1029 3683 1087 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 3979 3723 4037 3729
rect 3979 3720 3991 3723
rect 3936 3692 3991 3720
rect 3936 3680 3942 3692
rect 3979 3689 3991 3692
rect 4025 3689 4037 3723
rect 3979 3683 4037 3689
rect 4338 3680 4344 3732
rect 4396 3720 4402 3732
rect 4396 3692 5764 3720
rect 4396 3680 4402 3692
rect 5736 3664 5764 3692
rect 5810 3680 5816 3732
rect 5868 3720 5874 3732
rect 6730 3720 6736 3732
rect 5868 3692 6736 3720
rect 5868 3680 5874 3692
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 7834 3680 7840 3732
rect 7892 3680 7898 3732
rect 8389 3723 8447 3729
rect 8389 3689 8401 3723
rect 8435 3720 8447 3723
rect 8570 3720 8576 3732
rect 8435 3692 8576 3720
rect 8435 3689 8447 3692
rect 8389 3683 8447 3689
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 9131 3723 9189 3729
rect 9131 3689 9143 3723
rect 9177 3720 9189 3723
rect 9398 3720 9404 3732
rect 9177 3692 9404 3720
rect 9177 3689 9189 3692
rect 9131 3683 9189 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 11606 3680 11612 3732
rect 11664 3720 11670 3732
rect 12075 3723 12133 3729
rect 12075 3720 12087 3723
rect 11664 3692 12087 3720
rect 11664 3680 11670 3692
rect 12075 3689 12087 3692
rect 12121 3689 12133 3723
rect 12075 3683 12133 3689
rect 16206 3680 16212 3732
rect 16264 3720 16270 3732
rect 16482 3720 16488 3732
rect 16264 3692 16488 3720
rect 16264 3680 16270 3692
rect 16482 3680 16488 3692
rect 16540 3680 16546 3732
rect 16583 3723 16641 3729
rect 16583 3689 16595 3723
rect 16629 3720 16641 3723
rect 16850 3720 16856 3732
rect 16629 3692 16856 3720
rect 16629 3689 16641 3692
rect 16583 3683 16641 3689
rect 16850 3680 16856 3692
rect 16908 3680 16914 3732
rect 20349 3723 20407 3729
rect 17512 3692 20300 3720
rect 5718 3612 5724 3664
rect 5776 3612 5782 3664
rect 1670 3593 1676 3596
rect 1213 3587 1271 3593
rect 1213 3553 1225 3587
rect 1259 3553 1271 3587
rect 1213 3547 1271 3553
rect 1632 3587 1676 3593
rect 1632 3553 1644 3587
rect 1632 3547 1676 3553
rect 1026 3476 1032 3528
rect 1084 3516 1090 3528
rect 1228 3516 1256 3547
rect 1670 3544 1676 3547
rect 1728 3544 1734 3596
rect 3528 3584 3648 3588
rect 7852 3584 7880 3680
rect 8113 3655 8171 3661
rect 8113 3621 8125 3655
rect 8159 3652 8171 3655
rect 8478 3652 8484 3664
rect 8159 3624 8484 3652
rect 8159 3621 8171 3624
rect 8113 3615 8171 3621
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 10781 3655 10839 3661
rect 10781 3621 10793 3655
rect 10827 3652 10839 3655
rect 10827 3624 11744 3652
rect 10827 3621 10839 3624
rect 10781 3615 10839 3621
rect 1826 3560 7880 3584
rect 1826 3556 3556 3560
rect 3620 3556 7880 3560
rect 8573 3587 8631 3593
rect 1826 3525 1854 3556
rect 8573 3553 8585 3587
rect 8619 3553 8631 3587
rect 8573 3547 8631 3553
rect 1084 3488 1256 3516
rect 1305 3519 1363 3525
rect 1084 3476 1090 3488
rect 1305 3485 1317 3519
rect 1351 3485 1363 3519
rect 1305 3479 1363 3485
rect 1811 3519 1869 3525
rect 1811 3485 1823 3519
rect 1857 3485 1869 3519
rect 1811 3479 1869 3485
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3516 2099 3519
rect 2406 3516 2412 3528
rect 2087 3488 2412 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 1326 3380 1354 3479
rect 2406 3476 2412 3488
rect 2464 3476 2470 3528
rect 3510 3516 3516 3528
rect 2700 3488 3516 3516
rect 2700 3380 2728 3488
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 3970 3476 3976 3528
rect 4028 3476 4034 3528
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 4890 3516 4896 3528
rect 4295 3488 4896 3516
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 6362 3525 6368 3528
rect 5997 3519 6055 3525
rect 5997 3516 6009 3519
rect 5316 3488 6009 3516
rect 5316 3476 5322 3488
rect 5997 3485 6009 3488
rect 6043 3485 6055 3519
rect 5997 3479 6055 3485
rect 6324 3519 6368 3525
rect 6324 3485 6336 3519
rect 6324 3479 6368 3485
rect 6362 3476 6368 3479
rect 6420 3476 6426 3528
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6512 3488 6557 3516
rect 6512 3476 6518 3488
rect 6730 3476 6736 3528
rect 6788 3476 6794 3528
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 8588 3516 8616 3547
rect 8938 3544 8944 3596
rect 8996 3584 9002 3596
rect 9401 3587 9459 3593
rect 8996 3556 9352 3584
rect 8996 3544 9002 3556
rect 6972 3488 8616 3516
rect 8665 3519 8723 3525
rect 6972 3476 6978 3488
rect 8665 3485 8677 3519
rect 8711 3516 8723 3519
rect 9030 3516 9036 3528
rect 8711 3488 9036 3516
rect 8711 3485 8723 3488
rect 8665 3479 8723 3485
rect 9030 3476 9036 3488
rect 9088 3476 9094 3528
rect 9214 3525 9220 3528
rect 9171 3519 9220 3525
rect 9171 3485 9183 3519
rect 9217 3485 9220 3519
rect 9171 3479 9220 3485
rect 9214 3476 9220 3479
rect 9272 3476 9278 3528
rect 9324 3516 9352 3556
rect 9401 3553 9413 3587
rect 9447 3584 9459 3587
rect 9490 3584 9496 3596
rect 9447 3556 9496 3584
rect 9447 3553 9459 3556
rect 9401 3547 9459 3553
rect 9490 3544 9496 3556
rect 9548 3544 9554 3596
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3584 11115 3587
rect 11238 3584 11244 3596
rect 11103 3556 11244 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 11072 3516 11100 3547
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 11422 3544 11428 3596
rect 11480 3584 11486 3596
rect 11609 3587 11667 3593
rect 11609 3584 11621 3587
rect 11480 3556 11621 3584
rect 11480 3544 11486 3556
rect 11609 3553 11621 3556
rect 11655 3553 11667 3587
rect 11609 3547 11667 3553
rect 9324 3488 11100 3516
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3485 11391 3519
rect 11716 3516 11744 3624
rect 12158 3544 12164 3596
rect 12216 3584 12222 3596
rect 12345 3587 12403 3593
rect 12345 3584 12357 3587
rect 12216 3556 12357 3584
rect 12216 3544 12222 3556
rect 12345 3553 12357 3556
rect 12391 3553 12403 3587
rect 12345 3547 12403 3553
rect 13725 3587 13783 3593
rect 13725 3553 13737 3587
rect 13771 3584 13783 3587
rect 15933 3587 15991 3593
rect 13771 3556 14323 3584
rect 13771 3553 13783 3556
rect 13725 3547 13783 3553
rect 12072 3519 12130 3525
rect 12072 3516 12084 3519
rect 11716 3488 12084 3516
rect 11333 3479 11391 3485
rect 12072 3485 12084 3488
rect 12118 3485 12130 3519
rect 12072 3479 12130 3485
rect 5810 3448 5816 3460
rect 5460 3420 5816 3448
rect 1326 3352 2728 3380
rect 3329 3383 3387 3389
rect 3329 3349 3341 3383
rect 3375 3380 3387 3383
rect 5460 3380 5488 3420
rect 5810 3408 5816 3420
rect 5868 3408 5874 3460
rect 3375 3352 5488 3380
rect 5537 3383 5595 3389
rect 3375 3349 3387 3352
rect 3329 3343 3387 3349
rect 5537 3349 5549 3383
rect 5583 3380 5595 3383
rect 6454 3380 6460 3392
rect 5583 3352 6460 3380
rect 5583 3349 5595 3352
rect 5537 3343 5595 3349
rect 6454 3340 6460 3352
rect 6512 3340 6518 3392
rect 11348 3380 11376 3479
rect 13814 3476 13820 3528
rect 13872 3476 13878 3528
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14295 3527 14323 3556
rect 15933 3553 15945 3587
rect 15979 3584 15991 3587
rect 15979 3556 16623 3584
rect 15979 3553 15991 3556
rect 15933 3547 15991 3553
rect 14144 3519 14202 3525
rect 14144 3516 14156 3519
rect 14056 3488 14156 3516
rect 14056 3476 14062 3488
rect 14144 3485 14156 3488
rect 14190 3485 14202 3519
rect 14144 3479 14202 3485
rect 14280 3521 14338 3527
rect 14280 3487 14292 3521
rect 14326 3487 14338 3521
rect 14280 3481 14338 3487
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 14553 3519 14611 3525
rect 14553 3516 14565 3519
rect 14424 3488 14565 3516
rect 14424 3476 14430 3488
rect 14553 3485 14565 3488
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 16117 3519 16175 3525
rect 16117 3485 16129 3519
rect 16163 3516 16175 3519
rect 16390 3516 16396 3528
rect 16163 3488 16396 3516
rect 16163 3485 16175 3488
rect 16117 3479 16175 3485
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 16595 3527 16623 3556
rect 16666 3544 16672 3596
rect 16724 3584 16730 3596
rect 17512 3584 17540 3692
rect 20272 3652 20300 3692
rect 20349 3689 20361 3723
rect 20395 3720 20407 3723
rect 20806 3720 20812 3732
rect 20395 3692 20812 3720
rect 20395 3689 20407 3692
rect 20349 3683 20407 3689
rect 20806 3680 20812 3692
rect 20864 3680 20870 3732
rect 21082 3680 21088 3732
rect 21140 3680 21146 3732
rect 22554 3680 22560 3732
rect 22612 3720 22618 3732
rect 22747 3723 22805 3729
rect 22747 3720 22759 3723
rect 22612 3692 22759 3720
rect 22612 3680 22618 3692
rect 22747 3689 22759 3692
rect 22793 3720 22805 3723
rect 24210 3720 24216 3732
rect 22793 3692 24216 3720
rect 22793 3689 22805 3692
rect 22747 3683 22805 3689
rect 24210 3680 24216 3692
rect 24268 3680 24274 3732
rect 24854 3680 24860 3732
rect 24912 3720 24918 3732
rect 26053 3723 26111 3729
rect 26053 3720 26065 3723
rect 24912 3692 26065 3720
rect 24912 3680 24918 3692
rect 26053 3689 26065 3692
rect 26099 3689 26111 3723
rect 26053 3683 26111 3689
rect 26142 3680 26148 3732
rect 26200 3720 26206 3732
rect 29178 3720 29184 3732
rect 26200 3692 26740 3720
rect 26200 3680 26206 3692
rect 21100 3652 21128 3680
rect 20272 3624 21128 3652
rect 21542 3612 21548 3664
rect 21600 3612 21606 3664
rect 24302 3612 24308 3664
rect 24360 3652 24366 3664
rect 25041 3655 25099 3661
rect 25041 3652 25053 3655
rect 24360 3624 25053 3652
rect 24360 3612 24366 3624
rect 25041 3621 25053 3624
rect 25087 3621 25099 3655
rect 25041 3615 25099 3621
rect 16724 3556 17540 3584
rect 18233 3587 18291 3593
rect 16724 3544 16730 3556
rect 18233 3553 18245 3587
rect 18279 3584 18291 3587
rect 18279 3556 18831 3584
rect 18279 3553 18291 3556
rect 18233 3547 18291 3553
rect 16580 3521 16638 3527
rect 16580 3487 16592 3521
rect 16626 3487 16638 3521
rect 16580 3481 16638 3487
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3516 16911 3519
rect 17954 3516 17960 3528
rect 16899 3488 17960 3516
rect 16899 3485 16911 3488
rect 16853 3479 16911 3485
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 18322 3476 18328 3528
rect 18380 3476 18386 3528
rect 18690 3525 18696 3528
rect 18652 3519 18696 3525
rect 18652 3485 18664 3519
rect 18652 3479 18696 3485
rect 18690 3476 18696 3479
rect 18748 3476 18754 3528
rect 18803 3527 18831 3556
rect 19058 3544 19064 3596
rect 19116 3544 19122 3596
rect 19886 3544 19892 3596
rect 19944 3544 19950 3596
rect 20625 3587 20683 3593
rect 20625 3553 20637 3587
rect 20671 3584 20683 3587
rect 20714 3584 20720 3596
rect 20671 3556 20720 3584
rect 20671 3553 20683 3556
rect 20625 3547 20683 3553
rect 20714 3544 20720 3556
rect 20772 3544 20778 3596
rect 21269 3587 21327 3593
rect 21269 3553 21281 3587
rect 21315 3553 21327 3587
rect 21269 3547 21327 3553
rect 22005 3587 22063 3593
rect 22005 3553 22017 3587
rect 22051 3553 22063 3587
rect 22005 3547 22063 3553
rect 18788 3521 18846 3527
rect 18788 3487 18800 3521
rect 18834 3487 18846 3521
rect 19904 3516 19932 3544
rect 21284 3516 21312 3547
rect 19904 3488 21312 3516
rect 18788 3481 18846 3487
rect 21358 3476 21364 3528
rect 21416 3516 21422 3528
rect 21726 3516 21732 3528
rect 21416 3488 21732 3516
rect 21416 3476 21422 3488
rect 21726 3476 21732 3488
rect 21784 3516 21790 3528
rect 22020 3516 22048 3547
rect 22186 3544 22192 3596
rect 22244 3584 22250 3596
rect 22281 3587 22339 3593
rect 22281 3584 22293 3587
rect 22244 3556 22293 3584
rect 22244 3544 22250 3556
rect 22281 3553 22293 3556
rect 22327 3553 22339 3587
rect 22281 3547 22339 3553
rect 23014 3544 23020 3596
rect 23072 3544 23078 3596
rect 23750 3544 23756 3596
rect 23808 3584 23814 3596
rect 24765 3587 24823 3593
rect 24765 3584 24777 3587
rect 23808 3556 24777 3584
rect 23808 3544 23814 3556
rect 24765 3553 24777 3556
rect 24811 3553 24823 3587
rect 24765 3547 24823 3553
rect 25501 3587 25559 3593
rect 25501 3553 25513 3587
rect 25547 3553 25559 3587
rect 25501 3547 25559 3553
rect 21784 3488 22048 3516
rect 21784 3476 21790 3488
rect 22462 3476 22468 3528
rect 22520 3516 22526 3528
rect 22744 3521 22802 3527
rect 22744 3516 22756 3521
rect 22520 3488 22756 3516
rect 22520 3476 22526 3488
rect 22744 3487 22756 3488
rect 22790 3487 22802 3521
rect 22744 3481 22802 3487
rect 23474 3476 23480 3528
rect 23532 3516 23538 3528
rect 25516 3516 25544 3547
rect 25682 3544 25688 3596
rect 25740 3584 25746 3596
rect 26712 3593 26740 3692
rect 27448 3692 29184 3720
rect 26878 3612 26884 3664
rect 26936 3652 26942 3664
rect 26973 3655 27031 3661
rect 26973 3652 26985 3655
rect 26936 3624 26985 3652
rect 26936 3612 26942 3624
rect 26973 3621 26985 3624
rect 27019 3621 27031 3655
rect 26973 3615 27031 3621
rect 25777 3587 25835 3593
rect 25777 3584 25789 3587
rect 25740 3556 25789 3584
rect 25740 3544 25746 3556
rect 25777 3553 25789 3556
rect 25823 3553 25835 3587
rect 25777 3547 25835 3553
rect 26605 3587 26663 3593
rect 26605 3553 26617 3587
rect 26651 3553 26663 3587
rect 26605 3547 26663 3553
rect 26697 3587 26755 3593
rect 26697 3553 26709 3587
rect 26743 3584 26755 3587
rect 27341 3587 27399 3593
rect 27341 3584 27353 3587
rect 26743 3556 27353 3584
rect 26743 3553 26755 3556
rect 26697 3547 26755 3553
rect 27341 3553 27353 3556
rect 27387 3553 27399 3587
rect 27341 3547 27399 3553
rect 26620 3516 26648 3547
rect 27448 3516 27476 3692
rect 29178 3680 29184 3692
rect 29236 3680 29242 3732
rect 29822 3680 29828 3732
rect 29880 3680 29886 3732
rect 27890 3544 27896 3596
rect 27948 3584 27954 3596
rect 27985 3587 28043 3593
rect 27985 3584 27997 3587
rect 27948 3556 27997 3584
rect 27948 3544 27954 3556
rect 27985 3553 27997 3556
rect 28031 3553 28043 3587
rect 27985 3547 28043 3553
rect 28721 3587 28779 3593
rect 28721 3553 28733 3587
rect 28767 3584 28779 3587
rect 28810 3584 28816 3596
rect 28767 3556 28816 3584
rect 28767 3553 28779 3556
rect 28721 3547 28779 3553
rect 28810 3544 28816 3556
rect 28868 3544 28874 3596
rect 30098 3584 30104 3596
rect 29012 3556 30104 3584
rect 23532 3488 27476 3516
rect 23532 3476 23538 3488
rect 27614 3476 27620 3528
rect 27672 3476 27678 3528
rect 28166 3476 28172 3528
rect 28224 3516 28230 3528
rect 28312 3519 28370 3525
rect 28312 3516 28324 3519
rect 28224 3488 28324 3516
rect 28224 3476 28230 3488
rect 28312 3485 28324 3488
rect 28358 3485 28370 3519
rect 28312 3479 28370 3485
rect 28442 3476 28448 3528
rect 28500 3476 28506 3528
rect 28534 3476 28540 3528
rect 28592 3516 28598 3528
rect 29012 3516 29040 3556
rect 30098 3544 30104 3556
rect 30156 3544 30162 3596
rect 28592 3488 29040 3516
rect 28592 3476 28598 3488
rect 29086 3476 29092 3528
rect 29144 3516 29150 3528
rect 30377 3519 30435 3525
rect 30377 3516 30389 3519
rect 29144 3488 30389 3516
rect 29144 3476 29150 3488
rect 30377 3485 30389 3488
rect 30423 3485 30435 3519
rect 30377 3479 30435 3485
rect 13998 3380 14004 3392
rect 11348 3352 14004 3380
rect 13998 3340 14004 3352
rect 14056 3380 14062 3392
rect 14458 3380 14464 3392
rect 14056 3352 14464 3380
rect 14056 3340 14062 3352
rect 14458 3340 14464 3352
rect 14516 3340 14522 3392
rect 15930 3340 15936 3392
rect 15988 3380 15994 3392
rect 18046 3380 18052 3392
rect 15988 3352 18052 3380
rect 15988 3340 15994 3352
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 18340 3380 18368 3476
rect 19886 3408 19892 3460
rect 19944 3448 19950 3460
rect 26421 3451 26479 3457
rect 26421 3448 26433 3451
rect 19944 3420 22094 3448
rect 19944 3408 19950 3420
rect 19242 3380 19248 3392
rect 18340 3352 19248 3380
rect 19242 3340 19248 3352
rect 19300 3380 19306 3392
rect 20717 3383 20775 3389
rect 20717 3380 20729 3383
rect 19300 3352 20729 3380
rect 19300 3340 19306 3352
rect 20717 3349 20729 3352
rect 20763 3349 20775 3383
rect 20717 3343 20775 3349
rect 21818 3340 21824 3392
rect 21876 3340 21882 3392
rect 22066 3380 22094 3420
rect 23676 3420 26433 3448
rect 23676 3380 23704 3420
rect 26421 3417 26433 3420
rect 26467 3417 26479 3451
rect 26421 3411 26479 3417
rect 22066 3352 23704 3380
rect 24305 3383 24363 3389
rect 24305 3349 24317 3383
rect 24351 3380 24363 3383
rect 24578 3380 24584 3392
rect 24351 3352 24584 3380
rect 24351 3349 24363 3352
rect 24305 3343 24363 3349
rect 24578 3340 24584 3352
rect 24636 3340 24642 3392
rect 25314 3340 25320 3392
rect 25372 3340 25378 3392
rect 25590 3340 25596 3392
rect 25648 3340 25654 3392
rect 25682 3340 25688 3392
rect 25740 3380 25746 3392
rect 29546 3380 29552 3392
rect 25740 3352 29552 3380
rect 25740 3340 25746 3352
rect 29546 3340 29552 3352
rect 29604 3340 29610 3392
rect 552 3290 30912 3312
rect 552 3238 4193 3290
rect 4245 3238 4257 3290
rect 4309 3238 4321 3290
rect 4373 3238 4385 3290
rect 4437 3238 4449 3290
rect 4501 3238 11783 3290
rect 11835 3238 11847 3290
rect 11899 3238 11911 3290
rect 11963 3238 11975 3290
rect 12027 3238 12039 3290
rect 12091 3238 19373 3290
rect 19425 3238 19437 3290
rect 19489 3238 19501 3290
rect 19553 3238 19565 3290
rect 19617 3238 19629 3290
rect 19681 3238 26963 3290
rect 27015 3238 27027 3290
rect 27079 3238 27091 3290
rect 27143 3238 27155 3290
rect 27207 3238 27219 3290
rect 27271 3238 30912 3290
rect 552 3216 30912 3238
rect 3234 3136 3240 3188
rect 3292 3136 3298 3188
rect 5626 3176 5632 3188
rect 3620 3148 5632 3176
rect 3620 3117 3648 3148
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 5718 3136 5724 3188
rect 5776 3136 5782 3188
rect 8113 3179 8171 3185
rect 8113 3145 8125 3179
rect 8159 3176 8171 3179
rect 9214 3176 9220 3188
rect 8159 3148 9220 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 9674 3136 9680 3188
rect 9732 3176 9738 3188
rect 15930 3176 15936 3188
rect 9732 3148 15936 3176
rect 9732 3136 9738 3148
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 16390 3176 16396 3188
rect 16040 3148 16396 3176
rect 3605 3111 3663 3117
rect 3605 3077 3617 3111
rect 3651 3077 3663 3111
rect 3605 3071 3663 3077
rect 5810 3068 5816 3120
rect 5868 3108 5874 3120
rect 5994 3108 6000 3120
rect 5868 3080 6000 3108
rect 5868 3068 5874 3080
rect 5994 3068 6000 3080
rect 6052 3068 6058 3120
rect 13170 3068 13176 3120
rect 13228 3068 13234 3120
rect 1443 3043 1501 3049
rect 1443 3009 1455 3043
rect 1489 3040 1501 3043
rect 4246 3040 4252 3052
rect 1489 3012 4252 3040
rect 1489 3009 1501 3012
rect 1443 3003 1501 3009
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 5534 3040 5540 3052
rect 4362 3025 5540 3040
rect 4362 2994 4389 3025
rect 4377 2991 4389 2994
rect 4423 3012 5540 3025
rect 4423 2991 4435 3012
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 6595 3041 6653 3047
rect 6595 3007 6607 3041
rect 6641 3040 6653 3041
rect 7650 3040 7656 3052
rect 6641 3012 7656 3040
rect 6641 3007 6653 3012
rect 6595 3001 6653 3007
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 9398 3049 9404 3052
rect 9360 3043 9404 3049
rect 7892 3012 9168 3040
rect 7892 3000 7898 3012
rect 4377 2985 4435 2991
rect 937 2975 995 2981
rect 937 2941 949 2975
rect 983 2972 995 2975
rect 1578 2972 1584 2984
rect 983 2944 1584 2972
rect 983 2941 995 2944
rect 937 2935 995 2941
rect 1578 2932 1584 2944
rect 1636 2932 1642 2984
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2972 1731 2975
rect 2130 2972 2136 2984
rect 1719 2944 2136 2972
rect 1719 2941 1731 2944
rect 1673 2935 1731 2941
rect 2130 2932 2136 2944
rect 2188 2932 2194 2984
rect 3421 2975 3479 2981
rect 3421 2941 3433 2975
rect 3467 2972 3479 2975
rect 3467 2944 3556 2972
rect 3467 2941 3479 2944
rect 3421 2935 3479 2941
rect 3528 2916 3556 2944
rect 3694 2932 3700 2984
rect 3752 2932 3758 2984
rect 3789 2975 3847 2981
rect 3789 2941 3801 2975
rect 3835 2941 3847 2975
rect 3789 2935 3847 2941
rect 3050 2864 3056 2916
rect 3108 2864 3114 2916
rect 3510 2864 3516 2916
rect 3568 2864 3574 2916
rect 1403 2839 1461 2845
rect 1403 2805 1415 2839
rect 1449 2836 1461 2839
rect 3712 2836 3740 2932
rect 3804 2904 3832 2935
rect 3878 2932 3884 2984
rect 3936 2932 3942 2984
rect 4614 2932 4620 2984
rect 4672 2932 4678 2984
rect 6086 2932 6092 2984
rect 6144 2932 6150 2984
rect 6178 2932 6184 2984
rect 6236 2972 6242 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6236 2944 6837 2972
rect 6236 2932 6242 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 8478 2972 8484 2984
rect 6825 2935 6883 2941
rect 7668 2944 8484 2972
rect 3804 2876 3924 2904
rect 3896 2848 3924 2876
rect 1449 2808 3740 2836
rect 1449 2805 1461 2808
rect 1403 2799 1461 2805
rect 3878 2796 3884 2848
rect 3936 2796 3942 2848
rect 4154 2796 4160 2848
rect 4212 2836 4218 2848
rect 4347 2839 4405 2845
rect 4347 2836 4359 2839
rect 4212 2808 4359 2836
rect 4212 2796 4218 2808
rect 4347 2805 4359 2808
rect 4393 2805 4405 2839
rect 4347 2799 4405 2805
rect 6546 2796 6552 2848
rect 6604 2845 6610 2848
rect 6604 2836 6613 2845
rect 7668 2836 7696 2944
rect 8478 2932 8484 2944
rect 8536 2972 8542 2984
rect 8662 2972 8668 2984
rect 8536 2944 8668 2972
rect 8536 2932 8542 2944
rect 8662 2932 8668 2944
rect 8720 2932 8726 2984
rect 9030 2972 9036 2984
rect 8772 2944 9036 2972
rect 8573 2907 8631 2913
rect 8573 2873 8585 2907
rect 8619 2904 8631 2907
rect 8772 2904 8800 2944
rect 9030 2932 9036 2944
rect 9088 2932 9094 2984
rect 9140 2972 9168 3012
rect 9360 3009 9372 3043
rect 9360 3003 9404 3009
rect 9398 3000 9404 3003
rect 9456 3000 9462 3052
rect 9582 3047 9588 3052
rect 9539 3041 9588 3047
rect 9539 3007 9551 3041
rect 9585 3007 9588 3041
rect 9539 3001 9588 3007
rect 9582 3000 9588 3001
rect 9640 3000 9646 3052
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 11704 3043 11762 3049
rect 11704 3040 11716 3043
rect 11195 3012 11716 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 11704 3009 11716 3012
rect 11750 3009 11762 3043
rect 11704 3003 11762 3009
rect 9769 2975 9827 2981
rect 9769 2972 9781 2975
rect 9140 2944 9781 2972
rect 9769 2941 9781 2944
rect 9815 2941 9827 2975
rect 9769 2935 9827 2941
rect 11241 2975 11299 2981
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 11330 2972 11336 2984
rect 11287 2944 11336 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 11514 2932 11520 2984
rect 11572 2972 11578 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11572 2944 11989 2972
rect 11572 2932 11578 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 13188 2972 13216 3068
rect 13357 3043 13415 3049
rect 13357 3009 13369 3043
rect 13403 3040 13415 3043
rect 14464 3043 14522 3049
rect 14464 3040 14476 3043
rect 13403 3012 14476 3040
rect 13403 3009 13415 3012
rect 13357 3003 13415 3009
rect 14464 3009 14476 3012
rect 14510 3009 14522 3043
rect 14464 3003 14522 3009
rect 16040 2984 16068 3148
rect 16390 3136 16396 3148
rect 16448 3176 16454 3188
rect 19794 3176 19800 3188
rect 16448 3148 19800 3176
rect 16448 3136 16454 3148
rect 19794 3136 19800 3148
rect 19852 3136 19858 3188
rect 21818 3176 21824 3188
rect 20640 3148 21824 3176
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3040 16175 3043
rect 16672 3043 16730 3049
rect 16672 3040 16684 3043
rect 16163 3012 16684 3040
rect 16163 3009 16175 3012
rect 16117 3003 16175 3009
rect 16672 3009 16684 3012
rect 16718 3009 16730 3043
rect 16672 3003 16730 3009
rect 18325 3043 18383 3049
rect 18325 3009 18337 3043
rect 18371 3040 18383 3043
rect 19156 3043 19214 3049
rect 19156 3040 19168 3043
rect 18371 3012 19168 3040
rect 18371 3009 18383 3012
rect 18325 3003 18383 3009
rect 19156 3009 19168 3012
rect 19202 3009 19214 3043
rect 19156 3003 19214 3009
rect 19242 3000 19248 3052
rect 19300 3000 19306 3052
rect 19334 3000 19340 3052
rect 19392 3000 19398 3052
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3040 19487 3043
rect 20640 3040 20668 3148
rect 21818 3136 21824 3148
rect 21876 3136 21882 3188
rect 22278 3136 22284 3188
rect 22336 3176 22342 3188
rect 23385 3179 23443 3185
rect 23385 3176 23397 3179
rect 22336 3148 23397 3176
rect 22336 3136 22342 3148
rect 23385 3145 23397 3148
rect 23431 3145 23443 3179
rect 23385 3139 23443 3145
rect 19475 3012 20668 3040
rect 19475 3009 19487 3012
rect 19429 3003 19487 3009
rect 20714 3000 20720 3052
rect 20772 3000 20778 3052
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 21364 3043 21422 3049
rect 21364 3040 21376 3043
rect 20855 3012 21376 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 21364 3009 21376 3012
rect 21410 3009 21422 3043
rect 21364 3003 21422 3009
rect 21450 3000 21456 3052
rect 21508 3040 21514 3052
rect 21637 3043 21695 3049
rect 21637 3040 21649 3043
rect 21508 3012 21649 3040
rect 21508 3000 21514 3012
rect 21637 3009 21649 3012
rect 21683 3009 21695 3043
rect 23400 3040 23428 3139
rect 23566 3136 23572 3188
rect 23624 3176 23630 3188
rect 23842 3176 23848 3188
rect 23624 3148 23848 3176
rect 23624 3136 23630 3148
rect 23842 3136 23848 3148
rect 23900 3176 23906 3188
rect 25774 3176 25780 3188
rect 23900 3148 25780 3176
rect 23900 3136 23906 3148
rect 25774 3136 25780 3148
rect 25832 3136 25838 3188
rect 28534 3176 28540 3188
rect 26068 3148 28540 3176
rect 26068 3108 26096 3148
rect 28534 3136 28540 3148
rect 28592 3136 28598 3188
rect 30190 3136 30196 3188
rect 30248 3136 30254 3188
rect 25240 3080 26096 3108
rect 25240 3052 25268 3080
rect 23842 3040 23848 3052
rect 23400 3012 23848 3040
rect 21637 3003 21695 3009
rect 23842 3000 23848 3012
rect 23900 3000 23906 3052
rect 24026 3000 24032 3052
rect 24084 3040 24090 3052
rect 24308 3043 24366 3049
rect 24308 3040 24320 3043
rect 24084 3012 24320 3040
rect 24084 3000 24090 3012
rect 24308 3009 24320 3012
rect 24354 3009 24366 3043
rect 24308 3003 24366 3009
rect 25222 3000 25228 3052
rect 25280 3000 25286 3052
rect 26326 3000 26332 3052
rect 26384 3040 26390 3052
rect 26516 3043 26574 3049
rect 26516 3040 26528 3043
rect 26384 3012 26528 3040
rect 26384 3000 26390 3012
rect 26516 3009 26528 3012
rect 26562 3009 26574 3043
rect 26516 3003 26574 3009
rect 26602 3000 26608 3052
rect 26660 3040 26666 3052
rect 26789 3043 26847 3049
rect 26789 3040 26801 3043
rect 26660 3012 26801 3040
rect 26660 3000 26666 3012
rect 26789 3009 26801 3012
rect 26835 3009 26847 3043
rect 26789 3003 26847 3009
rect 27706 3000 27712 3052
rect 27764 3040 27770 3052
rect 29273 3043 29331 3049
rect 29273 3040 29285 3043
rect 27764 3012 29285 3040
rect 27764 3000 27770 3012
rect 29273 3009 29285 3012
rect 29319 3009 29331 3043
rect 29273 3003 29331 3009
rect 29914 3000 29920 3052
rect 29972 3000 29978 3052
rect 13725 2975 13783 2981
rect 13725 2972 13737 2975
rect 13188 2944 13737 2972
rect 11977 2935 12035 2941
rect 13725 2941 13737 2944
rect 13771 2941 13783 2975
rect 13725 2935 13783 2941
rect 13906 2932 13912 2984
rect 13964 2972 13970 2984
rect 14001 2975 14059 2981
rect 14001 2972 14013 2975
rect 13964 2944 14013 2972
rect 13964 2932 13970 2944
rect 14001 2941 14013 2944
rect 14047 2941 14059 2975
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14001 2935 14059 2941
rect 14108 2944 14749 2972
rect 8619 2876 8800 2904
rect 8619 2873 8631 2876
rect 8573 2867 8631 2873
rect 13170 2864 13176 2916
rect 13228 2904 13234 2916
rect 14108 2904 14136 2944
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 14737 2935 14795 2941
rect 16022 2932 16028 2984
rect 16080 2972 16086 2984
rect 16209 2975 16267 2981
rect 16209 2972 16221 2975
rect 16080 2944 16221 2972
rect 16080 2932 16086 2944
rect 16209 2941 16221 2944
rect 16255 2941 16267 2975
rect 16945 2975 17003 2981
rect 16945 2972 16957 2975
rect 16209 2935 16267 2941
rect 16316 2944 16957 2972
rect 13228 2876 14136 2904
rect 13228 2864 13234 2876
rect 6604 2808 7696 2836
rect 6604 2799 6613 2808
rect 6604 2796 6610 2799
rect 7742 2796 7748 2848
rect 7800 2836 7806 2848
rect 8665 2839 8723 2845
rect 8665 2836 8677 2839
rect 7800 2808 8677 2836
rect 7800 2796 7806 2808
rect 8665 2805 8677 2808
rect 8711 2805 8723 2839
rect 8665 2799 8723 2805
rect 8938 2796 8944 2848
rect 8996 2836 9002 2848
rect 11330 2836 11336 2848
rect 8996 2808 11336 2836
rect 8996 2796 9002 2808
rect 11330 2796 11336 2808
rect 11388 2796 11394 2848
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 11707 2839 11765 2845
rect 11707 2836 11719 2839
rect 11664 2808 11719 2836
rect 11664 2796 11670 2808
rect 11707 2805 11719 2808
rect 11753 2805 11765 2839
rect 11707 2799 11765 2805
rect 13541 2839 13599 2845
rect 13541 2805 13553 2839
rect 13587 2836 13599 2839
rect 14366 2836 14372 2848
rect 13587 2808 14372 2836
rect 13587 2805 13599 2808
rect 13541 2799 13599 2805
rect 14366 2796 14372 2808
rect 14424 2796 14430 2848
rect 14458 2796 14464 2848
rect 14516 2845 14522 2848
rect 14516 2836 14525 2845
rect 14516 2808 14561 2836
rect 14516 2799 14525 2808
rect 14516 2796 14522 2799
rect 15102 2796 15108 2848
rect 15160 2836 15166 2848
rect 16316 2836 16344 2944
rect 16945 2941 16957 2944
rect 16991 2941 17003 2975
rect 16945 2935 17003 2941
rect 18506 2932 18512 2984
rect 18564 2972 18570 2984
rect 18693 2975 18751 2981
rect 18693 2972 18705 2975
rect 18564 2944 18705 2972
rect 18564 2932 18570 2944
rect 18693 2941 18705 2944
rect 18739 2972 18751 2975
rect 19260 2972 19288 3000
rect 18739 2944 19288 2972
rect 19352 2972 19380 3000
rect 20732 2972 20760 3000
rect 20901 2975 20959 2981
rect 20901 2972 20913 2975
rect 19352 2944 20116 2972
rect 20732 2944 20913 2972
rect 18739 2941 18751 2944
rect 18693 2935 18751 2941
rect 18782 2864 18788 2916
rect 18840 2864 18846 2916
rect 15160 2808 16344 2836
rect 16675 2839 16733 2845
rect 15160 2796 15166 2808
rect 16675 2805 16687 2839
rect 16721 2836 16733 2839
rect 16850 2836 16856 2848
rect 16721 2808 16856 2836
rect 16721 2805 16733 2808
rect 16675 2799 16733 2805
rect 16850 2796 16856 2808
rect 16908 2796 16914 2848
rect 18800 2836 18828 2864
rect 19159 2839 19217 2845
rect 19159 2836 19171 2839
rect 18800 2808 19171 2836
rect 19159 2805 19171 2808
rect 19205 2805 19217 2839
rect 20088 2836 20116 2944
rect 20901 2941 20913 2944
rect 20947 2941 20959 2975
rect 20901 2935 20959 2941
rect 21228 2975 21286 2981
rect 21228 2941 21240 2975
rect 21274 2972 21286 2975
rect 21542 2972 21548 2984
rect 21274 2944 21548 2972
rect 21274 2941 21286 2944
rect 21228 2935 21286 2941
rect 21542 2932 21548 2944
rect 21600 2932 21606 2984
rect 23658 2972 23664 2984
rect 22940 2944 23664 2972
rect 22940 2836 22968 2944
rect 23658 2932 23664 2944
rect 23716 2932 23722 2984
rect 24486 2932 24492 2984
rect 24544 2972 24550 2984
rect 24581 2975 24639 2981
rect 24581 2972 24593 2975
rect 24544 2944 24593 2972
rect 24544 2932 24550 2944
rect 24581 2941 24593 2944
rect 24627 2941 24639 2975
rect 24581 2935 24639 2941
rect 26053 2975 26111 2981
rect 26053 2941 26065 2975
rect 26099 2972 26111 2975
rect 26418 2972 26424 2984
rect 26099 2944 26424 2972
rect 26099 2941 26111 2944
rect 26053 2935 26111 2941
rect 26418 2932 26424 2944
rect 26476 2932 26482 2984
rect 28166 2932 28172 2984
rect 28224 2972 28230 2984
rect 28997 2975 29055 2981
rect 28997 2972 29009 2975
rect 28224 2944 29009 2972
rect 28224 2932 28230 2944
rect 28997 2941 29009 2944
rect 29043 2972 29055 2975
rect 29932 2972 29960 3000
rect 29043 2944 29960 2972
rect 29043 2941 29055 2944
rect 28997 2935 29055 2941
rect 23017 2907 23075 2913
rect 23017 2873 23029 2907
rect 23063 2873 23075 2907
rect 23017 2867 23075 2873
rect 23293 2907 23351 2913
rect 23293 2873 23305 2907
rect 23339 2904 23351 2907
rect 23566 2904 23572 2916
rect 23339 2876 23572 2904
rect 23339 2873 23351 2876
rect 23293 2867 23351 2873
rect 20088 2808 22968 2836
rect 23032 2836 23060 2867
rect 23566 2864 23572 2876
rect 23624 2864 23630 2916
rect 29914 2864 29920 2916
rect 29972 2904 29978 2916
rect 30374 2904 30380 2916
rect 29972 2876 30380 2904
rect 29972 2864 29978 2876
rect 30374 2864 30380 2876
rect 30432 2864 30438 2916
rect 23934 2836 23940 2848
rect 23032 2808 23940 2836
rect 19159 2799 19217 2805
rect 23934 2796 23940 2808
rect 23992 2796 23998 2848
rect 24210 2796 24216 2848
rect 24268 2836 24274 2848
rect 24311 2839 24369 2845
rect 24311 2836 24323 2839
rect 24268 2808 24323 2836
rect 24268 2796 24274 2808
rect 24311 2805 24323 2808
rect 24357 2805 24369 2839
rect 24311 2799 24369 2805
rect 24670 2796 24676 2848
rect 24728 2836 24734 2848
rect 25685 2839 25743 2845
rect 25685 2836 25697 2839
rect 24728 2808 25697 2836
rect 24728 2796 24734 2808
rect 25685 2805 25697 2808
rect 25731 2805 25743 2839
rect 25685 2799 25743 2805
rect 26050 2796 26056 2848
rect 26108 2836 26114 2848
rect 26519 2839 26577 2845
rect 26519 2836 26531 2839
rect 26108 2808 26531 2836
rect 26108 2796 26114 2808
rect 26519 2805 26531 2808
rect 26565 2836 26577 2839
rect 26878 2836 26884 2848
rect 26565 2808 26884 2836
rect 26565 2805 26577 2808
rect 26519 2799 26577 2805
rect 26878 2796 26884 2808
rect 26936 2796 26942 2848
rect 28074 2796 28080 2848
rect 28132 2796 28138 2848
rect 552 2746 31072 2768
rect 552 2694 7988 2746
rect 8040 2694 8052 2746
rect 8104 2694 8116 2746
rect 8168 2694 8180 2746
rect 8232 2694 8244 2746
rect 8296 2694 15578 2746
rect 15630 2694 15642 2746
rect 15694 2694 15706 2746
rect 15758 2694 15770 2746
rect 15822 2694 15834 2746
rect 15886 2694 23168 2746
rect 23220 2694 23232 2746
rect 23284 2694 23296 2746
rect 23348 2694 23360 2746
rect 23412 2694 23424 2746
rect 23476 2694 30758 2746
rect 30810 2694 30822 2746
rect 30874 2694 30886 2746
rect 30938 2694 30950 2746
rect 31002 2694 31014 2746
rect 31066 2694 31072 2746
rect 552 2672 31072 2694
rect 934 2592 940 2644
rect 992 2592 998 2644
rect 1762 2592 1768 2644
rect 1820 2641 1826 2644
rect 1820 2632 1829 2641
rect 3329 2635 3387 2641
rect 1820 2604 1865 2632
rect 1820 2595 1829 2604
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 3510 2632 3516 2644
rect 3375 2604 3516 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 1820 2592 1826 2595
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 3979 2635 4037 2641
rect 3979 2601 3991 2635
rect 4025 2632 4037 2635
rect 4154 2632 4160 2644
rect 4025 2604 4160 2632
rect 4025 2601 4037 2604
rect 3979 2595 4037 2601
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 5534 2592 5540 2644
rect 5592 2592 5598 2644
rect 6362 2632 6368 2644
rect 6420 2641 6426 2644
rect 5736 2604 6368 2632
rect 5736 2508 5764 2604
rect 6362 2592 6368 2604
rect 6420 2595 6429 2641
rect 7300 2604 9536 2632
rect 6420 2592 6426 2595
rect 750 2456 756 2508
rect 808 2456 814 2508
rect 1121 2499 1179 2505
rect 1121 2465 1133 2499
rect 1167 2496 1179 2499
rect 3142 2496 3148 2508
rect 1167 2468 1716 2496
rect 1167 2465 1179 2468
rect 1121 2459 1179 2465
rect 768 2428 796 2456
rect 1688 2440 1716 2468
rect 1964 2468 3148 2496
rect 1305 2431 1363 2437
rect 1305 2428 1317 2431
rect 768 2400 1317 2428
rect 1305 2397 1317 2400
rect 1351 2397 1363 2431
rect 1305 2391 1363 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 1811 2431 1869 2437
rect 1811 2397 1823 2431
rect 1857 2428 1869 2431
rect 1964 2428 1992 2468
rect 3142 2456 3148 2468
rect 3200 2456 3206 2508
rect 4246 2456 4252 2508
rect 4304 2456 4310 2508
rect 5718 2456 5724 2508
rect 5776 2456 5782 2508
rect 5828 2468 6598 2496
rect 1857 2400 1992 2428
rect 2041 2431 2099 2437
rect 1857 2397 1869 2400
rect 1811 2391 1869 2397
rect 2041 2397 2053 2431
rect 2087 2428 2099 2431
rect 3513 2431 3571 2437
rect 2087 2400 2774 2428
rect 2087 2397 2099 2400
rect 2041 2391 2099 2397
rect 1670 2252 1676 2304
rect 1728 2292 1734 2304
rect 2130 2292 2136 2304
rect 1728 2264 2136 2292
rect 1728 2252 1734 2264
rect 2130 2252 2136 2264
rect 2188 2252 2194 2304
rect 2746 2292 2774 2400
rect 3513 2397 3525 2431
rect 3559 2428 3571 2431
rect 3786 2428 3792 2440
rect 3559 2400 3792 2428
rect 3559 2397 3571 2400
rect 3513 2391 3571 2397
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 4019 2433 4077 2439
rect 4019 2399 4031 2433
rect 4065 2428 4077 2433
rect 5828 2428 5856 2468
rect 4065 2400 5856 2428
rect 5905 2431 5963 2437
rect 4065 2399 4077 2400
rect 4019 2393 4077 2399
rect 5905 2397 5917 2431
rect 5951 2428 5963 2431
rect 6270 2428 6276 2440
rect 5951 2400 6276 2428
rect 5951 2397 5963 2400
rect 5905 2391 5963 2397
rect 5258 2320 5264 2372
rect 5316 2360 5322 2372
rect 5442 2360 5448 2372
rect 5316 2332 5448 2360
rect 5316 2320 5322 2332
rect 5442 2320 5448 2332
rect 5500 2360 5506 2372
rect 5920 2360 5948 2391
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 6454 2439 6460 2440
rect 6411 2433 6460 2439
rect 6411 2399 6423 2433
rect 6457 2399 6460 2433
rect 6411 2393 6460 2399
rect 6454 2388 6460 2393
rect 6512 2388 6518 2440
rect 6570 2428 6598 2468
rect 6638 2456 6644 2508
rect 6696 2456 6702 2508
rect 7300 2428 7328 2604
rect 9508 2564 9536 2604
rect 9582 2592 9588 2644
rect 9640 2632 9646 2644
rect 9953 2635 10011 2641
rect 9953 2632 9965 2635
rect 9640 2604 9965 2632
rect 9640 2592 9646 2604
rect 9953 2601 9965 2604
rect 9999 2601 10011 2635
rect 9953 2595 10011 2601
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 12986 2632 12992 2644
rect 10100 2604 12992 2632
rect 10100 2592 10106 2604
rect 9508 2536 10548 2564
rect 8478 2505 8484 2508
rect 8021 2499 8079 2505
rect 8021 2465 8033 2499
rect 8067 2496 8079 2499
rect 8440 2499 8484 2505
rect 8067 2468 8248 2496
rect 8067 2465 8079 2468
rect 8021 2459 8079 2465
rect 6570 2400 7328 2428
rect 7374 2388 7380 2440
rect 7432 2428 7438 2440
rect 7742 2428 7748 2440
rect 7432 2400 7748 2428
rect 7432 2388 7438 2400
rect 7742 2388 7748 2400
rect 7800 2428 7806 2440
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7800 2400 8125 2428
rect 7800 2388 7806 2400
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8220 2428 8248 2468
rect 8440 2465 8452 2499
rect 8440 2459 8484 2465
rect 8478 2456 8484 2459
rect 8536 2456 8542 2508
rect 8849 2499 8907 2505
rect 8849 2465 8861 2499
rect 8895 2496 8907 2499
rect 10318 2496 10324 2508
rect 8895 2468 10324 2496
rect 8895 2465 8907 2468
rect 8849 2459 8907 2465
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 10413 2499 10471 2505
rect 10413 2465 10425 2499
rect 10459 2465 10471 2499
rect 10413 2459 10471 2465
rect 8576 2431 8634 2437
rect 8576 2428 8588 2431
rect 8220 2400 8588 2428
rect 8113 2391 8171 2397
rect 8576 2397 8588 2400
rect 8622 2397 8634 2431
rect 8576 2391 8634 2397
rect 5500 2332 5948 2360
rect 5500 2320 5506 2332
rect 7558 2320 7564 2372
rect 7616 2320 7622 2372
rect 10428 2360 10456 2459
rect 10520 2440 10548 2536
rect 11072 2505 11100 2604
rect 12986 2592 12992 2604
rect 13044 2592 13050 2644
rect 14274 2592 14280 2644
rect 14332 2641 14338 2644
rect 14332 2632 14341 2641
rect 14458 2632 14464 2644
rect 14332 2604 14464 2632
rect 14332 2595 14341 2604
rect 14332 2592 14338 2595
rect 14458 2592 14464 2604
rect 14516 2592 14522 2644
rect 16583 2635 16641 2641
rect 16583 2601 16595 2635
rect 16629 2632 16641 2635
rect 16850 2632 16856 2644
rect 16629 2604 16856 2632
rect 16629 2601 16641 2604
rect 16583 2595 16641 2601
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 18782 2592 18788 2644
rect 18840 2641 18846 2644
rect 18840 2632 18849 2641
rect 18840 2604 18885 2632
rect 18840 2595 18849 2604
rect 18840 2592 18846 2595
rect 20714 2592 20720 2644
rect 20772 2632 20778 2644
rect 20809 2635 20867 2641
rect 20809 2632 20821 2635
rect 20772 2604 20821 2632
rect 20772 2592 20778 2604
rect 20809 2601 20821 2604
rect 20855 2601 20867 2635
rect 20809 2595 20867 2601
rect 21542 2592 21548 2644
rect 21600 2632 21606 2644
rect 21735 2635 21793 2641
rect 21735 2632 21747 2635
rect 21600 2604 21747 2632
rect 21600 2592 21606 2604
rect 21735 2601 21747 2604
rect 21781 2601 21793 2635
rect 21735 2595 21793 2601
rect 23477 2635 23535 2641
rect 23477 2601 23489 2635
rect 23523 2632 23535 2635
rect 24026 2632 24032 2644
rect 23523 2604 24032 2632
rect 23523 2601 23535 2604
rect 23477 2595 23535 2601
rect 24026 2592 24032 2604
rect 24084 2592 24090 2644
rect 25682 2632 25688 2644
rect 24228 2604 25688 2632
rect 11333 2567 11391 2573
rect 11333 2533 11345 2567
rect 11379 2564 11391 2567
rect 11606 2564 11612 2576
rect 11379 2536 11612 2564
rect 11379 2533 11391 2536
rect 11333 2527 11391 2533
rect 11606 2524 11612 2536
rect 11664 2524 11670 2576
rect 24228 2564 24256 2604
rect 25682 2592 25688 2604
rect 25740 2592 25746 2644
rect 25774 2592 25780 2644
rect 25832 2632 25838 2644
rect 26605 2635 26663 2641
rect 26605 2632 26617 2635
rect 25832 2604 26617 2632
rect 25832 2592 25838 2604
rect 26605 2601 26617 2604
rect 26651 2601 26663 2635
rect 26605 2595 26663 2601
rect 27338 2592 27344 2644
rect 27396 2632 27402 2644
rect 27706 2632 27712 2644
rect 27396 2604 27712 2632
rect 27396 2592 27402 2604
rect 27706 2592 27712 2604
rect 27764 2592 27770 2644
rect 27982 2592 27988 2644
rect 28040 2632 28046 2644
rect 28040 2604 28120 2632
rect 28040 2592 28046 2604
rect 23676 2536 24256 2564
rect 25516 2536 27660 2564
rect 11057 2499 11115 2505
rect 11057 2465 11069 2499
rect 11103 2465 11115 2499
rect 11057 2459 11115 2465
rect 11422 2456 11428 2508
rect 11480 2456 11486 2508
rect 11624 2496 11652 2524
rect 11936 2499 11994 2505
rect 11936 2496 11948 2499
rect 11624 2468 11948 2496
rect 11936 2465 11948 2468
rect 11982 2465 11994 2499
rect 11936 2459 11994 2465
rect 13725 2499 13783 2505
rect 13725 2465 13737 2499
rect 13771 2496 13783 2499
rect 13771 2468 14320 2496
rect 13771 2465 13783 2468
rect 13725 2459 13783 2465
rect 10502 2388 10508 2440
rect 10560 2388 10566 2440
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2428 10747 2431
rect 11238 2428 11244 2440
rect 10735 2400 11244 2428
rect 10735 2397 10747 2400
rect 10689 2391 10747 2397
rect 11238 2388 11244 2400
rect 11296 2428 11302 2440
rect 11440 2428 11468 2456
rect 11609 2431 11667 2437
rect 11609 2428 11621 2431
rect 11296 2400 11621 2428
rect 11296 2388 11302 2400
rect 11609 2397 11621 2400
rect 11655 2397 11667 2431
rect 11609 2391 11667 2397
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 12072 2431 12130 2437
rect 12072 2428 12084 2431
rect 11848 2400 12084 2428
rect 11848 2388 11854 2400
rect 12072 2397 12084 2400
rect 12118 2397 12130 2431
rect 12072 2391 12130 2397
rect 12342 2388 12348 2440
rect 12400 2388 12406 2440
rect 13814 2388 13820 2440
rect 13872 2388 13878 2440
rect 14292 2437 14320 2468
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 14553 2499 14611 2505
rect 14553 2496 14565 2499
rect 14516 2468 14565 2496
rect 14516 2456 14522 2468
rect 14553 2465 14565 2468
rect 14599 2465 14611 2499
rect 14553 2459 14611 2465
rect 15933 2499 15991 2505
rect 15933 2465 15945 2499
rect 15979 2496 15991 2499
rect 18233 2499 18291 2505
rect 15979 2468 16620 2496
rect 15979 2465 15991 2468
rect 15933 2459 15991 2465
rect 14280 2431 14338 2437
rect 14280 2397 14292 2431
rect 14326 2397 14338 2431
rect 14280 2391 14338 2397
rect 16022 2388 16028 2440
rect 16080 2428 16086 2440
rect 16592 2437 16620 2468
rect 18233 2465 18245 2499
rect 18279 2496 18291 2499
rect 20717 2499 20775 2505
rect 18279 2468 18828 2496
rect 18279 2465 18291 2468
rect 18233 2459 18291 2465
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 16080 2400 16129 2428
rect 16080 2388 16086 2400
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 16580 2431 16638 2437
rect 16580 2397 16592 2431
rect 16626 2397 16638 2431
rect 16580 2391 16638 2397
rect 16853 2431 16911 2437
rect 16853 2397 16865 2431
rect 16899 2428 16911 2431
rect 16899 2400 18276 2428
rect 16899 2397 16911 2400
rect 16853 2391 16911 2397
rect 10428 2332 11468 2360
rect 7576 2292 7604 2320
rect 2746 2264 7604 2292
rect 8110 2252 8116 2304
rect 8168 2292 8174 2304
rect 10962 2292 10968 2304
rect 8168 2264 10968 2292
rect 8168 2252 8174 2264
rect 10962 2252 10968 2264
rect 11020 2292 11026 2304
rect 11146 2292 11152 2304
rect 11020 2264 11152 2292
rect 11020 2252 11026 2264
rect 11146 2252 11152 2264
rect 11204 2252 11210 2304
rect 11440 2292 11468 2332
rect 13832 2292 13860 2388
rect 11440 2264 13860 2292
rect 18248 2292 18276 2400
rect 18322 2388 18328 2440
rect 18380 2388 18386 2440
rect 18800 2437 18828 2468
rect 20717 2465 20729 2499
rect 20763 2496 20775 2499
rect 22278 2496 22284 2508
rect 20763 2480 21410 2496
rect 21468 2480 22284 2496
rect 20763 2468 22284 2480
rect 20763 2465 20775 2468
rect 20717 2459 20775 2465
rect 21382 2452 21496 2468
rect 22278 2456 22284 2468
rect 22336 2456 22342 2508
rect 23676 2505 23704 2536
rect 25516 2508 25544 2536
rect 23661 2499 23719 2505
rect 23661 2465 23673 2499
rect 23707 2465 23719 2499
rect 23661 2459 23719 2465
rect 23750 2456 23756 2508
rect 23808 2496 23814 2508
rect 23937 2499 23995 2505
rect 23937 2496 23949 2499
rect 23808 2468 23949 2496
rect 23808 2456 23814 2468
rect 23937 2465 23949 2468
rect 23983 2465 23995 2499
rect 23937 2459 23995 2465
rect 24857 2499 24915 2505
rect 24857 2465 24869 2499
rect 24903 2496 24915 2499
rect 25314 2496 25320 2508
rect 24903 2468 25320 2496
rect 24903 2465 24915 2468
rect 24857 2459 24915 2465
rect 25314 2456 25320 2468
rect 25372 2456 25378 2508
rect 25498 2456 25504 2508
rect 25556 2456 25562 2508
rect 26418 2456 26424 2508
rect 26476 2496 26482 2508
rect 26513 2499 26571 2505
rect 26513 2496 26525 2499
rect 26476 2468 26525 2496
rect 26476 2456 26482 2468
rect 26513 2465 26525 2468
rect 26559 2465 26571 2499
rect 26513 2459 26571 2465
rect 27341 2499 27399 2505
rect 27341 2465 27353 2499
rect 27387 2496 27399 2499
rect 27522 2496 27528 2508
rect 27387 2468 27528 2496
rect 27387 2465 27399 2468
rect 27341 2459 27399 2465
rect 27522 2456 27528 2468
rect 27580 2456 27586 2508
rect 18788 2431 18846 2437
rect 18788 2397 18800 2431
rect 18834 2397 18846 2431
rect 18788 2391 18846 2397
rect 19061 2431 19119 2437
rect 19061 2397 19073 2431
rect 19107 2428 19119 2431
rect 21269 2431 21327 2437
rect 19107 2400 20668 2428
rect 19107 2397 19119 2400
rect 19061 2391 19119 2397
rect 20346 2320 20352 2372
rect 20404 2320 20410 2372
rect 20530 2292 20536 2304
rect 18248 2264 20536 2292
rect 20530 2252 20536 2264
rect 20588 2252 20594 2304
rect 20640 2292 20668 2400
rect 21269 2397 21281 2431
rect 21315 2397 21327 2431
rect 21269 2391 21327 2397
rect 20714 2320 20720 2372
rect 20772 2360 20778 2372
rect 21284 2360 21312 2391
rect 21634 2388 21640 2440
rect 21692 2428 21698 2440
rect 21732 2431 21790 2437
rect 21732 2428 21744 2431
rect 21692 2400 21744 2428
rect 21692 2388 21698 2400
rect 21732 2397 21744 2400
rect 21778 2397 21790 2431
rect 21732 2391 21790 2397
rect 22005 2431 22063 2437
rect 22005 2397 22017 2431
rect 22051 2428 22063 2431
rect 23474 2428 23480 2440
rect 22051 2400 23480 2428
rect 22051 2397 22063 2400
rect 22005 2391 22063 2397
rect 23474 2388 23480 2400
rect 23532 2388 23538 2440
rect 23566 2388 23572 2440
rect 23624 2428 23630 2440
rect 24118 2428 24124 2440
rect 23624 2400 24124 2428
rect 23624 2388 23630 2400
rect 24118 2388 24124 2400
rect 24176 2388 24182 2440
rect 24302 2388 24308 2440
rect 24360 2428 24366 2440
rect 24448 2431 24506 2437
rect 24448 2428 24460 2431
rect 24360 2400 24460 2428
rect 24360 2388 24366 2400
rect 24448 2397 24460 2400
rect 24494 2397 24506 2431
rect 24448 2391 24506 2397
rect 24578 2388 24584 2440
rect 24636 2428 24642 2440
rect 24636 2400 24681 2428
rect 24636 2388 24642 2400
rect 24762 2388 24768 2440
rect 24820 2428 24826 2440
rect 27632 2428 27660 2536
rect 27890 2456 27896 2508
rect 27948 2496 27954 2508
rect 27985 2499 28043 2505
rect 27985 2496 27997 2499
rect 27948 2468 27997 2496
rect 27948 2456 27954 2468
rect 27985 2465 27997 2468
rect 28031 2465 28043 2499
rect 28092 2496 28120 2604
rect 30006 2592 30012 2644
rect 30064 2592 30070 2644
rect 28312 2499 28370 2505
rect 28312 2496 28324 2499
rect 28092 2468 28324 2496
rect 27985 2459 28043 2465
rect 28312 2465 28324 2468
rect 28358 2465 28370 2499
rect 28312 2459 28370 2465
rect 28721 2499 28779 2505
rect 28721 2465 28733 2499
rect 28767 2496 28779 2499
rect 29730 2496 29736 2508
rect 28767 2468 29736 2496
rect 28767 2465 28779 2468
rect 28721 2459 28779 2465
rect 29730 2456 29736 2468
rect 29788 2456 29794 2508
rect 28166 2428 28172 2440
rect 24820 2400 27568 2428
rect 27632 2400 28172 2428
rect 24820 2388 24826 2400
rect 20772 2332 21312 2360
rect 20772 2320 20778 2332
rect 21910 2292 21916 2304
rect 20640 2264 21916 2292
rect 21910 2252 21916 2264
rect 21968 2252 21974 2304
rect 22186 2252 22192 2304
rect 22244 2292 22250 2304
rect 23109 2295 23167 2301
rect 23109 2292 23121 2295
rect 22244 2264 23121 2292
rect 22244 2252 22250 2264
rect 23109 2261 23121 2264
rect 23155 2261 23167 2295
rect 23109 2255 23167 2261
rect 23753 2295 23811 2301
rect 23753 2261 23765 2295
rect 23799 2292 23811 2295
rect 24486 2292 24492 2304
rect 23799 2264 24492 2292
rect 23799 2261 23811 2264
rect 23753 2255 23811 2261
rect 24486 2252 24492 2264
rect 24544 2252 24550 2304
rect 25958 2252 25964 2304
rect 26016 2252 26022 2304
rect 26418 2252 26424 2304
rect 26476 2292 26482 2304
rect 27433 2295 27491 2301
rect 27433 2292 27445 2295
rect 26476 2264 27445 2292
rect 26476 2252 26482 2264
rect 27433 2261 27445 2264
rect 27479 2261 27491 2295
rect 27540 2292 27568 2400
rect 28166 2388 28172 2400
rect 28224 2388 28230 2440
rect 28448 2433 28506 2439
rect 28448 2399 28460 2433
rect 28494 2428 28506 2433
rect 28534 2428 28540 2440
rect 28494 2400 28540 2428
rect 28494 2399 28506 2400
rect 28448 2393 28506 2399
rect 28534 2388 28540 2400
rect 28592 2388 28598 2440
rect 30377 2363 30435 2369
rect 30377 2329 30389 2363
rect 30423 2329 30435 2363
rect 30377 2323 30435 2329
rect 30392 2292 30420 2323
rect 27540 2264 30420 2292
rect 27433 2255 27491 2261
rect 552 2202 30912 2224
rect 552 2150 4193 2202
rect 4245 2150 4257 2202
rect 4309 2150 4321 2202
rect 4373 2150 4385 2202
rect 4437 2150 4449 2202
rect 4501 2150 11783 2202
rect 11835 2150 11847 2202
rect 11899 2150 11911 2202
rect 11963 2150 11975 2202
rect 12027 2150 12039 2202
rect 12091 2150 19373 2202
rect 19425 2150 19437 2202
rect 19489 2150 19501 2202
rect 19553 2150 19565 2202
rect 19617 2150 19629 2202
rect 19681 2150 26963 2202
rect 27015 2150 27027 2202
rect 27079 2150 27091 2202
rect 27143 2150 27155 2202
rect 27207 2150 27219 2202
rect 27271 2150 30912 2202
rect 552 2128 30912 2150
rect 1118 2048 1124 2100
rect 1176 2088 1182 2100
rect 3237 2091 3295 2097
rect 1176 2060 3188 2088
rect 1176 2048 1182 2060
rect 1443 1955 1501 1961
rect 1443 1921 1455 1955
rect 1489 1952 1501 1955
rect 2774 1952 2780 1964
rect 1489 1924 2780 1952
rect 1489 1921 1501 1924
rect 1443 1915 1501 1921
rect 2774 1912 2780 1924
rect 2832 1912 2838 1964
rect 937 1887 995 1893
rect 937 1853 949 1887
rect 983 1884 995 1887
rect 1302 1884 1308 1896
rect 983 1856 1308 1884
rect 983 1853 995 1856
rect 937 1847 995 1853
rect 1302 1844 1308 1856
rect 1360 1844 1366 1896
rect 1673 1887 1731 1893
rect 1673 1853 1685 1887
rect 1719 1884 1731 1887
rect 2498 1884 2504 1896
rect 1719 1856 2504 1884
rect 1719 1853 1731 1856
rect 1673 1847 1731 1853
rect 2498 1844 2504 1856
rect 2556 1844 2562 1896
rect 3160 1884 3188 2060
rect 3237 2057 3249 2091
rect 3283 2088 3295 2091
rect 3602 2088 3608 2100
rect 3283 2060 3608 2088
rect 3283 2057 3295 2060
rect 3237 2051 3295 2057
rect 3602 2048 3608 2060
rect 3660 2048 3666 2100
rect 4522 2048 4528 2100
rect 4580 2088 4586 2100
rect 5445 2091 5503 2097
rect 5445 2088 5457 2091
rect 4580 2060 5457 2088
rect 4580 2048 4586 2060
rect 5445 2057 5457 2060
rect 5491 2057 5503 2091
rect 5445 2051 5503 2057
rect 5626 2048 5632 2100
rect 5684 2088 5690 2100
rect 5684 2060 7604 2088
rect 5684 2048 5690 2060
rect 3605 1955 3663 1961
rect 3605 1921 3617 1955
rect 3651 1952 3663 1955
rect 3786 1952 3792 1964
rect 3651 1924 3792 1952
rect 3651 1921 3663 1924
rect 3605 1915 3663 1921
rect 3786 1912 3792 1924
rect 3844 1912 3850 1964
rect 3970 1961 3976 1964
rect 3932 1955 3976 1961
rect 3932 1921 3944 1955
rect 3932 1915 3976 1921
rect 3970 1912 3976 1915
rect 4028 1912 4034 1964
rect 4062 1912 4068 1964
rect 4120 1959 4126 1964
rect 4120 1953 4169 1959
rect 4120 1919 4123 1953
rect 4157 1919 4169 1953
rect 4120 1913 4169 1919
rect 4120 1912 4126 1913
rect 4338 1912 4344 1964
rect 4396 1912 4402 1964
rect 5994 1912 6000 1964
rect 6052 1952 6058 1964
rect 6276 1955 6334 1961
rect 6276 1952 6288 1955
rect 6052 1924 6288 1952
rect 6052 1912 6058 1924
rect 6276 1921 6288 1924
rect 6322 1921 6334 1955
rect 6276 1915 6334 1921
rect 6362 1912 6368 1964
rect 6420 1952 6426 1964
rect 7576 1952 7604 2060
rect 7650 2048 7656 2100
rect 7708 2048 7714 2100
rect 7834 2048 7840 2100
rect 7892 2088 7898 2100
rect 8021 2091 8079 2097
rect 8021 2088 8033 2091
rect 7892 2060 8033 2088
rect 7892 2048 7898 2060
rect 8021 2057 8033 2060
rect 8067 2057 8079 2091
rect 8021 2051 8079 2057
rect 8757 2091 8815 2097
rect 8757 2057 8769 2091
rect 8803 2088 8815 2091
rect 8846 2088 8852 2100
rect 8803 2060 8852 2088
rect 8803 2057 8815 2060
rect 8757 2051 8815 2057
rect 8846 2048 8852 2060
rect 8904 2048 8910 2100
rect 12342 2088 12348 2100
rect 8956 2060 12348 2088
rect 7742 1980 7748 2032
rect 7800 2020 7806 2032
rect 8956 2020 8984 2060
rect 12342 2048 12348 2060
rect 12400 2048 12406 2100
rect 13633 2091 13691 2097
rect 13633 2057 13645 2091
rect 13679 2088 13691 2091
rect 15102 2088 15108 2100
rect 13679 2060 15108 2088
rect 13679 2057 13691 2060
rect 13633 2051 13691 2057
rect 15102 2048 15108 2060
rect 15160 2048 15166 2100
rect 15948 2060 17908 2088
rect 7800 1992 8984 2020
rect 7800 1980 7806 1992
rect 6420 1924 6684 1952
rect 7576 1924 8340 1952
rect 6420 1912 6426 1924
rect 3421 1887 3479 1893
rect 3421 1884 3433 1887
rect 3160 1856 3433 1884
rect 3421 1853 3433 1856
rect 3467 1853 3479 1887
rect 3421 1847 3479 1853
rect 3050 1776 3056 1828
rect 3108 1776 3114 1828
rect 1403 1751 1461 1757
rect 1403 1717 1415 1751
rect 1449 1748 1461 1751
rect 1762 1748 1768 1760
rect 1449 1720 1768 1748
rect 1449 1717 1461 1720
rect 1403 1711 1461 1717
rect 1762 1708 1768 1720
rect 1820 1708 1826 1760
rect 3436 1748 3464 1847
rect 4430 1844 4436 1896
rect 4488 1884 4494 1896
rect 5442 1884 5448 1896
rect 4488 1856 5448 1884
rect 4488 1844 4494 1856
rect 5442 1844 5448 1856
rect 5500 1884 5506 1896
rect 5813 1887 5871 1893
rect 5813 1884 5825 1887
rect 5500 1856 5825 1884
rect 5500 1844 5506 1856
rect 5813 1853 5825 1856
rect 5859 1853 5871 1887
rect 6549 1887 6607 1893
rect 6549 1884 6561 1887
rect 5813 1847 5871 1853
rect 5920 1856 6561 1884
rect 5626 1776 5632 1828
rect 5684 1816 5690 1828
rect 5920 1816 5948 1856
rect 6549 1853 6561 1856
rect 6595 1853 6607 1887
rect 6656 1884 6684 1924
rect 6656 1856 7236 1884
rect 6549 1847 6607 1853
rect 5684 1788 5948 1816
rect 7208 1816 7236 1856
rect 8110 1844 8116 1896
rect 8168 1884 8174 1896
rect 8205 1887 8263 1893
rect 8205 1884 8217 1887
rect 8168 1856 8217 1884
rect 8168 1844 8174 1856
rect 8205 1853 8217 1856
rect 8251 1853 8263 1887
rect 8312 1884 8340 1924
rect 8846 1912 8852 1964
rect 8904 1952 8910 1964
rect 9496 1955 9554 1961
rect 9496 1952 9508 1955
rect 8904 1924 9508 1952
rect 8904 1912 8910 1924
rect 9496 1921 9508 1924
rect 9542 1921 9554 1955
rect 9496 1915 9554 1921
rect 11149 1955 11207 1961
rect 11149 1921 11161 1955
rect 11195 1952 11207 1955
rect 11704 1955 11762 1961
rect 11704 1952 11716 1955
rect 11195 1924 11716 1952
rect 11195 1921 11207 1924
rect 11149 1915 11207 1921
rect 11704 1921 11716 1924
rect 11750 1921 11762 1955
rect 11704 1915 11762 1921
rect 13357 1955 13415 1961
rect 13357 1921 13369 1955
rect 13403 1952 13415 1955
rect 14372 1955 14430 1961
rect 14372 1952 14384 1955
rect 13403 1924 14384 1952
rect 13403 1921 13415 1924
rect 13357 1915 13415 1921
rect 14372 1921 14384 1924
rect 14418 1921 14430 1955
rect 14372 1915 14430 1921
rect 8312 1856 8984 1884
rect 8205 1847 8263 1853
rect 8481 1819 8539 1825
rect 8481 1816 8493 1819
rect 7208 1788 8493 1816
rect 5684 1776 5690 1788
rect 8481 1785 8493 1788
rect 8527 1785 8539 1819
rect 8956 1816 8984 1856
rect 9030 1844 9036 1896
rect 9088 1844 9094 1896
rect 9769 1887 9827 1893
rect 9769 1884 9781 1887
rect 9140 1856 9781 1884
rect 9140 1816 9168 1856
rect 9769 1853 9781 1856
rect 9815 1853 9827 1887
rect 9769 1847 9827 1853
rect 11238 1844 11244 1896
rect 11296 1844 11302 1896
rect 11606 1893 11612 1896
rect 11568 1887 11612 1893
rect 11568 1853 11580 1887
rect 11568 1847 11612 1853
rect 11606 1844 11612 1847
rect 11664 1844 11670 1896
rect 11974 1844 11980 1896
rect 12032 1844 12038 1896
rect 13817 1887 13875 1893
rect 13817 1853 13829 1887
rect 13863 1853 13875 1887
rect 13817 1847 13875 1853
rect 8956 1788 9168 1816
rect 8481 1779 8539 1785
rect 5350 1748 5356 1760
rect 3436 1720 5356 1748
rect 5350 1708 5356 1720
rect 5408 1708 5414 1760
rect 5718 1708 5724 1760
rect 5776 1748 5782 1760
rect 6279 1751 6337 1757
rect 6279 1748 6291 1751
rect 5776 1720 6291 1748
rect 5776 1708 5782 1720
rect 6279 1717 6291 1720
rect 6325 1717 6337 1751
rect 6279 1711 6337 1717
rect 9030 1708 9036 1760
rect 9088 1748 9094 1760
rect 9398 1748 9404 1760
rect 9088 1720 9404 1748
rect 9088 1708 9094 1720
rect 9398 1708 9404 1720
rect 9456 1748 9462 1760
rect 9499 1751 9557 1757
rect 9499 1748 9511 1751
rect 9456 1720 9511 1748
rect 9456 1708 9462 1720
rect 9499 1717 9511 1720
rect 9545 1717 9557 1751
rect 9499 1711 9557 1717
rect 9674 1708 9680 1760
rect 9732 1748 9738 1760
rect 11974 1748 11980 1760
rect 9732 1720 11980 1748
rect 9732 1708 9738 1720
rect 11974 1708 11980 1720
rect 12032 1708 12038 1760
rect 13832 1748 13860 1847
rect 13906 1844 13912 1896
rect 13964 1844 13970 1896
rect 14274 1893 14280 1896
rect 14236 1887 14280 1893
rect 14236 1853 14248 1887
rect 14236 1847 14280 1853
rect 14274 1844 14280 1847
rect 14332 1844 14338 1896
rect 14642 1844 14648 1896
rect 14700 1844 14706 1896
rect 15948 1748 15976 2060
rect 17880 2020 17908 2060
rect 17954 2048 17960 2100
rect 18012 2088 18018 2100
rect 18325 2091 18383 2097
rect 18325 2088 18337 2091
rect 18012 2060 18337 2088
rect 18012 2048 18018 2060
rect 18325 2057 18337 2060
rect 18371 2057 18383 2091
rect 21726 2088 21732 2100
rect 18325 2051 18383 2057
rect 18708 2060 21732 2088
rect 18708 2020 18736 2060
rect 21726 2048 21732 2060
rect 21784 2048 21790 2100
rect 24026 2048 24032 2100
rect 24084 2088 24090 2100
rect 24762 2088 24768 2100
rect 24084 2060 24768 2088
rect 24084 2048 24090 2060
rect 24762 2048 24768 2060
rect 24820 2048 24826 2100
rect 27798 2048 27804 2100
rect 27856 2088 27862 2100
rect 28077 2091 28135 2097
rect 28077 2088 28089 2091
rect 27856 2060 28089 2088
rect 27856 2048 27862 2060
rect 28077 2057 28089 2060
rect 28123 2057 28135 2091
rect 29181 2091 29239 2097
rect 28077 2051 28135 2057
rect 28190 2060 28994 2088
rect 23109 2023 23167 2029
rect 23109 2020 23121 2023
rect 17880 1992 18736 2020
rect 22296 1992 23121 2020
rect 16022 1912 16028 1964
rect 16080 1952 16086 1964
rect 16117 1955 16175 1961
rect 16117 1952 16129 1955
rect 16080 1924 16129 1952
rect 16080 1912 16086 1924
rect 16117 1921 16129 1924
rect 16163 1921 16175 1955
rect 16580 1955 16638 1961
rect 16580 1952 16592 1955
rect 16117 1915 16175 1921
rect 16224 1924 16592 1952
rect 16224 1884 16252 1924
rect 16580 1921 16592 1924
rect 16626 1921 16638 1955
rect 16580 1915 16638 1921
rect 18233 1955 18291 1961
rect 18233 1921 18245 1955
rect 18279 1952 18291 1955
rect 19156 1955 19214 1961
rect 19156 1952 19168 1955
rect 18279 1924 19168 1952
rect 18279 1921 18291 1924
rect 18233 1915 18291 1921
rect 19156 1921 19168 1924
rect 19202 1921 19214 1955
rect 19156 1915 19214 1921
rect 20714 1912 20720 1964
rect 20772 1912 20778 1964
rect 21266 1961 21272 1964
rect 21228 1955 21272 1961
rect 21228 1921 21240 1955
rect 21228 1915 21272 1921
rect 21266 1912 21272 1915
rect 21324 1912 21330 1964
rect 21380 1953 21438 1959
rect 21380 1919 21392 1953
rect 21426 1950 21438 1953
rect 21637 1955 21695 1961
rect 21468 1950 21588 1952
rect 21426 1924 21588 1950
rect 21426 1922 21496 1924
rect 21426 1919 21438 1922
rect 21380 1913 21438 1919
rect 16040 1856 16252 1884
rect 16040 1825 16068 1856
rect 16666 1844 16672 1896
rect 16724 1884 16730 1896
rect 16853 1887 16911 1893
rect 16853 1884 16865 1887
rect 16724 1856 16865 1884
rect 16724 1844 16730 1856
rect 16853 1853 16865 1856
rect 16899 1853 16911 1887
rect 16853 1847 16911 1853
rect 18322 1844 18328 1896
rect 18380 1844 18386 1896
rect 18506 1844 18512 1896
rect 18564 1844 18570 1896
rect 18693 1887 18751 1893
rect 18693 1853 18705 1887
rect 18739 1853 18751 1887
rect 18693 1847 18751 1853
rect 16025 1819 16083 1825
rect 16025 1785 16037 1819
rect 16071 1785 16083 1819
rect 18340 1816 18368 1844
rect 18708 1816 18736 1847
rect 18782 1844 18788 1896
rect 18840 1884 18846 1896
rect 19020 1887 19078 1893
rect 19020 1884 19032 1887
rect 18840 1856 19032 1884
rect 18840 1844 18846 1856
rect 19020 1853 19032 1856
rect 19066 1853 19078 1887
rect 19020 1847 19078 1853
rect 19426 1844 19432 1896
rect 19484 1844 19490 1896
rect 20732 1884 20760 1912
rect 20898 1884 20904 1896
rect 20732 1856 20904 1884
rect 20898 1844 20904 1856
rect 20956 1844 20962 1896
rect 21560 1884 21588 1924
rect 21637 1921 21649 1955
rect 21683 1952 21695 1955
rect 22296 1952 22324 1992
rect 23109 1989 23121 1992
rect 23155 1989 23167 2023
rect 23750 2020 23756 2032
rect 23109 1983 23167 1989
rect 23308 1992 23756 2020
rect 21683 1924 22324 1952
rect 21683 1921 21695 1924
rect 21637 1915 21695 1921
rect 21726 1884 21732 1896
rect 21560 1856 21732 1884
rect 21726 1844 21732 1856
rect 21784 1844 21790 1896
rect 23308 1893 23336 1992
rect 23750 1980 23756 1992
rect 23808 1980 23814 2032
rect 23382 1912 23388 1964
rect 23440 1912 23446 1964
rect 23842 1912 23848 1964
rect 23900 1912 23906 1964
rect 24210 1961 24216 1964
rect 24172 1955 24216 1961
rect 24172 1921 24184 1955
rect 24172 1915 24216 1921
rect 24210 1912 24216 1915
rect 24268 1912 24274 1964
rect 24308 1953 24366 1959
rect 24308 1919 24320 1953
rect 24354 1919 24366 1953
rect 24308 1913 24366 1919
rect 23293 1887 23351 1893
rect 23293 1884 23305 1887
rect 22480 1856 23305 1884
rect 22480 1828 22508 1856
rect 23293 1853 23305 1856
rect 23339 1853 23351 1887
rect 23400 1884 23428 1912
rect 23569 1887 23627 1893
rect 23569 1884 23581 1887
rect 23400 1856 23581 1884
rect 23293 1847 23351 1853
rect 23569 1853 23581 1856
rect 23615 1853 23627 1887
rect 23569 1847 23627 1853
rect 23958 1880 24215 1884
rect 24323 1880 24351 1913
rect 24486 1912 24492 1964
rect 24544 1952 24550 1964
rect 24581 1955 24639 1961
rect 24581 1952 24593 1955
rect 24544 1924 24593 1952
rect 24544 1912 24550 1924
rect 24581 1921 24593 1924
rect 24627 1921 24639 1955
rect 24581 1915 24639 1921
rect 24946 1912 24952 1964
rect 25004 1952 25010 1964
rect 26237 1955 26295 1961
rect 26237 1952 26249 1955
rect 25004 1924 26249 1952
rect 25004 1912 25010 1924
rect 26237 1921 26249 1924
rect 26283 1952 26295 1955
rect 26418 1952 26424 1964
rect 26283 1924 26424 1952
rect 26283 1921 26295 1924
rect 26237 1915 26295 1921
rect 26418 1912 26424 1924
rect 26476 1912 26482 1964
rect 26733 1937 26791 1943
rect 26733 1903 26745 1937
rect 26779 1903 26791 1937
rect 26878 1912 26884 1964
rect 26936 1952 26942 1964
rect 26973 1955 27031 1961
rect 26973 1952 26985 1955
rect 26936 1924 26985 1952
rect 26936 1912 26942 1924
rect 26973 1921 26985 1924
rect 27019 1921 27031 1955
rect 26973 1915 27031 1921
rect 27430 1912 27436 1964
rect 27488 1952 27494 1964
rect 28190 1952 28218 2060
rect 28966 2020 28994 2060
rect 29181 2057 29193 2091
rect 29227 2088 29239 2091
rect 29362 2088 29368 2100
rect 29227 2060 29368 2088
rect 29227 2057 29239 2060
rect 29181 2051 29239 2057
rect 29362 2048 29368 2060
rect 29420 2048 29426 2100
rect 29454 2048 29460 2100
rect 29512 2088 29518 2100
rect 29641 2091 29699 2097
rect 29641 2088 29653 2091
rect 29512 2060 29653 2088
rect 29512 2048 29518 2060
rect 29641 2057 29653 2060
rect 29687 2057 29699 2091
rect 29641 2051 29699 2057
rect 30101 2023 30159 2029
rect 30101 2020 30113 2023
rect 28966 1992 30113 2020
rect 30101 1989 30113 1992
rect 30147 1989 30159 2023
rect 30101 1983 30159 1989
rect 27488 1924 28218 1952
rect 27488 1912 27494 1924
rect 28258 1912 28264 1964
rect 28316 1912 28322 1964
rect 28552 1924 28764 1952
rect 26733 1897 26791 1903
rect 23958 1856 24351 1880
rect 18340 1788 18736 1816
rect 20809 1819 20867 1825
rect 16025 1779 16083 1785
rect 20809 1785 20821 1819
rect 20855 1816 20867 1819
rect 20990 1816 20996 1828
rect 20855 1788 20996 1816
rect 20855 1785 20867 1788
rect 20809 1779 20867 1785
rect 20990 1776 20996 1788
rect 21048 1776 21054 1828
rect 22462 1776 22468 1828
rect 22520 1776 22526 1828
rect 22922 1816 22928 1828
rect 22664 1788 22928 1816
rect 13832 1720 15976 1748
rect 16583 1751 16641 1757
rect 16583 1717 16595 1751
rect 16629 1748 16641 1751
rect 16850 1748 16856 1760
rect 16629 1720 16856 1748
rect 16629 1717 16641 1720
rect 16583 1711 16641 1717
rect 16850 1708 16856 1720
rect 16908 1708 16914 1760
rect 17126 1708 17132 1760
rect 17184 1748 17190 1760
rect 19242 1748 19248 1760
rect 17184 1720 19248 1748
rect 17184 1708 17190 1720
rect 19242 1708 19248 1720
rect 19300 1708 19306 1760
rect 20070 1708 20076 1760
rect 20128 1748 20134 1760
rect 22664 1748 22692 1788
rect 22922 1776 22928 1788
rect 22980 1776 22986 1828
rect 23017 1819 23075 1825
rect 23017 1785 23029 1819
rect 23063 1816 23075 1819
rect 23958 1816 23986 1856
rect 24187 1852 24351 1856
rect 26050 1844 26056 1896
rect 26108 1884 26114 1896
rect 26564 1887 26622 1893
rect 26564 1884 26576 1887
rect 26108 1856 26576 1884
rect 26108 1844 26114 1856
rect 26564 1853 26576 1856
rect 26610 1853 26622 1887
rect 26763 1884 26791 1897
rect 28276 1884 28304 1912
rect 26763 1856 28304 1884
rect 26564 1847 26622 1853
rect 23063 1788 23986 1816
rect 23063 1785 23075 1788
rect 23017 1779 23075 1785
rect 27706 1776 27712 1828
rect 27764 1816 27770 1828
rect 28552 1816 28580 1924
rect 28629 1887 28687 1893
rect 28629 1853 28641 1887
rect 28675 1853 28687 1887
rect 28736 1884 28764 1924
rect 28989 1887 29047 1893
rect 28736 1880 28948 1884
rect 28989 1880 29001 1887
rect 28736 1856 29001 1880
rect 28629 1847 28687 1853
rect 28920 1853 29001 1856
rect 29035 1853 29047 1887
rect 28920 1852 29047 1853
rect 28989 1847 29047 1852
rect 27764 1788 28580 1816
rect 27764 1776 27770 1788
rect 28644 1760 28672 1847
rect 28718 1776 28724 1828
rect 28776 1816 28782 1828
rect 30377 1819 30435 1825
rect 30377 1816 30389 1819
rect 28776 1788 30389 1816
rect 28776 1776 28782 1788
rect 30377 1785 30389 1788
rect 30423 1785 30435 1819
rect 30377 1779 30435 1785
rect 20128 1720 22692 1748
rect 20128 1708 20134 1720
rect 22738 1708 22744 1760
rect 22796 1748 22802 1760
rect 23385 1751 23443 1757
rect 23385 1748 23397 1751
rect 22796 1720 23397 1748
rect 22796 1708 22802 1720
rect 23385 1717 23397 1720
rect 23431 1717 23443 1751
rect 23385 1711 23443 1717
rect 23474 1708 23480 1760
rect 23532 1748 23538 1760
rect 23658 1748 23664 1760
rect 23532 1720 23664 1748
rect 23532 1708 23538 1720
rect 23658 1708 23664 1720
rect 23716 1708 23722 1760
rect 24486 1708 24492 1760
rect 24544 1748 24550 1760
rect 24854 1748 24860 1760
rect 24544 1720 24860 1748
rect 24544 1708 24550 1720
rect 24854 1708 24860 1720
rect 24912 1708 24918 1760
rect 24946 1708 24952 1760
rect 25004 1748 25010 1760
rect 25685 1751 25743 1757
rect 25685 1748 25697 1751
rect 25004 1720 25697 1748
rect 25004 1708 25010 1720
rect 25685 1717 25697 1720
rect 25731 1717 25743 1751
rect 25685 1711 25743 1717
rect 26602 1708 26608 1760
rect 26660 1748 26666 1760
rect 28626 1748 28632 1760
rect 26660 1720 28632 1748
rect 26660 1708 26666 1720
rect 28626 1708 28632 1720
rect 28684 1708 28690 1760
rect 28810 1708 28816 1760
rect 28868 1748 28874 1760
rect 29086 1748 29092 1760
rect 28868 1720 29092 1748
rect 28868 1708 28874 1720
rect 29086 1708 29092 1720
rect 29144 1708 29150 1760
rect 552 1658 31072 1680
rect 552 1606 7988 1658
rect 8040 1606 8052 1658
rect 8104 1606 8116 1658
rect 8168 1606 8180 1658
rect 8232 1606 8244 1658
rect 8296 1606 15578 1658
rect 15630 1606 15642 1658
rect 15694 1606 15706 1658
rect 15758 1606 15770 1658
rect 15822 1606 15834 1658
rect 15886 1606 23168 1658
rect 23220 1606 23232 1658
rect 23284 1606 23296 1658
rect 23348 1606 23360 1658
rect 23412 1606 23424 1658
rect 23476 1606 30758 1658
rect 30810 1606 30822 1658
rect 30874 1606 30886 1658
rect 30938 1606 30950 1658
rect 31002 1606 31014 1658
rect 31066 1606 31072 1658
rect 552 1584 31072 1606
rect 1029 1547 1087 1553
rect 1029 1513 1041 1547
rect 1075 1544 1087 1547
rect 1210 1544 1216 1556
rect 1075 1516 1216 1544
rect 1075 1513 1087 1516
rect 1029 1507 1087 1513
rect 1210 1504 1216 1516
rect 1268 1504 1274 1556
rect 1762 1504 1768 1556
rect 1820 1553 1826 1556
rect 1820 1507 1829 1553
rect 1820 1504 1826 1507
rect 3050 1504 3056 1556
rect 3108 1544 3114 1556
rect 3108 1516 5488 1544
rect 3108 1504 3114 1516
rect 5460 1476 5488 1516
rect 5534 1504 5540 1556
rect 5592 1504 5598 1556
rect 5902 1504 5908 1556
rect 5960 1504 5966 1556
rect 6923 1547 6981 1553
rect 6018 1516 6183 1544
rect 6018 1476 6046 1516
rect 5460 1448 6046 1476
rect 6155 1476 6183 1516
rect 6923 1513 6935 1547
rect 6969 1544 6981 1547
rect 8481 1547 8539 1553
rect 6969 1516 8432 1544
rect 6969 1513 6981 1516
rect 6923 1507 6981 1513
rect 8404 1476 8432 1516
rect 8481 1513 8493 1547
rect 8527 1544 8539 1547
rect 8527 1516 11376 1544
rect 8527 1513 8539 1516
rect 8481 1507 8539 1513
rect 11057 1479 11115 1485
rect 6155 1448 6598 1476
rect 8404 1448 8800 1476
rect 1026 1368 1032 1420
rect 1084 1408 1090 1420
rect 1213 1411 1271 1417
rect 1213 1408 1225 1411
rect 1084 1380 1225 1408
rect 1084 1368 1090 1380
rect 1213 1377 1225 1380
rect 1259 1377 1271 1411
rect 1213 1371 1271 1377
rect 1302 1368 1308 1420
rect 1360 1368 1366 1420
rect 2130 1408 2136 1420
rect 1964 1380 2136 1408
rect 1801 1361 1859 1367
rect 1801 1358 1813 1361
rect 1780 1327 1813 1358
rect 1847 1340 1859 1361
rect 1964 1340 1992 1380
rect 2130 1368 2136 1380
rect 2188 1368 2194 1420
rect 3421 1411 3479 1417
rect 3421 1377 3433 1411
rect 3467 1408 3479 1411
rect 5810 1408 5816 1420
rect 3467 1380 5816 1408
rect 3467 1377 3479 1380
rect 3421 1371 3479 1377
rect 5810 1368 5816 1380
rect 5868 1368 5874 1420
rect 5994 1368 6000 1420
rect 6052 1408 6058 1420
rect 6089 1411 6147 1417
rect 6089 1408 6101 1411
rect 6052 1380 6101 1408
rect 6052 1368 6058 1380
rect 6089 1377 6101 1380
rect 6135 1377 6147 1411
rect 6089 1371 6147 1377
rect 6178 1368 6184 1420
rect 6236 1408 6242 1420
rect 6365 1411 6423 1417
rect 6236 1380 6316 1408
rect 6236 1368 6242 1380
rect 1847 1327 1992 1340
rect 1780 1312 1992 1327
rect 2038 1300 2044 1352
rect 2096 1300 2102 1352
rect 3510 1300 3516 1352
rect 3568 1300 3574 1352
rect 3878 1349 3884 1352
rect 3840 1343 3884 1349
rect 3840 1309 3852 1343
rect 3840 1303 3884 1309
rect 3878 1300 3884 1303
rect 3936 1300 3942 1352
rect 4062 1349 4068 1352
rect 4019 1343 4068 1349
rect 4019 1309 4031 1343
rect 4065 1309 4068 1343
rect 4019 1303 4068 1309
rect 4062 1300 4068 1303
rect 4120 1300 4126 1352
rect 4246 1300 4252 1352
rect 4304 1300 4310 1352
rect 4338 1300 4344 1352
rect 4396 1340 4402 1352
rect 6288 1340 6316 1380
rect 6365 1377 6377 1411
rect 6411 1377 6423 1411
rect 6570 1408 6598 1448
rect 8665 1411 8723 1417
rect 6570 1380 6979 1408
rect 6365 1371 6423 1377
rect 4396 1312 6132 1340
rect 4396 1300 4402 1312
rect 5626 1232 5632 1284
rect 5684 1232 5690 1284
rect 1670 1164 1676 1216
rect 1728 1204 1734 1216
rect 4430 1204 4436 1216
rect 1728 1176 4436 1204
rect 1728 1164 1734 1176
rect 4430 1164 4436 1176
rect 4488 1164 4494 1216
rect 4614 1164 4620 1216
rect 4672 1204 4678 1216
rect 5644 1204 5672 1232
rect 4672 1176 5672 1204
rect 6104 1204 6132 1312
rect 6196 1312 6316 1340
rect 6196 1281 6224 1312
rect 6181 1275 6239 1281
rect 6181 1241 6193 1275
rect 6227 1241 6239 1275
rect 6181 1235 6239 1241
rect 6380 1204 6408 1371
rect 6951 1367 6979 1380
rect 8665 1377 8677 1411
rect 8711 1377 8723 1411
rect 8665 1371 8723 1377
rect 8772 1392 8800 1448
rect 11057 1445 11069 1479
rect 11103 1476 11115 1479
rect 11238 1476 11244 1488
rect 11103 1448 11244 1476
rect 11103 1445 11115 1448
rect 11057 1439 11115 1445
rect 11238 1436 11244 1448
rect 11296 1436 11302 1488
rect 11348 1476 11376 1516
rect 11606 1504 11612 1556
rect 11664 1544 11670 1556
rect 12075 1547 12133 1553
rect 12075 1544 12087 1547
rect 11664 1516 12087 1544
rect 11664 1504 11670 1516
rect 12075 1513 12087 1516
rect 12121 1513 12133 1547
rect 12075 1507 12133 1513
rect 14274 1504 14280 1556
rect 14332 1553 14338 1556
rect 14332 1544 14341 1553
rect 16583 1547 16641 1553
rect 14332 1516 14377 1544
rect 14332 1507 14341 1516
rect 16583 1513 16595 1547
rect 16629 1544 16641 1547
rect 16850 1544 16856 1556
rect 16629 1516 16856 1544
rect 16629 1513 16641 1516
rect 16583 1507 16641 1513
rect 14332 1504 14338 1507
rect 16850 1504 16856 1516
rect 16908 1504 16914 1556
rect 18782 1504 18788 1556
rect 18840 1553 18846 1556
rect 18840 1544 18849 1553
rect 18840 1516 18885 1544
rect 18840 1507 18849 1516
rect 18840 1504 18846 1507
rect 19426 1504 19432 1556
rect 19484 1544 19490 1556
rect 20809 1547 20867 1553
rect 20809 1544 20821 1547
rect 19484 1516 20821 1544
rect 19484 1504 19490 1516
rect 20809 1513 20821 1516
rect 20855 1513 20867 1547
rect 20809 1507 20867 1513
rect 20898 1504 20904 1556
rect 20956 1544 20962 1556
rect 20956 1516 21312 1544
rect 20956 1504 20962 1516
rect 11698 1476 11704 1488
rect 11348 1448 11704 1476
rect 11698 1436 11704 1448
rect 11756 1436 11762 1488
rect 20070 1436 20076 1488
rect 20128 1436 20134 1488
rect 20441 1479 20499 1485
rect 20441 1445 20453 1479
rect 20487 1476 20499 1479
rect 20487 1448 21120 1476
rect 20487 1445 20499 1448
rect 20441 1439 20499 1445
rect 11425 1411 11483 1417
rect 11425 1408 11437 1411
rect 6951 1361 7011 1367
rect 8680 1364 8714 1371
rect 8772 1364 8846 1392
rect 6457 1343 6515 1349
rect 6457 1309 6469 1343
rect 6503 1309 6515 1343
rect 6951 1330 6965 1361
rect 6953 1327 6965 1330
rect 6999 1327 7011 1361
rect 6953 1321 7011 1327
rect 6457 1303 6515 1309
rect 6104 1176 6408 1204
rect 6472 1204 6500 1303
rect 7190 1300 7196 1352
rect 7248 1300 7254 1352
rect 8686 1204 8714 1364
rect 8818 1340 8846 1364
rect 10704 1380 11437 1408
rect 9030 1349 9036 1352
rect 8992 1343 9036 1349
rect 8992 1340 9004 1343
rect 8818 1312 9004 1340
rect 8992 1309 9004 1312
rect 8992 1303 9036 1309
rect 9030 1300 9036 1303
rect 9088 1300 9094 1352
rect 9122 1300 9128 1352
rect 9180 1340 9186 1352
rect 9401 1343 9459 1349
rect 9180 1312 9225 1340
rect 9180 1300 9186 1312
rect 9401 1309 9413 1343
rect 9447 1340 9459 1343
rect 10134 1340 10140 1352
rect 9447 1312 10140 1340
rect 9447 1309 9459 1312
rect 9401 1303 9459 1309
rect 10134 1300 10140 1312
rect 10192 1300 10198 1352
rect 8938 1204 8944 1216
rect 6472 1176 8944 1204
rect 4672 1164 4678 1176
rect 8938 1164 8944 1176
rect 8996 1204 9002 1216
rect 10704 1204 10732 1380
rect 11425 1377 11437 1380
rect 11471 1377 11483 1411
rect 13725 1411 13783 1417
rect 11425 1371 11483 1377
rect 11532 1380 11744 1408
rect 10781 1343 10839 1349
rect 10781 1309 10793 1343
rect 10827 1340 10839 1343
rect 11532 1340 11560 1380
rect 10827 1312 11560 1340
rect 11609 1343 11667 1349
rect 10827 1309 10839 1312
rect 10781 1303 10839 1309
rect 11609 1309 11621 1343
rect 11655 1309 11667 1343
rect 11716 1340 11744 1380
rect 13725 1377 13737 1411
rect 13771 1408 13783 1411
rect 15933 1411 15991 1417
rect 13771 1380 14320 1408
rect 13771 1377 13783 1380
rect 13725 1371 13783 1377
rect 12072 1361 12130 1367
rect 12072 1340 12084 1361
rect 11716 1327 12084 1340
rect 12118 1327 12130 1361
rect 11716 1321 12130 1327
rect 11716 1312 12112 1321
rect 11609 1303 11667 1309
rect 11238 1232 11244 1284
rect 11296 1272 11302 1284
rect 11624 1272 11652 1303
rect 12158 1300 12164 1352
rect 12216 1340 12222 1352
rect 12345 1343 12403 1349
rect 12345 1340 12357 1343
rect 12216 1312 12357 1340
rect 12216 1300 12222 1312
rect 12345 1309 12357 1312
rect 12391 1309 12403 1343
rect 12345 1303 12403 1309
rect 13814 1300 13820 1352
rect 13872 1300 13878 1352
rect 14292 1349 14320 1380
rect 15933 1377 15945 1411
rect 15979 1408 15991 1411
rect 18233 1411 18291 1417
rect 15979 1380 16620 1408
rect 15979 1377 15991 1380
rect 15933 1371 15991 1377
rect 14280 1343 14338 1349
rect 14280 1309 14292 1343
rect 14326 1309 14338 1343
rect 14280 1303 14338 1309
rect 14366 1300 14372 1352
rect 14424 1340 14430 1352
rect 14553 1343 14611 1349
rect 14553 1340 14565 1343
rect 14424 1312 14565 1340
rect 14424 1300 14430 1312
rect 14553 1309 14565 1312
rect 14599 1309 14611 1343
rect 14553 1303 14611 1309
rect 16022 1300 16028 1352
rect 16080 1340 16086 1352
rect 16592 1349 16620 1380
rect 18233 1377 18245 1411
rect 18279 1408 18291 1411
rect 20088 1408 20116 1436
rect 20717 1411 20775 1417
rect 20717 1408 20729 1411
rect 18279 1380 18828 1408
rect 20088 1380 20729 1408
rect 18279 1377 18291 1380
rect 18233 1371 18291 1377
rect 16117 1343 16175 1349
rect 16117 1340 16129 1343
rect 16080 1312 16129 1340
rect 16080 1300 16086 1312
rect 16117 1309 16129 1312
rect 16163 1309 16175 1343
rect 16117 1303 16175 1309
rect 16580 1343 16638 1349
rect 16580 1309 16592 1343
rect 16626 1309 16638 1343
rect 16580 1303 16638 1309
rect 16850 1300 16856 1352
rect 16908 1300 16914 1352
rect 18322 1300 18328 1352
rect 18380 1300 18386 1352
rect 18800 1349 18828 1380
rect 20717 1377 20729 1380
rect 20763 1377 20775 1411
rect 20717 1371 20775 1377
rect 20993 1411 21051 1417
rect 20993 1377 21005 1411
rect 21039 1377 21051 1411
rect 20993 1371 21051 1377
rect 18788 1343 18846 1349
rect 18788 1309 18800 1343
rect 18834 1309 18846 1343
rect 18788 1303 18846 1309
rect 19061 1343 19119 1349
rect 19061 1309 19073 1343
rect 19107 1340 19119 1343
rect 20898 1340 20904 1352
rect 19107 1312 20904 1340
rect 19107 1309 19119 1312
rect 19061 1303 19119 1309
rect 20898 1300 20904 1312
rect 20956 1300 20962 1352
rect 11296 1244 11652 1272
rect 11296 1232 11302 1244
rect 13354 1232 13360 1284
rect 13412 1232 13418 1284
rect 20530 1232 20536 1284
rect 20588 1232 20594 1284
rect 21008 1272 21036 1371
rect 21092 1340 21120 1448
rect 21284 1417 21312 1516
rect 21542 1504 21548 1556
rect 21600 1544 21606 1556
rect 21735 1547 21793 1553
rect 21735 1544 21747 1547
rect 21600 1516 21747 1544
rect 21600 1504 21606 1516
rect 21735 1513 21747 1516
rect 21781 1513 21793 1547
rect 21735 1507 21793 1513
rect 21910 1504 21916 1556
rect 21968 1544 21974 1556
rect 21968 1516 22692 1544
rect 21968 1504 21974 1516
rect 21269 1411 21327 1417
rect 21269 1377 21281 1411
rect 21315 1377 21327 1411
rect 21269 1371 21327 1377
rect 21358 1368 21364 1420
rect 21416 1408 21422 1420
rect 22462 1408 22468 1420
rect 21416 1380 22468 1408
rect 21416 1368 21422 1380
rect 22462 1368 22468 1380
rect 22520 1368 22526 1420
rect 22664 1408 22692 1516
rect 22922 1504 22928 1556
rect 22980 1504 22986 1556
rect 23477 1547 23535 1553
rect 23477 1513 23489 1547
rect 23523 1513 23535 1547
rect 23477 1507 23535 1513
rect 22940 1408 22968 1504
rect 23106 1436 23112 1488
rect 23164 1476 23170 1488
rect 23492 1476 23520 1507
rect 23658 1504 23664 1556
rect 23716 1544 23722 1556
rect 23753 1547 23811 1553
rect 23753 1544 23765 1547
rect 23716 1516 23765 1544
rect 23716 1504 23722 1516
rect 23753 1513 23765 1516
rect 23799 1513 23811 1547
rect 23753 1507 23811 1513
rect 24854 1504 24860 1556
rect 24912 1544 24918 1556
rect 26881 1547 26939 1553
rect 26881 1544 26893 1547
rect 24912 1516 26893 1544
rect 24912 1504 24918 1516
rect 26881 1513 26893 1516
rect 26927 1513 26939 1547
rect 26881 1507 26939 1513
rect 27249 1547 27307 1553
rect 27249 1513 27261 1547
rect 27295 1513 27307 1547
rect 27249 1507 27307 1513
rect 24210 1476 24216 1488
rect 23164 1448 23520 1476
rect 23768 1448 24216 1476
rect 23164 1436 23170 1448
rect 23768 1420 23796 1448
rect 24210 1436 24216 1448
rect 24268 1436 24274 1488
rect 26326 1436 26332 1488
rect 26384 1476 26390 1488
rect 27264 1476 27292 1507
rect 27522 1504 27528 1556
rect 27580 1504 27586 1556
rect 28166 1544 28172 1556
rect 27632 1516 28172 1544
rect 27632 1476 27660 1516
rect 28166 1504 28172 1516
rect 28224 1504 28230 1556
rect 28994 1504 29000 1556
rect 29052 1544 29058 1556
rect 29457 1547 29515 1553
rect 29457 1544 29469 1547
rect 29052 1516 29469 1544
rect 29052 1504 29058 1516
rect 29457 1513 29469 1516
rect 29503 1513 29515 1547
rect 29457 1507 29515 1513
rect 26384 1448 27292 1476
rect 27356 1448 27660 1476
rect 26384 1436 26390 1448
rect 23661 1411 23719 1417
rect 23661 1408 23673 1411
rect 22664 1380 22876 1408
rect 22940 1380 23673 1408
rect 21732 1343 21790 1349
rect 21732 1340 21744 1343
rect 21092 1312 21744 1340
rect 21732 1309 21744 1312
rect 21778 1309 21790 1343
rect 21732 1303 21790 1309
rect 22005 1343 22063 1349
rect 22005 1309 22017 1343
rect 22051 1340 22063 1343
rect 22738 1340 22744 1352
rect 22051 1312 22744 1340
rect 22051 1309 22063 1312
rect 22005 1303 22063 1309
rect 22738 1300 22744 1312
rect 22796 1300 22802 1352
rect 21266 1272 21272 1284
rect 21008 1244 21272 1272
rect 8996 1176 10732 1204
rect 8996 1164 9002 1176
rect 11146 1164 11152 1216
rect 11204 1204 11210 1216
rect 13372 1204 13400 1232
rect 11204 1176 13400 1204
rect 11204 1164 11210 1176
rect 13814 1164 13820 1216
rect 13872 1204 13878 1216
rect 14642 1204 14648 1216
rect 13872 1176 14648 1204
rect 13872 1164 13878 1176
rect 14642 1164 14648 1176
rect 14700 1164 14706 1216
rect 16298 1164 16304 1216
rect 16356 1204 16362 1216
rect 17770 1204 17776 1216
rect 16356 1176 17776 1204
rect 16356 1164 16362 1176
rect 17770 1164 17776 1176
rect 17828 1204 17834 1216
rect 21008 1204 21036 1244
rect 21266 1232 21272 1244
rect 21324 1232 21330 1284
rect 22848 1272 22876 1380
rect 23661 1377 23673 1380
rect 23707 1377 23719 1411
rect 23661 1371 23719 1377
rect 23676 1340 23704 1371
rect 23750 1368 23756 1420
rect 23808 1368 23814 1420
rect 23934 1368 23940 1420
rect 23992 1368 23998 1420
rect 24121 1411 24179 1417
rect 24121 1408 24133 1411
rect 24044 1380 24133 1408
rect 23952 1340 23980 1368
rect 24044 1352 24072 1380
rect 24121 1377 24133 1380
rect 24167 1377 24179 1411
rect 24228 1408 24256 1436
rect 24448 1411 24506 1417
rect 24448 1408 24460 1411
rect 24228 1380 24460 1408
rect 24121 1371 24179 1377
rect 24448 1377 24460 1380
rect 24494 1377 24506 1411
rect 24448 1371 24506 1377
rect 25314 1368 25320 1420
rect 25372 1408 25378 1420
rect 25372 1380 26562 1408
rect 25372 1368 25378 1380
rect 24617 1361 24675 1367
rect 24617 1358 24629 1361
rect 23676 1312 23980 1340
rect 24026 1300 24032 1352
rect 24084 1300 24090 1352
rect 24302 1340 24308 1352
rect 24136 1312 24308 1340
rect 23106 1272 23112 1284
rect 22848 1244 23112 1272
rect 23106 1232 23112 1244
rect 23164 1232 23170 1284
rect 23293 1275 23351 1281
rect 23293 1241 23305 1275
rect 23339 1272 23351 1275
rect 24136 1272 24164 1312
rect 24302 1300 24308 1312
rect 24360 1300 24366 1352
rect 24596 1327 24629 1358
rect 24663 1352 24675 1361
rect 24663 1327 24676 1352
rect 24596 1312 24676 1327
rect 24670 1300 24676 1312
rect 24728 1300 24734 1352
rect 24857 1343 24915 1349
rect 24857 1309 24869 1343
rect 24903 1340 24915 1343
rect 25590 1340 25596 1352
rect 24903 1312 25596 1340
rect 24903 1309 24915 1312
rect 24857 1303 24915 1309
rect 25590 1300 25596 1312
rect 25648 1300 25654 1352
rect 26534 1340 26562 1380
rect 26602 1368 26608 1420
rect 26660 1368 26666 1420
rect 27356 1417 27384 1448
rect 26697 1411 26755 1417
rect 26697 1377 26709 1411
rect 26743 1408 26755 1411
rect 27065 1411 27123 1417
rect 27065 1408 27077 1411
rect 26743 1380 27077 1408
rect 26743 1377 26755 1380
rect 26697 1371 26755 1377
rect 27065 1377 27077 1380
rect 27111 1377 27123 1411
rect 27065 1371 27123 1377
rect 27341 1411 27399 1417
rect 27341 1377 27353 1411
rect 27387 1377 27399 1411
rect 27341 1371 27399 1377
rect 26712 1340 26740 1371
rect 26534 1312 26740 1340
rect 27080 1340 27108 1371
rect 27430 1368 27436 1420
rect 27488 1408 27494 1420
rect 27617 1411 27675 1417
rect 27617 1408 27629 1411
rect 27488 1380 27629 1408
rect 27488 1368 27494 1380
rect 27617 1377 27629 1380
rect 27663 1377 27675 1411
rect 27617 1371 27675 1377
rect 27706 1368 27712 1420
rect 27764 1368 27770 1420
rect 27944 1411 28002 1417
rect 27944 1408 27956 1411
rect 27816 1380 27956 1408
rect 27724 1340 27752 1368
rect 27816 1352 27844 1380
rect 27944 1377 27956 1380
rect 27990 1377 28002 1411
rect 27944 1371 28002 1377
rect 29454 1368 29460 1420
rect 29512 1408 29518 1420
rect 30009 1411 30067 1417
rect 30009 1408 30021 1411
rect 29512 1380 30021 1408
rect 29512 1368 29518 1380
rect 30009 1377 30021 1380
rect 30055 1377 30067 1411
rect 30009 1371 30067 1377
rect 27080 1312 27752 1340
rect 27798 1300 27804 1352
rect 27856 1300 27862 1352
rect 28074 1300 28080 1352
rect 28132 1340 28138 1352
rect 28132 1312 28177 1340
rect 28132 1300 28138 1312
rect 28350 1300 28356 1352
rect 28408 1300 28414 1352
rect 29914 1300 29920 1352
rect 29972 1340 29978 1352
rect 30377 1343 30435 1349
rect 30377 1340 30389 1343
rect 29972 1312 30389 1340
rect 29972 1300 29978 1312
rect 30377 1309 30389 1312
rect 30423 1309 30435 1343
rect 30377 1303 30435 1309
rect 23339 1244 24164 1272
rect 25961 1275 26019 1281
rect 23339 1241 23351 1244
rect 23293 1235 23351 1241
rect 25961 1241 25973 1275
rect 26007 1241 26019 1275
rect 25961 1235 26019 1241
rect 17828 1176 21036 1204
rect 17828 1164 17834 1176
rect 21082 1164 21088 1216
rect 21140 1204 21146 1216
rect 25976 1204 26004 1235
rect 21140 1176 26004 1204
rect 21140 1164 21146 1176
rect 26418 1164 26424 1216
rect 26476 1164 26482 1216
rect 552 1114 30912 1136
rect 552 1062 4193 1114
rect 4245 1062 4257 1114
rect 4309 1062 4321 1114
rect 4373 1062 4385 1114
rect 4437 1062 4449 1114
rect 4501 1062 11783 1114
rect 11835 1062 11847 1114
rect 11899 1062 11911 1114
rect 11963 1062 11975 1114
rect 12027 1062 12039 1114
rect 12091 1062 19373 1114
rect 19425 1062 19437 1114
rect 19489 1062 19501 1114
rect 19553 1062 19565 1114
rect 19617 1062 19629 1114
rect 19681 1062 26963 1114
rect 27015 1062 27027 1114
rect 27079 1062 27091 1114
rect 27143 1062 27155 1114
rect 27207 1062 27219 1114
rect 27271 1062 30912 1114
rect 552 1040 30912 1062
rect 2590 960 2596 1012
rect 2648 960 2654 1012
rect 2774 960 2780 1012
rect 2832 960 2838 1012
rect 3237 1003 3295 1009
rect 3237 969 3249 1003
rect 3283 1000 3295 1003
rect 3326 1000 3332 1012
rect 3283 972 3332 1000
rect 3283 969 3295 972
rect 3237 963 3295 969
rect 3326 960 3332 972
rect 3384 960 3390 1012
rect 3605 1003 3663 1009
rect 3605 969 3617 1003
rect 3651 1000 3663 1003
rect 4614 1000 4620 1012
rect 3651 972 4620 1000
rect 3651 969 3663 972
rect 3605 963 3663 969
rect 4614 960 4620 972
rect 4672 960 4678 1012
rect 4709 1003 4767 1009
rect 4709 969 4721 1003
rect 4755 1000 4767 1003
rect 4982 1000 4988 1012
rect 4755 972 4988 1000
rect 4755 969 4767 972
rect 4709 963 4767 969
rect 4982 960 4988 972
rect 5040 960 5046 1012
rect 5074 960 5080 1012
rect 5132 960 5138 1012
rect 5166 960 5172 1012
rect 5224 960 5230 1012
rect 7282 1000 7288 1012
rect 6012 972 7288 1000
rect 2608 932 2636 960
rect 3881 935 3939 941
rect 3881 932 3893 935
rect 2608 904 3893 932
rect 3881 901 3893 904
rect 3927 901 3939 935
rect 3881 895 3939 901
rect 4157 935 4215 941
rect 4157 901 4169 935
rect 4203 932 4215 935
rect 4798 932 4804 944
rect 4203 904 4804 932
rect 4203 901 4215 904
rect 4157 895 4215 901
rect 4798 892 4804 904
rect 4856 892 4862 944
rect 5810 892 5816 944
rect 5868 892 5874 944
rect 934 824 940 876
rect 992 824 998 876
rect 1443 867 1501 873
rect 1443 833 1455 867
rect 1489 864 1501 867
rect 1489 836 1624 864
rect 1489 833 1501 836
rect 1443 827 1501 833
rect 1596 796 1624 836
rect 1670 824 1676 876
rect 1728 824 1734 876
rect 1762 824 1768 876
rect 1820 864 1826 876
rect 5442 864 5448 876
rect 1820 836 5448 864
rect 1820 824 1826 836
rect 3436 805 3464 836
rect 5442 824 5448 836
rect 5500 824 5506 876
rect 3421 799 3479 805
rect 1596 768 3188 796
rect 1403 663 1461 669
rect 1403 629 1415 663
rect 1449 660 1461 663
rect 3050 660 3056 672
rect 1449 632 3056 660
rect 1449 629 1461 632
rect 1403 623 1461 629
rect 3050 620 3056 632
rect 3108 620 3114 672
rect 3160 660 3188 768
rect 3421 765 3433 799
rect 3467 765 3479 799
rect 3421 759 3479 765
rect 3602 756 3608 808
rect 3660 796 3666 808
rect 3789 799 3847 805
rect 3789 796 3801 799
rect 3660 768 3801 796
rect 3660 756 3666 768
rect 3789 765 3801 768
rect 3835 765 3847 799
rect 3789 759 3847 765
rect 4065 799 4123 805
rect 4065 765 4077 799
rect 4111 796 4123 799
rect 4246 796 4252 808
rect 4111 768 4252 796
rect 4111 765 4123 768
rect 4065 759 4123 765
rect 3694 688 3700 740
rect 3752 728 3758 740
rect 4080 728 4108 759
rect 4246 756 4252 768
rect 4304 756 4310 808
rect 4341 799 4399 805
rect 4341 765 4353 799
rect 4387 765 4399 799
rect 4341 759 4399 765
rect 3752 700 4108 728
rect 4356 728 4384 759
rect 4430 756 4436 808
rect 4488 796 4494 808
rect 5353 799 5411 805
rect 5353 796 5365 799
rect 4488 768 5365 796
rect 4488 756 4494 768
rect 5353 765 5365 768
rect 5399 796 5411 799
rect 5534 796 5540 808
rect 5399 768 5540 796
rect 5399 765 5411 768
rect 5353 759 5411 765
rect 5534 756 5540 768
rect 5592 756 5598 808
rect 6012 805 6040 972
rect 7282 960 7288 972
rect 7340 960 7346 1012
rect 8389 1003 8447 1009
rect 8389 969 8401 1003
rect 8435 1000 8447 1003
rect 8662 1000 8668 1012
rect 8435 972 8668 1000
rect 8435 969 8447 972
rect 8389 963 8447 969
rect 8662 960 8668 972
rect 8720 960 8726 1012
rect 10502 960 10508 1012
rect 10560 960 10566 1012
rect 11330 960 11336 1012
rect 11388 1000 11394 1012
rect 11517 1003 11575 1009
rect 11517 1000 11529 1003
rect 11388 972 11529 1000
rect 11388 960 11394 972
rect 11517 969 11529 972
rect 11563 969 11575 1003
rect 11517 963 11575 969
rect 11977 1003 12035 1009
rect 11977 969 11989 1003
rect 12023 1000 12035 1003
rect 12250 1000 12256 1012
rect 12023 972 12256 1000
rect 12023 969 12035 972
rect 11977 963 12035 969
rect 12250 960 12256 972
rect 12308 960 12314 1012
rect 13170 960 13176 1012
rect 13228 960 13234 1012
rect 13541 1003 13599 1009
rect 13541 969 13553 1003
rect 13587 1000 13599 1003
rect 14182 1000 14188 1012
rect 13587 972 14188 1000
rect 13587 969 13599 972
rect 13541 963 13599 969
rect 14182 960 14188 972
rect 14240 960 14246 1012
rect 16117 1003 16175 1009
rect 16117 969 16129 1003
rect 16163 1000 16175 1003
rect 16666 1000 16672 1012
rect 16163 972 16672 1000
rect 16163 969 16175 972
rect 16117 963 16175 969
rect 16666 960 16672 972
rect 16724 960 16730 1012
rect 16850 960 16856 1012
rect 16908 1000 16914 1012
rect 18693 1003 18751 1009
rect 18693 1000 18705 1003
rect 16908 972 18705 1000
rect 16908 960 16914 972
rect 18693 969 18705 972
rect 18739 969 18751 1003
rect 18693 963 18751 969
rect 20806 960 20812 1012
rect 20864 960 20870 1012
rect 20898 960 20904 1012
rect 20956 1000 20962 1012
rect 21269 1003 21327 1009
rect 21269 1000 21281 1003
rect 20956 972 21281 1000
rect 20956 960 20962 972
rect 21269 969 21281 972
rect 21315 969 21327 1003
rect 21269 963 21327 969
rect 21542 960 21548 1012
rect 21600 1000 21606 1012
rect 23014 1000 23020 1012
rect 21600 972 23020 1000
rect 21600 960 21606 972
rect 23014 960 23020 972
rect 23072 960 23078 1012
rect 23474 960 23480 1012
rect 23532 1000 23538 1012
rect 23569 1003 23627 1009
rect 23569 1000 23581 1003
rect 23532 972 23581 1000
rect 23532 960 23538 972
rect 23569 969 23581 972
rect 23615 969 23627 1003
rect 26418 1000 26424 1012
rect 23569 963 23627 969
rect 23676 972 26424 1000
rect 10778 892 10784 944
rect 10836 932 10842 944
rect 11241 935 11299 941
rect 11241 932 11253 935
rect 10836 904 11253 932
rect 10836 892 10842 904
rect 11241 901 11253 904
rect 11287 932 11299 935
rect 12710 932 12716 944
rect 11287 904 12716 932
rect 11287 901 11299 904
rect 11241 895 11299 901
rect 12710 892 12716 904
rect 12768 892 12774 944
rect 12897 935 12955 941
rect 12897 901 12909 935
rect 12943 932 12955 935
rect 13722 932 13728 944
rect 12943 904 13728 932
rect 12943 901 12955 904
rect 12897 895 12955 901
rect 13722 892 13728 904
rect 13780 892 13786 944
rect 16390 892 16396 944
rect 16448 892 16454 944
rect 18417 935 18475 941
rect 18417 901 18429 935
rect 18463 932 18475 935
rect 18966 932 18972 944
rect 18463 904 18972 932
rect 18463 901 18475 904
rect 18417 895 18475 901
rect 18966 892 18972 904
rect 19024 892 19030 944
rect 23676 932 23704 972
rect 26418 960 26424 972
rect 26476 960 26482 1012
rect 26602 960 26608 1012
rect 26660 960 26666 1012
rect 28534 960 28540 1012
rect 28592 960 28598 1012
rect 29454 960 29460 1012
rect 29512 1000 29518 1012
rect 29825 1003 29883 1009
rect 29825 1000 29837 1003
rect 29512 972 29837 1000
rect 29512 960 29518 972
rect 29825 969 29837 972
rect 29871 1000 29883 1003
rect 30193 1003 30251 1009
rect 30193 1000 30205 1003
rect 29871 972 30205 1000
rect 29871 969 29883 972
rect 29825 963 29883 969
rect 30193 969 30205 972
rect 30239 969 30251 1003
rect 30193 963 30251 969
rect 23492 904 23704 932
rect 6270 824 6276 876
rect 6328 864 6334 876
rect 6416 867 6474 873
rect 6638 871 6644 876
rect 6416 864 6428 867
rect 6328 836 6428 864
rect 6328 824 6334 836
rect 6416 833 6428 836
rect 6462 833 6474 867
rect 6416 827 6474 833
rect 6595 865 6644 871
rect 6595 831 6607 865
rect 6641 831 6644 865
rect 6595 825 6644 831
rect 6638 824 6644 825
rect 6696 824 6702 876
rect 6730 824 6736 876
rect 6788 864 6794 876
rect 6825 867 6883 873
rect 6825 864 6837 867
rect 6788 836 6837 864
rect 6788 824 6794 836
rect 6825 833 6837 836
rect 6871 833 6883 867
rect 6825 827 6883 833
rect 8205 867 8263 873
rect 8205 833 8217 867
rect 8251 864 8263 867
rect 8846 864 8852 876
rect 8251 836 8852 864
rect 8251 833 8263 836
rect 8205 827 8263 833
rect 8846 824 8852 836
rect 8904 824 8910 876
rect 9214 871 9220 876
rect 9171 865 9220 871
rect 9171 831 9183 865
rect 9217 831 9220 865
rect 9171 825 9220 831
rect 9214 824 9220 825
rect 9272 824 9278 876
rect 11146 864 11152 876
rect 9324 836 11152 864
rect 5629 799 5687 805
rect 5629 765 5641 799
rect 5675 796 5687 799
rect 5997 799 6055 805
rect 5997 796 6009 799
rect 5675 768 6009 796
rect 5675 765 5687 768
rect 5629 759 5687 765
rect 5997 765 6009 768
rect 6043 765 6055 799
rect 5997 759 6055 765
rect 6086 756 6092 808
rect 6144 756 6150 808
rect 8294 756 8300 808
rect 8352 796 8358 808
rect 9030 805 9036 808
rect 8573 799 8631 805
rect 8573 796 8585 799
rect 8352 768 8585 796
rect 8352 756 8358 768
rect 8573 765 8585 768
rect 8619 765 8631 799
rect 8573 759 8631 765
rect 8665 799 8723 805
rect 8665 765 8677 799
rect 8711 765 8723 799
rect 8665 759 8723 765
rect 8992 799 9036 805
rect 8992 765 9004 799
rect 9088 796 9094 808
rect 9324 796 9352 836
rect 11146 824 11152 836
rect 11204 824 11210 876
rect 11514 824 11520 876
rect 11572 864 11578 876
rect 13817 867 13875 873
rect 13817 864 13829 867
rect 11572 836 13829 864
rect 11572 824 11578 836
rect 13817 833 13829 836
rect 13863 833 13875 867
rect 13817 827 13875 833
rect 9088 768 9352 796
rect 9401 799 9459 805
rect 8992 759 9036 765
rect 5902 728 5908 740
rect 4356 700 5908 728
rect 3752 688 3758 700
rect 5902 688 5908 700
rect 5960 688 5966 740
rect 8386 688 8392 740
rect 8444 728 8450 740
rect 8680 728 8708 759
rect 9030 756 9036 759
rect 9088 756 9094 768
rect 9401 765 9413 799
rect 9447 796 9459 799
rect 10778 796 10784 808
rect 9447 768 10784 796
rect 9447 765 9459 768
rect 9401 759 9459 765
rect 10778 756 10784 768
rect 10836 756 10842 808
rect 11422 756 11428 808
rect 11480 796 11486 808
rect 12250 796 12256 808
rect 11480 768 12256 796
rect 11480 756 11486 768
rect 12250 756 12256 768
rect 12308 756 12314 808
rect 12434 756 12440 808
rect 12492 796 12498 808
rect 13081 799 13139 805
rect 13081 796 13093 799
rect 12492 768 13093 796
rect 12492 756 12498 768
rect 13081 765 13093 768
rect 13127 765 13139 799
rect 13081 759 13139 765
rect 13354 756 13360 808
rect 13412 756 13418 808
rect 13538 756 13544 808
rect 13596 796 13602 808
rect 13725 799 13783 805
rect 13725 796 13737 799
rect 13596 768 13737 796
rect 13596 756 13602 768
rect 13725 765 13737 768
rect 13771 765 13783 799
rect 13832 796 13860 827
rect 14274 824 14280 876
rect 14332 871 14338 876
rect 14332 865 14381 871
rect 14332 831 14335 865
rect 14369 831 14381 865
rect 16408 864 16436 892
rect 16856 867 16914 873
rect 16856 864 16868 867
rect 16408 836 16868 864
rect 14332 825 14381 831
rect 16856 833 16868 836
rect 16902 833 16914 867
rect 16856 827 16914 833
rect 14332 824 14338 825
rect 17126 824 17132 876
rect 17184 824 17190 876
rect 17862 824 17868 876
rect 17920 824 17926 876
rect 19334 873 19340 876
rect 19296 867 19340 873
rect 19296 833 19308 867
rect 19296 827 19340 833
rect 19334 824 19340 827
rect 19392 824 19398 876
rect 19475 867 19533 873
rect 19475 833 19487 867
rect 19521 864 19533 867
rect 19521 836 19656 864
rect 19521 833 19533 836
rect 19475 827 19533 833
rect 14458 796 14464 808
rect 13832 768 14464 796
rect 13725 759 13783 765
rect 14458 756 14464 768
rect 14516 756 14522 808
rect 14550 756 14556 808
rect 14608 756 14614 808
rect 16298 756 16304 808
rect 16356 756 16362 808
rect 16390 756 16396 808
rect 16448 756 16454 808
rect 17880 796 17908 824
rect 16500 768 17908 796
rect 18877 799 18935 805
rect 8444 700 8708 728
rect 8444 688 8450 700
rect 10962 688 10968 740
rect 11020 728 11026 740
rect 12158 728 12164 740
rect 11020 700 12164 728
rect 11020 688 11026 700
rect 12158 688 12164 700
rect 12216 688 12222 740
rect 16500 728 16528 768
rect 18877 765 18889 799
rect 18923 765 18935 799
rect 18877 759 18935 765
rect 18969 799 19027 805
rect 18969 765 18981 799
rect 19015 796 19027 799
rect 19628 796 19656 836
rect 19702 824 19708 876
rect 19760 824 19766 876
rect 21358 824 21364 876
rect 21416 824 21422 876
rect 21545 867 21603 873
rect 21545 833 21557 867
rect 21591 864 21603 867
rect 22051 867 22109 873
rect 21591 836 21680 864
rect 21591 833 21603 836
rect 21545 827 21603 833
rect 21376 796 21404 824
rect 19015 768 19104 796
rect 19628 768 21404 796
rect 21453 799 21511 805
rect 19015 765 19027 768
rect 18969 759 19027 765
rect 12268 700 12940 728
rect 4706 660 4712 672
rect 3160 632 4712 660
rect 4706 620 4712 632
rect 4764 620 4770 672
rect 5445 663 5503 669
rect 5445 629 5457 663
rect 5491 660 5503 663
rect 10778 660 10784 672
rect 5491 632 10784 660
rect 5491 629 5503 632
rect 5445 623 5503 629
rect 10778 620 10784 632
rect 10836 620 10842 672
rect 11146 620 11152 672
rect 11204 660 11210 672
rect 12268 660 12296 700
rect 11204 632 12296 660
rect 11204 620 11210 632
rect 12802 620 12808 672
rect 12860 620 12866 672
rect 12912 660 12940 700
rect 15212 700 16528 728
rect 14283 663 14341 669
rect 14283 660 14295 663
rect 12912 632 14295 660
rect 14283 629 14295 632
rect 14329 660 14341 663
rect 15212 660 15240 700
rect 14329 632 15240 660
rect 14329 629 14341 632
rect 14283 623 14341 629
rect 15286 620 15292 672
rect 15344 660 15350 672
rect 15657 663 15715 669
rect 15657 660 15669 663
rect 15344 632 15669 660
rect 15344 620 15350 632
rect 15657 629 15669 632
rect 15703 629 15715 663
rect 15657 623 15715 629
rect 16758 620 16764 672
rect 16816 660 16822 672
rect 16859 663 16917 669
rect 16859 660 16871 663
rect 16816 632 16871 660
rect 16816 620 16822 632
rect 16859 629 16871 632
rect 16905 660 16917 663
rect 17862 660 17868 672
rect 16905 632 17868 660
rect 16905 629 16917 632
rect 16859 623 16917 629
rect 17862 620 17868 632
rect 17920 620 17926 672
rect 18892 660 18920 759
rect 19076 740 19104 768
rect 21453 765 21465 799
rect 21499 765 21511 799
rect 21453 759 21511 765
rect 19058 688 19064 740
rect 19116 688 19122 740
rect 21468 728 21496 759
rect 21542 728 21548 740
rect 21379 700 21548 728
rect 21379 660 21407 700
rect 21542 688 21548 700
rect 21600 688 21606 740
rect 18892 632 21407 660
rect 21652 660 21680 836
rect 22051 833 22063 867
rect 22097 864 22109 867
rect 22186 864 22192 876
rect 22097 836 22192 864
rect 22097 833 22109 836
rect 22051 827 22109 833
rect 22186 824 22192 836
rect 22244 824 22250 876
rect 22281 867 22339 873
rect 22281 833 22293 867
rect 22327 864 22339 867
rect 23492 864 23520 904
rect 26694 892 26700 944
rect 26752 892 26758 944
rect 22327 836 23520 864
rect 22327 833 22339 836
rect 22281 827 22339 833
rect 23842 824 23848 876
rect 23900 824 23906 876
rect 24302 824 24308 876
rect 24360 864 24366 876
rect 24581 867 24639 873
rect 24360 836 24405 864
rect 24360 824 24366 836
rect 24581 833 24593 867
rect 24627 833 24639 867
rect 24581 827 24639 833
rect 21872 799 21930 805
rect 21872 765 21884 799
rect 21918 796 21930 799
rect 21918 768 23980 796
rect 21918 765 21930 768
rect 21872 759 21930 765
rect 23842 688 23848 740
rect 23900 688 23906 740
rect 23860 660 23888 688
rect 21652 632 23888 660
rect 23952 660 23980 768
rect 24394 756 24400 808
rect 24452 796 24458 808
rect 24596 796 24624 827
rect 25222 824 25228 876
rect 25280 864 25286 876
rect 26712 864 26740 892
rect 27160 867 27218 873
rect 27160 864 27172 867
rect 25280 836 26280 864
rect 26712 836 27172 864
rect 25280 824 25286 836
rect 26252 805 26280 836
rect 27160 833 27172 836
rect 27206 833 27218 867
rect 27160 827 27218 833
rect 27338 824 27344 876
rect 27396 824 27402 876
rect 27433 867 27491 873
rect 27433 833 27445 867
rect 27479 864 27491 867
rect 29270 864 29276 876
rect 27479 836 29276 864
rect 27479 833 27491 836
rect 27433 827 27491 833
rect 29270 824 29276 836
rect 29328 824 29334 876
rect 24452 768 24624 796
rect 26237 799 26295 805
rect 24452 756 24458 768
rect 26237 765 26249 799
rect 26283 765 26295 799
rect 26237 759 26295 765
rect 26421 799 26479 805
rect 26421 765 26433 799
rect 26467 796 26479 799
rect 26510 796 26516 808
rect 26467 768 26516 796
rect 26467 765 26479 768
rect 26421 759 26479 765
rect 26510 756 26516 768
rect 26568 756 26574 808
rect 26697 799 26755 805
rect 26697 765 26709 799
rect 26743 796 26755 799
rect 27356 796 27384 824
rect 26743 768 27384 796
rect 26743 765 26755 768
rect 26697 759 26755 765
rect 28626 756 28632 808
rect 28684 796 28690 808
rect 28997 799 29055 805
rect 28997 796 29009 799
rect 28684 768 29009 796
rect 28684 756 28690 768
rect 28997 765 29009 768
rect 29043 765 29055 799
rect 28997 759 29055 765
rect 24118 660 24124 672
rect 23952 632 24124 660
rect 24118 620 24124 632
rect 24176 660 24182 672
rect 24311 663 24369 669
rect 24311 660 24323 663
rect 24176 632 24323 660
rect 24176 620 24182 632
rect 24311 629 24323 632
rect 24357 629 24369 663
rect 24311 623 24369 629
rect 25682 620 25688 672
rect 25740 620 25746 672
rect 26050 620 26056 672
rect 26108 620 26114 672
rect 26234 620 26240 672
rect 26292 660 26298 672
rect 27163 663 27221 669
rect 27163 660 27175 663
rect 26292 632 27175 660
rect 26292 620 26298 632
rect 27163 629 27175 632
rect 27209 660 27221 663
rect 27798 660 27804 672
rect 27209 632 27804 660
rect 27209 629 27221 632
rect 27163 623 27221 629
rect 27798 620 27804 632
rect 27856 620 27862 672
rect 29178 620 29184 672
rect 29236 620 29242 672
rect 552 570 31072 592
rect 552 518 7988 570
rect 8040 518 8052 570
rect 8104 518 8116 570
rect 8168 518 8180 570
rect 8232 518 8244 570
rect 8296 518 15578 570
rect 15630 518 15642 570
rect 15694 518 15706 570
rect 15758 518 15770 570
rect 15822 518 15834 570
rect 15886 518 23168 570
rect 23220 518 23232 570
rect 23284 518 23296 570
rect 23348 518 23360 570
rect 23412 518 23424 570
rect 23476 518 30758 570
rect 30810 518 30822 570
rect 30874 518 30886 570
rect 30938 518 30950 570
rect 31002 518 31014 570
rect 31066 518 31072 570
rect 552 496 31072 518
rect 3050 416 3056 468
rect 3108 456 3114 468
rect 5718 456 5724 468
rect 3108 428 5724 456
rect 3108 416 3114 428
rect 5718 416 5724 428
rect 5776 416 5782 468
rect 5810 416 5816 468
rect 5868 456 5874 468
rect 14366 456 14372 468
rect 5868 428 14372 456
rect 5868 416 5874 428
rect 14366 416 14372 428
rect 14424 416 14430 468
rect 14550 416 14556 468
rect 14608 456 14614 468
rect 26050 456 26056 468
rect 14608 428 26056 456
rect 14608 416 14614 428
rect 26050 416 26056 428
rect 26108 416 26114 468
rect 3510 348 3516 400
rect 3568 388 3574 400
rect 8386 388 8392 400
rect 3568 360 8392 388
rect 3568 348 3574 360
rect 8386 348 8392 360
rect 8444 388 8450 400
rect 8444 360 11100 388
rect 8444 348 8450 360
rect 3878 280 3884 332
rect 3936 320 3942 332
rect 9030 320 9036 332
rect 3936 292 9036 320
rect 3936 280 3942 292
rect 9030 280 9036 292
rect 9088 280 9094 332
rect 11072 320 11100 360
rect 12802 348 12808 400
rect 12860 388 12866 400
rect 19058 388 19064 400
rect 12860 360 19064 388
rect 12860 348 12866 360
rect 19058 348 19064 360
rect 19116 388 19122 400
rect 24486 388 24492 400
rect 19116 360 24492 388
rect 19116 348 19122 360
rect 24486 348 24492 360
rect 24544 348 24550 400
rect 25682 348 25688 400
rect 25740 348 25746 400
rect 11514 320 11520 332
rect 11072 292 11520 320
rect 11514 280 11520 292
rect 11572 280 11578 332
rect 14274 280 14280 332
rect 14332 320 14338 332
rect 25700 320 25728 348
rect 14332 292 25728 320
rect 14332 280 14338 292
rect 11330 212 11336 264
rect 11388 212 11394 264
rect 12710 212 12716 264
rect 12768 252 12774 264
rect 15562 252 15568 264
rect 12768 224 15568 252
rect 12768 212 12774 224
rect 15562 212 15568 224
rect 15620 212 15626 264
rect 24026 252 24032 264
rect 16592 224 24032 252
rect 1302 144 1308 196
rect 1360 184 1366 196
rect 6086 184 6092 196
rect 1360 156 6092 184
rect 1360 144 1366 156
rect 6086 144 6092 156
rect 6144 144 6150 196
rect 11348 116 11376 212
rect 12250 144 12256 196
rect 12308 184 12314 196
rect 12308 156 13768 184
rect 12308 144 12314 156
rect 13740 116 13768 156
rect 14458 144 14464 196
rect 14516 184 14522 196
rect 16592 184 16620 224
rect 24026 212 24032 224
rect 24084 212 24090 264
rect 14516 156 16620 184
rect 14516 144 14522 156
rect 17862 144 17868 196
rect 17920 184 17926 196
rect 26234 184 26240 196
rect 17920 156 26240 184
rect 17920 144 17926 156
rect 26234 144 26240 156
rect 26292 144 26298 196
rect 15470 116 15476 128
rect 11348 88 13676 116
rect 13740 88 15476 116
rect 5534 8 5540 60
rect 5592 48 5598 60
rect 12434 48 12440 60
rect 5592 20 12440 48
rect 5592 8 5598 20
rect 12434 8 12440 20
rect 12492 8 12498 60
rect 13648 48 13676 88
rect 15470 76 15476 88
rect 15528 76 15534 128
rect 16390 48 16396 60
rect 13648 20 16396 48
rect 16390 8 16396 20
rect 16448 8 16454 60
<< via1 >>
rect 7656 22244 7708 22296
rect 7748 22244 7800 22296
rect 14924 22244 14976 22296
rect 22284 22244 22336 22296
rect 22376 22244 22428 22296
rect 23664 22244 23716 22296
rect 23756 22244 23808 22296
rect 28540 22244 28592 22296
rect 5356 22176 5408 22228
rect 5448 22176 5500 22228
rect 14372 22176 14424 22228
rect 18972 22176 19024 22228
rect 21732 22176 21784 22228
rect 30380 22176 30432 22228
rect 1768 22108 1820 22160
rect 7288 22108 7340 22160
rect 7656 22108 7708 22160
rect 9956 22108 10008 22160
rect 13176 22108 13228 22160
rect 22468 22108 22520 22160
rect 22744 22108 22796 22160
rect 25596 22108 25648 22160
rect 3608 22040 3660 22092
rect 1952 21972 2004 22024
rect 7748 21972 7800 22024
rect 3976 21904 4028 21956
rect 12716 21972 12768 22024
rect 12900 21972 12952 22024
rect 13084 21972 13136 22024
rect 18512 22040 18564 22092
rect 18604 22040 18656 22092
rect 23756 22040 23808 22092
rect 25044 22040 25096 22092
rect 14004 21972 14056 22024
rect 16672 21972 16724 22024
rect 21824 21972 21876 22024
rect 1676 21836 1728 21888
rect 4988 21836 5040 21888
rect 6828 21836 6880 21888
rect 17316 21904 17368 21956
rect 20812 21904 20864 21956
rect 21364 21904 21416 21956
rect 27896 21972 27948 22024
rect 31208 21972 31260 22024
rect 22836 21904 22888 21956
rect 25780 21904 25832 21956
rect 8392 21836 8444 21888
rect 10692 21836 10744 21888
rect 10968 21836 11020 21888
rect 20720 21836 20772 21888
rect 21456 21836 21508 21888
rect 22376 21836 22428 21888
rect 22560 21836 22612 21888
rect 25872 21836 25924 21888
rect 4193 21734 4245 21786
rect 4257 21734 4309 21786
rect 4321 21734 4373 21786
rect 4385 21734 4437 21786
rect 4449 21734 4501 21786
rect 11783 21734 11835 21786
rect 11847 21734 11899 21786
rect 11911 21734 11963 21786
rect 11975 21734 12027 21786
rect 12039 21734 12091 21786
rect 19373 21734 19425 21786
rect 19437 21734 19489 21786
rect 19501 21734 19553 21786
rect 19565 21734 19617 21786
rect 19629 21734 19681 21786
rect 26963 21734 27015 21786
rect 27027 21734 27079 21786
rect 27091 21734 27143 21786
rect 27155 21734 27207 21786
rect 27219 21734 27271 21786
rect 8576 21632 8628 21684
rect 7288 21564 7340 21616
rect 10140 21632 10192 21684
rect 10232 21632 10284 21684
rect 13176 21675 13228 21684
rect 13176 21641 13185 21675
rect 13185 21641 13219 21675
rect 13219 21641 13228 21675
rect 13176 21632 13228 21641
rect 3148 21496 3200 21548
rect 4068 21496 4120 21548
rect 5356 21496 5408 21548
rect 1216 21428 1268 21480
rect 1676 21471 1728 21480
rect 1676 21437 1685 21471
rect 1685 21437 1719 21471
rect 1719 21437 1728 21471
rect 1676 21428 1728 21437
rect 2780 21428 2832 21480
rect 5264 21428 5316 21480
rect 6000 21496 6052 21548
rect 9128 21539 9180 21548
rect 9128 21505 9140 21539
rect 9140 21505 9174 21539
rect 9174 21505 9180 21539
rect 9128 21496 9180 21505
rect 10784 21496 10836 21548
rect 5540 21428 5592 21480
rect 6552 21471 6604 21480
rect 6552 21437 6561 21471
rect 6561 21437 6595 21471
rect 6595 21437 6604 21471
rect 6552 21428 6604 21437
rect 7196 21428 7248 21480
rect 8300 21428 8352 21480
rect 3056 21403 3108 21412
rect 3056 21369 3065 21403
rect 3065 21369 3099 21403
rect 3099 21369 3108 21403
rect 3056 21360 3108 21369
rect 5356 21360 5408 21412
rect 2320 21292 2372 21344
rect 5908 21360 5960 21412
rect 7288 21292 7340 21344
rect 7840 21335 7892 21344
rect 7840 21301 7849 21335
rect 7849 21301 7883 21335
rect 7883 21301 7892 21335
rect 7840 21292 7892 21301
rect 8392 21360 8444 21412
rect 8668 21471 8720 21480
rect 8668 21437 8677 21471
rect 8677 21437 8711 21471
rect 8711 21437 8720 21471
rect 8668 21428 8720 21437
rect 9220 21428 9272 21480
rect 10048 21428 10100 21480
rect 10968 21471 11020 21480
rect 10968 21437 10977 21471
rect 10977 21437 11011 21471
rect 11011 21437 11020 21471
rect 10968 21428 11020 21437
rect 12992 21496 13044 21548
rect 14188 21496 14240 21548
rect 8760 21360 8812 21412
rect 10600 21360 10652 21412
rect 11704 21471 11756 21480
rect 11704 21437 11713 21471
rect 11713 21437 11747 21471
rect 11747 21437 11756 21471
rect 11704 21428 11756 21437
rect 13084 21428 13136 21480
rect 13544 21471 13596 21480
rect 13544 21437 13553 21471
rect 13553 21437 13587 21471
rect 13587 21437 13596 21471
rect 13544 21428 13596 21437
rect 13268 21360 13320 21412
rect 15752 21632 15804 21684
rect 21916 21632 21968 21684
rect 15384 21496 15436 21548
rect 17960 21564 18012 21616
rect 18604 21564 18656 21616
rect 20720 21607 20772 21616
rect 20720 21573 20729 21607
rect 20729 21573 20763 21607
rect 20763 21573 20772 21607
rect 20720 21564 20772 21573
rect 20812 21564 20864 21616
rect 25596 21632 25648 21684
rect 25964 21632 26016 21684
rect 15016 21428 15068 21480
rect 15752 21471 15804 21480
rect 15752 21437 15761 21471
rect 15761 21437 15795 21471
rect 15795 21437 15804 21471
rect 15752 21428 15804 21437
rect 16120 21471 16172 21480
rect 16120 21437 16129 21471
rect 16129 21437 16163 21471
rect 16163 21437 16172 21471
rect 16120 21428 16172 21437
rect 17684 21428 17736 21480
rect 18328 21428 18380 21480
rect 19064 21428 19116 21480
rect 19340 21428 19392 21480
rect 20444 21428 20496 21480
rect 16212 21360 16264 21412
rect 17960 21403 18012 21412
rect 17960 21369 17969 21403
rect 17969 21369 18003 21403
rect 18003 21369 18012 21403
rect 17960 21360 18012 21369
rect 8944 21292 8996 21344
rect 10324 21292 10376 21344
rect 10508 21335 10560 21344
rect 10508 21301 10517 21335
rect 10517 21301 10551 21335
rect 10551 21301 10560 21335
rect 10508 21292 10560 21301
rect 10968 21292 11020 21344
rect 12808 21335 12860 21344
rect 12808 21301 12817 21335
rect 12817 21301 12851 21335
rect 12851 21301 12860 21335
rect 12808 21292 12860 21301
rect 14004 21335 14056 21344
rect 14004 21301 14019 21335
rect 14019 21301 14053 21335
rect 14053 21301 14056 21335
rect 14004 21292 14056 21301
rect 15476 21292 15528 21344
rect 17592 21292 17644 21344
rect 18236 21292 18288 21344
rect 20076 21335 20128 21344
rect 20076 21301 20085 21335
rect 20085 21301 20119 21335
rect 20119 21301 20128 21335
rect 20076 21292 20128 21301
rect 20812 21292 20864 21344
rect 21456 21539 21508 21548
rect 21456 21505 21465 21539
rect 21465 21505 21499 21539
rect 21499 21505 21508 21539
rect 21456 21496 21508 21505
rect 22008 21496 22060 21548
rect 23296 21496 23348 21548
rect 24492 21539 24544 21548
rect 24492 21505 24501 21539
rect 24501 21505 24535 21539
rect 24535 21505 24544 21539
rect 24492 21496 24544 21505
rect 25504 21564 25556 21616
rect 29460 21632 29512 21684
rect 30380 21675 30432 21684
rect 30380 21641 30389 21675
rect 30389 21641 30423 21675
rect 30423 21641 30432 21675
rect 30380 21632 30432 21641
rect 22192 21471 22244 21480
rect 22192 21437 22201 21471
rect 22201 21437 22235 21471
rect 22235 21437 22244 21471
rect 22192 21428 22244 21437
rect 22309 21471 22361 21480
rect 22309 21437 22318 21471
rect 22318 21437 22352 21471
rect 22352 21437 22361 21471
rect 22309 21428 22361 21437
rect 23112 21428 23164 21480
rect 23572 21428 23624 21480
rect 23848 21471 23900 21480
rect 23848 21437 23857 21471
rect 23857 21437 23891 21471
rect 23891 21437 23900 21471
rect 23848 21428 23900 21437
rect 23940 21428 23992 21480
rect 24768 21471 24820 21480
rect 24768 21437 24777 21471
rect 24777 21437 24811 21471
rect 24811 21437 24820 21471
rect 24768 21428 24820 21437
rect 24952 21428 25004 21480
rect 25044 21471 25096 21480
rect 25044 21437 25053 21471
rect 25053 21437 25087 21471
rect 25087 21437 25096 21471
rect 25044 21428 25096 21437
rect 25780 21471 25832 21480
rect 25780 21437 25789 21471
rect 25789 21437 25823 21471
rect 25823 21437 25832 21471
rect 25780 21428 25832 21437
rect 26056 21428 26108 21480
rect 26700 21471 26752 21480
rect 26700 21437 26709 21471
rect 26709 21437 26743 21471
rect 26743 21437 26752 21471
rect 26700 21428 26752 21437
rect 29092 21471 29144 21480
rect 29092 21437 29101 21471
rect 29101 21437 29135 21471
rect 29135 21437 29144 21471
rect 29092 21428 29144 21437
rect 29276 21471 29328 21480
rect 29276 21437 29285 21471
rect 29285 21437 29319 21471
rect 29319 21437 29328 21471
rect 29276 21428 29328 21437
rect 29828 21496 29880 21548
rect 31116 21496 31168 21548
rect 28448 21360 28500 21412
rect 22008 21292 22060 21344
rect 23112 21335 23164 21344
rect 23112 21301 23121 21335
rect 23121 21301 23155 21335
rect 23155 21301 23164 21335
rect 23112 21292 23164 21301
rect 23756 21292 23808 21344
rect 23940 21292 23992 21344
rect 25320 21292 25372 21344
rect 25688 21335 25740 21344
rect 25688 21301 25697 21335
rect 25697 21301 25731 21335
rect 25731 21301 25740 21335
rect 25688 21292 25740 21301
rect 27804 21335 27856 21344
rect 27804 21301 27813 21335
rect 27813 21301 27847 21335
rect 27847 21301 27856 21335
rect 27804 21292 27856 21301
rect 28356 21335 28408 21344
rect 28356 21301 28365 21335
rect 28365 21301 28399 21335
rect 28399 21301 28408 21335
rect 28356 21292 28408 21301
rect 30104 21292 30156 21344
rect 7988 21190 8040 21242
rect 8052 21190 8104 21242
rect 8116 21190 8168 21242
rect 8180 21190 8232 21242
rect 8244 21190 8296 21242
rect 15578 21190 15630 21242
rect 15642 21190 15694 21242
rect 15706 21190 15758 21242
rect 15770 21190 15822 21242
rect 15834 21190 15886 21242
rect 23168 21190 23220 21242
rect 23232 21190 23284 21242
rect 23296 21190 23348 21242
rect 23360 21190 23412 21242
rect 23424 21190 23476 21242
rect 30758 21190 30810 21242
rect 30822 21190 30874 21242
rect 30886 21190 30938 21242
rect 30950 21190 31002 21242
rect 31014 21190 31066 21242
rect 1768 21131 1820 21140
rect 1768 21097 1783 21131
rect 1783 21097 1817 21131
rect 1817 21097 1820 21131
rect 1768 21088 1820 21097
rect 5816 21088 5868 21140
rect 5908 21088 5960 21140
rect 5264 21020 5316 21072
rect 8668 21088 8720 21140
rect 9496 21088 9548 21140
rect 9772 21088 9824 21140
rect 11520 21088 11572 21140
rect 11612 21088 11664 21140
rect 14924 21088 14976 21140
rect 16672 21088 16724 21140
rect 19064 21088 19116 21140
rect 20168 21088 20220 21140
rect 20812 21131 20864 21140
rect 20812 21097 20821 21131
rect 20821 21097 20855 21131
rect 20855 21097 20864 21131
rect 20812 21088 20864 21097
rect 22192 21088 22244 21140
rect 23388 21088 23440 21140
rect 25044 21088 25096 21140
rect 25320 21131 25372 21140
rect 25320 21097 25329 21131
rect 25329 21097 25363 21131
rect 25363 21097 25372 21131
rect 25320 21088 25372 21097
rect 25504 21088 25556 21140
rect 27896 21088 27948 21140
rect 10232 21020 10284 21072
rect 10416 21063 10468 21072
rect 10416 21029 10425 21063
rect 10425 21029 10459 21063
rect 10459 21029 10468 21063
rect 10416 21020 10468 21029
rect 10876 21020 10928 21072
rect 12900 21020 12952 21072
rect 756 20884 808 20936
rect 5540 20952 5592 21004
rect 1492 20884 1544 20936
rect 2412 20884 2464 20936
rect 3700 20884 3752 20936
rect 3976 20927 4028 20936
rect 3976 20893 3988 20927
rect 3988 20893 4022 20927
rect 4022 20893 4028 20927
rect 3976 20884 4028 20893
rect 4252 20927 4304 20936
rect 4252 20893 4261 20927
rect 4261 20893 4295 20927
rect 4295 20893 4304 20927
rect 4252 20884 4304 20893
rect 5816 20995 5868 21004
rect 5816 20961 5825 20995
rect 5825 20961 5859 20995
rect 5859 20961 5868 20995
rect 5816 20952 5868 20961
rect 6460 20884 6512 20936
rect 6736 20884 6788 20936
rect 7472 20952 7524 21004
rect 8576 20952 8628 21004
rect 9588 20952 9640 21004
rect 10692 20952 10744 21004
rect 7840 20884 7892 20936
rect 8392 20884 8444 20936
rect 8852 20884 8904 20936
rect 9496 20884 9548 20936
rect 11152 20884 11204 20936
rect 11244 20927 11296 20936
rect 11244 20893 11253 20927
rect 11253 20893 11287 20927
rect 11287 20893 11296 20927
rect 11244 20884 11296 20893
rect 11520 20884 11572 20936
rect 11796 20884 11848 20936
rect 14004 20952 14056 21004
rect 15108 20952 15160 21004
rect 15752 20995 15804 21004
rect 15752 20961 15761 20995
rect 15761 20961 15795 20995
rect 15795 20961 15804 20995
rect 15752 20952 15804 20961
rect 16028 20952 16080 21004
rect 16488 20952 16540 21004
rect 18328 21020 18380 21072
rect 19340 21020 19392 21072
rect 20260 21020 20312 21072
rect 25228 21020 25280 21072
rect 26148 21020 26200 21072
rect 18788 20952 18840 21004
rect 18972 20995 19024 21004
rect 18972 20961 18981 20995
rect 18981 20961 19015 20995
rect 19015 20961 19024 20995
rect 18972 20952 19024 20961
rect 13360 20884 13412 20936
rect 848 20748 900 20800
rect 2688 20748 2740 20800
rect 4712 20748 4764 20800
rect 7656 20791 7708 20800
rect 7656 20757 7665 20791
rect 7665 20757 7699 20791
rect 7699 20757 7708 20791
rect 7656 20748 7708 20757
rect 12992 20816 13044 20868
rect 14096 20884 14148 20936
rect 14280 20884 14332 20936
rect 15016 20884 15068 20936
rect 16120 20927 16172 20936
rect 16120 20893 16129 20927
rect 16129 20893 16163 20927
rect 16163 20893 16172 20927
rect 16120 20884 16172 20893
rect 19248 20927 19300 20936
rect 19248 20893 19257 20927
rect 19257 20893 19291 20927
rect 19291 20893 19300 20927
rect 22560 20952 22612 21004
rect 19248 20884 19300 20893
rect 21180 20884 21232 20936
rect 17684 20859 17736 20868
rect 17684 20825 17693 20859
rect 17693 20825 17727 20859
rect 17727 20825 17736 20859
rect 17684 20816 17736 20825
rect 11796 20748 11848 20800
rect 18052 20791 18104 20800
rect 18052 20757 18061 20791
rect 18061 20757 18095 20791
rect 18095 20757 18104 20791
rect 18052 20748 18104 20757
rect 18696 20748 18748 20800
rect 22652 20816 22704 20868
rect 25780 20995 25832 21004
rect 25780 20961 25789 20995
rect 25789 20961 25823 20995
rect 25823 20961 25832 20995
rect 25780 20952 25832 20961
rect 25872 20952 25924 21004
rect 27344 20952 27396 21004
rect 26056 20884 26108 20936
rect 26424 20927 26476 20936
rect 26424 20893 26433 20927
rect 26433 20893 26467 20927
rect 26467 20893 26476 20927
rect 26424 20884 26476 20893
rect 26792 20884 26844 20936
rect 28632 20927 28684 20936
rect 28632 20893 28644 20927
rect 28644 20893 28678 20927
rect 28678 20893 28684 20927
rect 28632 20884 28684 20893
rect 30472 20884 30524 20936
rect 25964 20859 26016 20868
rect 25964 20825 25973 20859
rect 25973 20825 26007 20859
rect 26007 20825 26016 20859
rect 25964 20816 26016 20825
rect 23572 20748 23624 20800
rect 24124 20748 24176 20800
rect 29736 20816 29788 20868
rect 26608 20748 26660 20800
rect 4193 20646 4245 20698
rect 4257 20646 4309 20698
rect 4321 20646 4373 20698
rect 4385 20646 4437 20698
rect 4449 20646 4501 20698
rect 11783 20646 11835 20698
rect 11847 20646 11899 20698
rect 11911 20646 11963 20698
rect 11975 20646 12027 20698
rect 12039 20646 12091 20698
rect 19373 20646 19425 20698
rect 19437 20646 19489 20698
rect 19501 20646 19553 20698
rect 19565 20646 19617 20698
rect 19629 20646 19681 20698
rect 26963 20646 27015 20698
rect 27027 20646 27079 20698
rect 27091 20646 27143 20698
rect 27155 20646 27207 20698
rect 27219 20646 27271 20698
rect 6000 20544 6052 20596
rect 7104 20587 7156 20596
rect 7104 20553 7113 20587
rect 7113 20553 7147 20587
rect 7147 20553 7156 20587
rect 7104 20544 7156 20553
rect 9588 20544 9640 20596
rect 10876 20544 10928 20596
rect 13360 20544 13412 20596
rect 3516 20519 3568 20528
rect 3516 20485 3525 20519
rect 3525 20485 3559 20519
rect 3559 20485 3568 20519
rect 3516 20476 3568 20485
rect 3700 20476 3752 20528
rect 5264 20476 5316 20528
rect 7748 20476 7800 20528
rect 8484 20476 8536 20528
rect 10692 20476 10744 20528
rect 11060 20476 11112 20528
rect 1308 20340 1360 20392
rect 1676 20383 1728 20392
rect 1676 20349 1685 20383
rect 1685 20349 1719 20383
rect 1719 20349 1728 20383
rect 1676 20340 1728 20349
rect 3792 20340 3844 20392
rect 4896 20340 4948 20392
rect 5264 20383 5316 20392
rect 5264 20349 5273 20383
rect 5273 20349 5307 20383
rect 5307 20349 5316 20383
rect 5264 20340 5316 20349
rect 8852 20408 8904 20460
rect 8944 20408 8996 20460
rect 9404 20408 9456 20460
rect 9588 20408 9640 20460
rect 10232 20408 10284 20460
rect 10324 20408 10376 20460
rect 6000 20383 6052 20392
rect 6000 20349 6009 20383
rect 6009 20349 6043 20383
rect 6043 20349 6052 20383
rect 6000 20340 6052 20349
rect 6460 20340 6512 20392
rect 8300 20340 8352 20392
rect 8392 20340 8444 20392
rect 8576 20340 8628 20392
rect 10968 20383 11020 20392
rect 10968 20349 10977 20383
rect 10977 20349 11011 20383
rect 11011 20349 11020 20383
rect 10968 20340 11020 20349
rect 11244 20383 11296 20392
rect 11244 20349 11253 20383
rect 11253 20349 11287 20383
rect 11287 20349 11296 20383
rect 11244 20340 11296 20349
rect 11428 20408 11480 20460
rect 11612 20408 11664 20460
rect 12808 20408 12860 20460
rect 13820 20408 13872 20460
rect 14004 20433 14056 20460
rect 14004 20408 14049 20433
rect 14049 20408 14056 20433
rect 12072 20340 12124 20392
rect 12624 20340 12676 20392
rect 12900 20340 12952 20392
rect 14648 20340 14700 20392
rect 21916 20544 21968 20596
rect 22008 20544 22060 20596
rect 24308 20544 24360 20596
rect 25136 20544 25188 20596
rect 15200 20408 15252 20460
rect 16120 20340 16172 20392
rect 19064 20408 19116 20460
rect 18604 20340 18656 20392
rect 26240 20476 26292 20528
rect 19248 20451 19300 20460
rect 19248 20417 19257 20451
rect 19257 20417 19291 20451
rect 19291 20417 19300 20451
rect 19248 20408 19300 20417
rect 21180 20408 21232 20460
rect 7564 20272 7616 20324
rect 1584 20204 1636 20256
rect 3332 20204 3384 20256
rect 3884 20247 3936 20256
rect 3884 20213 3893 20247
rect 3893 20213 3927 20247
rect 3927 20213 3936 20247
rect 3884 20204 3936 20213
rect 4436 20247 4488 20256
rect 4436 20213 4445 20247
rect 4445 20213 4479 20247
rect 4479 20213 4488 20247
rect 4436 20204 4488 20213
rect 5356 20204 5408 20256
rect 5540 20204 5592 20256
rect 5908 20204 5960 20256
rect 11152 20272 11204 20324
rect 11336 20272 11388 20324
rect 15108 20272 15160 20324
rect 11520 20204 11572 20256
rect 14372 20204 14424 20256
rect 15384 20247 15436 20256
rect 15384 20213 15393 20247
rect 15393 20213 15427 20247
rect 15427 20213 15436 20247
rect 15384 20204 15436 20213
rect 18696 20272 18748 20324
rect 19156 20272 19208 20324
rect 21548 20383 21600 20392
rect 21548 20349 21557 20383
rect 21557 20349 21591 20383
rect 21591 20349 21600 20383
rect 21548 20340 21600 20349
rect 23388 20340 23440 20392
rect 25228 20340 25280 20392
rect 16764 20204 16816 20256
rect 17224 20204 17276 20256
rect 17960 20204 18012 20256
rect 20260 20272 20312 20324
rect 21824 20272 21876 20324
rect 22560 20272 22612 20324
rect 22192 20204 22244 20256
rect 26424 20340 26476 20392
rect 26792 20340 26844 20392
rect 29276 20340 29328 20392
rect 29368 20340 29420 20392
rect 29828 20383 29880 20392
rect 29828 20349 29837 20383
rect 29837 20349 29871 20383
rect 29871 20349 29880 20383
rect 29828 20340 29880 20349
rect 30196 20340 30248 20392
rect 29092 20315 29144 20324
rect 29092 20281 29101 20315
rect 29101 20281 29135 20315
rect 29135 20281 29144 20315
rect 29092 20272 29144 20281
rect 24768 20204 24820 20256
rect 26148 20204 26200 20256
rect 26792 20204 26844 20256
rect 27344 20204 27396 20256
rect 27804 20204 27856 20256
rect 29920 20247 29972 20256
rect 29920 20213 29929 20247
rect 29929 20213 29963 20247
rect 29963 20213 29972 20247
rect 29920 20204 29972 20213
rect 30104 20315 30156 20324
rect 30104 20281 30113 20315
rect 30113 20281 30147 20315
rect 30147 20281 30156 20315
rect 30104 20272 30156 20281
rect 30656 20272 30708 20324
rect 7988 20102 8040 20154
rect 8052 20102 8104 20154
rect 8116 20102 8168 20154
rect 8180 20102 8232 20154
rect 8244 20102 8296 20154
rect 15578 20102 15630 20154
rect 15642 20102 15694 20154
rect 15706 20102 15758 20154
rect 15770 20102 15822 20154
rect 15834 20102 15886 20154
rect 23168 20102 23220 20154
rect 23232 20102 23284 20154
rect 23296 20102 23348 20154
rect 23360 20102 23412 20154
rect 23424 20102 23476 20154
rect 30758 20102 30810 20154
rect 30822 20102 30874 20154
rect 30886 20102 30938 20154
rect 30950 20102 31002 20154
rect 31014 20102 31066 20154
rect 1584 20000 1636 20052
rect 1308 19907 1360 19916
rect 1308 19873 1317 19907
rect 1317 19873 1351 19907
rect 1351 19873 1360 19907
rect 1308 19864 1360 19873
rect 3332 20043 3384 20052
rect 3332 20009 3341 20043
rect 3341 20009 3375 20043
rect 3375 20009 3384 20043
rect 3332 20000 3384 20009
rect 3608 19975 3660 19984
rect 3608 19941 3617 19975
rect 3617 19941 3651 19975
rect 3651 19941 3660 19975
rect 3608 19932 3660 19941
rect 4528 19975 4580 19984
rect 4528 19941 4537 19975
rect 4537 19941 4571 19975
rect 4571 19941 4580 19975
rect 4528 19932 4580 19941
rect 4712 19975 4764 19984
rect 4712 19941 4721 19975
rect 4721 19941 4755 19975
rect 4755 19941 4764 19975
rect 4712 19932 4764 19941
rect 5080 19975 5132 19984
rect 5080 19941 5089 19975
rect 5089 19941 5123 19975
rect 5123 19941 5132 19975
rect 5080 19932 5132 19941
rect 5264 19975 5316 19984
rect 5264 19941 5273 19975
rect 5273 19941 5307 19975
rect 5307 19941 5316 19975
rect 5264 19932 5316 19941
rect 5908 19932 5960 19984
rect 8576 19932 8628 19984
rect 3700 19864 3752 19916
rect 3884 19864 3936 19916
rect 5632 19864 5684 19916
rect 5816 19907 5868 19916
rect 5816 19873 5825 19907
rect 5825 19873 5859 19907
rect 5859 19873 5868 19907
rect 5816 19864 5868 19873
rect 6828 19864 6880 19916
rect 7012 19907 7064 19916
rect 7012 19873 7021 19907
rect 7021 19873 7055 19907
rect 7055 19873 7064 19907
rect 7012 19864 7064 19873
rect 7840 19864 7892 19916
rect 1584 19796 1636 19848
rect 1952 19796 2004 19848
rect 2044 19839 2096 19848
rect 2044 19805 2053 19839
rect 2053 19805 2087 19839
rect 2087 19805 2096 19839
rect 2044 19796 2096 19805
rect 3332 19796 3384 19848
rect 8392 19796 8444 19848
rect 8944 19839 8996 19848
rect 8944 19805 8956 19839
rect 8956 19805 8990 19839
rect 8990 19805 8996 19839
rect 8944 19796 8996 19805
rect 11612 19932 11664 19984
rect 9312 19796 9364 19848
rect 9404 19796 9456 19848
rect 9588 19796 9640 19848
rect 5264 19728 5316 19780
rect 5724 19728 5776 19780
rect 11888 19864 11940 19916
rect 12440 19864 12492 19916
rect 11612 19796 11664 19848
rect 12164 19839 12216 19848
rect 12164 19805 12166 19839
rect 12166 19805 12216 19839
rect 12164 19796 12216 19805
rect 14188 19907 14240 19916
rect 14188 19873 14197 19907
rect 14197 19873 14231 19907
rect 14231 19873 14240 19907
rect 14188 19864 14240 19873
rect 15752 19932 15804 19984
rect 18880 20000 18932 20052
rect 19064 20000 19116 20052
rect 20720 20000 20772 20052
rect 15476 19864 15528 19916
rect 4068 19660 4120 19712
rect 5540 19703 5592 19712
rect 5540 19669 5549 19703
rect 5549 19669 5583 19703
rect 5583 19669 5592 19703
rect 5540 19660 5592 19669
rect 6460 19660 6512 19712
rect 11336 19728 11388 19780
rect 11428 19728 11480 19780
rect 11704 19728 11756 19780
rect 13912 19728 13964 19780
rect 14096 19728 14148 19780
rect 15292 19796 15344 19848
rect 16304 19932 16356 19984
rect 17684 19932 17736 19984
rect 19800 19975 19852 19984
rect 19800 19941 19809 19975
rect 19809 19941 19843 19975
rect 19843 19941 19852 19975
rect 19800 19932 19852 19941
rect 20628 19932 20680 19984
rect 20076 19864 20128 19916
rect 20168 19907 20220 19916
rect 20168 19873 20177 19907
rect 20177 19873 20211 19907
rect 20211 19873 20220 19907
rect 20168 19864 20220 19873
rect 20260 19864 20312 19916
rect 9036 19660 9088 19712
rect 9128 19660 9180 19712
rect 9404 19660 9456 19712
rect 12256 19660 12308 19712
rect 12440 19660 12492 19712
rect 13268 19660 13320 19712
rect 13636 19703 13688 19712
rect 13636 19669 13645 19703
rect 13645 19669 13679 19703
rect 13679 19669 13688 19703
rect 13636 19660 13688 19669
rect 14464 19660 14516 19712
rect 16028 19660 16080 19712
rect 16488 19796 16540 19848
rect 17960 19839 18012 19848
rect 17960 19805 17969 19839
rect 17969 19805 18003 19839
rect 18003 19805 18012 19839
rect 17960 19796 18012 19805
rect 21088 19907 21140 19916
rect 21088 19873 21097 19907
rect 21097 19873 21131 19907
rect 21131 19873 21140 19907
rect 21088 19864 21140 19873
rect 22560 20000 22612 20052
rect 21548 19932 21600 19984
rect 16764 19660 16816 19712
rect 18972 19660 19024 19712
rect 20168 19660 20220 19712
rect 20628 19703 20680 19712
rect 20628 19669 20637 19703
rect 20637 19669 20671 19703
rect 20671 19669 20680 19703
rect 20628 19660 20680 19669
rect 22008 19907 22060 19916
rect 22008 19873 22017 19907
rect 22017 19873 22051 19907
rect 22051 19873 22060 19907
rect 22008 19864 22060 19873
rect 22652 19932 22704 19984
rect 23848 20000 23900 20052
rect 25228 20000 25280 20052
rect 26240 20000 26292 20052
rect 29276 20000 29328 20052
rect 30564 20000 30616 20052
rect 23388 19728 23440 19780
rect 24308 19839 24360 19848
rect 24308 19805 24317 19839
rect 24317 19805 24351 19839
rect 24351 19805 24360 19839
rect 24308 19796 24360 19805
rect 26332 19864 26384 19916
rect 27620 19864 27672 19916
rect 27988 19864 28040 19916
rect 28540 19864 28592 19916
rect 26332 19728 26384 19780
rect 22100 19660 22152 19712
rect 22192 19660 22244 19712
rect 26056 19703 26108 19712
rect 26056 19669 26065 19703
rect 26065 19669 26099 19703
rect 26099 19669 26108 19703
rect 26056 19660 26108 19669
rect 26148 19660 26200 19712
rect 27804 19796 27856 19848
rect 28264 19796 28316 19848
rect 28816 19839 28868 19848
rect 28816 19805 28818 19839
rect 28818 19805 28868 19839
rect 28816 19796 28868 19805
rect 29000 19796 29052 19848
rect 29552 19796 29604 19848
rect 30012 19660 30064 19712
rect 30288 19660 30340 19712
rect 4193 19558 4245 19610
rect 4257 19558 4309 19610
rect 4321 19558 4373 19610
rect 4385 19558 4437 19610
rect 4449 19558 4501 19610
rect 11783 19558 11835 19610
rect 11847 19558 11899 19610
rect 11911 19558 11963 19610
rect 11975 19558 12027 19610
rect 12039 19558 12091 19610
rect 19373 19558 19425 19610
rect 19437 19558 19489 19610
rect 19501 19558 19553 19610
rect 19565 19558 19617 19610
rect 19629 19558 19681 19610
rect 26963 19558 27015 19610
rect 27027 19558 27079 19610
rect 27091 19558 27143 19610
rect 27155 19558 27207 19610
rect 27219 19558 27271 19610
rect 1216 19456 1268 19508
rect 3792 19456 3844 19508
rect 8208 19456 8260 19508
rect 8300 19456 8352 19508
rect 5172 19388 5224 19440
rect 1308 19320 1360 19372
rect 1584 19320 1636 19372
rect 2228 19320 2280 19372
rect 3792 19320 3844 19372
rect 848 19295 900 19304
rect 848 19261 857 19295
rect 857 19261 891 19295
rect 891 19261 900 19295
rect 848 19252 900 19261
rect 664 19184 716 19236
rect 2504 19295 2556 19304
rect 2504 19261 2513 19295
rect 2513 19261 2547 19295
rect 2547 19261 2556 19295
rect 2504 19252 2556 19261
rect 3976 19252 4028 19304
rect 5172 19252 5224 19304
rect 5816 19388 5868 19440
rect 7656 19388 7708 19440
rect 10232 19499 10284 19508
rect 10232 19465 10241 19499
rect 10241 19465 10275 19499
rect 10275 19465 10284 19499
rect 10232 19456 10284 19465
rect 11244 19456 11296 19508
rect 11796 19456 11848 19508
rect 12624 19456 12676 19508
rect 14096 19456 14148 19508
rect 11152 19388 11204 19440
rect 5632 19320 5684 19372
rect 8392 19363 8444 19372
rect 8392 19329 8401 19363
rect 8401 19329 8435 19363
rect 8435 19329 8444 19363
rect 8392 19320 8444 19329
rect 8576 19320 8628 19372
rect 9036 19320 9088 19372
rect 9312 19320 9364 19372
rect 11428 19320 11480 19372
rect 2964 19184 3016 19236
rect 6552 19295 6604 19304
rect 6552 19261 6561 19295
rect 6561 19261 6595 19295
rect 6595 19261 6604 19295
rect 6552 19252 6604 19261
rect 7196 19252 7248 19304
rect 8668 19252 8720 19304
rect 9864 19252 9916 19304
rect 10140 19252 10192 19304
rect 10232 19184 10284 19236
rect 11244 19295 11296 19304
rect 11244 19261 11253 19295
rect 11253 19261 11287 19295
rect 11287 19261 11296 19295
rect 11244 19252 11296 19261
rect 12900 19320 12952 19372
rect 15936 19388 15988 19440
rect 14924 19252 14976 19304
rect 15108 19295 15160 19304
rect 15108 19261 15117 19295
rect 15117 19261 15151 19295
rect 15151 19261 15160 19295
rect 15108 19252 15160 19261
rect 12992 19184 13044 19236
rect 14556 19184 14608 19236
rect 16488 19456 16540 19508
rect 16856 19456 16908 19508
rect 17684 19456 17736 19508
rect 17960 19456 18012 19508
rect 19156 19456 19208 19508
rect 21916 19456 21968 19508
rect 22100 19456 22152 19508
rect 22836 19456 22888 19508
rect 23572 19499 23624 19508
rect 23572 19465 23581 19499
rect 23581 19465 23615 19499
rect 23615 19465 23624 19499
rect 23572 19456 23624 19465
rect 26516 19456 26568 19508
rect 18144 19363 18196 19372
rect 18144 19329 18153 19363
rect 18153 19329 18187 19363
rect 18187 19329 18196 19363
rect 18144 19320 18196 19329
rect 18236 19320 18288 19372
rect 17316 19252 17368 19304
rect 17408 19252 17460 19304
rect 18420 19252 18472 19304
rect 18512 19295 18564 19304
rect 18512 19261 18521 19295
rect 18521 19261 18555 19295
rect 18555 19261 18564 19295
rect 18512 19252 18564 19261
rect 18696 19295 18748 19304
rect 18696 19261 18705 19295
rect 18705 19261 18739 19295
rect 18739 19261 18748 19295
rect 18696 19252 18748 19261
rect 15384 19184 15436 19236
rect 16212 19184 16264 19236
rect 19340 19320 19392 19372
rect 22836 19320 22888 19372
rect 30288 19431 30340 19440
rect 30288 19397 30297 19431
rect 30297 19397 30331 19431
rect 30331 19397 30340 19431
rect 30288 19388 30340 19397
rect 27252 19320 27304 19372
rect 27344 19320 27396 19372
rect 19892 19252 19944 19304
rect 20076 19252 20128 19304
rect 20444 19295 20496 19304
rect 20444 19261 20453 19295
rect 20453 19261 20487 19295
rect 20487 19261 20496 19295
rect 20444 19252 20496 19261
rect 20168 19184 20220 19236
rect 20812 19252 20864 19304
rect 3240 19159 3292 19168
rect 3240 19125 3249 19159
rect 3249 19125 3283 19159
rect 3283 19125 3292 19159
rect 3240 19116 3292 19125
rect 4988 19159 5040 19168
rect 4988 19125 4997 19159
rect 4997 19125 5031 19159
rect 5031 19125 5040 19159
rect 4988 19116 5040 19125
rect 5448 19116 5500 19168
rect 5724 19116 5776 19168
rect 8668 19116 8720 19168
rect 9220 19116 9272 19168
rect 11244 19116 11296 19168
rect 11520 19116 11572 19168
rect 14004 19116 14056 19168
rect 14280 19116 14332 19168
rect 14832 19116 14884 19168
rect 14924 19159 14976 19168
rect 14924 19125 14933 19159
rect 14933 19125 14967 19159
rect 14967 19125 14976 19159
rect 14924 19116 14976 19125
rect 15108 19116 15160 19168
rect 16396 19116 16448 19168
rect 16764 19116 16816 19168
rect 18328 19116 18380 19168
rect 20260 19116 20312 19168
rect 20444 19116 20496 19168
rect 22652 19252 22704 19304
rect 22468 19227 22520 19236
rect 22468 19193 22477 19227
rect 22477 19193 22511 19227
rect 22511 19193 22520 19227
rect 22468 19184 22520 19193
rect 23664 19184 23716 19236
rect 24492 19295 24544 19304
rect 24492 19261 24501 19295
rect 24501 19261 24535 19295
rect 24535 19261 24544 19295
rect 24492 19252 24544 19261
rect 25136 19252 25188 19304
rect 25504 19252 25556 19304
rect 26700 19295 26752 19304
rect 26700 19261 26709 19295
rect 26709 19261 26743 19295
rect 26743 19261 26752 19295
rect 26700 19252 26752 19261
rect 27528 19252 27580 19304
rect 29184 19252 29236 19304
rect 29828 19320 29880 19372
rect 29644 19252 29696 19304
rect 24492 19116 24544 19168
rect 28172 19184 28224 19236
rect 26332 19159 26384 19168
rect 26332 19125 26341 19159
rect 26341 19125 26375 19159
rect 26375 19125 26384 19159
rect 26332 19116 26384 19125
rect 26792 19116 26844 19168
rect 26976 19116 27028 19168
rect 28816 19184 28868 19236
rect 29368 19116 29420 19168
rect 7988 19014 8040 19066
rect 8052 19014 8104 19066
rect 8116 19014 8168 19066
rect 8180 19014 8232 19066
rect 8244 19014 8296 19066
rect 15578 19014 15630 19066
rect 15642 19014 15694 19066
rect 15706 19014 15758 19066
rect 15770 19014 15822 19066
rect 15834 19014 15886 19066
rect 23168 19014 23220 19066
rect 23232 19014 23284 19066
rect 23296 19014 23348 19066
rect 23360 19014 23412 19066
rect 23424 19014 23476 19066
rect 30758 19014 30810 19066
rect 30822 19014 30874 19066
rect 30886 19014 30938 19066
rect 30950 19014 31002 19066
rect 31014 19014 31066 19066
rect 1584 18912 1636 18964
rect 3056 18912 3108 18964
rect 3240 18912 3292 18964
rect 1216 18819 1268 18828
rect 1216 18785 1225 18819
rect 1225 18785 1259 18819
rect 1259 18785 1268 18819
rect 1216 18776 1268 18785
rect 1308 18751 1360 18760
rect 1308 18717 1317 18751
rect 1317 18717 1351 18751
rect 1351 18717 1360 18751
rect 1308 18708 1360 18717
rect 2872 18776 2924 18828
rect 2964 18776 3016 18828
rect 3424 18887 3476 18896
rect 3424 18853 3433 18887
rect 3433 18853 3467 18887
rect 3467 18853 3476 18887
rect 3424 18844 3476 18853
rect 5632 18887 5684 18896
rect 5632 18853 5641 18887
rect 5641 18853 5675 18887
rect 5675 18853 5684 18887
rect 5632 18844 5684 18853
rect 5816 18844 5868 18896
rect 2504 18708 2556 18760
rect 3424 18572 3476 18624
rect 3700 18708 3752 18760
rect 6184 18776 6236 18828
rect 4988 18708 5040 18760
rect 6092 18708 6144 18760
rect 6368 18751 6420 18760
rect 6368 18717 6380 18751
rect 6380 18717 6414 18751
rect 6414 18717 6420 18751
rect 6368 18708 6420 18717
rect 6644 18751 6696 18760
rect 6644 18717 6653 18751
rect 6653 18717 6687 18751
rect 6687 18717 6696 18751
rect 6644 18708 6696 18717
rect 5540 18640 5592 18692
rect 8484 18912 8536 18964
rect 7472 18844 7524 18896
rect 9036 18912 9088 18964
rect 9128 18955 9180 18964
rect 9128 18921 9143 18955
rect 9143 18921 9177 18955
rect 9177 18921 9180 18955
rect 9128 18912 9180 18921
rect 11060 18912 11112 18964
rect 11428 18912 11480 18964
rect 14924 18912 14976 18964
rect 15016 18912 15068 18964
rect 15936 18912 15988 18964
rect 7380 18776 7432 18828
rect 7748 18776 7800 18828
rect 8484 18708 8536 18760
rect 8944 18708 8996 18760
rect 13452 18819 13504 18828
rect 13452 18785 13461 18819
rect 13461 18785 13495 18819
rect 13495 18785 13504 18819
rect 13452 18776 13504 18785
rect 15936 18819 15988 18828
rect 15936 18785 15945 18819
rect 15945 18785 15979 18819
rect 15979 18785 15988 18819
rect 15936 18776 15988 18785
rect 16488 18912 16540 18964
rect 17776 18912 17828 18964
rect 20628 18912 20680 18964
rect 19800 18844 19852 18896
rect 21272 18844 21324 18896
rect 23020 18912 23072 18964
rect 25688 18912 25740 18964
rect 26976 18912 27028 18964
rect 28816 18955 28868 18964
rect 28816 18921 28831 18955
rect 28831 18921 28865 18955
rect 28865 18921 28868 18955
rect 28816 18912 28868 18921
rect 29092 18912 29144 18964
rect 29368 18912 29420 18964
rect 30196 18955 30248 18964
rect 30196 18921 30205 18955
rect 30205 18921 30239 18955
rect 30239 18921 30248 18955
rect 30196 18912 30248 18921
rect 24216 18844 24268 18896
rect 10968 18751 11020 18760
rect 10968 18717 10977 18751
rect 10977 18717 11011 18751
rect 11011 18717 11020 18751
rect 10968 18708 11020 18717
rect 11250 18708 11302 18760
rect 11520 18708 11572 18760
rect 11704 18751 11756 18760
rect 11704 18717 11713 18751
rect 11713 18717 11747 18751
rect 11747 18717 11756 18751
rect 11704 18708 11756 18717
rect 11796 18708 11848 18760
rect 12716 18640 12768 18692
rect 5172 18572 5224 18624
rect 13084 18572 13136 18624
rect 13268 18615 13320 18624
rect 13268 18581 13277 18615
rect 13277 18581 13311 18615
rect 13311 18581 13320 18615
rect 13268 18572 13320 18581
rect 14372 18708 14424 18760
rect 16764 18708 16816 18760
rect 17684 18708 17736 18760
rect 14740 18572 14792 18624
rect 16488 18572 16540 18624
rect 18144 18615 18196 18624
rect 18144 18581 18153 18615
rect 18153 18581 18187 18615
rect 18187 18581 18196 18615
rect 18144 18572 18196 18581
rect 18972 18776 19024 18828
rect 20444 18776 20496 18828
rect 18696 18708 18748 18760
rect 18788 18708 18840 18760
rect 22284 18776 22336 18828
rect 20812 18708 20864 18760
rect 21456 18708 21508 18760
rect 22008 18708 22060 18760
rect 22652 18708 22704 18760
rect 22928 18708 22980 18760
rect 23848 18776 23900 18828
rect 24492 18819 24544 18828
rect 24492 18785 24494 18819
rect 24494 18785 24544 18819
rect 24492 18776 24544 18785
rect 27896 18844 27948 18896
rect 25872 18776 25924 18828
rect 26884 18776 26936 18828
rect 28264 18776 28316 18828
rect 23756 18572 23808 18624
rect 23848 18615 23900 18624
rect 23848 18581 23857 18615
rect 23857 18581 23891 18615
rect 23891 18581 23900 18615
rect 23848 18572 23900 18581
rect 26056 18708 26108 18760
rect 26148 18708 26200 18760
rect 24400 18572 24452 18624
rect 25596 18572 25648 18624
rect 27896 18640 27948 18692
rect 29368 18776 29420 18828
rect 28816 18751 28868 18760
rect 28816 18717 28828 18751
rect 28828 18717 28862 18751
rect 28862 18717 28868 18751
rect 28816 18708 28868 18717
rect 29000 18708 29052 18760
rect 29092 18751 29144 18760
rect 29092 18717 29101 18751
rect 29101 18717 29135 18751
rect 29135 18717 29144 18751
rect 29092 18708 29144 18717
rect 26424 18572 26476 18624
rect 26700 18572 26752 18624
rect 28172 18572 28224 18624
rect 28540 18572 28592 18624
rect 31300 18572 31352 18624
rect 4193 18470 4245 18522
rect 4257 18470 4309 18522
rect 4321 18470 4373 18522
rect 4385 18470 4437 18522
rect 4449 18470 4501 18522
rect 11783 18470 11835 18522
rect 11847 18470 11899 18522
rect 11911 18470 11963 18522
rect 11975 18470 12027 18522
rect 12039 18470 12091 18522
rect 19373 18470 19425 18522
rect 19437 18470 19489 18522
rect 19501 18470 19553 18522
rect 19565 18470 19617 18522
rect 19629 18470 19681 18522
rect 26963 18470 27015 18522
rect 27027 18470 27079 18522
rect 27091 18470 27143 18522
rect 27155 18470 27207 18522
rect 27219 18470 27271 18522
rect 1216 18368 1268 18420
rect 3608 18368 3660 18420
rect 3700 18368 3752 18420
rect 5724 18368 5776 18420
rect 6368 18368 6420 18420
rect 6920 18368 6972 18420
rect 13636 18368 13688 18420
rect 17868 18368 17920 18420
rect 18052 18368 18104 18420
rect 21272 18368 21324 18420
rect 21456 18368 21508 18420
rect 23756 18368 23808 18420
rect 3056 18232 3108 18284
rect 4252 18232 4304 18284
rect 5540 18232 5592 18284
rect 5632 18232 5684 18284
rect 1676 18207 1728 18216
rect 1676 18173 1685 18207
rect 1685 18173 1719 18207
rect 1719 18173 1728 18207
rect 1676 18164 1728 18173
rect 1216 18028 1268 18080
rect 1584 18028 1636 18080
rect 1768 18028 1820 18080
rect 3608 18164 3660 18216
rect 4528 18164 4580 18216
rect 4712 18164 4764 18216
rect 5448 18164 5500 18216
rect 6092 18207 6144 18216
rect 6092 18173 6101 18207
rect 6101 18173 6135 18207
rect 6135 18173 6144 18207
rect 6092 18164 6144 18173
rect 8392 18232 8444 18284
rect 8944 18232 8996 18284
rect 9128 18232 9180 18284
rect 9312 18275 9364 18284
rect 9312 18241 9321 18275
rect 9321 18241 9355 18275
rect 9355 18241 9364 18275
rect 9312 18232 9364 18241
rect 15936 18300 15988 18352
rect 16212 18300 16264 18352
rect 19248 18300 19300 18352
rect 12256 18232 12308 18284
rect 14188 18275 14240 18284
rect 7472 18164 7524 18216
rect 8484 18164 8536 18216
rect 3700 18028 3752 18080
rect 3884 18028 3936 18080
rect 5080 18028 5132 18080
rect 5908 18028 5960 18080
rect 6184 18028 6236 18080
rect 6736 18028 6788 18080
rect 6828 18028 6880 18080
rect 8484 18028 8536 18080
rect 10692 18096 10744 18148
rect 13544 18164 13596 18216
rect 13728 18164 13780 18216
rect 13820 18207 13872 18216
rect 13820 18173 13829 18207
rect 13829 18173 13863 18207
rect 13863 18173 13872 18207
rect 13820 18164 13872 18173
rect 14188 18241 14190 18275
rect 14190 18241 14240 18275
rect 14188 18232 14240 18241
rect 17040 18232 17092 18284
rect 17132 18275 17184 18284
rect 17132 18241 17141 18275
rect 17141 18241 17175 18275
rect 17175 18241 17184 18275
rect 17132 18232 17184 18241
rect 17316 18232 17368 18284
rect 16856 18207 16908 18216
rect 16856 18173 16865 18207
rect 16865 18173 16899 18207
rect 16899 18173 16908 18207
rect 16856 18164 16908 18173
rect 18328 18232 18380 18284
rect 19892 18300 19944 18352
rect 24400 18343 24452 18352
rect 24400 18309 24409 18343
rect 24409 18309 24443 18343
rect 24443 18309 24452 18343
rect 24400 18300 24452 18309
rect 9036 18071 9088 18080
rect 9036 18037 9051 18071
rect 9051 18037 9085 18071
rect 9085 18037 9088 18071
rect 9036 18028 9088 18037
rect 11060 18028 11112 18080
rect 12992 18028 13044 18080
rect 13176 18071 13228 18080
rect 13176 18037 13185 18071
rect 13185 18037 13219 18071
rect 13219 18037 13228 18071
rect 13176 18028 13228 18037
rect 13912 18028 13964 18080
rect 15844 18028 15896 18080
rect 16396 18028 16448 18080
rect 17132 18028 17184 18080
rect 20168 18164 20220 18216
rect 20536 18232 20588 18284
rect 24032 18232 24084 18284
rect 24216 18232 24268 18284
rect 24860 18232 24912 18284
rect 25596 18232 25648 18284
rect 26148 18300 26200 18352
rect 30104 18368 30156 18420
rect 30288 18411 30340 18420
rect 30288 18377 30297 18411
rect 30297 18377 30331 18411
rect 30331 18377 30340 18411
rect 30288 18368 30340 18377
rect 28724 18300 28776 18352
rect 29736 18300 29788 18352
rect 30380 18300 30432 18352
rect 21732 18164 21784 18216
rect 19616 18096 19668 18148
rect 19800 18139 19852 18148
rect 19800 18105 19809 18139
rect 19809 18105 19843 18139
rect 19843 18105 19852 18139
rect 19800 18096 19852 18105
rect 17960 18028 18012 18080
rect 19984 18071 20036 18080
rect 19984 18037 19993 18071
rect 19993 18037 20027 18071
rect 20027 18037 20036 18071
rect 19984 18028 20036 18037
rect 20812 18071 20864 18080
rect 20812 18037 20827 18071
rect 20827 18037 20861 18071
rect 20861 18037 20864 18071
rect 20812 18028 20864 18037
rect 20996 18028 21048 18080
rect 22468 18096 22520 18148
rect 22836 18096 22888 18148
rect 24584 18207 24636 18216
rect 24584 18173 24593 18207
rect 24593 18173 24627 18207
rect 24627 18173 24636 18207
rect 24584 18164 24636 18173
rect 26056 18164 26108 18216
rect 26516 18164 26568 18216
rect 22192 18071 22244 18080
rect 22192 18037 22201 18071
rect 22201 18037 22235 18071
rect 22235 18037 22244 18071
rect 22192 18028 22244 18037
rect 23572 18139 23624 18148
rect 23572 18105 23581 18139
rect 23581 18105 23615 18139
rect 23615 18105 23624 18139
rect 23572 18096 23624 18105
rect 23756 18096 23808 18148
rect 24124 18096 24176 18148
rect 28540 18164 28592 18216
rect 29736 18164 29788 18216
rect 27896 18096 27948 18148
rect 24952 18028 25004 18080
rect 25320 18028 25372 18080
rect 28356 18028 28408 18080
rect 28908 18096 28960 18148
rect 29828 18028 29880 18080
rect 30012 18028 30064 18080
rect 7988 17926 8040 17978
rect 8052 17926 8104 17978
rect 8116 17926 8168 17978
rect 8180 17926 8232 17978
rect 8244 17926 8296 17978
rect 15578 17926 15630 17978
rect 15642 17926 15694 17978
rect 15706 17926 15758 17978
rect 15770 17926 15822 17978
rect 15834 17926 15886 17978
rect 23168 17926 23220 17978
rect 23232 17926 23284 17978
rect 23296 17926 23348 17978
rect 23360 17926 23412 17978
rect 23424 17926 23476 17978
rect 30758 17926 30810 17978
rect 30822 17926 30874 17978
rect 30886 17926 30938 17978
rect 30950 17926 31002 17978
rect 31014 17926 31066 17978
rect 1308 17824 1360 17876
rect 1768 17867 1820 17876
rect 1768 17833 1783 17867
rect 1783 17833 1817 17867
rect 1817 17833 1820 17867
rect 1768 17824 1820 17833
rect 3148 17867 3200 17876
rect 3148 17833 3157 17867
rect 3157 17833 3191 17867
rect 3191 17833 3200 17867
rect 3148 17824 3200 17833
rect 3424 17824 3476 17876
rect 8760 17824 8812 17876
rect 8944 17824 8996 17876
rect 9680 17824 9732 17876
rect 10692 17824 10744 17876
rect 11152 17824 11204 17876
rect 12164 17824 12216 17876
rect 1216 17484 1268 17536
rect 1676 17620 1728 17672
rect 3148 17688 3200 17740
rect 3516 17731 3568 17740
rect 3516 17697 3525 17731
rect 3525 17697 3559 17731
rect 3559 17697 3568 17731
rect 3516 17688 3568 17697
rect 5632 17799 5684 17808
rect 5632 17765 5641 17799
rect 5641 17765 5675 17799
rect 5675 17765 5684 17799
rect 5632 17756 5684 17765
rect 5724 17756 5776 17808
rect 3240 17620 3292 17672
rect 3884 17663 3936 17672
rect 3884 17629 3886 17663
rect 3886 17629 3936 17663
rect 3884 17620 3936 17629
rect 5816 17731 5868 17740
rect 5816 17697 5825 17731
rect 5825 17697 5859 17731
rect 5859 17697 5868 17731
rect 5816 17688 5868 17697
rect 8576 17799 8628 17808
rect 8576 17765 8585 17799
rect 8585 17765 8619 17799
rect 8619 17765 8628 17799
rect 8576 17756 8628 17765
rect 8668 17756 8720 17808
rect 10784 17799 10836 17808
rect 10784 17765 10793 17799
rect 10793 17765 10827 17799
rect 10827 17765 10836 17799
rect 10784 17756 10836 17765
rect 6736 17688 6788 17740
rect 11336 17756 11388 17808
rect 13544 17756 13596 17808
rect 5448 17620 5500 17672
rect 5632 17620 5684 17672
rect 6092 17620 6144 17672
rect 6644 17620 6696 17672
rect 7012 17620 7064 17672
rect 9220 17688 9272 17740
rect 9496 17688 9548 17740
rect 11152 17688 11204 17740
rect 11244 17688 11296 17740
rect 11612 17688 11664 17740
rect 8208 17620 8260 17672
rect 8392 17552 8444 17604
rect 8852 17620 8904 17672
rect 12256 17663 12308 17672
rect 12256 17629 12265 17663
rect 12265 17629 12299 17663
rect 12299 17629 12308 17663
rect 12256 17620 12308 17629
rect 13176 17688 13228 17740
rect 15292 17824 15344 17876
rect 16212 17824 16264 17876
rect 16580 17824 16632 17876
rect 16672 17824 16724 17876
rect 15568 17756 15620 17808
rect 16028 17756 16080 17808
rect 17316 17824 17368 17876
rect 16304 17731 16356 17740
rect 16304 17697 16313 17731
rect 16313 17697 16347 17731
rect 16347 17697 16356 17731
rect 16304 17688 16356 17697
rect 5816 17484 5868 17536
rect 10416 17484 10468 17536
rect 12256 17484 12308 17536
rect 12716 17484 12768 17536
rect 13820 17663 13872 17672
rect 13820 17629 13829 17663
rect 13829 17629 13863 17663
rect 13863 17629 13872 17663
rect 13820 17620 13872 17629
rect 14188 17663 14240 17672
rect 14188 17629 14190 17663
rect 14190 17629 14240 17663
rect 14188 17620 14240 17629
rect 16212 17663 16264 17672
rect 16212 17629 16221 17663
rect 16221 17629 16255 17663
rect 16255 17629 16264 17663
rect 16212 17620 16264 17629
rect 16304 17552 16356 17604
rect 15384 17484 15436 17536
rect 16672 17620 16724 17672
rect 16856 17620 16908 17672
rect 18788 17688 18840 17740
rect 20076 17688 20128 17740
rect 20260 17688 20312 17740
rect 19524 17620 19576 17672
rect 21272 17663 21324 17672
rect 21272 17629 21281 17663
rect 21281 17629 21315 17663
rect 21315 17629 21324 17663
rect 21272 17620 21324 17629
rect 21456 17620 21508 17672
rect 23020 17688 23072 17740
rect 23940 17824 23992 17876
rect 24032 17824 24084 17876
rect 26792 17824 26844 17876
rect 27068 17824 27120 17876
rect 28540 17824 28592 17876
rect 28724 17824 28776 17876
rect 29276 17824 29328 17876
rect 29644 17824 29696 17876
rect 28264 17756 28316 17808
rect 23848 17688 23900 17740
rect 24216 17688 24268 17740
rect 24400 17688 24452 17740
rect 24952 17688 25004 17740
rect 25228 17688 25280 17740
rect 25872 17688 25924 17740
rect 18328 17484 18380 17536
rect 18788 17527 18840 17536
rect 18788 17493 18797 17527
rect 18797 17493 18831 17527
rect 18831 17493 18840 17527
rect 18788 17484 18840 17493
rect 19156 17484 19208 17536
rect 21180 17552 21232 17604
rect 24768 17620 24820 17672
rect 25596 17620 25648 17672
rect 26148 17620 26200 17672
rect 26424 17663 26476 17672
rect 26424 17629 26433 17663
rect 26433 17629 26467 17663
rect 26467 17629 26476 17663
rect 26424 17620 26476 17629
rect 26884 17663 26936 17672
rect 26884 17629 26896 17663
rect 26896 17629 26930 17663
rect 26930 17629 26936 17663
rect 26884 17620 26936 17629
rect 21548 17484 21600 17536
rect 23940 17595 23992 17604
rect 23940 17561 23949 17595
rect 23949 17561 23983 17595
rect 23983 17561 23992 17595
rect 23940 17552 23992 17561
rect 25780 17484 25832 17536
rect 28540 17620 28592 17672
rect 29000 17620 29052 17672
rect 29276 17620 29328 17672
rect 30380 17595 30432 17604
rect 30380 17561 30389 17595
rect 30389 17561 30423 17595
rect 30423 17561 30432 17595
rect 30380 17552 30432 17561
rect 30656 17484 30708 17536
rect 4193 17382 4245 17434
rect 4257 17382 4309 17434
rect 4321 17382 4373 17434
rect 4385 17382 4437 17434
rect 4449 17382 4501 17434
rect 11783 17382 11835 17434
rect 11847 17382 11899 17434
rect 11911 17382 11963 17434
rect 11975 17382 12027 17434
rect 12039 17382 12091 17434
rect 19373 17382 19425 17434
rect 19437 17382 19489 17434
rect 19501 17382 19553 17434
rect 19565 17382 19617 17434
rect 19629 17382 19681 17434
rect 26963 17382 27015 17434
rect 27027 17382 27079 17434
rect 27091 17382 27143 17434
rect 27155 17382 27207 17434
rect 27219 17382 27271 17434
rect 5724 17280 5776 17332
rect 5816 17323 5868 17332
rect 5816 17289 5825 17323
rect 5825 17289 5859 17323
rect 5859 17289 5868 17323
rect 5816 17280 5868 17289
rect 9220 17280 9272 17332
rect 9312 17280 9364 17332
rect 1216 17144 1268 17196
rect 2136 17144 2188 17196
rect 3332 17187 3384 17196
rect 3332 17153 3341 17187
rect 3341 17153 3375 17187
rect 3375 17153 3384 17187
rect 3332 17144 3384 17153
rect 3516 17144 3568 17196
rect 2964 17076 3016 17128
rect 3976 17076 4028 17128
rect 4528 17076 4580 17128
rect 5264 17144 5316 17196
rect 6828 17187 6880 17196
rect 6828 17153 6837 17187
rect 6837 17153 6871 17187
rect 6871 17153 6880 17187
rect 6828 17144 6880 17153
rect 8484 17212 8536 17264
rect 10600 17212 10652 17264
rect 10876 17212 10928 17264
rect 1768 16940 1820 16992
rect 3884 16940 3936 16992
rect 5080 16940 5132 16992
rect 5724 16940 5776 16992
rect 6092 17119 6144 17128
rect 6092 17085 6101 17119
rect 6101 17085 6135 17119
rect 6135 17085 6144 17119
rect 6092 17076 6144 17085
rect 6184 17076 6236 17128
rect 7104 17076 7156 17128
rect 8392 17076 8444 17128
rect 8576 17119 8628 17128
rect 8576 17085 8585 17119
rect 8585 17085 8619 17119
rect 8619 17085 8628 17119
rect 8576 17076 8628 17085
rect 6920 16940 6972 16992
rect 9220 17144 9272 17196
rect 12164 17280 12216 17332
rect 12348 17280 12400 17332
rect 14096 17280 14148 17332
rect 15016 17280 15068 17332
rect 18052 17280 18104 17332
rect 18604 17280 18656 17332
rect 20260 17280 20312 17332
rect 12808 17144 12860 17196
rect 9036 17076 9088 17128
rect 9312 17076 9364 17128
rect 9496 17076 9548 17128
rect 10508 17076 10560 17128
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 11244 17119 11296 17128
rect 11244 17085 11253 17119
rect 11253 17085 11287 17119
rect 11287 17085 11296 17119
rect 11244 17076 11296 17085
rect 10968 17008 11020 17060
rect 12256 17076 12308 17128
rect 13544 17212 13596 17264
rect 13084 17144 13136 17196
rect 16212 17212 16264 17264
rect 22376 17280 22428 17332
rect 23204 17280 23256 17332
rect 15568 17144 15620 17196
rect 9680 16940 9732 16992
rect 10140 16940 10192 16992
rect 11336 16940 11388 16992
rect 11888 16940 11940 16992
rect 13636 16940 13688 16992
rect 14924 17076 14976 17128
rect 14648 17008 14700 17060
rect 16672 17076 16724 17128
rect 17132 17187 17184 17196
rect 17132 17153 17141 17187
rect 17141 17153 17175 17187
rect 17175 17153 17184 17187
rect 17132 17144 17184 17153
rect 19984 17144 20036 17196
rect 18696 17119 18748 17128
rect 18696 17085 18705 17119
rect 18705 17085 18739 17119
rect 18739 17085 18748 17119
rect 18696 17076 18748 17085
rect 22008 17212 22060 17264
rect 25780 17323 25832 17332
rect 25780 17289 25789 17323
rect 25789 17289 25823 17323
rect 25823 17289 25832 17323
rect 25780 17280 25832 17289
rect 25964 17280 26016 17332
rect 28448 17280 28500 17332
rect 28724 17323 28776 17332
rect 28724 17289 28733 17323
rect 28733 17289 28767 17323
rect 28767 17289 28776 17323
rect 28724 17280 28776 17289
rect 29828 17280 29880 17332
rect 21088 17144 21140 17196
rect 21180 17187 21232 17196
rect 21180 17153 21189 17187
rect 21189 17153 21223 17187
rect 21223 17153 21232 17187
rect 21180 17144 21232 17153
rect 20536 17076 20588 17128
rect 20812 17119 20864 17128
rect 20812 17085 20814 17119
rect 20814 17085 20864 17119
rect 20812 17076 20864 17085
rect 21456 17076 21508 17128
rect 22560 17076 22612 17128
rect 23204 17119 23256 17128
rect 23204 17085 23213 17119
rect 23213 17085 23247 17119
rect 23247 17085 23256 17119
rect 23204 17076 23256 17085
rect 25872 17212 25924 17264
rect 27712 17212 27764 17264
rect 24216 17144 24268 17196
rect 26332 17144 26384 17196
rect 26148 17119 26200 17128
rect 26148 17085 26157 17119
rect 26157 17085 26191 17119
rect 26191 17085 26200 17119
rect 26148 17076 26200 17085
rect 26516 17076 26568 17128
rect 28080 17076 28132 17128
rect 29276 17076 29328 17128
rect 29644 17119 29696 17128
rect 29644 17085 29653 17119
rect 29653 17085 29687 17119
rect 29687 17085 29696 17119
rect 29644 17076 29696 17085
rect 16856 16983 16908 16992
rect 16856 16949 16871 16983
rect 16871 16949 16905 16983
rect 16905 16949 16908 16983
rect 16856 16940 16908 16949
rect 17040 16940 17092 16992
rect 18420 16940 18472 16992
rect 20076 16983 20128 16992
rect 20076 16949 20085 16983
rect 20085 16949 20119 16983
rect 20119 16949 20128 16983
rect 20076 16940 20128 16949
rect 24400 16983 24452 16992
rect 24400 16949 24415 16983
rect 24415 16949 24449 16983
rect 24449 16949 24452 16983
rect 24400 16940 24452 16949
rect 26424 16940 26476 16992
rect 26792 16940 26844 16992
rect 28540 16940 28592 16992
rect 29460 16940 29512 16992
rect 30012 17076 30064 17128
rect 31116 17076 31168 17128
rect 30012 16940 30064 16992
rect 31024 16940 31076 16992
rect 7988 16838 8040 16890
rect 8052 16838 8104 16890
rect 8116 16838 8168 16890
rect 8180 16838 8232 16890
rect 8244 16838 8296 16890
rect 15578 16838 15630 16890
rect 15642 16838 15694 16890
rect 15706 16838 15758 16890
rect 15770 16838 15822 16890
rect 15834 16838 15886 16890
rect 23168 16838 23220 16890
rect 23232 16838 23284 16890
rect 23296 16838 23348 16890
rect 23360 16838 23412 16890
rect 23424 16838 23476 16890
rect 30758 16838 30810 16890
rect 30822 16838 30874 16890
rect 30886 16838 30938 16890
rect 30950 16838 31002 16890
rect 31014 16838 31066 16890
rect 1216 16736 1268 16788
rect 2320 16736 2372 16788
rect 3056 16779 3108 16788
rect 3056 16745 3065 16779
rect 3065 16745 3099 16779
rect 3099 16745 3108 16779
rect 3056 16736 3108 16745
rect 3332 16736 3384 16788
rect 3608 16600 3660 16652
rect 4528 16600 4580 16652
rect 5540 16779 5592 16788
rect 5540 16745 5549 16779
rect 5549 16745 5583 16779
rect 5583 16745 5592 16779
rect 5540 16736 5592 16745
rect 5080 16668 5132 16720
rect 7012 16736 7064 16788
rect 8668 16736 8720 16788
rect 8944 16736 8996 16788
rect 10508 16779 10560 16788
rect 10508 16745 10517 16779
rect 10517 16745 10551 16779
rect 10551 16745 10560 16779
rect 10508 16736 10560 16745
rect 7288 16668 7340 16720
rect 11888 16736 11940 16788
rect 12808 16736 12860 16788
rect 16120 16779 16172 16788
rect 16120 16745 16129 16779
rect 16129 16745 16163 16779
rect 16163 16745 16172 16779
rect 16120 16736 16172 16745
rect 17040 16736 17092 16788
rect 17960 16736 18012 16788
rect 19156 16736 19208 16788
rect 5908 16600 5960 16652
rect 1032 16532 1084 16584
rect 1584 16575 1636 16584
rect 1584 16541 1586 16575
rect 1586 16541 1636 16575
rect 1584 16532 1636 16541
rect 1768 16532 1820 16584
rect 940 16439 992 16448
rect 940 16405 949 16439
rect 949 16405 983 16439
rect 983 16405 992 16439
rect 940 16396 992 16405
rect 3700 16532 3752 16584
rect 3884 16575 3936 16584
rect 3884 16541 3886 16575
rect 3886 16541 3936 16575
rect 3884 16532 3936 16541
rect 4068 16532 4120 16584
rect 6552 16643 6604 16652
rect 6552 16609 6561 16643
rect 6561 16609 6595 16643
rect 6595 16609 6604 16643
rect 6552 16600 6604 16609
rect 9404 16643 9456 16652
rect 9404 16609 9413 16643
rect 9413 16609 9447 16643
rect 9447 16609 9456 16643
rect 9404 16600 9456 16609
rect 13912 16668 13964 16720
rect 8668 16575 8720 16584
rect 8668 16541 8677 16575
rect 8677 16541 8711 16575
rect 8711 16541 8720 16575
rect 8668 16532 8720 16541
rect 11060 16643 11112 16652
rect 11060 16609 11069 16643
rect 11069 16609 11103 16643
rect 11103 16609 11112 16643
rect 11060 16600 11112 16609
rect 10324 16532 10376 16584
rect 14188 16643 14240 16652
rect 11244 16532 11296 16584
rect 11796 16532 11848 16584
rect 11980 16575 12032 16584
rect 11980 16541 11982 16575
rect 11982 16541 12032 16575
rect 11980 16532 12032 16541
rect 14188 16609 14190 16643
rect 14190 16609 14240 16643
rect 14188 16600 14240 16609
rect 13820 16575 13872 16584
rect 13820 16541 13829 16575
rect 13829 16541 13863 16575
rect 13863 16541 13872 16575
rect 13820 16532 13872 16541
rect 15476 16600 15528 16652
rect 16212 16600 16264 16652
rect 14464 16534 14516 16586
rect 17040 16600 17092 16652
rect 21180 16736 21232 16788
rect 16672 16532 16724 16584
rect 17132 16532 17184 16584
rect 18420 16532 18472 16584
rect 20076 16600 20128 16652
rect 21088 16643 21140 16652
rect 21088 16609 21097 16643
rect 21097 16609 21131 16643
rect 21131 16609 21140 16643
rect 21088 16600 21140 16609
rect 23848 16779 23900 16788
rect 23848 16745 23857 16779
rect 23857 16745 23891 16779
rect 23891 16745 23900 16779
rect 23848 16736 23900 16745
rect 21364 16600 21416 16652
rect 22376 16600 22428 16652
rect 23940 16600 23992 16652
rect 24216 16736 24268 16788
rect 24400 16736 24452 16788
rect 27896 16736 27948 16788
rect 28356 16736 28408 16788
rect 29920 16736 29972 16788
rect 30380 16779 30432 16788
rect 30380 16745 30389 16779
rect 30389 16745 30423 16779
rect 30423 16745 30432 16779
rect 30380 16736 30432 16745
rect 31024 16736 31076 16788
rect 27988 16668 28040 16720
rect 26056 16600 26108 16652
rect 27252 16600 27304 16652
rect 27620 16600 27672 16652
rect 10784 16464 10836 16516
rect 5264 16396 5316 16448
rect 5540 16396 5592 16448
rect 10140 16396 10192 16448
rect 11336 16507 11388 16516
rect 11336 16473 11345 16507
rect 11345 16473 11379 16507
rect 11379 16473 11388 16507
rect 11336 16464 11388 16473
rect 12716 16396 12768 16448
rect 13452 16439 13504 16448
rect 13452 16405 13461 16439
rect 13461 16405 13495 16439
rect 13495 16405 13504 16439
rect 13452 16396 13504 16405
rect 14280 16396 14332 16448
rect 15476 16464 15528 16516
rect 15936 16396 15988 16448
rect 19432 16464 19484 16516
rect 20536 16532 20588 16584
rect 20904 16532 20956 16584
rect 21272 16575 21324 16584
rect 21272 16541 21281 16575
rect 21281 16541 21315 16575
rect 21315 16541 21324 16575
rect 21272 16532 21324 16541
rect 21456 16532 21508 16584
rect 22744 16464 22796 16516
rect 18420 16396 18472 16448
rect 19156 16439 19208 16448
rect 19156 16405 19165 16439
rect 19165 16405 19199 16439
rect 19199 16405 19208 16439
rect 19156 16396 19208 16405
rect 19248 16396 19300 16448
rect 21088 16396 21140 16448
rect 21180 16396 21232 16448
rect 22468 16396 22520 16448
rect 25044 16532 25096 16584
rect 26148 16532 26200 16584
rect 26792 16575 26844 16584
rect 26792 16541 26794 16575
rect 26794 16541 26844 16575
rect 26792 16532 26844 16541
rect 27896 16532 27948 16584
rect 28172 16532 28224 16584
rect 28448 16532 28500 16584
rect 29276 16532 29328 16584
rect 29552 16532 29604 16584
rect 29644 16532 29696 16584
rect 26792 16396 26844 16448
rect 28264 16439 28316 16448
rect 28264 16405 28273 16439
rect 28273 16405 28307 16439
rect 28307 16405 28316 16439
rect 28264 16396 28316 16405
rect 29368 16396 29420 16448
rect 4193 16294 4245 16346
rect 4257 16294 4309 16346
rect 4321 16294 4373 16346
rect 4385 16294 4437 16346
rect 4449 16294 4501 16346
rect 11783 16294 11835 16346
rect 11847 16294 11899 16346
rect 11911 16294 11963 16346
rect 11975 16294 12027 16346
rect 12039 16294 12091 16346
rect 19373 16294 19425 16346
rect 19437 16294 19489 16346
rect 19501 16294 19553 16346
rect 19565 16294 19617 16346
rect 19629 16294 19681 16346
rect 26963 16294 27015 16346
rect 27027 16294 27079 16346
rect 27091 16294 27143 16346
rect 27155 16294 27207 16346
rect 27219 16294 27271 16346
rect 2964 16235 3016 16244
rect 2964 16201 2973 16235
rect 2973 16201 3007 16235
rect 3007 16201 3016 16235
rect 2964 16192 3016 16201
rect 5540 16192 5592 16244
rect 5632 16235 5684 16244
rect 5632 16201 5641 16235
rect 5641 16201 5675 16235
rect 5675 16201 5684 16235
rect 5632 16192 5684 16201
rect 10324 16192 10376 16244
rect 10140 16124 10192 16176
rect 8300 16056 8352 16108
rect 8392 16056 8444 16108
rect 1032 15988 1084 16040
rect 3332 15963 3384 15972
rect 3332 15929 3341 15963
rect 3341 15929 3375 15963
rect 3375 15929 3384 15963
rect 3332 15920 3384 15929
rect 3700 15988 3752 16040
rect 4436 15988 4488 16040
rect 4896 15988 4948 16040
rect 6184 15988 6236 16040
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 7104 15988 7156 16040
rect 8484 15988 8536 16040
rect 8668 16031 8720 16040
rect 8668 15997 8677 16031
rect 8677 15997 8711 16031
rect 8711 15997 8720 16031
rect 8668 15988 8720 15997
rect 13452 16192 13504 16244
rect 13728 16192 13780 16244
rect 9680 15988 9732 16040
rect 11244 16099 11296 16108
rect 11244 16065 11253 16099
rect 11253 16065 11287 16099
rect 11287 16065 11296 16099
rect 11244 16056 11296 16065
rect 11428 16056 11480 16108
rect 16488 16192 16540 16244
rect 14464 16167 14516 16176
rect 14464 16133 14473 16167
rect 14473 16133 14507 16167
rect 14507 16133 14516 16167
rect 14464 16124 14516 16133
rect 11612 15988 11664 16040
rect 14740 16056 14792 16108
rect 14832 15988 14884 16040
rect 14924 15988 14976 16040
rect 18420 16192 18472 16244
rect 20536 16192 20588 16244
rect 15292 16031 15344 16040
rect 15292 15997 15301 16031
rect 15301 15997 15335 16031
rect 15335 15997 15344 16031
rect 15292 15988 15344 15997
rect 16856 16031 16908 16040
rect 16856 15997 16865 16031
rect 16865 15997 16899 16031
rect 16899 15997 16908 16031
rect 16856 15988 16908 15997
rect 17500 15988 17552 16040
rect 22100 16192 22152 16244
rect 22836 16192 22888 16244
rect 20720 16167 20772 16176
rect 20720 16133 20729 16167
rect 20729 16133 20763 16167
rect 20763 16133 20772 16167
rect 20720 16124 20772 16133
rect 22652 16124 22704 16176
rect 25320 16124 25372 16176
rect 27160 16192 27212 16244
rect 28356 16192 28408 16244
rect 28448 16235 28500 16244
rect 28448 16201 28457 16235
rect 28457 16201 28491 16235
rect 28491 16201 28500 16235
rect 28448 16192 28500 16201
rect 28908 16192 28960 16244
rect 27620 16124 27672 16176
rect 29000 16124 29052 16176
rect 29552 16124 29604 16176
rect 21272 16099 21324 16108
rect 21272 16065 21274 16099
rect 21274 16065 21324 16099
rect 21272 16056 21324 16065
rect 1676 15852 1728 15904
rect 3516 15852 3568 15904
rect 3700 15852 3752 15904
rect 3884 15852 3936 15904
rect 4436 15852 4488 15904
rect 6092 15852 6144 15904
rect 6460 15852 6512 15904
rect 8576 15852 8628 15904
rect 8944 15852 8996 15904
rect 11704 15895 11756 15904
rect 11704 15861 11719 15895
rect 11719 15861 11753 15895
rect 11753 15861 11756 15895
rect 11704 15852 11756 15861
rect 11888 15852 11940 15904
rect 13452 15920 13504 15972
rect 13544 15920 13596 15972
rect 14004 15920 14056 15972
rect 14280 15963 14332 15972
rect 14280 15929 14289 15963
rect 14289 15929 14323 15963
rect 14323 15929 14332 15963
rect 14280 15920 14332 15929
rect 13084 15895 13136 15904
rect 13084 15861 13093 15895
rect 13093 15861 13127 15895
rect 13127 15861 13136 15895
rect 13084 15852 13136 15861
rect 14188 15852 14240 15904
rect 15016 15895 15068 15904
rect 15016 15861 15031 15895
rect 15031 15861 15065 15895
rect 15065 15861 15068 15895
rect 15016 15852 15068 15861
rect 17132 15852 17184 15904
rect 20812 15988 20864 16040
rect 20904 16031 20956 16040
rect 20904 15997 20913 16031
rect 20913 15997 20947 16031
rect 20947 15997 20956 16031
rect 20904 15988 20956 15997
rect 20168 15920 20220 15972
rect 22928 15988 22980 16040
rect 19064 15852 19116 15904
rect 22744 15895 22796 15904
rect 22744 15861 22753 15895
rect 22753 15861 22787 15895
rect 22787 15861 22796 15895
rect 22744 15852 22796 15861
rect 23848 16099 23900 16108
rect 23848 16065 23857 16099
rect 23857 16065 23891 16099
rect 23891 16065 23900 16099
rect 23848 16056 23900 16065
rect 24216 16099 24268 16108
rect 24216 16065 24218 16099
rect 24218 16065 24268 16099
rect 24216 16056 24268 16065
rect 25964 16056 26016 16108
rect 26424 16099 26476 16108
rect 26424 16065 26426 16099
rect 26426 16065 26476 16099
rect 26424 16056 26476 16065
rect 29276 16056 29328 16108
rect 30012 16124 30064 16176
rect 23940 15988 23992 16040
rect 26148 15988 26200 16040
rect 26608 15988 26660 16040
rect 27160 15988 27212 16040
rect 28172 15988 28224 16040
rect 28724 15988 28776 16040
rect 28908 15988 28960 16040
rect 29000 15988 29052 16040
rect 27528 15920 27580 15972
rect 24124 15852 24176 15904
rect 24308 15852 24360 15904
rect 29276 15852 29328 15904
rect 29552 15852 29604 15904
rect 30012 15852 30064 15904
rect 30380 15920 30432 15972
rect 31024 15852 31076 15904
rect 7988 15750 8040 15802
rect 8052 15750 8104 15802
rect 8116 15750 8168 15802
rect 8180 15750 8232 15802
rect 8244 15750 8296 15802
rect 15578 15750 15630 15802
rect 15642 15750 15694 15802
rect 15706 15750 15758 15802
rect 15770 15750 15822 15802
rect 15834 15750 15886 15802
rect 23168 15750 23220 15802
rect 23232 15750 23284 15802
rect 23296 15750 23348 15802
rect 23360 15750 23412 15802
rect 23424 15750 23476 15802
rect 30758 15750 30810 15802
rect 30822 15750 30874 15802
rect 30886 15750 30938 15802
rect 30950 15750 31002 15802
rect 31014 15750 31066 15802
rect 3148 15691 3200 15700
rect 3148 15657 3157 15691
rect 3157 15657 3191 15691
rect 3191 15657 3200 15691
rect 3148 15648 3200 15657
rect 4988 15648 5040 15700
rect 11888 15648 11940 15700
rect 11980 15648 12032 15700
rect 13084 15648 13136 15700
rect 14188 15648 14240 15700
rect 14832 15648 14884 15700
rect 18236 15648 18288 15700
rect 6460 15580 6512 15632
rect 11704 15580 11756 15632
rect 16948 15580 17000 15632
rect 1676 15487 1728 15496
rect 1676 15453 1678 15487
rect 1678 15453 1728 15487
rect 848 15351 900 15360
rect 848 15317 857 15351
rect 857 15317 891 15351
rect 891 15317 900 15351
rect 848 15308 900 15317
rect 1124 15308 1176 15360
rect 1676 15444 1728 15453
rect 2044 15487 2096 15496
rect 2044 15453 2053 15487
rect 2053 15453 2087 15487
rect 2087 15453 2096 15487
rect 2044 15444 2096 15453
rect 3516 15487 3568 15496
rect 3516 15453 3525 15487
rect 3525 15453 3559 15487
rect 3559 15453 3568 15487
rect 3516 15444 3568 15453
rect 3884 15487 3936 15496
rect 3884 15453 3886 15487
rect 3886 15453 3936 15487
rect 3884 15444 3936 15453
rect 3976 15487 4028 15496
rect 3976 15453 3988 15487
rect 3988 15453 4022 15487
rect 4022 15453 4028 15487
rect 3976 15444 4028 15453
rect 4620 15444 4672 15496
rect 5724 15444 5776 15496
rect 3792 15308 3844 15360
rect 6184 15351 6236 15360
rect 6184 15317 6193 15351
rect 6193 15317 6227 15351
rect 6227 15317 6236 15351
rect 7196 15487 7248 15496
rect 7196 15453 7205 15487
rect 7205 15453 7239 15487
rect 7239 15453 7248 15487
rect 7196 15444 7248 15453
rect 7656 15444 7708 15496
rect 7840 15444 7892 15496
rect 8668 15487 8720 15496
rect 8668 15453 8677 15487
rect 8677 15453 8711 15487
rect 8711 15453 8720 15487
rect 8668 15444 8720 15453
rect 8852 15444 8904 15496
rect 9128 15487 9180 15496
rect 9128 15453 9140 15487
rect 9140 15453 9174 15487
rect 9174 15453 9180 15487
rect 9128 15444 9180 15453
rect 9312 15444 9364 15496
rect 6184 15308 6236 15317
rect 8300 15351 8352 15360
rect 8300 15317 8309 15351
rect 8309 15317 8343 15351
rect 8343 15317 8352 15351
rect 8300 15308 8352 15317
rect 11244 15512 11296 15564
rect 12716 15444 12768 15496
rect 13452 15512 13504 15564
rect 13820 15555 13872 15564
rect 13820 15521 13829 15555
rect 13829 15521 13863 15555
rect 13863 15521 13872 15555
rect 13820 15512 13872 15521
rect 14464 15512 14516 15564
rect 15936 15512 15988 15564
rect 11980 15308 12032 15360
rect 13452 15351 13504 15360
rect 13452 15317 13461 15351
rect 13461 15317 13495 15351
rect 13495 15317 13504 15351
rect 13452 15308 13504 15317
rect 14740 15444 14792 15496
rect 17040 15555 17092 15564
rect 17040 15521 17049 15555
rect 17049 15521 17083 15555
rect 17083 15521 17092 15555
rect 17040 15512 17092 15521
rect 19156 15512 19208 15564
rect 17132 15487 17184 15496
rect 17132 15453 17141 15487
rect 17141 15453 17175 15487
rect 17175 15453 17184 15487
rect 17132 15444 17184 15453
rect 17316 15444 17368 15496
rect 23756 15648 23808 15700
rect 24216 15648 24268 15700
rect 21364 15512 21416 15564
rect 21548 15512 21600 15564
rect 23848 15512 23900 15564
rect 27528 15648 27580 15700
rect 28264 15648 28316 15700
rect 29000 15648 29052 15700
rect 26424 15580 26476 15632
rect 29644 15648 29696 15700
rect 31024 15648 31076 15700
rect 31208 15648 31260 15700
rect 29736 15580 29788 15632
rect 30932 15580 30984 15632
rect 18604 15376 18656 15428
rect 19248 15376 19300 15428
rect 19800 15444 19852 15496
rect 20904 15444 20956 15496
rect 21272 15487 21324 15496
rect 21272 15453 21281 15487
rect 21281 15453 21315 15487
rect 21315 15453 21324 15487
rect 21272 15444 21324 15453
rect 21824 15444 21876 15496
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22008 15444 22060 15453
rect 23664 15444 23716 15496
rect 24032 15446 24084 15498
rect 24124 15444 24176 15496
rect 15384 15308 15436 15360
rect 16028 15308 16080 15360
rect 16672 15308 16724 15360
rect 16856 15351 16908 15360
rect 16856 15317 16865 15351
rect 16865 15317 16899 15351
rect 16899 15317 16908 15351
rect 16856 15308 16908 15317
rect 18972 15351 19024 15360
rect 18972 15317 18981 15351
rect 18981 15317 19015 15351
rect 19015 15317 19024 15351
rect 18972 15308 19024 15317
rect 19800 15308 19852 15360
rect 20996 15351 21048 15360
rect 20996 15317 21005 15351
rect 21005 15317 21039 15351
rect 21039 15317 21048 15351
rect 20996 15308 21048 15317
rect 22008 15308 22060 15360
rect 22652 15308 22704 15360
rect 24032 15308 24084 15360
rect 26332 15512 26384 15564
rect 26792 15512 26844 15564
rect 26976 15512 27028 15564
rect 27620 15555 27672 15564
rect 27620 15521 27629 15555
rect 27629 15521 27663 15555
rect 27663 15521 27672 15555
rect 27620 15512 27672 15521
rect 26148 15444 26200 15496
rect 26332 15308 26384 15360
rect 26424 15308 26476 15360
rect 26792 15308 26844 15360
rect 26976 15308 27028 15360
rect 27988 15487 28040 15496
rect 27988 15453 27997 15487
rect 27997 15453 28031 15487
rect 28031 15453 28040 15487
rect 27988 15444 28040 15453
rect 28172 15444 28224 15496
rect 28540 15444 28592 15496
rect 28724 15487 28776 15496
rect 28724 15453 28733 15487
rect 28733 15453 28767 15487
rect 28767 15453 28776 15487
rect 28724 15444 28776 15453
rect 30012 15512 30064 15564
rect 31208 15376 31260 15428
rect 28356 15308 28408 15360
rect 4193 15206 4245 15258
rect 4257 15206 4309 15258
rect 4321 15206 4373 15258
rect 4385 15206 4437 15258
rect 4449 15206 4501 15258
rect 11783 15206 11835 15258
rect 11847 15206 11899 15258
rect 11911 15206 11963 15258
rect 11975 15206 12027 15258
rect 12039 15206 12091 15258
rect 19373 15206 19425 15258
rect 19437 15206 19489 15258
rect 19501 15206 19553 15258
rect 19565 15206 19617 15258
rect 19629 15206 19681 15258
rect 26963 15206 27015 15258
rect 27027 15206 27079 15258
rect 27091 15206 27143 15258
rect 27155 15206 27207 15258
rect 27219 15206 27271 15258
rect 1400 15104 1452 15156
rect 2872 15104 2924 15156
rect 5724 15104 5776 15156
rect 5908 15104 5960 15156
rect 1124 14968 1176 15020
rect 1308 14968 1360 15020
rect 3056 14968 3108 15020
rect 3792 15011 3844 15020
rect 3792 14977 3801 15011
rect 3801 14977 3835 15011
rect 3835 14977 3844 15011
rect 3792 14968 3844 14977
rect 8300 15104 8352 15156
rect 13268 15104 13320 15156
rect 14464 15104 14516 15156
rect 10968 15079 11020 15088
rect 10968 15045 10977 15079
rect 10977 15045 11011 15079
rect 11011 15045 11020 15079
rect 10968 15036 11020 15045
rect 14004 15036 14056 15088
rect 15844 15104 15896 15156
rect 8852 14968 8904 15020
rect 10784 14968 10836 15020
rect 11244 15011 11296 15020
rect 11244 14977 11253 15011
rect 11253 14977 11287 15011
rect 11287 14977 11296 15011
rect 11244 14968 11296 14977
rect 3884 14900 3936 14952
rect 4528 14943 4580 14952
rect 4528 14909 4537 14943
rect 4537 14909 4571 14943
rect 4571 14909 4580 14943
rect 4528 14900 4580 14909
rect 5632 14900 5684 14952
rect 6184 14900 6236 14952
rect 6460 14943 6512 14952
rect 6460 14909 6462 14943
rect 6462 14909 6512 14943
rect 6460 14900 6512 14909
rect 6736 14900 6788 14952
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 6920 14900 6972 14952
rect 8392 14900 8444 14952
rect 8668 14943 8720 14952
rect 8668 14909 8677 14943
rect 8677 14909 8711 14943
rect 8711 14909 8720 14943
rect 8668 14900 8720 14909
rect 1676 14764 1728 14816
rect 7564 14832 7616 14884
rect 8484 14832 8536 14884
rect 4068 14764 4120 14816
rect 11336 14900 11388 14952
rect 11980 14943 12032 14952
rect 11980 14909 11989 14943
rect 11989 14909 12023 14943
rect 12023 14909 12032 14943
rect 11980 14900 12032 14909
rect 12808 14900 12860 14952
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 15016 15011 15068 15020
rect 15016 14977 15018 15011
rect 15018 14977 15068 15011
rect 15016 14968 15068 14977
rect 14464 14832 14516 14884
rect 15292 14900 15344 14952
rect 15384 14943 15436 14952
rect 15384 14909 15393 14943
rect 15393 14909 15427 14943
rect 15427 14909 15436 14943
rect 15384 14900 15436 14909
rect 14740 14832 14792 14884
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 17316 14968 17368 15020
rect 19064 14968 19116 15020
rect 19708 15011 19760 15020
rect 16948 14900 17000 14952
rect 17592 14900 17644 14952
rect 18788 14900 18840 14952
rect 19708 14977 19717 15011
rect 19717 14977 19751 15011
rect 19751 14977 19760 15011
rect 19708 14968 19760 14977
rect 20904 14968 20956 15020
rect 21364 15104 21416 15156
rect 23848 15104 23900 15156
rect 26056 15147 26108 15156
rect 26056 15113 26065 15147
rect 26065 15113 26099 15147
rect 26099 15113 26108 15147
rect 26056 15104 26108 15113
rect 27068 15104 27120 15156
rect 27436 15104 27488 15156
rect 28080 15104 28132 15156
rect 28632 15104 28684 15156
rect 29644 15104 29696 15156
rect 30380 15104 30432 15156
rect 31116 15104 31168 15156
rect 23664 14968 23716 15020
rect 24032 14968 24084 15020
rect 24216 15011 24268 15020
rect 24216 14977 24218 15011
rect 24218 14977 24268 15011
rect 24216 14968 24268 14977
rect 24768 14968 24820 15020
rect 9772 14764 9824 14816
rect 10416 14764 10468 14816
rect 10508 14807 10560 14816
rect 10508 14773 10517 14807
rect 10517 14773 10551 14807
rect 10551 14773 10560 14807
rect 10508 14764 10560 14773
rect 10968 14764 11020 14816
rect 11704 14807 11756 14816
rect 11704 14773 11719 14807
rect 11719 14773 11753 14807
rect 11753 14773 11756 14807
rect 11704 14764 11756 14773
rect 13820 14807 13872 14816
rect 13820 14773 13829 14807
rect 13829 14773 13863 14807
rect 13863 14773 13872 14807
rect 13820 14764 13872 14773
rect 16488 14807 16540 14816
rect 16488 14773 16497 14807
rect 16497 14773 16531 14807
rect 16531 14773 16540 14807
rect 16488 14764 16540 14773
rect 16764 14764 16816 14816
rect 19064 14764 19116 14816
rect 19248 14807 19300 14816
rect 19248 14773 19257 14807
rect 19257 14773 19291 14807
rect 19291 14773 19300 14807
rect 19248 14764 19300 14773
rect 21456 14900 21508 14952
rect 22376 14900 22428 14952
rect 23020 14832 23072 14884
rect 25044 14900 25096 14952
rect 26424 14968 26476 15020
rect 29920 15036 29972 15088
rect 27068 15011 27120 15020
rect 26332 14943 26384 14952
rect 26332 14909 26341 14943
rect 26341 14909 26375 14943
rect 26375 14909 26384 14943
rect 26332 14900 26384 14909
rect 25504 14832 25556 14884
rect 26148 14832 26200 14884
rect 26700 14943 26752 14952
rect 26700 14909 26709 14943
rect 26709 14909 26743 14943
rect 26743 14909 26752 14943
rect 26700 14900 26752 14909
rect 27068 14977 27070 15011
rect 27070 14977 27120 15011
rect 27068 14968 27120 14977
rect 27252 14968 27304 15020
rect 27620 14968 27672 15020
rect 27896 14900 27948 14952
rect 20076 14764 20128 14816
rect 20812 14764 20864 14816
rect 20904 14764 20956 14816
rect 21824 14764 21876 14816
rect 22284 14764 22336 14816
rect 26240 14764 26292 14816
rect 26424 14764 26476 14816
rect 28356 14900 28408 14952
rect 29460 14900 29512 14952
rect 30288 14900 30340 14952
rect 28908 14832 28960 14884
rect 29000 14764 29052 14816
rect 30288 14764 30340 14816
rect 30748 14900 30800 14952
rect 30932 14764 30984 14816
rect 7988 14662 8040 14714
rect 8052 14662 8104 14714
rect 8116 14662 8168 14714
rect 8180 14662 8232 14714
rect 8244 14662 8296 14714
rect 15578 14662 15630 14714
rect 15642 14662 15694 14714
rect 15706 14662 15758 14714
rect 15770 14662 15822 14714
rect 15834 14662 15886 14714
rect 23168 14662 23220 14714
rect 23232 14662 23284 14714
rect 23296 14662 23348 14714
rect 23360 14662 23412 14714
rect 23424 14662 23476 14714
rect 30758 14662 30810 14714
rect 30822 14662 30874 14714
rect 30886 14662 30938 14714
rect 30950 14662 31002 14714
rect 31014 14662 31066 14714
rect 940 14560 992 14612
rect 1216 14535 1268 14544
rect 1216 14501 1225 14535
rect 1225 14501 1259 14535
rect 1259 14501 1268 14535
rect 1216 14492 1268 14501
rect 1400 14492 1452 14544
rect 2228 14560 2280 14612
rect 3792 14560 3844 14612
rect 3608 14492 3660 14544
rect 4436 14560 4488 14612
rect 4528 14560 4580 14612
rect 4712 14560 4764 14612
rect 5448 14603 5500 14612
rect 5448 14569 5457 14603
rect 5457 14569 5491 14603
rect 5491 14569 5500 14603
rect 5448 14560 5500 14569
rect 6184 14560 6236 14612
rect 6828 14560 6880 14612
rect 7380 14560 7432 14612
rect 8300 14560 8352 14612
rect 9312 14560 9364 14612
rect 9404 14603 9456 14612
rect 9404 14569 9413 14603
rect 9413 14569 9447 14603
rect 9447 14569 9456 14603
rect 9404 14560 9456 14569
rect 10416 14560 10468 14612
rect 1400 14356 1452 14408
rect 1676 14356 1728 14408
rect 1952 14356 2004 14408
rect 2136 14356 2188 14408
rect 2596 14356 2648 14408
rect 4988 14424 5040 14476
rect 5540 14492 5592 14544
rect 5908 14424 5960 14476
rect 6279 14424 6331 14476
rect 6644 14492 6696 14544
rect 4804 14288 4856 14340
rect 4896 14331 4948 14340
rect 4896 14297 4905 14331
rect 4905 14297 4939 14331
rect 4939 14297 4948 14331
rect 4896 14288 4948 14297
rect 6276 14288 6328 14340
rect 1768 14220 1820 14272
rect 3332 14220 3384 14272
rect 3516 14263 3568 14272
rect 3516 14229 3525 14263
rect 3525 14229 3559 14263
rect 3559 14229 3568 14263
rect 3516 14220 3568 14229
rect 4620 14220 4672 14272
rect 4988 14220 5040 14272
rect 5724 14220 5776 14272
rect 6828 14399 6880 14408
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 7196 14399 7248 14408
rect 7196 14365 7198 14399
rect 7198 14365 7248 14399
rect 7196 14356 7248 14365
rect 7288 14399 7340 14408
rect 7288 14365 7300 14399
rect 7300 14365 7334 14399
rect 7334 14365 7340 14399
rect 7288 14356 7340 14365
rect 7564 14399 7616 14408
rect 7564 14365 7573 14399
rect 7573 14365 7607 14399
rect 7607 14365 7616 14399
rect 7564 14356 7616 14365
rect 8576 14424 8628 14476
rect 9772 14492 9824 14544
rect 10048 14535 10100 14544
rect 10048 14501 10057 14535
rect 10057 14501 10091 14535
rect 10091 14501 10100 14535
rect 10048 14492 10100 14501
rect 11152 14492 11204 14544
rect 11980 14560 12032 14612
rect 12072 14603 12124 14612
rect 12072 14569 12087 14603
rect 12087 14569 12121 14603
rect 12121 14569 12124 14603
rect 12072 14560 12124 14569
rect 12992 14560 13044 14612
rect 11612 14492 11664 14544
rect 10968 14424 11020 14476
rect 16488 14560 16540 14612
rect 16764 14560 16816 14612
rect 19248 14560 19300 14612
rect 20812 14560 20864 14612
rect 22284 14560 22336 14612
rect 26148 14560 26200 14612
rect 15292 14492 15344 14544
rect 18328 14492 18380 14544
rect 19156 14492 19208 14544
rect 6644 14220 6696 14272
rect 7012 14220 7064 14272
rect 8208 14220 8260 14272
rect 8760 14220 8812 14272
rect 8852 14263 8904 14272
rect 8852 14229 8861 14263
rect 8861 14229 8895 14263
rect 8895 14229 8904 14263
rect 8852 14220 8904 14229
rect 11336 14356 11388 14408
rect 13912 14424 13964 14476
rect 15200 14424 15252 14476
rect 16120 14467 16172 14476
rect 16120 14433 16129 14467
rect 16129 14433 16163 14467
rect 16163 14433 16172 14467
rect 16120 14424 16172 14433
rect 16764 14424 16816 14476
rect 17316 14424 17368 14476
rect 21640 14492 21692 14544
rect 23756 14535 23808 14544
rect 23756 14501 23765 14535
rect 23765 14501 23799 14535
rect 23799 14501 23808 14535
rect 23756 14492 23808 14501
rect 11152 14288 11204 14340
rect 11244 14288 11296 14340
rect 12348 14399 12400 14408
rect 12348 14365 12357 14399
rect 12357 14365 12391 14399
rect 12391 14365 12400 14399
rect 12348 14356 12400 14365
rect 13452 14356 13504 14408
rect 14004 14356 14056 14408
rect 14188 14399 14240 14408
rect 14188 14365 14190 14399
rect 14190 14365 14240 14399
rect 14188 14356 14240 14365
rect 14464 14356 14516 14408
rect 14556 14399 14608 14408
rect 14556 14365 14565 14399
rect 14565 14365 14599 14399
rect 14599 14365 14608 14399
rect 14556 14356 14608 14365
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 9864 14220 9916 14272
rect 14096 14220 14148 14272
rect 14648 14220 14700 14272
rect 14740 14220 14792 14272
rect 16304 14263 16356 14272
rect 16304 14229 16313 14263
rect 16313 14229 16347 14263
rect 16347 14229 16356 14263
rect 16304 14220 16356 14229
rect 18972 14288 19024 14340
rect 19156 14288 19208 14340
rect 19708 14399 19760 14408
rect 19708 14365 19717 14399
rect 19717 14365 19751 14399
rect 19751 14365 19760 14399
rect 19708 14356 19760 14365
rect 21272 14424 21324 14476
rect 22836 14424 22888 14476
rect 23664 14424 23716 14476
rect 24216 14467 24268 14476
rect 24216 14433 24218 14467
rect 24218 14433 24268 14467
rect 24216 14424 24268 14433
rect 24676 14424 24728 14476
rect 26240 14467 26292 14476
rect 26240 14433 26241 14467
rect 26241 14433 26275 14467
rect 26275 14433 26292 14467
rect 26240 14424 26292 14433
rect 26792 14492 26844 14544
rect 27068 14492 27120 14544
rect 27252 14492 27304 14544
rect 27896 14492 27948 14544
rect 22284 14356 22336 14408
rect 24308 14383 24353 14408
rect 24353 14383 24360 14408
rect 24308 14356 24360 14383
rect 24492 14356 24544 14408
rect 24952 14356 25004 14408
rect 27988 14467 28040 14476
rect 27988 14433 27997 14467
rect 27997 14433 28031 14467
rect 28031 14433 28040 14467
rect 27988 14424 28040 14433
rect 28264 14560 28316 14612
rect 29184 14560 29236 14612
rect 29920 14560 29972 14612
rect 30748 14560 30800 14612
rect 29460 14492 29512 14544
rect 28356 14356 28408 14408
rect 29920 14356 29972 14408
rect 21548 14220 21600 14272
rect 27896 14288 27948 14340
rect 22744 14220 22796 14272
rect 23296 14220 23348 14272
rect 25044 14220 25096 14272
rect 26056 14263 26108 14272
rect 26056 14229 26065 14263
rect 26065 14229 26099 14263
rect 26099 14229 26108 14263
rect 26056 14220 26108 14229
rect 26700 14220 26752 14272
rect 26792 14220 26844 14272
rect 27068 14220 27120 14272
rect 27160 14220 27212 14272
rect 27620 14220 27672 14272
rect 4193 14118 4245 14170
rect 4257 14118 4309 14170
rect 4321 14118 4373 14170
rect 4385 14118 4437 14170
rect 4449 14118 4501 14170
rect 11783 14118 11835 14170
rect 11847 14118 11899 14170
rect 11911 14118 11963 14170
rect 11975 14118 12027 14170
rect 12039 14118 12091 14170
rect 19373 14118 19425 14170
rect 19437 14118 19489 14170
rect 19501 14118 19553 14170
rect 19565 14118 19617 14170
rect 19629 14118 19681 14170
rect 26963 14118 27015 14170
rect 27027 14118 27079 14170
rect 27091 14118 27143 14170
rect 27155 14118 27207 14170
rect 27219 14118 27271 14170
rect 3516 14016 3568 14068
rect 4160 14016 4212 14068
rect 7288 14016 7340 14068
rect 756 13880 808 13932
rect 2780 13880 2832 13932
rect 4160 13880 4212 13932
rect 5632 13880 5684 13932
rect 2596 13812 2648 13864
rect 3056 13855 3108 13864
rect 3056 13821 3065 13855
rect 3065 13821 3099 13855
rect 3099 13821 3108 13855
rect 3056 13812 3108 13821
rect 3424 13812 3476 13864
rect 3516 13855 3568 13864
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 5816 13812 5868 13864
rect 6276 13880 6328 13932
rect 6460 13923 6512 13932
rect 6460 13889 6462 13923
rect 6462 13889 6512 13923
rect 6460 13880 6512 13889
rect 9864 14016 9916 14068
rect 9956 14016 10008 14068
rect 11612 14016 11664 14068
rect 12348 14016 12400 14068
rect 12532 14016 12584 14068
rect 13268 14016 13320 14068
rect 14556 14016 14608 14068
rect 8392 13948 8444 14000
rect 6920 13812 6972 13864
rect 8208 13812 8260 13864
rect 8392 13855 8444 13864
rect 8392 13821 8401 13855
rect 8401 13821 8435 13855
rect 8435 13821 8444 13855
rect 8392 13812 8444 13821
rect 9128 13948 9180 14000
rect 11152 13948 11204 14000
rect 11336 13880 11388 13932
rect 11704 13880 11756 13932
rect 12716 13991 12768 14000
rect 12716 13957 12725 13991
rect 12725 13957 12759 13991
rect 12759 13957 12768 13991
rect 12716 13948 12768 13957
rect 14004 13948 14056 14000
rect 9312 13812 9364 13864
rect 9404 13812 9456 13864
rect 9496 13812 9548 13864
rect 10048 13855 10100 13864
rect 10048 13821 10050 13855
rect 10050 13821 10100 13855
rect 10048 13812 10100 13821
rect 10416 13855 10468 13864
rect 10416 13821 10425 13855
rect 10425 13821 10459 13855
rect 10459 13821 10468 13855
rect 10416 13812 10468 13821
rect 10508 13812 10560 13864
rect 11060 13812 11112 13864
rect 11888 13855 11940 13864
rect 11888 13821 11897 13855
rect 11897 13821 11931 13855
rect 11931 13821 11940 13855
rect 11888 13812 11940 13821
rect 5540 13744 5592 13796
rect 7840 13744 7892 13796
rect 11428 13744 11480 13796
rect 11796 13787 11848 13796
rect 11796 13753 11805 13787
rect 11805 13753 11839 13787
rect 11839 13753 11848 13787
rect 11796 13744 11848 13753
rect 1952 13676 2004 13728
rect 3332 13719 3384 13728
rect 3332 13685 3341 13719
rect 3341 13685 3375 13719
rect 3375 13685 3384 13719
rect 3332 13676 3384 13685
rect 3700 13676 3752 13728
rect 3792 13676 3844 13728
rect 3976 13676 4028 13728
rect 4528 13676 4580 13728
rect 6460 13676 6512 13728
rect 6644 13676 6696 13728
rect 8668 13676 8720 13728
rect 12256 13676 12308 13728
rect 13452 13880 13504 13932
rect 13728 13880 13780 13932
rect 13912 13880 13964 13932
rect 13728 13744 13780 13796
rect 14740 13880 14792 13932
rect 16856 14016 16908 14068
rect 18236 14059 18288 14068
rect 18236 14025 18245 14059
rect 18245 14025 18279 14059
rect 18279 14025 18288 14059
rect 18236 14016 18288 14025
rect 19064 14059 19116 14068
rect 19064 14025 19073 14059
rect 19073 14025 19107 14059
rect 19107 14025 19116 14059
rect 19064 14016 19116 14025
rect 16028 13991 16080 14000
rect 16028 13957 16037 13991
rect 16037 13957 16071 13991
rect 16071 13957 16080 13991
rect 16028 13948 16080 13957
rect 18696 13948 18748 14000
rect 16764 13923 16816 13932
rect 16764 13889 16766 13923
rect 16766 13889 16816 13923
rect 16764 13880 16816 13889
rect 21916 14016 21968 14068
rect 24860 14016 24912 14068
rect 26056 14016 26108 14068
rect 26516 14059 26568 14068
rect 26516 14025 26525 14059
rect 26525 14025 26559 14059
rect 26559 14025 26568 14059
rect 26516 14016 26568 14025
rect 26608 14016 26660 14068
rect 27436 14016 27488 14068
rect 27528 14016 27580 14068
rect 29092 14016 29144 14068
rect 29552 14059 29604 14068
rect 29552 14025 29561 14059
rect 29561 14025 29595 14059
rect 29595 14025 29604 14059
rect 29552 14016 29604 14025
rect 29828 14059 29880 14068
rect 29828 14025 29837 14059
rect 29837 14025 29871 14059
rect 29871 14025 29880 14059
rect 29828 14016 29880 14025
rect 31116 14016 31168 14068
rect 21456 13948 21508 14000
rect 24492 13948 24544 14000
rect 20536 13880 20588 13932
rect 24216 13880 24268 13932
rect 14832 13812 14884 13864
rect 13084 13676 13136 13728
rect 14188 13676 14240 13728
rect 14924 13676 14976 13728
rect 16672 13676 16724 13728
rect 17132 13676 17184 13728
rect 19340 13676 19392 13728
rect 19984 13855 20036 13864
rect 19984 13821 19993 13855
rect 19993 13821 20027 13855
rect 20027 13821 20036 13855
rect 19984 13812 20036 13821
rect 20628 13812 20680 13864
rect 20720 13855 20772 13864
rect 20720 13821 20729 13855
rect 20729 13821 20763 13855
rect 20763 13821 20772 13855
rect 20720 13812 20772 13821
rect 22928 13855 22980 13864
rect 22560 13744 22612 13796
rect 20352 13676 20404 13728
rect 20812 13676 20864 13728
rect 21916 13676 21968 13728
rect 22928 13821 22937 13855
rect 22937 13821 22971 13855
rect 22971 13821 22980 13855
rect 22928 13812 22980 13821
rect 22744 13744 22796 13796
rect 23296 13812 23348 13864
rect 23388 13855 23440 13864
rect 23388 13821 23397 13855
rect 23397 13821 23431 13855
rect 23431 13821 23440 13855
rect 23388 13812 23440 13821
rect 23020 13719 23072 13728
rect 23020 13685 23029 13719
rect 23029 13685 23063 13719
rect 23063 13685 23072 13719
rect 23020 13676 23072 13685
rect 23756 13812 23808 13864
rect 23940 13812 23992 13864
rect 24032 13855 24084 13864
rect 24032 13821 24041 13855
rect 24041 13821 24075 13855
rect 24075 13821 24084 13855
rect 24400 13880 24452 13932
rect 24032 13812 24084 13821
rect 24768 13812 24820 13864
rect 26424 13880 26476 13932
rect 27344 13880 27396 13932
rect 29184 13948 29236 14000
rect 30748 13948 30800 14000
rect 29552 13880 29604 13932
rect 29644 13880 29696 13932
rect 25688 13812 25740 13864
rect 26976 13812 27028 13864
rect 27528 13812 27580 13864
rect 28908 13812 28960 13864
rect 29092 13812 29144 13864
rect 24584 13744 24636 13796
rect 24124 13719 24176 13728
rect 24124 13685 24133 13719
rect 24133 13685 24167 13719
rect 24167 13685 24176 13719
rect 24124 13676 24176 13685
rect 26516 13676 26568 13728
rect 27160 13719 27212 13728
rect 27160 13685 27175 13719
rect 27175 13685 27209 13719
rect 27209 13685 27212 13719
rect 29276 13812 29328 13864
rect 31392 13880 31444 13932
rect 30380 13855 30432 13864
rect 30380 13821 30389 13855
rect 30389 13821 30423 13855
rect 30423 13821 30432 13855
rect 30380 13812 30432 13821
rect 29644 13744 29696 13796
rect 30288 13744 30340 13796
rect 27160 13676 27212 13685
rect 29828 13676 29880 13728
rect 7988 13574 8040 13626
rect 8052 13574 8104 13626
rect 8116 13574 8168 13626
rect 8180 13574 8232 13626
rect 8244 13574 8296 13626
rect 15578 13574 15630 13626
rect 15642 13574 15694 13626
rect 15706 13574 15758 13626
rect 15770 13574 15822 13626
rect 15834 13574 15886 13626
rect 23168 13574 23220 13626
rect 23232 13574 23284 13626
rect 23296 13574 23348 13626
rect 23360 13574 23412 13626
rect 23424 13574 23476 13626
rect 30758 13574 30810 13626
rect 30822 13574 30874 13626
rect 30886 13574 30938 13626
rect 30950 13574 31002 13626
rect 31014 13574 31066 13626
rect 1676 13472 1728 13524
rect 3424 13472 3476 13524
rect 3976 13515 4028 13524
rect 3976 13481 3991 13515
rect 3991 13481 4025 13515
rect 4025 13481 4028 13515
rect 3976 13472 4028 13481
rect 5816 13515 5868 13524
rect 5816 13481 5825 13515
rect 5825 13481 5859 13515
rect 5859 13481 5868 13515
rect 5816 13472 5868 13481
rect 6092 13515 6144 13524
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 6920 13472 6972 13524
rect 7196 13472 7248 13524
rect 7840 13472 7892 13524
rect 9220 13472 9272 13524
rect 848 13336 900 13388
rect 1216 13379 1268 13388
rect 1216 13345 1225 13379
rect 1225 13345 1259 13379
rect 1259 13345 1268 13379
rect 1216 13336 1268 13345
rect 1308 13379 1360 13388
rect 1308 13345 1317 13379
rect 1317 13345 1351 13379
rect 1351 13345 1360 13379
rect 1308 13336 1360 13345
rect 5816 13336 5868 13388
rect 6184 13336 6236 13388
rect 6460 13336 6512 13388
rect 6828 13379 6880 13388
rect 6828 13345 6837 13379
rect 6837 13345 6871 13379
rect 6871 13345 6880 13379
rect 6828 13336 6880 13345
rect 8484 13404 8536 13456
rect 9128 13404 9180 13456
rect 8852 13336 8904 13388
rect 9312 13379 9364 13388
rect 9312 13345 9321 13379
rect 9321 13345 9355 13379
rect 9355 13345 9364 13379
rect 9312 13336 9364 13345
rect 9588 13447 9640 13456
rect 9588 13413 9597 13447
rect 9597 13413 9631 13447
rect 9631 13413 9640 13447
rect 9588 13404 9640 13413
rect 11152 13515 11204 13524
rect 11152 13481 11161 13515
rect 11161 13481 11195 13515
rect 11195 13481 11204 13515
rect 11152 13472 11204 13481
rect 11796 13472 11848 13524
rect 9864 13379 9916 13388
rect 9864 13345 9873 13379
rect 9873 13345 9907 13379
rect 9907 13345 9916 13379
rect 9864 13336 9916 13345
rect 10968 13379 11020 13388
rect 10968 13345 10977 13379
rect 10977 13345 11011 13379
rect 11011 13345 11020 13379
rect 10968 13336 11020 13345
rect 11428 13336 11480 13388
rect 11612 13336 11664 13388
rect 11704 13336 11756 13388
rect 14464 13472 14516 13524
rect 14924 13404 14976 13456
rect 15384 13472 15436 13524
rect 20352 13472 20404 13524
rect 20720 13472 20772 13524
rect 21916 13472 21968 13524
rect 16764 13404 16816 13456
rect 2228 13268 2280 13320
rect 3792 13268 3844 13320
rect 3976 13311 4028 13320
rect 3976 13277 3988 13311
rect 3988 13277 4022 13311
rect 4022 13277 4028 13311
rect 3976 13268 4028 13277
rect 5080 13268 5132 13320
rect 7196 13268 7248 13320
rect 7288 13311 7340 13320
rect 7288 13277 7300 13311
rect 7300 13277 7334 13311
rect 7334 13277 7340 13311
rect 7288 13268 7340 13277
rect 8760 13268 8812 13320
rect 9128 13268 9180 13320
rect 5356 13200 5408 13252
rect 6276 13200 6328 13252
rect 6368 13200 6420 13252
rect 6736 13200 6788 13252
rect 9496 13200 9548 13252
rect 10140 13200 10192 13252
rect 10692 13268 10744 13320
rect 11060 13268 11112 13320
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 11336 13268 11388 13320
rect 12348 13268 12400 13320
rect 12440 13311 12492 13320
rect 12440 13277 12449 13311
rect 12449 13277 12483 13311
rect 12483 13277 12492 13311
rect 12440 13268 12492 13277
rect 12808 13311 12860 13320
rect 12808 13277 12810 13311
rect 12810 13277 12860 13311
rect 12808 13268 12860 13277
rect 13084 13336 13136 13388
rect 12992 13268 13044 13320
rect 15108 13336 15160 13388
rect 15476 13336 15528 13388
rect 16304 13379 16356 13388
rect 16304 13345 16313 13379
rect 16313 13345 16347 13379
rect 16347 13345 16356 13379
rect 16304 13336 16356 13345
rect 1584 13132 1636 13184
rect 3148 13132 3200 13184
rect 3516 13132 3568 13184
rect 6092 13132 6144 13184
rect 7104 13132 7156 13184
rect 7656 13132 7708 13184
rect 9220 13132 9272 13184
rect 9312 13132 9364 13184
rect 10600 13175 10652 13184
rect 10600 13141 10609 13175
rect 10609 13141 10643 13175
rect 10643 13141 10652 13175
rect 10600 13132 10652 13141
rect 13360 13132 13412 13184
rect 13820 13132 13872 13184
rect 14004 13132 14056 13184
rect 14740 13200 14792 13252
rect 16580 13336 16632 13388
rect 18696 13336 18748 13388
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 20904 13336 20956 13388
rect 21272 13336 21324 13388
rect 21640 13336 21692 13388
rect 23940 13515 23992 13524
rect 23940 13481 23949 13515
rect 23949 13481 23983 13515
rect 23983 13481 23992 13515
rect 23940 13472 23992 13481
rect 24124 13472 24176 13524
rect 26976 13472 27028 13524
rect 27436 13472 27488 13524
rect 29276 13472 29328 13524
rect 29736 13472 29788 13524
rect 23848 13404 23900 13456
rect 24216 13404 24268 13456
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 19892 13268 19944 13320
rect 22100 13268 22152 13320
rect 22376 13311 22428 13320
rect 22376 13277 22388 13311
rect 22388 13277 22422 13311
rect 22422 13277 22428 13311
rect 22376 13268 22428 13277
rect 22652 13311 22704 13320
rect 22652 13277 22661 13311
rect 22661 13277 22695 13311
rect 22695 13277 22704 13311
rect 22652 13268 22704 13277
rect 24308 13268 24360 13320
rect 24860 13379 24912 13388
rect 24860 13345 24869 13379
rect 24869 13345 24903 13379
rect 24903 13345 24912 13379
rect 24860 13336 24912 13345
rect 24768 13268 24820 13320
rect 26424 13311 26476 13320
rect 26424 13277 26433 13311
rect 26433 13277 26467 13311
rect 26467 13277 26476 13311
rect 26424 13268 26476 13277
rect 26608 13268 26660 13320
rect 26792 13311 26844 13320
rect 26792 13277 26794 13311
rect 26794 13277 26844 13311
rect 26792 13268 26844 13277
rect 26976 13336 27028 13388
rect 16212 13132 16264 13184
rect 16672 13175 16724 13184
rect 16672 13141 16681 13175
rect 16681 13141 16715 13175
rect 16715 13141 16724 13175
rect 16672 13132 16724 13141
rect 17408 13132 17460 13184
rect 19708 13132 19760 13184
rect 20168 13132 20220 13184
rect 24032 13200 24084 13252
rect 22284 13132 22336 13184
rect 23020 13132 23072 13184
rect 26792 13132 26844 13184
rect 28632 13311 28684 13320
rect 28632 13277 28641 13311
rect 28641 13277 28675 13311
rect 28675 13277 28684 13311
rect 28632 13268 28684 13277
rect 29828 13268 29880 13320
rect 28908 13132 28960 13184
rect 30288 13132 30340 13184
rect 4193 13030 4245 13082
rect 4257 13030 4309 13082
rect 4321 13030 4373 13082
rect 4385 13030 4437 13082
rect 4449 13030 4501 13082
rect 11783 13030 11835 13082
rect 11847 13030 11899 13082
rect 11911 13030 11963 13082
rect 11975 13030 12027 13082
rect 12039 13030 12091 13082
rect 19373 13030 19425 13082
rect 19437 13030 19489 13082
rect 19501 13030 19553 13082
rect 19565 13030 19617 13082
rect 19629 13030 19681 13082
rect 26963 13030 27015 13082
rect 27027 13030 27079 13082
rect 27091 13030 27143 13082
rect 27155 13030 27207 13082
rect 27219 13030 27271 13082
rect 1216 12928 1268 12980
rect 1308 12792 1360 12844
rect 1584 12792 1636 12844
rect 4252 12928 4304 12980
rect 7288 12928 7340 12980
rect 8760 12971 8812 12980
rect 8760 12937 8769 12971
rect 8769 12937 8803 12971
rect 8803 12937 8812 12971
rect 8760 12928 8812 12937
rect 3424 12860 3476 12912
rect 8392 12860 8444 12912
rect 2320 12724 2372 12776
rect 2964 12724 3016 12776
rect 3424 12767 3476 12776
rect 3424 12733 3433 12767
rect 3433 12733 3467 12767
rect 3467 12733 3476 12767
rect 3424 12724 3476 12733
rect 3608 12724 3660 12776
rect 4252 12792 4304 12844
rect 5632 12792 5684 12844
rect 6736 12792 6788 12844
rect 6644 12724 6696 12776
rect 1676 12588 1728 12640
rect 3516 12588 3568 12640
rect 4528 12588 4580 12640
rect 6920 12588 6972 12640
rect 7840 12724 7892 12776
rect 8576 12724 8628 12776
rect 8760 12724 8812 12776
rect 9220 12928 9272 12980
rect 11244 12928 11296 12980
rect 12072 12971 12124 12980
rect 12072 12937 12081 12971
rect 12081 12937 12115 12971
rect 12115 12937 12124 12971
rect 12072 12928 12124 12937
rect 12348 12928 12400 12980
rect 9404 12860 9456 12912
rect 9956 12792 10008 12844
rect 10876 12792 10928 12844
rect 11704 12792 11756 12844
rect 13360 12860 13412 12912
rect 11244 12724 11296 12776
rect 9680 12588 9732 12640
rect 9956 12588 10008 12640
rect 10692 12588 10744 12640
rect 11336 12588 11388 12640
rect 12900 12724 12952 12776
rect 11796 12656 11848 12708
rect 13176 12724 13228 12776
rect 13452 12724 13504 12776
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 13820 12792 13872 12844
rect 15108 12928 15160 12980
rect 17316 12928 17368 12980
rect 21640 12928 21692 12980
rect 22652 12928 22704 12980
rect 19340 12860 19392 12912
rect 19708 12903 19760 12912
rect 19708 12869 19717 12903
rect 19717 12869 19751 12903
rect 19751 12869 19760 12903
rect 19708 12860 19760 12869
rect 19892 12860 19944 12912
rect 22376 12860 22428 12912
rect 22560 12860 22612 12912
rect 16396 12767 16448 12776
rect 16396 12733 16405 12767
rect 16405 12733 16439 12767
rect 16439 12733 16448 12767
rect 16396 12724 16448 12733
rect 16028 12656 16080 12708
rect 19064 12767 19116 12776
rect 19064 12733 19073 12767
rect 19073 12733 19107 12767
rect 19107 12733 19116 12767
rect 19064 12724 19116 12733
rect 20168 12792 20220 12844
rect 20628 12792 20680 12844
rect 23756 12928 23808 12980
rect 24952 12928 25004 12980
rect 25596 12928 25648 12980
rect 25688 12971 25740 12980
rect 25688 12937 25697 12971
rect 25697 12937 25731 12971
rect 25731 12937 25740 12971
rect 25688 12928 25740 12937
rect 27160 12928 27212 12980
rect 29920 12971 29972 12980
rect 29920 12937 29929 12971
rect 29929 12937 29963 12971
rect 29963 12937 29972 12971
rect 29920 12928 29972 12937
rect 30380 12971 30432 12980
rect 30380 12937 30389 12971
rect 30389 12937 30423 12971
rect 30423 12937 30432 12971
rect 30380 12928 30432 12937
rect 27712 12860 27764 12912
rect 19432 12724 19484 12776
rect 20076 12724 20128 12776
rect 20260 12724 20312 12776
rect 22928 12767 22980 12776
rect 22928 12733 22937 12767
rect 22937 12733 22971 12767
rect 22971 12733 22980 12767
rect 22928 12724 22980 12733
rect 23756 12724 23808 12776
rect 23848 12767 23900 12776
rect 23848 12733 23857 12767
rect 23857 12733 23891 12767
rect 23891 12733 23900 12767
rect 23848 12724 23900 12733
rect 24032 12792 24084 12844
rect 25596 12792 25648 12844
rect 26700 12792 26752 12844
rect 27160 12792 27212 12844
rect 30288 12792 30340 12844
rect 24860 12724 24912 12776
rect 25872 12724 25924 12776
rect 26424 12724 26476 12776
rect 27988 12724 28040 12776
rect 23572 12656 23624 12708
rect 23940 12656 23992 12708
rect 26148 12656 26200 12708
rect 27528 12656 27580 12708
rect 11980 12588 12032 12640
rect 13084 12588 13136 12640
rect 14188 12588 14240 12640
rect 16856 12631 16908 12640
rect 16856 12597 16871 12631
rect 16871 12597 16905 12631
rect 16905 12597 16908 12631
rect 16856 12588 16908 12597
rect 17408 12588 17460 12640
rect 18788 12588 18840 12640
rect 18880 12631 18932 12640
rect 18880 12597 18889 12631
rect 18889 12597 18923 12631
rect 18923 12597 18932 12631
rect 18880 12588 18932 12597
rect 19340 12588 19392 12640
rect 19800 12588 19852 12640
rect 19984 12588 20036 12640
rect 20812 12588 20864 12640
rect 22008 12588 22060 12640
rect 22836 12588 22888 12640
rect 24124 12588 24176 12640
rect 24308 12631 24360 12640
rect 24308 12597 24323 12631
rect 24323 12597 24357 12631
rect 24357 12597 24360 12631
rect 24308 12588 24360 12597
rect 26884 12588 26936 12640
rect 27436 12588 27488 12640
rect 29000 12656 29052 12708
rect 29184 12656 29236 12708
rect 30380 12724 30432 12776
rect 29644 12699 29696 12708
rect 29644 12665 29653 12699
rect 29653 12665 29687 12699
rect 29687 12665 29696 12699
rect 29644 12656 29696 12665
rect 29460 12588 29512 12640
rect 29736 12631 29788 12640
rect 29736 12597 29745 12631
rect 29745 12597 29779 12631
rect 29779 12597 29788 12631
rect 29736 12588 29788 12597
rect 7988 12486 8040 12538
rect 8052 12486 8104 12538
rect 8116 12486 8168 12538
rect 8180 12486 8232 12538
rect 8244 12486 8296 12538
rect 15578 12486 15630 12538
rect 15642 12486 15694 12538
rect 15706 12486 15758 12538
rect 15770 12486 15822 12538
rect 15834 12486 15886 12538
rect 23168 12486 23220 12538
rect 23232 12486 23284 12538
rect 23296 12486 23348 12538
rect 23360 12486 23412 12538
rect 23424 12486 23476 12538
rect 30758 12486 30810 12538
rect 30822 12486 30874 12538
rect 30886 12486 30938 12538
rect 30950 12486 31002 12538
rect 31014 12486 31066 12538
rect 3148 12384 3200 12436
rect 3240 12384 3292 12436
rect 3792 12384 3844 12436
rect 3976 12427 4028 12436
rect 3976 12393 3991 12427
rect 3991 12393 4025 12427
rect 4025 12393 4028 12427
rect 3976 12384 4028 12393
rect 4528 12384 4580 12436
rect 5632 12384 5684 12436
rect 5724 12384 5776 12436
rect 5908 12384 5960 12436
rect 6276 12384 6328 12436
rect 8300 12384 8352 12436
rect 8484 12384 8536 12436
rect 1308 12291 1360 12300
rect 1308 12257 1317 12291
rect 1317 12257 1351 12291
rect 1351 12257 1360 12291
rect 1308 12248 1360 12257
rect 1676 12291 1728 12300
rect 1676 12257 1678 12291
rect 1678 12257 1728 12291
rect 1676 12248 1728 12257
rect 11244 12427 11296 12436
rect 11244 12393 11253 12427
rect 11253 12393 11287 12427
rect 11287 12393 11296 12427
rect 11244 12384 11296 12393
rect 12164 12384 12216 12436
rect 12900 12384 12952 12436
rect 13268 12384 13320 12436
rect 14188 12384 14240 12436
rect 15200 12384 15252 12436
rect 15936 12384 15988 12436
rect 16580 12384 16632 12436
rect 1768 12207 1813 12232
rect 1813 12207 1820 12232
rect 1768 12180 1820 12207
rect 1952 12180 2004 12232
rect 3240 12180 3292 12232
rect 3516 12223 3568 12232
rect 3516 12189 3525 12223
rect 3525 12189 3559 12223
rect 3559 12189 3568 12223
rect 3516 12180 3568 12189
rect 3884 12180 3936 12232
rect 4068 12180 4120 12232
rect 5080 12180 5132 12232
rect 6368 12248 6420 12300
rect 6460 12291 6512 12300
rect 6460 12257 6469 12291
rect 6469 12257 6503 12291
rect 6503 12257 6512 12291
rect 6460 12248 6512 12257
rect 3332 12112 3384 12164
rect 6644 12180 6696 12232
rect 6828 12223 6880 12232
rect 6828 12189 6830 12223
rect 6830 12189 6880 12223
rect 6828 12180 6880 12189
rect 6920 12223 6972 12232
rect 6920 12189 6932 12223
rect 6932 12189 6966 12223
rect 6966 12189 6972 12223
rect 6920 12180 6972 12189
rect 7104 12248 7156 12300
rect 7472 12248 7524 12300
rect 9864 12248 9916 12300
rect 11152 12291 11204 12300
rect 11152 12257 11161 12291
rect 11161 12257 11195 12291
rect 11195 12257 11204 12291
rect 11152 12248 11204 12257
rect 11796 12248 11848 12300
rect 8576 12180 8628 12232
rect 6184 12112 6236 12164
rect 1952 12044 2004 12096
rect 4068 12044 4120 12096
rect 6092 12087 6144 12096
rect 6092 12053 6101 12087
rect 6101 12053 6135 12087
rect 6135 12053 6144 12087
rect 6092 12044 6144 12053
rect 8024 12044 8076 12096
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 8852 12180 8904 12232
rect 9128 12223 9180 12232
rect 9128 12189 9140 12223
rect 9140 12189 9174 12223
rect 9174 12189 9180 12223
rect 9128 12180 9180 12189
rect 12072 12248 12124 12300
rect 12440 12291 12492 12300
rect 12440 12257 12449 12291
rect 12449 12257 12483 12291
rect 12483 12257 12492 12291
rect 12440 12248 12492 12257
rect 12808 12291 12860 12300
rect 12808 12257 12810 12291
rect 12810 12257 12860 12291
rect 12808 12248 12860 12257
rect 10692 12155 10744 12164
rect 10692 12121 10701 12155
rect 10701 12121 10735 12155
rect 10735 12121 10744 12155
rect 10692 12112 10744 12121
rect 12624 12180 12676 12232
rect 13452 12248 13504 12300
rect 14832 12248 14884 12300
rect 19064 12384 19116 12436
rect 20168 12384 20220 12436
rect 20260 12427 20312 12436
rect 20260 12393 20269 12427
rect 20269 12393 20303 12427
rect 20303 12393 20312 12427
rect 20260 12384 20312 12393
rect 20628 12384 20680 12436
rect 22008 12384 22060 12436
rect 23112 12427 23164 12436
rect 23112 12393 23121 12427
rect 23121 12393 23155 12427
rect 23155 12393 23164 12427
rect 23112 12384 23164 12393
rect 17408 12291 17460 12300
rect 17408 12257 17417 12291
rect 17417 12257 17451 12291
rect 17451 12257 17460 12291
rect 17408 12248 17460 12257
rect 13268 12180 13320 12232
rect 13360 12180 13412 12232
rect 9404 12044 9456 12096
rect 10600 12044 10652 12096
rect 11060 12044 11112 12096
rect 14280 12180 14332 12232
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 16580 12180 16632 12232
rect 17868 12180 17920 12232
rect 17960 12223 18012 12232
rect 17960 12189 17969 12223
rect 17969 12189 18003 12223
rect 18003 12189 18012 12223
rect 17960 12180 18012 12189
rect 18420 12223 18472 12232
rect 18420 12189 18432 12223
rect 18432 12189 18466 12223
rect 18466 12189 18472 12223
rect 18420 12180 18472 12189
rect 18696 12291 18748 12300
rect 18696 12257 18705 12291
rect 18705 12257 18739 12291
rect 18739 12257 18748 12291
rect 18696 12248 18748 12257
rect 21180 12248 21232 12300
rect 23848 12384 23900 12436
rect 25596 12384 25648 12436
rect 25780 12384 25832 12436
rect 27528 12384 27580 12436
rect 27620 12384 27672 12436
rect 28448 12384 28500 12436
rect 19064 12180 19116 12232
rect 19892 12180 19944 12232
rect 21548 12180 21600 12232
rect 21824 12180 21876 12232
rect 23940 12223 23992 12232
rect 23940 12189 23952 12223
rect 23952 12189 23986 12223
rect 23986 12189 23992 12223
rect 23940 12180 23992 12189
rect 24124 12248 24176 12300
rect 25780 12291 25832 12300
rect 25780 12257 25789 12291
rect 25789 12257 25823 12291
rect 25823 12257 25832 12291
rect 25780 12248 25832 12257
rect 26516 12248 26568 12300
rect 24308 12180 24360 12232
rect 14096 12044 14148 12096
rect 17040 12087 17092 12096
rect 17040 12053 17049 12087
rect 17049 12053 17083 12087
rect 17083 12053 17092 12087
rect 17040 12044 17092 12053
rect 18328 12044 18380 12096
rect 19432 12044 19484 12096
rect 20996 12044 21048 12096
rect 25780 12044 25832 12096
rect 26332 12044 26384 12096
rect 26884 12223 26936 12232
rect 26884 12189 26896 12223
rect 26896 12189 26930 12223
rect 26930 12189 26936 12223
rect 26884 12180 26936 12189
rect 27160 12291 27212 12300
rect 27160 12257 27169 12291
rect 27169 12257 27203 12291
rect 27203 12257 27212 12291
rect 27160 12248 27212 12257
rect 27988 12248 28040 12300
rect 28908 12291 28960 12300
rect 28908 12257 28917 12291
rect 28917 12257 28951 12291
rect 28951 12257 28960 12291
rect 28908 12248 28960 12257
rect 29736 12248 29788 12300
rect 27804 12180 27856 12232
rect 28264 12112 28316 12164
rect 27620 12044 27672 12096
rect 28908 12044 28960 12096
rect 4193 11942 4245 11994
rect 4257 11942 4309 11994
rect 4321 11942 4373 11994
rect 4385 11942 4437 11994
rect 4449 11942 4501 11994
rect 11783 11942 11835 11994
rect 11847 11942 11899 11994
rect 11911 11942 11963 11994
rect 11975 11942 12027 11994
rect 12039 11942 12091 11994
rect 19373 11942 19425 11994
rect 19437 11942 19489 11994
rect 19501 11942 19553 11994
rect 19565 11942 19617 11994
rect 19629 11942 19681 11994
rect 26963 11942 27015 11994
rect 27027 11942 27079 11994
rect 27091 11942 27143 11994
rect 27155 11942 27207 11994
rect 27219 11942 27271 11994
rect 1400 11840 1452 11892
rect 2872 11840 2924 11892
rect 2044 11704 2096 11756
rect 3516 11704 3568 11756
rect 6092 11840 6144 11892
rect 6920 11840 6972 11892
rect 7564 11840 7616 11892
rect 8576 11840 8628 11892
rect 9036 11840 9088 11892
rect 940 11679 992 11688
rect 940 11645 949 11679
rect 949 11645 983 11679
rect 983 11645 992 11679
rect 940 11636 992 11645
rect 1676 11679 1728 11688
rect 1676 11645 1685 11679
rect 1685 11645 1719 11679
rect 1719 11645 1728 11679
rect 1676 11636 1728 11645
rect 3240 11636 3292 11688
rect 3608 11636 3660 11688
rect 4712 11636 4764 11688
rect 5540 11679 5592 11688
rect 5540 11645 5549 11679
rect 5549 11645 5583 11679
rect 5583 11645 5592 11679
rect 5540 11636 5592 11645
rect 6092 11704 6144 11756
rect 11520 11883 11572 11892
rect 11520 11849 11529 11883
rect 11529 11849 11563 11883
rect 11563 11849 11572 11883
rect 11520 11840 11572 11849
rect 12348 11883 12400 11892
rect 12348 11849 12357 11883
rect 12357 11849 12391 11883
rect 12391 11849 12400 11883
rect 12348 11840 12400 11849
rect 12992 11840 13044 11892
rect 13084 11840 13136 11892
rect 9680 11772 9732 11824
rect 11336 11772 11388 11824
rect 12716 11772 12768 11824
rect 7840 11704 7892 11756
rect 6276 11679 6328 11688
rect 6276 11645 6285 11679
rect 6285 11645 6319 11679
rect 6319 11645 6328 11679
rect 6276 11636 6328 11645
rect 6644 11636 6696 11688
rect 8024 11636 8076 11688
rect 2872 11500 2924 11552
rect 3976 11500 4028 11552
rect 4068 11500 4120 11552
rect 5632 11500 5684 11552
rect 6736 11500 6788 11552
rect 7012 11500 7064 11552
rect 7564 11500 7616 11552
rect 8300 11636 8352 11688
rect 8484 11704 8536 11756
rect 10600 11704 10652 11756
rect 8760 11636 8812 11688
rect 9312 11636 9364 11688
rect 9404 11636 9456 11688
rect 10784 11636 10836 11688
rect 12256 11636 12308 11688
rect 13176 11772 13228 11824
rect 13268 11704 13320 11756
rect 14188 11704 14240 11756
rect 14280 11747 14332 11756
rect 14280 11713 14289 11747
rect 14289 11713 14323 11747
rect 14323 11713 14332 11747
rect 14280 11704 14332 11713
rect 13084 11636 13136 11688
rect 13544 11679 13596 11688
rect 13544 11645 13553 11679
rect 13553 11645 13587 11679
rect 13587 11645 13596 11679
rect 13544 11636 13596 11645
rect 13636 11636 13688 11688
rect 8852 11500 8904 11552
rect 9956 11500 10008 11552
rect 10048 11500 10100 11552
rect 10324 11500 10376 11552
rect 15844 11636 15896 11688
rect 18328 11840 18380 11892
rect 18420 11883 18472 11892
rect 18420 11849 18429 11883
rect 18429 11849 18463 11883
rect 18463 11849 18472 11883
rect 18420 11840 18472 11849
rect 17868 11772 17920 11824
rect 20536 11883 20588 11892
rect 20536 11849 20545 11883
rect 20545 11849 20579 11883
rect 20579 11849 20588 11883
rect 20536 11840 20588 11849
rect 21548 11840 21600 11892
rect 20996 11772 21048 11824
rect 16672 11636 16724 11688
rect 17040 11704 17092 11756
rect 17960 11704 18012 11756
rect 18696 11747 18748 11756
rect 18696 11713 18705 11747
rect 18705 11713 18739 11747
rect 18739 11713 18748 11747
rect 18696 11704 18748 11713
rect 17868 11636 17920 11688
rect 19340 11704 19392 11756
rect 23940 11840 23992 11892
rect 25688 11840 25740 11892
rect 26884 11840 26936 11892
rect 26976 11840 27028 11892
rect 24308 11704 24360 11756
rect 28448 11772 28500 11824
rect 28816 11840 28868 11892
rect 29552 11772 29604 11824
rect 26516 11704 26568 11756
rect 19892 11636 19944 11688
rect 21180 11636 21232 11688
rect 22284 11679 22336 11688
rect 22284 11645 22293 11679
rect 22293 11645 22327 11679
rect 22327 11645 22336 11679
rect 22284 11636 22336 11645
rect 22928 11636 22980 11688
rect 23940 11679 23992 11688
rect 23940 11645 23949 11679
rect 23949 11645 23983 11679
rect 23983 11645 23992 11679
rect 23940 11636 23992 11645
rect 24860 11636 24912 11688
rect 25228 11679 25280 11688
rect 25228 11645 25237 11679
rect 25237 11645 25271 11679
rect 25271 11645 25280 11679
rect 25228 11636 25280 11645
rect 25504 11636 25556 11688
rect 28724 11704 28776 11756
rect 15200 11500 15252 11552
rect 15936 11543 15988 11552
rect 15936 11509 15945 11543
rect 15945 11509 15979 11543
rect 15979 11509 15988 11543
rect 15936 11500 15988 11509
rect 16120 11543 16172 11552
rect 16120 11509 16129 11543
rect 16129 11509 16163 11543
rect 16163 11509 16172 11543
rect 16120 11500 16172 11509
rect 17132 11500 17184 11552
rect 18788 11500 18840 11552
rect 19064 11500 19116 11552
rect 28540 11568 28592 11620
rect 29000 11568 29052 11620
rect 21088 11543 21140 11552
rect 21088 11509 21097 11543
rect 21097 11509 21131 11543
rect 21131 11509 21140 11543
rect 21088 11500 21140 11509
rect 21640 11500 21692 11552
rect 22008 11543 22060 11552
rect 22008 11509 22023 11543
rect 22023 11509 22057 11543
rect 22057 11509 22060 11543
rect 22008 11500 22060 11509
rect 26976 11500 27028 11552
rect 27528 11500 27580 11552
rect 27712 11500 27764 11552
rect 29644 11636 29696 11688
rect 30380 11636 30432 11688
rect 31300 11636 31352 11688
rect 29644 11500 29696 11552
rect 30288 11500 30340 11552
rect 7988 11398 8040 11450
rect 8052 11398 8104 11450
rect 8116 11398 8168 11450
rect 8180 11398 8232 11450
rect 8244 11398 8296 11450
rect 15578 11398 15630 11450
rect 15642 11398 15694 11450
rect 15706 11398 15758 11450
rect 15770 11398 15822 11450
rect 15834 11398 15886 11450
rect 23168 11398 23220 11450
rect 23232 11398 23284 11450
rect 23296 11398 23348 11450
rect 23360 11398 23412 11450
rect 23424 11398 23476 11450
rect 30758 11398 30810 11450
rect 30822 11398 30874 11450
rect 30886 11398 30938 11450
rect 30950 11398 31002 11450
rect 31014 11398 31066 11450
rect 1400 11339 1452 11348
rect 1400 11305 1409 11339
rect 1409 11305 1443 11339
rect 1443 11305 1452 11339
rect 1400 11296 1452 11305
rect 1768 11296 1820 11348
rect 2136 11296 2188 11348
rect 664 11228 716 11280
rect 3608 11296 3660 11348
rect 3884 11296 3936 11348
rect 4988 11296 5040 11348
rect 6000 11296 6052 11348
rect 6276 11296 6328 11348
rect 1308 11160 1360 11212
rect 2136 11160 2188 11212
rect 1952 11092 2004 11144
rect 3976 11271 4028 11280
rect 3976 11237 3985 11271
rect 3985 11237 4019 11271
rect 4019 11237 4028 11271
rect 3976 11228 4028 11237
rect 3608 11024 3660 11076
rect 4620 11160 4672 11212
rect 4712 11203 4764 11212
rect 4712 11169 4721 11203
rect 4721 11169 4755 11203
rect 4755 11169 4764 11203
rect 4712 11160 4764 11169
rect 3792 11092 3844 11144
rect 4068 11024 4120 11076
rect 1676 10956 1728 11008
rect 4528 10956 4580 11008
rect 5448 11160 5500 11212
rect 5724 11160 5776 11212
rect 5816 11160 5868 11212
rect 6736 11228 6788 11280
rect 9128 11296 9180 11348
rect 9404 11296 9456 11348
rect 10416 11296 10468 11348
rect 10692 11296 10744 11348
rect 6920 11160 6972 11212
rect 7564 11203 7616 11212
rect 7564 11169 7573 11203
rect 7573 11169 7607 11203
rect 7607 11169 7616 11203
rect 7564 11160 7616 11169
rect 7656 11160 7708 11212
rect 6644 11092 6696 11144
rect 7288 11137 7340 11144
rect 7288 11103 7300 11137
rect 7300 11103 7334 11137
rect 7334 11103 7340 11137
rect 7288 11092 7340 11103
rect 9312 11160 9364 11212
rect 9496 11160 9548 11212
rect 10784 11228 10836 11280
rect 10968 11228 11020 11280
rect 10048 11160 10100 11212
rect 10600 11160 10652 11212
rect 10692 11203 10744 11212
rect 10692 11169 10701 11203
rect 10701 11169 10735 11203
rect 10735 11169 10744 11203
rect 10692 11160 10744 11169
rect 5356 11024 5408 11076
rect 6460 10999 6512 11008
rect 6460 10965 6469 10999
rect 6469 10965 6503 10999
rect 6503 10965 6512 10999
rect 6460 10956 6512 10965
rect 9128 11024 9180 11076
rect 9312 11024 9364 11076
rect 10140 11092 10192 11144
rect 12164 11160 12216 11212
rect 14648 11296 14700 11348
rect 16120 11296 16172 11348
rect 18604 11296 18656 11348
rect 18788 11339 18840 11348
rect 18788 11305 18797 11339
rect 18797 11305 18831 11339
rect 18831 11305 18840 11339
rect 18788 11296 18840 11305
rect 10508 11067 10560 11076
rect 10508 11033 10517 11067
rect 10517 11033 10551 11067
rect 10551 11033 10560 11067
rect 10508 11024 10560 11033
rect 10968 11067 11020 11076
rect 10968 11033 10977 11067
rect 10977 11033 11011 11067
rect 11011 11033 11020 11067
rect 10968 11024 11020 11033
rect 11612 11024 11664 11076
rect 11152 10956 11204 11008
rect 12440 11135 12492 11144
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 12440 11092 12492 11101
rect 12808 11135 12860 11144
rect 12808 11101 12810 11135
rect 12810 11101 12860 11135
rect 12808 11092 12860 11101
rect 13084 11160 13136 11212
rect 14832 11203 14884 11212
rect 14832 11169 14841 11203
rect 14841 11169 14875 11203
rect 14875 11169 14884 11203
rect 14832 11160 14884 11169
rect 15476 11160 15528 11212
rect 16580 11092 16632 11144
rect 16672 11092 16724 11144
rect 16948 11092 17000 11144
rect 17132 11135 17184 11144
rect 17132 11101 17134 11135
rect 17134 11101 17184 11135
rect 17132 11092 17184 11101
rect 20536 11296 20588 11348
rect 21824 11296 21876 11348
rect 22928 11296 22980 11348
rect 19064 11228 19116 11280
rect 19524 11160 19576 11212
rect 20628 11160 20680 11212
rect 25504 11296 25556 11348
rect 26148 11296 26200 11348
rect 29000 11296 29052 11348
rect 29552 11296 29604 11348
rect 30380 11296 30432 11348
rect 11796 11067 11848 11076
rect 11796 11033 11805 11067
rect 11805 11033 11839 11067
rect 11839 11033 11848 11067
rect 11796 11024 11848 11033
rect 12256 11024 12308 11076
rect 14648 11067 14700 11076
rect 14648 11033 14657 11067
rect 14657 11033 14691 11067
rect 14691 11033 14700 11067
rect 14648 11024 14700 11033
rect 14924 11067 14976 11076
rect 14924 11033 14933 11067
rect 14933 11033 14967 11067
rect 14967 11033 14976 11067
rect 14924 11024 14976 11033
rect 15476 11067 15528 11076
rect 15476 11033 15485 11067
rect 15485 11033 15519 11067
rect 15519 11033 15528 11067
rect 15476 11024 15528 11033
rect 16212 11024 16264 11076
rect 18696 11024 18748 11076
rect 19156 11092 19208 11144
rect 21548 11092 21600 11144
rect 22008 11092 22060 11144
rect 22100 11092 22152 11144
rect 22376 11092 22428 11144
rect 23572 11092 23624 11144
rect 13544 10956 13596 11008
rect 14188 10956 14240 11008
rect 18972 10956 19024 11008
rect 21180 10956 21232 11008
rect 21272 10999 21324 11008
rect 21272 10965 21281 10999
rect 21281 10965 21315 10999
rect 21315 10965 21324 10999
rect 21272 10956 21324 10965
rect 21640 10956 21692 11008
rect 22100 10956 22152 11008
rect 22652 10956 22704 11008
rect 24124 11092 24176 11144
rect 28172 11160 28224 11212
rect 30196 11160 30248 11212
rect 24676 11135 24728 11144
rect 24676 11101 24685 11135
rect 24685 11101 24719 11135
rect 24719 11101 24728 11135
rect 24676 11092 24728 11101
rect 26424 11135 26476 11144
rect 26424 11101 26433 11135
rect 26433 11101 26467 11135
rect 26467 11101 26476 11135
rect 26424 11092 26476 11101
rect 26608 11092 26660 11144
rect 26884 11135 26936 11144
rect 26884 11101 26896 11135
rect 26896 11101 26930 11135
rect 26930 11101 26936 11135
rect 26884 11092 26936 11101
rect 27528 11092 27580 11144
rect 28448 11092 28500 11144
rect 28080 11024 28132 11076
rect 30012 11067 30064 11076
rect 30012 11033 30021 11067
rect 30021 11033 30055 11067
rect 30055 11033 30064 11067
rect 30012 11024 30064 11033
rect 23848 10956 23900 11008
rect 30104 10956 30156 11008
rect 4193 10854 4245 10906
rect 4257 10854 4309 10906
rect 4321 10854 4373 10906
rect 4385 10854 4437 10906
rect 4449 10854 4501 10906
rect 11783 10854 11835 10906
rect 11847 10854 11899 10906
rect 11911 10854 11963 10906
rect 11975 10854 12027 10906
rect 12039 10854 12091 10906
rect 19373 10854 19425 10906
rect 19437 10854 19489 10906
rect 19501 10854 19553 10906
rect 19565 10854 19617 10906
rect 19629 10854 19681 10906
rect 26963 10854 27015 10906
rect 27027 10854 27079 10906
rect 27091 10854 27143 10906
rect 27155 10854 27207 10906
rect 27219 10854 27271 10906
rect 1308 10616 1360 10668
rect 5080 10752 5132 10804
rect 6092 10752 6144 10804
rect 7748 10752 7800 10804
rect 8852 10752 8904 10804
rect 11152 10752 11204 10804
rect 848 10548 900 10600
rect 3240 10591 3292 10600
rect 3240 10557 3249 10591
rect 3249 10557 3283 10591
rect 3283 10557 3292 10591
rect 3240 10548 3292 10557
rect 4436 10616 4488 10668
rect 1768 10412 1820 10464
rect 2044 10412 2096 10464
rect 4620 10548 4672 10600
rect 5540 10591 5592 10600
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 5540 10548 5592 10557
rect 5816 10548 5868 10600
rect 5908 10548 5960 10600
rect 6276 10591 6328 10600
rect 6276 10557 6285 10591
rect 6285 10557 6319 10591
rect 6319 10557 6328 10591
rect 6276 10548 6328 10557
rect 8668 10548 8720 10600
rect 13360 10684 13412 10736
rect 9404 10616 9456 10668
rect 9864 10616 9916 10668
rect 10048 10659 10100 10668
rect 10048 10625 10050 10659
rect 10050 10625 10100 10659
rect 10048 10616 10100 10625
rect 9312 10548 9364 10600
rect 11060 10616 11112 10668
rect 13820 10616 13872 10668
rect 14188 10616 14240 10668
rect 16764 10752 16816 10804
rect 16948 10752 17000 10804
rect 19248 10795 19300 10804
rect 19248 10761 19257 10795
rect 19257 10761 19291 10795
rect 19291 10761 19300 10795
rect 19248 10752 19300 10761
rect 21548 10752 21600 10804
rect 22284 10752 22336 10804
rect 26792 10752 26844 10804
rect 30564 10752 30616 10804
rect 16764 10616 16816 10668
rect 17500 10616 17552 10668
rect 21272 10684 21324 10736
rect 21916 10684 21968 10736
rect 19892 10616 19944 10668
rect 20720 10616 20772 10668
rect 21456 10616 21508 10668
rect 21732 10616 21784 10668
rect 7656 10523 7708 10532
rect 7656 10489 7665 10523
rect 7665 10489 7699 10523
rect 7699 10489 7708 10523
rect 7656 10480 7708 10489
rect 7840 10480 7892 10532
rect 10324 10548 10376 10600
rect 12164 10548 12216 10600
rect 12348 10548 12400 10600
rect 12624 10548 12676 10600
rect 12900 10548 12952 10600
rect 13452 10548 13504 10600
rect 13544 10591 13596 10600
rect 13544 10557 13553 10591
rect 13553 10557 13587 10591
rect 13587 10557 13596 10591
rect 13544 10548 13596 10557
rect 3976 10412 4028 10464
rect 4436 10412 4488 10464
rect 4712 10412 4764 10464
rect 6184 10412 6236 10464
rect 8760 10412 8812 10464
rect 9404 10455 9456 10464
rect 9404 10421 9413 10455
rect 9413 10421 9447 10455
rect 9447 10421 9456 10455
rect 9404 10412 9456 10421
rect 10416 10412 10468 10464
rect 12072 10455 12124 10464
rect 12072 10421 12081 10455
rect 12081 10421 12115 10455
rect 12115 10421 12124 10455
rect 12072 10412 12124 10421
rect 12440 10412 12492 10464
rect 12624 10455 12676 10464
rect 12624 10421 12633 10455
rect 12633 10421 12667 10455
rect 12667 10421 12676 10455
rect 12624 10412 12676 10421
rect 13084 10412 13136 10464
rect 16488 10548 16540 10600
rect 19156 10548 19208 10600
rect 18696 10480 18748 10532
rect 18788 10523 18840 10532
rect 18788 10489 18797 10523
rect 18797 10489 18831 10523
rect 18831 10489 18840 10523
rect 18788 10480 18840 10489
rect 13912 10412 13964 10464
rect 15292 10412 15344 10464
rect 16672 10412 16724 10464
rect 16856 10455 16908 10464
rect 16856 10421 16871 10455
rect 16871 10421 16905 10455
rect 16905 10421 16908 10455
rect 16856 10412 16908 10421
rect 17040 10412 17092 10464
rect 20260 10591 20312 10600
rect 20260 10557 20269 10591
rect 20269 10557 20303 10591
rect 20303 10557 20312 10591
rect 20260 10548 20312 10557
rect 21824 10548 21876 10600
rect 22928 10616 22980 10668
rect 23480 10659 23532 10668
rect 23480 10625 23489 10659
rect 23489 10625 23523 10659
rect 23523 10625 23532 10659
rect 23480 10616 23532 10625
rect 24952 10659 25004 10668
rect 20996 10480 21048 10532
rect 21548 10480 21600 10532
rect 19616 10412 19668 10464
rect 23020 10548 23072 10600
rect 23848 10480 23900 10532
rect 22100 10412 22152 10464
rect 24308 10548 24360 10600
rect 24952 10625 24954 10659
rect 24954 10625 25004 10659
rect 24952 10616 25004 10625
rect 27804 10616 27856 10668
rect 29184 10616 29236 10668
rect 29736 10616 29788 10668
rect 25688 10548 25740 10600
rect 25780 10548 25832 10600
rect 29460 10548 29512 10600
rect 29552 10548 29604 10600
rect 24124 10480 24176 10532
rect 24032 10455 24084 10464
rect 24032 10421 24041 10455
rect 24041 10421 24075 10455
rect 24075 10421 24084 10455
rect 24032 10412 24084 10421
rect 25136 10412 25188 10464
rect 25412 10412 25464 10464
rect 29000 10412 29052 10464
rect 29368 10412 29420 10464
rect 30104 10412 30156 10464
rect 30288 10455 30340 10464
rect 30288 10421 30297 10455
rect 30297 10421 30331 10455
rect 30331 10421 30340 10455
rect 30288 10412 30340 10421
rect 7988 10310 8040 10362
rect 8052 10310 8104 10362
rect 8116 10310 8168 10362
rect 8180 10310 8232 10362
rect 8244 10310 8296 10362
rect 15578 10310 15630 10362
rect 15642 10310 15694 10362
rect 15706 10310 15758 10362
rect 15770 10310 15822 10362
rect 15834 10310 15886 10362
rect 23168 10310 23220 10362
rect 23232 10310 23284 10362
rect 23296 10310 23348 10362
rect 23360 10310 23412 10362
rect 23424 10310 23476 10362
rect 30758 10310 30810 10362
rect 30822 10310 30874 10362
rect 30886 10310 30938 10362
rect 30950 10310 31002 10362
rect 31014 10310 31066 10362
rect 1768 10208 1820 10260
rect 3976 10208 4028 10260
rect 5540 10208 5592 10260
rect 6460 10208 6512 10260
rect 5816 10140 5868 10192
rect 6184 10183 6236 10192
rect 6184 10149 6193 10183
rect 6193 10149 6227 10183
rect 6227 10149 6236 10183
rect 6828 10208 6880 10260
rect 7840 10208 7892 10260
rect 6184 10140 6236 10149
rect 1308 10004 1360 10056
rect 1400 10004 1452 10056
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 4528 10072 4580 10124
rect 5632 10072 5684 10124
rect 6736 10072 6788 10124
rect 9496 10208 9548 10260
rect 12072 10208 12124 10260
rect 13360 10251 13412 10260
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 13452 10208 13504 10260
rect 15476 10208 15528 10260
rect 16212 10208 16264 10260
rect 17132 10208 17184 10260
rect 5724 9936 5776 9988
rect 7104 10004 7156 10056
rect 7196 10047 7248 10056
rect 7196 10013 7205 10047
rect 7205 10013 7239 10047
rect 7239 10013 7248 10047
rect 7196 10004 7248 10013
rect 7288 10004 7340 10056
rect 8484 10004 8536 10056
rect 9036 10047 9088 10056
rect 9036 10013 9038 10047
rect 9038 10013 9088 10047
rect 9036 10004 9088 10013
rect 9404 10115 9456 10124
rect 9404 10081 9413 10115
rect 9413 10081 9447 10115
rect 9447 10081 9456 10115
rect 9404 10072 9456 10081
rect 9680 10072 9732 10124
rect 10232 10072 10284 10124
rect 10600 10072 10652 10124
rect 12900 10072 12952 10124
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 15476 10072 15528 10124
rect 10784 10004 10836 10056
rect 11336 10047 11388 10056
rect 11336 10013 11338 10047
rect 11338 10013 11388 10047
rect 11336 10004 11388 10013
rect 11428 10047 11480 10056
rect 11428 10013 11440 10047
rect 11440 10013 11474 10047
rect 11474 10013 11480 10047
rect 11428 10004 11480 10013
rect 13912 10047 13964 10056
rect 13912 10013 13914 10047
rect 13914 10013 13964 10047
rect 13912 10004 13964 10013
rect 14004 10049 14056 10056
rect 14004 10015 14032 10049
rect 14032 10015 14056 10049
rect 14004 10004 14056 10015
rect 15936 10115 15988 10124
rect 15936 10081 15953 10115
rect 15953 10081 15987 10115
rect 15987 10081 15988 10115
rect 15936 10072 15988 10081
rect 8576 9936 8628 9988
rect 16396 10004 16448 10056
rect 16948 10072 17000 10124
rect 17040 10115 17092 10124
rect 17040 10081 17049 10115
rect 17049 10081 17083 10115
rect 17083 10081 17092 10115
rect 17040 10072 17092 10081
rect 18696 10140 18748 10192
rect 19064 10208 19116 10260
rect 20260 10208 20312 10260
rect 20996 10251 21048 10260
rect 20996 10217 21005 10251
rect 21005 10217 21039 10251
rect 21039 10217 21048 10251
rect 20996 10208 21048 10217
rect 19616 10183 19668 10192
rect 19616 10149 19625 10183
rect 19625 10149 19659 10183
rect 19659 10149 19668 10183
rect 19616 10140 19668 10149
rect 17776 10004 17828 10056
rect 19524 10072 19576 10124
rect 19708 10072 19760 10124
rect 20628 10140 20680 10192
rect 20260 10072 20312 10124
rect 18788 10004 18840 10056
rect 22652 10208 22704 10260
rect 22836 10208 22888 10260
rect 23572 10208 23624 10260
rect 24676 10208 24728 10260
rect 24952 10208 25004 10260
rect 22928 10140 22980 10192
rect 26332 10208 26384 10260
rect 21640 10115 21692 10124
rect 21640 10081 21642 10115
rect 21642 10081 21692 10115
rect 21640 10072 21692 10081
rect 22008 10115 22060 10124
rect 22008 10081 22017 10115
rect 22017 10081 22051 10115
rect 22051 10081 22060 10115
rect 22008 10072 22060 10081
rect 21456 10004 21508 10056
rect 21916 10004 21968 10056
rect 23480 10004 23532 10056
rect 26516 10140 26568 10192
rect 30288 10140 30340 10192
rect 24492 10115 24544 10124
rect 24492 10081 24494 10115
rect 24494 10081 24544 10115
rect 24492 10072 24544 10081
rect 25136 10072 25188 10124
rect 11152 9868 11204 9920
rect 12164 9868 12216 9920
rect 15384 9911 15436 9920
rect 15384 9877 15393 9911
rect 15393 9877 15427 9911
rect 15427 9877 15436 9911
rect 15384 9868 15436 9877
rect 16120 9911 16172 9920
rect 16120 9877 16129 9911
rect 16129 9877 16163 9911
rect 16163 9877 16172 9911
rect 16120 9868 16172 9877
rect 16948 9868 17000 9920
rect 18052 9868 18104 9920
rect 19524 9868 19576 9920
rect 19984 9868 20036 9920
rect 23572 9936 23624 9988
rect 23664 9868 23716 9920
rect 24860 10047 24912 10056
rect 24860 10013 24869 10047
rect 24869 10013 24903 10047
rect 24903 10013 24912 10047
rect 24860 10004 24912 10013
rect 24952 10004 25004 10056
rect 26424 10047 26476 10056
rect 26424 10013 26433 10047
rect 26433 10013 26467 10047
rect 26467 10013 26476 10047
rect 26424 10004 26476 10013
rect 26608 10004 26660 10056
rect 28172 10072 28224 10124
rect 28908 10115 28960 10124
rect 28908 10081 28917 10115
rect 28917 10081 28951 10115
rect 28951 10081 28960 10115
rect 28908 10072 28960 10081
rect 28264 10004 28316 10056
rect 24308 9868 24360 9920
rect 26056 9868 26108 9920
rect 28172 9868 28224 9920
rect 30380 9911 30432 9920
rect 30380 9877 30389 9911
rect 30389 9877 30423 9911
rect 30423 9877 30432 9911
rect 30380 9868 30432 9877
rect 4193 9766 4245 9818
rect 4257 9766 4309 9818
rect 4321 9766 4373 9818
rect 4385 9766 4437 9818
rect 4449 9766 4501 9818
rect 11783 9766 11835 9818
rect 11847 9766 11899 9818
rect 11911 9766 11963 9818
rect 11975 9766 12027 9818
rect 12039 9766 12091 9818
rect 19373 9766 19425 9818
rect 19437 9766 19489 9818
rect 19501 9766 19553 9818
rect 19565 9766 19617 9818
rect 19629 9766 19681 9818
rect 26963 9766 27015 9818
rect 27027 9766 27079 9818
rect 27091 9766 27143 9818
rect 27155 9766 27207 9818
rect 27219 9766 27271 9818
rect 1400 9664 1452 9716
rect 2044 9664 2096 9716
rect 2596 9664 2648 9716
rect 5724 9664 5776 9716
rect 6276 9664 6328 9716
rect 6460 9664 6512 9716
rect 8760 9664 8812 9716
rect 8852 9664 8904 9716
rect 10324 9664 10376 9716
rect 1308 9528 1360 9580
rect 1032 9460 1084 9512
rect 4712 9528 4764 9580
rect 3424 9460 3476 9512
rect 3976 9503 4028 9512
rect 3976 9469 3978 9503
rect 3978 9469 4028 9503
rect 3976 9460 4028 9469
rect 5172 9460 5224 9512
rect 6460 9528 6512 9580
rect 7012 9528 7064 9580
rect 8484 9528 8536 9580
rect 10508 9528 10560 9580
rect 6736 9460 6788 9512
rect 8392 9460 8444 9512
rect 9220 9460 9272 9512
rect 1768 9324 1820 9376
rect 1952 9324 2004 9376
rect 3424 9324 3476 9376
rect 5080 9392 5132 9444
rect 5908 9392 5960 9444
rect 7840 9392 7892 9444
rect 5356 9324 5408 9376
rect 6368 9324 6420 9376
rect 8944 9324 8996 9376
rect 9036 9367 9088 9376
rect 9036 9333 9051 9367
rect 9051 9333 9085 9367
rect 9085 9333 9088 9367
rect 9036 9324 9088 9333
rect 9588 9324 9640 9376
rect 12808 9664 12860 9716
rect 12992 9664 13044 9716
rect 13452 9664 13504 9716
rect 15476 9664 15528 9716
rect 17776 9664 17828 9716
rect 19156 9664 19208 9716
rect 23756 9664 23808 9716
rect 20536 9639 20588 9648
rect 20536 9605 20545 9639
rect 20545 9605 20579 9639
rect 20579 9605 20588 9639
rect 20536 9596 20588 9605
rect 22376 9596 22428 9648
rect 23112 9596 23164 9648
rect 25228 9664 25280 9716
rect 25688 9707 25740 9716
rect 25688 9673 25697 9707
rect 25697 9673 25731 9707
rect 25731 9673 25740 9707
rect 25688 9664 25740 9673
rect 28264 9707 28316 9716
rect 28264 9673 28273 9707
rect 28273 9673 28307 9707
rect 28307 9673 28316 9707
rect 28264 9664 28316 9673
rect 27528 9596 27580 9648
rect 10784 9503 10836 9512
rect 10784 9469 10793 9503
rect 10793 9469 10827 9503
rect 10827 9469 10836 9503
rect 10784 9460 10836 9469
rect 11060 9528 11112 9580
rect 11244 9571 11296 9580
rect 11244 9537 11256 9571
rect 11256 9537 11290 9571
rect 11290 9537 11296 9571
rect 11244 9528 11296 9537
rect 11428 9528 11480 9580
rect 11520 9503 11572 9512
rect 11520 9469 11529 9503
rect 11529 9469 11563 9503
rect 11563 9469 11572 9503
rect 11520 9460 11572 9469
rect 13176 9528 13228 9580
rect 13268 9528 13320 9580
rect 13544 9571 13596 9580
rect 13544 9537 13553 9571
rect 13553 9537 13587 9571
rect 13587 9537 13596 9571
rect 13544 9528 13596 9537
rect 14096 9528 14148 9580
rect 14648 9528 14700 9580
rect 16764 9460 16816 9512
rect 17132 9503 17184 9512
rect 17132 9469 17141 9503
rect 17141 9469 17175 9503
rect 17175 9469 17184 9503
rect 17132 9460 17184 9469
rect 21180 9528 21232 9580
rect 21640 9571 21692 9580
rect 21640 9537 21649 9571
rect 21649 9537 21683 9571
rect 21683 9537 21692 9571
rect 21640 9528 21692 9537
rect 23848 9571 23900 9580
rect 23848 9537 23857 9571
rect 23857 9537 23891 9571
rect 23891 9537 23900 9571
rect 23848 9528 23900 9537
rect 24032 9528 24084 9580
rect 25320 9528 25372 9580
rect 18696 9503 18748 9512
rect 18696 9469 18705 9503
rect 18705 9469 18739 9503
rect 18739 9469 18748 9503
rect 18696 9460 18748 9469
rect 19340 9460 19392 9512
rect 19432 9503 19484 9512
rect 19432 9469 19441 9503
rect 19441 9469 19475 9503
rect 19475 9469 19484 9503
rect 19432 9460 19484 9469
rect 19892 9460 19944 9512
rect 11152 9324 11204 9376
rect 11336 9324 11388 9376
rect 12624 9367 12676 9376
rect 12624 9333 12633 9367
rect 12633 9333 12667 9367
rect 12667 9333 12676 9367
rect 12624 9324 12676 9333
rect 13176 9392 13228 9444
rect 13360 9392 13412 9444
rect 15936 9392 15988 9444
rect 13912 9324 13964 9376
rect 18604 9392 18656 9444
rect 17224 9324 17276 9376
rect 19064 9324 19116 9376
rect 19340 9324 19392 9376
rect 22560 9460 22612 9512
rect 22376 9392 22428 9444
rect 23480 9460 23532 9512
rect 24492 9460 24544 9512
rect 25688 9460 25740 9512
rect 26976 9528 27028 9580
rect 26056 9503 26108 9512
rect 26056 9469 26065 9503
rect 26065 9469 26099 9503
rect 26099 9469 26108 9503
rect 26056 9460 26108 9469
rect 26424 9460 26476 9512
rect 28908 9528 28960 9580
rect 29460 9664 29512 9716
rect 30288 9664 30340 9716
rect 30656 9596 30708 9648
rect 29092 9528 29144 9580
rect 27528 9392 27580 9444
rect 21364 9367 21416 9376
rect 21364 9333 21379 9367
rect 21379 9333 21413 9367
rect 21413 9333 21416 9367
rect 21364 9324 21416 9333
rect 23756 9324 23808 9376
rect 24492 9324 24544 9376
rect 25780 9324 25832 9376
rect 25872 9324 25924 9376
rect 26516 9367 26568 9376
rect 26516 9333 26531 9367
rect 26531 9333 26565 9367
rect 26565 9333 26568 9367
rect 26516 9324 26568 9333
rect 27896 9367 27948 9376
rect 27896 9333 27905 9367
rect 27905 9333 27939 9367
rect 27939 9333 27948 9367
rect 27896 9324 27948 9333
rect 29000 9367 29052 9376
rect 29000 9333 29009 9367
rect 29009 9333 29043 9367
rect 29043 9333 29052 9367
rect 29000 9324 29052 9333
rect 29368 9324 29420 9376
rect 30104 9324 30156 9376
rect 30288 9367 30340 9376
rect 30288 9333 30297 9367
rect 30297 9333 30331 9367
rect 30331 9333 30340 9367
rect 30288 9324 30340 9333
rect 7988 9222 8040 9274
rect 8052 9222 8104 9274
rect 8116 9222 8168 9274
rect 8180 9222 8232 9274
rect 8244 9222 8296 9274
rect 15578 9222 15630 9274
rect 15642 9222 15694 9274
rect 15706 9222 15758 9274
rect 15770 9222 15822 9274
rect 15834 9222 15886 9274
rect 23168 9222 23220 9274
rect 23232 9222 23284 9274
rect 23296 9222 23348 9274
rect 23360 9222 23412 9274
rect 23424 9222 23476 9274
rect 30758 9222 30810 9274
rect 30822 9222 30874 9274
rect 30886 9222 30938 9274
rect 30950 9222 31002 9274
rect 31014 9222 31066 9274
rect 1308 9163 1360 9172
rect 1308 9129 1317 9163
rect 1317 9129 1351 9163
rect 1351 9129 1360 9163
rect 1308 9120 1360 9129
rect 2872 9163 2924 9172
rect 2872 9129 2887 9163
rect 2887 9129 2921 9163
rect 2921 9129 2924 9163
rect 2872 9120 2924 9129
rect 4620 9163 4672 9172
rect 4620 9129 4629 9163
rect 4629 9129 4663 9163
rect 4663 9129 4672 9163
rect 4620 9120 4672 9129
rect 1952 9052 2004 9104
rect 7196 9120 7248 9172
rect 7564 9120 7616 9172
rect 7656 9120 7708 9172
rect 7840 9120 7892 9172
rect 9220 9120 9272 9172
rect 11520 9120 11572 9172
rect 1768 8984 1820 9036
rect 2412 9027 2464 9036
rect 2412 8993 2421 9027
rect 2421 8993 2455 9027
rect 2455 8993 2464 9027
rect 2412 8984 2464 8993
rect 2964 8916 3016 8968
rect 3332 8916 3384 8968
rect 1768 8848 1820 8900
rect 1952 8848 2004 8900
rect 1676 8780 1728 8832
rect 5080 8848 5132 8900
rect 4804 8780 4856 8832
rect 4896 8823 4948 8832
rect 4896 8789 4905 8823
rect 4905 8789 4939 8823
rect 4939 8789 4948 8823
rect 4896 8780 4948 8789
rect 4988 8780 5040 8832
rect 5356 8848 5408 8900
rect 5448 8891 5500 8900
rect 5448 8857 5457 8891
rect 5457 8857 5491 8891
rect 5491 8857 5500 8891
rect 5448 8848 5500 8857
rect 6092 8984 6144 9036
rect 6368 9027 6420 9036
rect 6368 8993 6377 9027
rect 6377 8993 6411 9027
rect 6411 8993 6420 9027
rect 6368 8984 6420 8993
rect 6644 9027 6696 9036
rect 6644 8993 6653 9027
rect 6653 8993 6687 9027
rect 6687 8993 6696 9027
rect 6644 8984 6696 8993
rect 7196 9027 7248 9036
rect 7196 8993 7205 9027
rect 7205 8993 7239 9027
rect 7239 8993 7248 9027
rect 7196 8984 7248 8993
rect 7472 9027 7524 9036
rect 7472 8993 7481 9027
rect 7481 8993 7515 9027
rect 7515 8993 7524 9027
rect 7472 8984 7524 8993
rect 6276 8848 6328 8900
rect 7012 8916 7064 8968
rect 13912 9120 13964 9172
rect 15660 9120 15712 9172
rect 16120 9120 16172 9172
rect 17132 9120 17184 9172
rect 17224 9120 17276 9172
rect 17868 9120 17920 9172
rect 19432 9120 19484 9172
rect 20444 9120 20496 9172
rect 21640 9120 21692 9172
rect 22008 9120 22060 9172
rect 23572 9120 23624 9172
rect 23664 9120 23716 9172
rect 19156 9052 19208 9104
rect 21364 9052 21416 9104
rect 8208 8984 8260 9036
rect 10508 9027 10560 9036
rect 10508 8993 10517 9027
rect 10517 8993 10551 9027
rect 10551 8993 10560 9027
rect 10508 8984 10560 8993
rect 11336 9027 11388 9036
rect 11336 8993 11338 9027
rect 11338 8993 11388 9027
rect 11336 8984 11388 8993
rect 11612 8984 11664 9036
rect 12348 8984 12400 9036
rect 12716 8984 12768 9036
rect 13544 9027 13596 9036
rect 13544 8993 13553 9027
rect 13553 8993 13587 9027
rect 13587 8993 13596 9027
rect 13544 8984 13596 8993
rect 14924 8984 14976 9036
rect 15476 8984 15528 9036
rect 16120 8984 16172 9036
rect 16488 8984 16540 9036
rect 16672 8984 16724 9036
rect 16948 8984 17000 9036
rect 18788 8984 18840 9036
rect 8300 8959 8352 8968
rect 8300 8925 8309 8959
rect 8309 8925 8343 8959
rect 8343 8925 8352 8959
rect 8300 8916 8352 8925
rect 8484 8916 8536 8968
rect 5816 8823 5868 8832
rect 5816 8789 5825 8823
rect 5825 8789 5859 8823
rect 5859 8789 5868 8823
rect 5816 8780 5868 8789
rect 6368 8780 6420 8832
rect 6460 8823 6512 8832
rect 6460 8789 6469 8823
rect 6469 8789 6503 8823
rect 6503 8789 6512 8823
rect 6460 8780 6512 8789
rect 7012 8823 7064 8832
rect 7012 8789 7021 8823
rect 7021 8789 7055 8823
rect 7055 8789 7064 8823
rect 7012 8780 7064 8789
rect 9404 8848 9456 8900
rect 8484 8780 8536 8832
rect 8668 8780 8720 8832
rect 10876 8916 10928 8968
rect 11152 8916 11204 8968
rect 11520 8916 11572 8968
rect 12808 8916 12860 8968
rect 13084 8916 13136 8968
rect 15200 8916 15252 8968
rect 17132 8916 17184 8968
rect 10600 8891 10652 8900
rect 10600 8857 10609 8891
rect 10609 8857 10643 8891
rect 10643 8857 10652 8891
rect 10600 8848 10652 8857
rect 15476 8848 15528 8900
rect 11336 8780 11388 8832
rect 12348 8780 12400 8832
rect 15568 8823 15620 8832
rect 15568 8789 15577 8823
rect 15577 8789 15611 8823
rect 15611 8789 15620 8823
rect 15568 8780 15620 8789
rect 16488 8780 16540 8832
rect 19248 8780 19300 8832
rect 19984 8984 20036 9036
rect 20536 8984 20588 9036
rect 22008 8984 22060 9036
rect 22284 8984 22336 9036
rect 20628 8916 20680 8968
rect 19708 8848 19760 8900
rect 20352 8848 20404 8900
rect 21916 8848 21968 8900
rect 22560 8984 22612 9036
rect 23756 8984 23808 9036
rect 24860 9120 24912 9172
rect 24952 9163 25004 9172
rect 24952 9129 24961 9163
rect 24961 9129 24995 9163
rect 24995 9129 25004 9163
rect 24952 9120 25004 9129
rect 25688 9163 25740 9172
rect 25688 9129 25697 9163
rect 25697 9129 25731 9163
rect 25731 9129 25740 9163
rect 25688 9120 25740 9129
rect 23572 8916 23624 8968
rect 22652 8891 22704 8900
rect 22652 8857 22661 8891
rect 22661 8857 22695 8891
rect 22695 8857 22704 8891
rect 22652 8848 22704 8857
rect 25596 9027 25648 9036
rect 25596 8993 25605 9027
rect 25605 8993 25639 9027
rect 25639 8993 25648 9027
rect 25596 8984 25648 8993
rect 25780 8984 25832 9036
rect 27528 9120 27580 9172
rect 27896 9120 27948 9172
rect 26148 9027 26200 9036
rect 26148 8993 26157 9027
rect 26157 8993 26191 9027
rect 26191 8993 26200 9027
rect 26148 8984 26200 8993
rect 26332 8984 26384 9036
rect 25504 8916 25556 8968
rect 26608 8916 26660 8968
rect 29000 9120 29052 9172
rect 29276 9120 29328 9172
rect 30472 9120 30524 9172
rect 29828 9052 29880 9104
rect 30196 9052 30248 9104
rect 28632 9027 28684 9036
rect 28632 8993 28641 9027
rect 28641 8993 28675 9027
rect 28675 8993 28684 9027
rect 28632 8984 28684 8993
rect 30012 8984 30064 9036
rect 29368 8916 29420 8968
rect 29552 8916 29604 8968
rect 20812 8780 20864 8832
rect 22192 8780 22244 8832
rect 25412 8823 25464 8832
rect 25412 8789 25421 8823
rect 25421 8789 25455 8823
rect 25455 8789 25464 8823
rect 25412 8780 25464 8789
rect 26884 8780 26936 8832
rect 28264 8823 28316 8832
rect 28264 8789 28273 8823
rect 28273 8789 28307 8823
rect 28307 8789 28316 8823
rect 28264 8780 28316 8789
rect 28908 8780 28960 8832
rect 29368 8780 29420 8832
rect 30012 8780 30064 8832
rect 30472 8780 30524 8832
rect 4193 8678 4245 8730
rect 4257 8678 4309 8730
rect 4321 8678 4373 8730
rect 4385 8678 4437 8730
rect 4449 8678 4501 8730
rect 11783 8678 11835 8730
rect 11847 8678 11899 8730
rect 11911 8678 11963 8730
rect 11975 8678 12027 8730
rect 12039 8678 12091 8730
rect 19373 8678 19425 8730
rect 19437 8678 19489 8730
rect 19501 8678 19553 8730
rect 19565 8678 19617 8730
rect 19629 8678 19681 8730
rect 26963 8678 27015 8730
rect 27027 8678 27079 8730
rect 27091 8678 27143 8730
rect 27155 8678 27207 8730
rect 27219 8678 27271 8730
rect 940 8576 992 8628
rect 2780 8619 2832 8628
rect 2780 8585 2789 8619
rect 2789 8585 2823 8619
rect 2823 8585 2832 8619
rect 2780 8576 2832 8585
rect 2412 8508 2464 8560
rect 3240 8508 3292 8560
rect 4712 8508 4764 8560
rect 756 8372 808 8424
rect 1584 8372 1636 8424
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 2964 8440 3016 8492
rect 3056 8440 3108 8492
rect 2688 8304 2740 8356
rect 3240 8415 3292 8424
rect 3240 8381 3249 8415
rect 3249 8381 3283 8415
rect 3283 8381 3292 8415
rect 3240 8372 3292 8381
rect 3608 8415 3660 8424
rect 3608 8381 3610 8415
rect 3610 8381 3660 8415
rect 3608 8372 3660 8381
rect 7104 8576 7156 8628
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 5816 8440 5868 8492
rect 5908 8440 5960 8492
rect 6736 8440 6788 8492
rect 8300 8576 8352 8628
rect 8392 8619 8444 8628
rect 8392 8585 8401 8619
rect 8401 8585 8435 8619
rect 8435 8585 8444 8619
rect 8392 8576 8444 8585
rect 8484 8576 8536 8628
rect 9128 8576 9180 8628
rect 6000 8279 6052 8288
rect 6000 8245 6015 8279
rect 6015 8245 6049 8279
rect 6049 8245 6052 8279
rect 6000 8236 6052 8245
rect 7840 8236 7892 8288
rect 8760 8508 8812 8560
rect 9312 8508 9364 8560
rect 8484 8440 8536 8492
rect 8668 8440 8720 8492
rect 9128 8440 9180 8492
rect 10968 8440 11020 8492
rect 11520 8619 11572 8628
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 11152 8508 11204 8560
rect 12532 8508 12584 8560
rect 13084 8551 13136 8560
rect 13084 8517 13093 8551
rect 13093 8517 13127 8551
rect 13127 8517 13136 8551
rect 13084 8508 13136 8517
rect 15108 8508 15160 8560
rect 15200 8508 15252 8560
rect 9220 8372 9272 8424
rect 9496 8415 9548 8424
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 9588 8372 9640 8424
rect 11336 8372 11388 8424
rect 11704 8372 11756 8424
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 13912 8483 13964 8492
rect 13912 8449 13914 8483
rect 13914 8449 13964 8483
rect 13912 8440 13964 8449
rect 16028 8576 16080 8628
rect 16672 8576 16724 8628
rect 15568 8508 15620 8560
rect 17592 8619 17644 8628
rect 17592 8585 17601 8619
rect 17601 8585 17635 8619
rect 17635 8585 17644 8619
rect 17592 8576 17644 8585
rect 18604 8576 18656 8628
rect 17960 8508 18012 8560
rect 17132 8440 17184 8492
rect 18696 8483 18748 8492
rect 9036 8236 9088 8288
rect 9128 8279 9180 8288
rect 9128 8245 9137 8279
rect 9137 8245 9171 8279
rect 9171 8245 9180 8279
rect 9128 8236 9180 8245
rect 11612 8236 11664 8288
rect 12072 8236 12124 8288
rect 14188 8372 14240 8424
rect 15660 8372 15712 8424
rect 17592 8372 17644 8424
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 19064 8483 19116 8492
rect 19064 8449 19066 8483
rect 19066 8449 19116 8483
rect 19064 8440 19116 8449
rect 19156 8483 19208 8492
rect 19156 8449 19168 8483
rect 19168 8449 19202 8483
rect 19202 8449 19208 8483
rect 19156 8440 19208 8449
rect 19340 8440 19392 8492
rect 20720 8619 20772 8628
rect 20720 8585 20729 8619
rect 20729 8585 20763 8619
rect 20763 8585 20772 8619
rect 20720 8576 20772 8585
rect 22284 8576 22336 8628
rect 25596 8576 25648 8628
rect 25872 8619 25924 8628
rect 25872 8585 25881 8619
rect 25881 8585 25915 8619
rect 25915 8585 25924 8619
rect 25872 8576 25924 8585
rect 26424 8576 26476 8628
rect 25412 8508 25464 8560
rect 20720 8440 20772 8492
rect 22008 8440 22060 8492
rect 22192 8440 22244 8492
rect 18420 8415 18472 8424
rect 18420 8381 18429 8415
rect 18429 8381 18463 8415
rect 18463 8381 18472 8415
rect 18420 8372 18472 8381
rect 21456 8372 21508 8424
rect 21916 8372 21968 8424
rect 22928 8372 22980 8424
rect 23756 8372 23808 8424
rect 23848 8415 23900 8424
rect 23848 8381 23857 8415
rect 23857 8381 23891 8415
rect 23891 8381 23900 8415
rect 23848 8372 23900 8381
rect 27804 8576 27856 8628
rect 28540 8619 28592 8628
rect 28540 8585 28549 8619
rect 28549 8585 28583 8619
rect 28583 8585 28592 8619
rect 28540 8576 28592 8585
rect 29184 8576 29236 8628
rect 28632 8508 28684 8560
rect 26516 8372 26568 8424
rect 28080 8440 28132 8492
rect 27344 8372 27396 8424
rect 30380 8440 30432 8492
rect 13636 8236 13688 8288
rect 14556 8236 14608 8288
rect 26792 8304 26844 8356
rect 28816 8304 28868 8356
rect 30196 8372 30248 8424
rect 31208 8304 31260 8356
rect 16028 8236 16080 8288
rect 19064 8236 19116 8288
rect 21640 8236 21692 8288
rect 21916 8236 21968 8288
rect 22560 8236 22612 8288
rect 25044 8236 25096 8288
rect 28080 8236 28132 8288
rect 29184 8279 29236 8288
rect 29184 8245 29193 8279
rect 29193 8245 29227 8279
rect 29227 8245 29236 8279
rect 29184 8236 29236 8245
rect 7988 8134 8040 8186
rect 8052 8134 8104 8186
rect 8116 8134 8168 8186
rect 8180 8134 8232 8186
rect 8244 8134 8296 8186
rect 15578 8134 15630 8186
rect 15642 8134 15694 8186
rect 15706 8134 15758 8186
rect 15770 8134 15822 8186
rect 15834 8134 15886 8186
rect 23168 8134 23220 8186
rect 23232 8134 23284 8186
rect 23296 8134 23348 8186
rect 23360 8134 23412 8186
rect 23424 8134 23476 8186
rect 30758 8134 30810 8186
rect 30822 8134 30874 8186
rect 30886 8134 30938 8186
rect 30950 8134 31002 8186
rect 31014 8134 31066 8186
rect 2228 8032 2280 8084
rect 1584 7896 1636 7948
rect 1768 7896 1820 7948
rect 1492 7828 1544 7880
rect 2044 7964 2096 8016
rect 5172 8075 5224 8084
rect 5172 8041 5181 8075
rect 5181 8041 5215 8075
rect 5215 8041 5224 8075
rect 5172 8032 5224 8041
rect 5724 8032 5776 8084
rect 6644 8032 6696 8084
rect 7656 8075 7708 8084
rect 7656 8041 7665 8075
rect 7665 8041 7699 8075
rect 7699 8041 7708 8075
rect 7656 8032 7708 8041
rect 1308 7760 1360 7812
rect 3240 7896 3292 7948
rect 5172 7896 5224 7948
rect 5816 7964 5868 8016
rect 1124 7692 1176 7744
rect 5540 7828 5592 7880
rect 5264 7760 5316 7812
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 6000 7828 6052 7880
rect 9680 8032 9732 8084
rect 11336 8032 11388 8084
rect 10324 7964 10376 8016
rect 7840 7760 7892 7812
rect 8392 7896 8444 7948
rect 9128 7896 9180 7948
rect 9312 7896 9364 7948
rect 8576 7828 8628 7880
rect 10600 7828 10652 7880
rect 11244 7896 11296 7948
rect 14832 8032 14884 8084
rect 16028 8032 16080 8084
rect 16672 8032 16724 8084
rect 11152 7828 11204 7880
rect 11336 7871 11388 7880
rect 11336 7837 11345 7871
rect 11345 7837 11379 7871
rect 11379 7837 11388 7871
rect 11336 7828 11388 7837
rect 11704 7871 11756 7880
rect 11704 7837 11706 7871
rect 11706 7837 11756 7871
rect 11704 7828 11756 7837
rect 11796 7871 11848 7880
rect 11796 7837 11841 7871
rect 11841 7837 11848 7871
rect 13728 7939 13780 7948
rect 13728 7905 13737 7939
rect 13737 7905 13771 7939
rect 13771 7905 13780 7939
rect 13728 7896 13780 7905
rect 16212 8007 16264 8016
rect 16212 7973 16221 8007
rect 16221 7973 16255 8007
rect 16255 7973 16264 8007
rect 16212 7964 16264 7973
rect 16304 7964 16356 8016
rect 17592 8075 17644 8084
rect 17592 8041 17601 8075
rect 17601 8041 17635 8075
rect 17635 8041 17644 8075
rect 17592 8032 17644 8041
rect 19064 8032 19116 8084
rect 19892 8075 19944 8084
rect 19892 8041 19901 8075
rect 19901 8041 19935 8075
rect 19935 8041 19944 8075
rect 19892 8032 19944 8041
rect 21916 8032 21968 8084
rect 16396 7896 16448 7948
rect 11796 7828 11848 7837
rect 8300 7760 8352 7812
rect 15384 7828 15436 7880
rect 3240 7692 3292 7744
rect 4068 7692 4120 7744
rect 6000 7692 6052 7744
rect 7564 7692 7616 7744
rect 8944 7692 8996 7744
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 10692 7735 10744 7744
rect 10692 7701 10701 7735
rect 10701 7701 10735 7735
rect 10735 7701 10744 7735
rect 10692 7692 10744 7701
rect 10784 7692 10836 7744
rect 13176 7735 13228 7744
rect 13176 7701 13185 7735
rect 13185 7701 13219 7735
rect 13219 7701 13228 7735
rect 13176 7692 13228 7701
rect 13820 7692 13872 7744
rect 14556 7692 14608 7744
rect 14740 7692 14792 7744
rect 18144 7896 18196 7948
rect 20536 7939 20588 7948
rect 20536 7905 20545 7939
rect 20545 7905 20579 7939
rect 20579 7905 20588 7939
rect 20536 7896 20588 7905
rect 20628 7896 20680 7948
rect 21272 7964 21324 8016
rect 18420 7828 18472 7880
rect 18880 7828 18932 7880
rect 23020 8032 23072 8084
rect 25320 8075 25372 8084
rect 25320 8041 25329 8075
rect 25329 8041 25363 8075
rect 25363 8041 25372 8075
rect 25320 8032 25372 8041
rect 27804 8032 27856 8084
rect 28356 8032 28408 8084
rect 25044 7964 25096 8016
rect 29368 7964 29420 8016
rect 24492 7896 24544 7948
rect 26424 7896 26476 7948
rect 27528 7896 27580 7948
rect 28080 7896 28132 7948
rect 28448 7939 28500 7948
rect 28448 7905 28457 7939
rect 28457 7905 28491 7939
rect 28491 7905 28500 7939
rect 28448 7896 28500 7905
rect 29552 7896 29604 7948
rect 29920 7896 29972 7948
rect 21456 7828 21508 7880
rect 21640 7871 21692 7880
rect 21640 7837 21642 7871
rect 21642 7837 21692 7871
rect 21640 7828 21692 7837
rect 15660 7735 15712 7744
rect 15660 7701 15669 7735
rect 15669 7701 15703 7735
rect 15703 7701 15712 7735
rect 15660 7692 15712 7701
rect 15752 7692 15804 7744
rect 16764 7692 16816 7744
rect 17500 7692 17552 7744
rect 20444 7692 20496 7744
rect 22192 7692 22244 7744
rect 22928 7828 22980 7880
rect 23664 7828 23716 7880
rect 24124 7828 24176 7880
rect 26608 7828 26660 7880
rect 27252 7828 27304 7880
rect 27712 7871 27764 7880
rect 27712 7837 27721 7871
rect 27721 7837 27755 7871
rect 27755 7837 27764 7871
rect 27712 7828 27764 7837
rect 28172 7871 28224 7880
rect 28172 7837 28184 7871
rect 28184 7837 28218 7871
rect 28218 7837 28224 7871
rect 28172 7828 28224 7837
rect 25228 7692 25280 7744
rect 27436 7735 27488 7744
rect 27436 7701 27445 7735
rect 27445 7701 27479 7735
rect 27479 7701 27488 7735
rect 27436 7692 27488 7701
rect 28816 7692 28868 7744
rect 30380 7735 30432 7744
rect 30380 7701 30389 7735
rect 30389 7701 30423 7735
rect 30423 7701 30432 7735
rect 30380 7692 30432 7701
rect 4193 7590 4245 7642
rect 4257 7590 4309 7642
rect 4321 7590 4373 7642
rect 4385 7590 4437 7642
rect 4449 7590 4501 7642
rect 11783 7590 11835 7642
rect 11847 7590 11899 7642
rect 11911 7590 11963 7642
rect 11975 7590 12027 7642
rect 12039 7590 12091 7642
rect 19373 7590 19425 7642
rect 19437 7590 19489 7642
rect 19501 7590 19553 7642
rect 19565 7590 19617 7642
rect 19629 7590 19681 7642
rect 26963 7590 27015 7642
rect 27027 7590 27079 7642
rect 27091 7590 27143 7642
rect 27155 7590 27207 7642
rect 27219 7590 27271 7642
rect 1124 7352 1176 7404
rect 756 7284 808 7336
rect 7656 7488 7708 7540
rect 7564 7420 7616 7472
rect 2044 7284 2096 7336
rect 3240 7327 3292 7336
rect 3240 7293 3249 7327
rect 3249 7293 3283 7327
rect 3283 7293 3292 7327
rect 3240 7284 3292 7293
rect 3332 7284 3384 7336
rect 3056 7259 3108 7268
rect 3056 7225 3065 7259
rect 3065 7225 3099 7259
rect 3099 7225 3108 7259
rect 3056 7216 3108 7225
rect 5264 7352 5316 7404
rect 5448 7352 5500 7404
rect 5908 7395 5960 7404
rect 5908 7361 5910 7395
rect 5910 7361 5960 7395
rect 5908 7352 5960 7361
rect 6736 7352 6788 7404
rect 8576 7352 8628 7404
rect 5080 7284 5132 7336
rect 7840 7284 7892 7336
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 8392 7284 8444 7293
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 13176 7488 13228 7540
rect 11244 7420 11296 7472
rect 12624 7352 12676 7404
rect 1492 7148 1544 7200
rect 1768 7148 1820 7200
rect 4436 7148 4488 7200
rect 4620 7148 4672 7200
rect 10968 7284 11020 7336
rect 11244 7327 11296 7336
rect 11244 7293 11253 7327
rect 11253 7293 11287 7327
rect 11287 7293 11296 7327
rect 11244 7284 11296 7293
rect 12440 7284 12492 7336
rect 13176 7352 13228 7404
rect 15752 7488 15804 7540
rect 16212 7531 16264 7540
rect 16212 7497 16221 7531
rect 16221 7497 16255 7531
rect 16255 7497 16264 7531
rect 16212 7488 16264 7497
rect 17776 7531 17828 7540
rect 17776 7497 17785 7531
rect 17785 7497 17819 7531
rect 17819 7497 17828 7531
rect 17776 7488 17828 7497
rect 18880 7488 18932 7540
rect 19892 7488 19944 7540
rect 20812 7488 20864 7540
rect 23572 7531 23624 7540
rect 23572 7497 23581 7531
rect 23581 7497 23615 7531
rect 23615 7497 23624 7531
rect 23572 7488 23624 7497
rect 24124 7488 24176 7540
rect 27528 7488 27580 7540
rect 12992 7284 13044 7336
rect 13268 7284 13320 7336
rect 14464 7284 14516 7336
rect 15292 7352 15344 7404
rect 15568 7352 15620 7404
rect 16580 7284 16632 7336
rect 16764 7284 16816 7336
rect 17132 7327 17184 7336
rect 17132 7293 17141 7327
rect 17141 7293 17175 7327
rect 17175 7293 17184 7327
rect 17132 7284 17184 7293
rect 17500 7284 17552 7336
rect 18512 7352 18564 7404
rect 19064 7395 19116 7404
rect 19064 7361 19066 7395
rect 19066 7361 19116 7395
rect 19064 7352 19116 7361
rect 21732 7352 21784 7404
rect 21916 7395 21968 7404
rect 21916 7361 21918 7395
rect 21918 7361 21968 7395
rect 21916 7352 21968 7361
rect 22008 7377 22060 7404
rect 22008 7352 22020 7377
rect 22020 7352 22054 7377
rect 22054 7352 22060 7377
rect 22192 7352 22244 7404
rect 22652 7352 22704 7404
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 24400 7352 24452 7404
rect 7656 7148 7708 7200
rect 10508 7148 10560 7200
rect 11704 7191 11756 7200
rect 11704 7157 11719 7191
rect 11719 7157 11753 7191
rect 11753 7157 11756 7191
rect 18420 7284 18472 7336
rect 11704 7148 11756 7157
rect 13084 7191 13136 7200
rect 13084 7157 13093 7191
rect 13093 7157 13127 7191
rect 13127 7157 13136 7191
rect 13084 7148 13136 7157
rect 14188 7148 14240 7200
rect 14832 7191 14884 7200
rect 14832 7157 14847 7191
rect 14847 7157 14881 7191
rect 14881 7157 14884 7191
rect 14832 7148 14884 7157
rect 15016 7148 15068 7200
rect 16764 7191 16816 7200
rect 16764 7157 16773 7191
rect 16773 7157 16807 7191
rect 16807 7157 16816 7191
rect 16764 7148 16816 7157
rect 18604 7216 18656 7268
rect 17592 7191 17644 7200
rect 17592 7157 17601 7191
rect 17601 7157 17635 7191
rect 17635 7157 17644 7191
rect 17592 7148 17644 7157
rect 17776 7148 17828 7200
rect 20444 7284 20496 7336
rect 20904 7284 20956 7336
rect 21548 7327 21600 7336
rect 21548 7293 21557 7327
rect 21557 7293 21591 7327
rect 21591 7293 21600 7327
rect 21548 7284 21600 7293
rect 22376 7148 22428 7200
rect 22560 7148 22612 7200
rect 24860 7327 24912 7336
rect 24860 7293 24869 7327
rect 24869 7293 24903 7327
rect 24903 7293 24912 7327
rect 24860 7284 24912 7293
rect 24492 7148 24544 7200
rect 24768 7148 24820 7200
rect 26148 7284 26200 7336
rect 25688 7216 25740 7268
rect 29276 7284 29328 7336
rect 29460 7327 29512 7336
rect 29460 7293 29469 7327
rect 29469 7293 29503 7327
rect 29503 7293 29512 7327
rect 29460 7284 29512 7293
rect 26608 7148 26660 7200
rect 26976 7148 27028 7200
rect 28540 7191 28592 7200
rect 28540 7157 28549 7191
rect 28549 7157 28583 7191
rect 28583 7157 28592 7191
rect 28540 7148 28592 7157
rect 28632 7148 28684 7200
rect 29736 7148 29788 7200
rect 7988 7046 8040 7098
rect 8052 7046 8104 7098
rect 8116 7046 8168 7098
rect 8180 7046 8232 7098
rect 8244 7046 8296 7098
rect 15578 7046 15630 7098
rect 15642 7046 15694 7098
rect 15706 7046 15758 7098
rect 15770 7046 15822 7098
rect 15834 7046 15886 7098
rect 23168 7046 23220 7098
rect 23232 7046 23284 7098
rect 23296 7046 23348 7098
rect 23360 7046 23412 7098
rect 23424 7046 23476 7098
rect 30758 7046 30810 7098
rect 30822 7046 30874 7098
rect 30886 7046 30938 7098
rect 30950 7046 31002 7098
rect 31014 7046 31066 7098
rect 756 6876 808 6928
rect 940 6647 992 6656
rect 940 6613 949 6647
rect 949 6613 983 6647
rect 983 6613 992 6647
rect 940 6604 992 6613
rect 1216 6647 1268 6656
rect 1216 6613 1225 6647
rect 1225 6613 1259 6647
rect 1259 6613 1268 6647
rect 1216 6604 1268 6613
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 3240 6944 3292 6996
rect 3424 6944 3476 6996
rect 5080 6944 5132 6996
rect 5448 6944 5500 6996
rect 5816 6944 5868 6996
rect 1768 6919 1820 6928
rect 1768 6885 1777 6919
rect 1777 6885 1811 6919
rect 1811 6885 1820 6919
rect 1768 6876 1820 6885
rect 2044 6876 2096 6928
rect 3608 6876 3660 6928
rect 3976 6876 4028 6928
rect 4620 6876 4672 6928
rect 1676 6740 1728 6792
rect 3240 6740 3292 6792
rect 4344 6808 4396 6860
rect 5080 6851 5132 6860
rect 3884 6740 3936 6792
rect 5080 6817 5089 6851
rect 5089 6817 5123 6851
rect 5123 6817 5132 6851
rect 5080 6808 5132 6817
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 5908 6808 5960 6860
rect 8576 6944 8628 6996
rect 11704 6944 11756 6996
rect 17776 6987 17828 6996
rect 17776 6953 17785 6987
rect 17785 6953 17819 6987
rect 17819 6953 17828 6987
rect 17776 6944 17828 6953
rect 18512 6987 18564 6996
rect 18512 6953 18527 6987
rect 18527 6953 18561 6987
rect 18561 6953 18564 6987
rect 18512 6944 18564 6953
rect 18696 6944 18748 6996
rect 20076 6944 20128 6996
rect 8484 6808 8536 6860
rect 1860 6672 1912 6724
rect 5448 6740 5500 6792
rect 6368 6740 6420 6792
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 3884 6647 3936 6656
rect 3884 6613 3893 6647
rect 3893 6613 3927 6647
rect 3927 6613 3936 6647
rect 3884 6604 3936 6613
rect 5356 6604 5408 6656
rect 5448 6647 5500 6656
rect 5448 6613 5457 6647
rect 5457 6613 5491 6647
rect 5491 6613 5500 6647
rect 5448 6604 5500 6613
rect 5816 6604 5868 6656
rect 7748 6604 7800 6656
rect 10416 6647 10468 6656
rect 10416 6613 10425 6647
rect 10425 6613 10459 6647
rect 10459 6613 10468 6647
rect 10416 6604 10468 6613
rect 11152 6808 11204 6860
rect 11244 6808 11296 6860
rect 11336 6851 11388 6860
rect 11336 6817 11345 6851
rect 11345 6817 11379 6851
rect 11379 6817 11388 6851
rect 11336 6808 11388 6817
rect 13820 6851 13872 6860
rect 13820 6817 13829 6851
rect 13829 6817 13863 6851
rect 13863 6817 13872 6851
rect 13820 6808 13872 6817
rect 13912 6808 13964 6860
rect 14188 6851 14240 6860
rect 14188 6817 14190 6851
rect 14190 6817 14240 6851
rect 14188 6808 14240 6817
rect 11060 6604 11112 6656
rect 12348 6740 12400 6792
rect 15936 6808 15988 6860
rect 16028 6808 16080 6860
rect 16396 6851 16448 6860
rect 16396 6817 16405 6851
rect 16405 6817 16439 6851
rect 16439 6817 16448 6851
rect 16396 6808 16448 6817
rect 17132 6876 17184 6928
rect 15660 6715 15712 6724
rect 15660 6681 15669 6715
rect 15669 6681 15703 6715
rect 15703 6681 15712 6715
rect 15660 6672 15712 6681
rect 16764 6740 16816 6792
rect 17316 6740 17368 6792
rect 16396 6672 16448 6724
rect 13268 6647 13320 6656
rect 13268 6613 13277 6647
rect 13277 6613 13311 6647
rect 13311 6613 13320 6647
rect 13268 6604 13320 6613
rect 13728 6604 13780 6656
rect 16212 6604 16264 6656
rect 16672 6604 16724 6656
rect 17592 6808 17644 6860
rect 17776 6808 17828 6860
rect 18420 6740 18472 6792
rect 18604 6740 18656 6792
rect 18696 6740 18748 6792
rect 19708 6808 19760 6860
rect 18972 6740 19024 6792
rect 20536 6808 20588 6860
rect 22100 6876 22152 6928
rect 23664 6944 23716 6996
rect 30012 6944 30064 6996
rect 22928 6808 22980 6860
rect 21088 6740 21140 6792
rect 22100 6783 22152 6792
rect 22100 6749 22109 6783
rect 22109 6749 22143 6783
rect 22143 6749 22152 6783
rect 22100 6740 22152 6749
rect 22468 6783 22520 6792
rect 22468 6749 22470 6783
rect 22470 6749 22520 6783
rect 22468 6740 22520 6749
rect 22744 6740 22796 6792
rect 23020 6740 23072 6792
rect 23664 6808 23716 6860
rect 24584 6851 24636 6860
rect 24584 6817 24593 6851
rect 24593 6817 24627 6851
rect 24627 6817 24636 6851
rect 24584 6808 24636 6817
rect 26148 6876 26200 6928
rect 27344 6876 27396 6928
rect 27620 6919 27672 6928
rect 27620 6885 27629 6919
rect 27629 6885 27663 6919
rect 27663 6885 27672 6919
rect 27620 6876 27672 6885
rect 27804 6876 27856 6928
rect 24952 6740 25004 6792
rect 17408 6647 17460 6656
rect 17408 6613 17417 6647
rect 17417 6613 17451 6647
rect 17451 6613 17460 6647
rect 17408 6604 17460 6613
rect 18052 6604 18104 6656
rect 18420 6604 18472 6656
rect 19156 6604 19208 6656
rect 20260 6647 20312 6656
rect 20260 6613 20269 6647
rect 20269 6613 20303 6647
rect 20303 6613 20312 6647
rect 20260 6604 20312 6613
rect 20352 6604 20404 6656
rect 21548 6604 21600 6656
rect 22376 6604 22428 6656
rect 23296 6604 23348 6656
rect 24124 6647 24176 6656
rect 24124 6613 24133 6647
rect 24133 6613 24167 6647
rect 24167 6613 24176 6647
rect 24124 6604 24176 6613
rect 24860 6604 24912 6656
rect 26240 6808 26292 6860
rect 26700 6808 26752 6860
rect 27712 6851 27764 6860
rect 27712 6817 27721 6851
rect 27721 6817 27755 6851
rect 27755 6817 27764 6851
rect 27712 6808 27764 6817
rect 30288 6808 30340 6860
rect 28264 6740 28316 6792
rect 27344 6672 27396 6724
rect 29552 6715 29604 6724
rect 29552 6681 29561 6715
rect 29561 6681 29595 6715
rect 29595 6681 29604 6715
rect 29552 6672 29604 6681
rect 28908 6604 28960 6656
rect 4193 6502 4245 6554
rect 4257 6502 4309 6554
rect 4321 6502 4373 6554
rect 4385 6502 4437 6554
rect 4449 6502 4501 6554
rect 11783 6502 11835 6554
rect 11847 6502 11899 6554
rect 11911 6502 11963 6554
rect 11975 6502 12027 6554
rect 12039 6502 12091 6554
rect 19373 6502 19425 6554
rect 19437 6502 19489 6554
rect 19501 6502 19553 6554
rect 19565 6502 19617 6554
rect 19629 6502 19681 6554
rect 26963 6502 27015 6554
rect 27027 6502 27079 6554
rect 27091 6502 27143 6554
rect 27155 6502 27207 6554
rect 27219 6502 27271 6554
rect 1216 6400 1268 6452
rect 2780 6443 2832 6452
rect 2780 6409 2789 6443
rect 2789 6409 2823 6443
rect 2823 6409 2832 6443
rect 2780 6400 2832 6409
rect 2136 6264 2188 6316
rect 4068 6264 4120 6316
rect 5724 6264 5776 6316
rect 5908 6307 5960 6316
rect 5908 6273 5910 6307
rect 5910 6273 5960 6307
rect 5908 6264 5960 6273
rect 6092 6264 6144 6316
rect 6460 6264 6512 6316
rect 756 6196 808 6248
rect 1584 6196 1636 6248
rect 2596 6196 2648 6248
rect 2872 6196 2924 6248
rect 3608 6196 3660 6248
rect 5264 6196 5316 6248
rect 7748 6128 7800 6180
rect 2136 6060 2188 6112
rect 4252 6060 4304 6112
rect 5080 6103 5132 6112
rect 5080 6069 5089 6103
rect 5089 6069 5123 6103
rect 5123 6069 5132 6103
rect 5080 6060 5132 6069
rect 5540 6060 5592 6112
rect 7656 6060 7708 6112
rect 9864 6400 9916 6452
rect 10600 6400 10652 6452
rect 13268 6400 13320 6452
rect 13452 6400 13504 6452
rect 14556 6400 14608 6452
rect 14648 6400 14700 6452
rect 16028 6400 16080 6452
rect 16212 6443 16264 6452
rect 16212 6409 16221 6443
rect 16221 6409 16255 6443
rect 16255 6409 16264 6443
rect 16212 6400 16264 6409
rect 8576 6264 8628 6316
rect 8484 6196 8536 6248
rect 10416 6196 10468 6248
rect 10508 6196 10560 6248
rect 11060 6307 11112 6316
rect 11060 6273 11072 6307
rect 11072 6273 11106 6307
rect 11106 6273 11112 6307
rect 11060 6264 11112 6273
rect 13084 6264 13136 6316
rect 11336 6239 11388 6248
rect 11336 6205 11345 6239
rect 11345 6205 11379 6239
rect 11379 6205 11388 6239
rect 11336 6196 11388 6205
rect 12716 6196 12768 6248
rect 13360 6264 13412 6316
rect 14372 6307 14424 6316
rect 14372 6273 14381 6307
rect 14381 6273 14415 6307
rect 14415 6273 14424 6307
rect 14372 6264 14424 6273
rect 14740 6264 14792 6316
rect 15200 6264 15252 6316
rect 15476 6264 15528 6316
rect 8944 6060 8996 6112
rect 11244 6060 11296 6112
rect 11796 6060 11848 6112
rect 13912 6128 13964 6180
rect 20628 6400 20680 6452
rect 20720 6443 20772 6452
rect 20720 6409 20729 6443
rect 20729 6409 20763 6443
rect 20763 6409 20772 6443
rect 20720 6400 20772 6409
rect 22744 6443 22796 6452
rect 22744 6409 22753 6443
rect 22753 6409 22787 6443
rect 22787 6409 22796 6443
rect 22744 6400 22796 6409
rect 17040 6332 17092 6384
rect 17776 6332 17828 6384
rect 17132 6239 17184 6248
rect 17132 6205 17141 6239
rect 17141 6205 17175 6239
rect 17175 6205 17184 6239
rect 17132 6196 17184 6205
rect 17500 6239 17552 6248
rect 17500 6205 17509 6239
rect 17509 6205 17543 6239
rect 17543 6205 17552 6239
rect 17500 6196 17552 6205
rect 17960 6239 18012 6248
rect 17960 6205 17969 6239
rect 17969 6205 18003 6239
rect 18003 6205 18012 6239
rect 17960 6196 18012 6205
rect 18144 6196 18196 6248
rect 18696 6332 18748 6384
rect 19248 6264 19300 6316
rect 18604 6196 18656 6248
rect 20536 6196 20588 6248
rect 21180 6196 21232 6248
rect 21548 6196 21600 6248
rect 21732 6196 21784 6248
rect 23296 6332 23348 6384
rect 24308 6264 24360 6316
rect 23848 6196 23900 6248
rect 25504 6196 25556 6248
rect 12440 6103 12492 6112
rect 12440 6069 12449 6103
rect 12449 6069 12483 6103
rect 12483 6069 12492 6103
rect 12440 6060 12492 6069
rect 12808 6103 12860 6112
rect 12808 6069 12817 6103
rect 12817 6069 12851 6103
rect 12851 6069 12860 6103
rect 12808 6060 12860 6069
rect 13084 6103 13136 6112
rect 13084 6069 13093 6103
rect 13093 6069 13127 6103
rect 13127 6069 13136 6103
rect 13084 6060 13136 6069
rect 13544 6103 13596 6112
rect 13544 6069 13553 6103
rect 13553 6069 13587 6103
rect 13587 6069 13596 6103
rect 13544 6060 13596 6069
rect 14464 6060 14516 6112
rect 14832 6103 14884 6112
rect 14832 6069 14847 6103
rect 14847 6069 14881 6103
rect 14881 6069 14884 6103
rect 14832 6060 14884 6069
rect 16856 6060 16908 6112
rect 16948 6103 17000 6112
rect 16948 6069 16957 6103
rect 16957 6069 16991 6103
rect 16991 6069 17000 6103
rect 16948 6060 17000 6069
rect 17224 6103 17276 6112
rect 17224 6069 17233 6103
rect 17233 6069 17267 6103
rect 17267 6069 17276 6103
rect 17224 6060 17276 6069
rect 18052 6060 18104 6112
rect 18972 6060 19024 6112
rect 19064 6060 19116 6112
rect 21548 6060 21600 6112
rect 22836 6060 22888 6112
rect 24400 6060 24452 6112
rect 25780 6060 25832 6112
rect 25872 6103 25924 6112
rect 25872 6069 25881 6103
rect 25881 6069 25915 6103
rect 25915 6069 25924 6103
rect 25872 6060 25924 6069
rect 26148 6264 26200 6316
rect 26700 6307 26752 6316
rect 26700 6273 26709 6307
rect 26709 6273 26743 6307
rect 26743 6273 26752 6307
rect 26700 6264 26752 6273
rect 26884 6264 26936 6316
rect 27436 6307 27488 6316
rect 27436 6273 27445 6307
rect 27445 6273 27479 6307
rect 27479 6273 27488 6307
rect 27436 6264 27488 6273
rect 26516 6196 26568 6248
rect 27896 6196 27948 6248
rect 26792 6128 26844 6180
rect 26332 6060 26384 6112
rect 26424 6103 26476 6112
rect 26424 6069 26433 6103
rect 26433 6069 26467 6103
rect 26467 6069 26476 6103
rect 26424 6060 26476 6069
rect 26608 6060 26660 6112
rect 29644 6060 29696 6112
rect 7988 5958 8040 6010
rect 8052 5958 8104 6010
rect 8116 5958 8168 6010
rect 8180 5958 8232 6010
rect 8244 5958 8296 6010
rect 15578 5958 15630 6010
rect 15642 5958 15694 6010
rect 15706 5958 15758 6010
rect 15770 5958 15822 6010
rect 15834 5958 15886 6010
rect 23168 5958 23220 6010
rect 23232 5958 23284 6010
rect 23296 5958 23348 6010
rect 23360 5958 23412 6010
rect 23424 5958 23476 6010
rect 30758 5958 30810 6010
rect 30822 5958 30874 6010
rect 30886 5958 30938 6010
rect 30950 5958 31002 6010
rect 31014 5958 31066 6010
rect 1032 5856 1084 5908
rect 1768 5899 1820 5908
rect 1768 5865 1783 5899
rect 1783 5865 1817 5899
rect 1817 5865 1820 5899
rect 1768 5856 1820 5865
rect 2136 5856 2188 5908
rect 664 5720 716 5772
rect 1400 5720 1452 5772
rect 3884 5856 3936 5908
rect 3976 5899 4028 5908
rect 3976 5865 3991 5899
rect 3991 5865 4025 5899
rect 4025 5865 4028 5899
rect 3976 5856 4028 5865
rect 5448 5856 5500 5908
rect 6092 5856 6144 5908
rect 7564 5856 7616 5908
rect 8668 5856 8720 5908
rect 10600 5856 10652 5908
rect 12716 5856 12768 5908
rect 13544 5856 13596 5908
rect 20352 5856 20404 5908
rect 21088 5856 21140 5908
rect 21548 5856 21600 5908
rect 22468 5856 22520 5908
rect 25688 5899 25740 5908
rect 25688 5865 25697 5899
rect 25697 5865 25731 5899
rect 25731 5865 25740 5899
rect 25688 5856 25740 5865
rect 25780 5856 25832 5908
rect 29276 5856 29328 5908
rect 29460 5856 29512 5908
rect 3516 5695 3568 5704
rect 3516 5661 3525 5695
rect 3525 5661 3559 5695
rect 3559 5661 3568 5695
rect 3516 5652 3568 5661
rect 4068 5652 4120 5704
rect 4620 5652 4672 5704
rect 4988 5652 5040 5704
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 6276 5695 6328 5704
rect 6276 5661 6288 5695
rect 6288 5661 6322 5695
rect 6322 5661 6328 5695
rect 6276 5652 6328 5661
rect 6736 5652 6788 5704
rect 7748 5652 7800 5704
rect 8484 5695 8536 5704
rect 8484 5661 8496 5695
rect 8496 5661 8530 5695
rect 8530 5661 8536 5695
rect 8484 5652 8536 5661
rect 8760 5695 8812 5704
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 11428 5763 11480 5772
rect 11428 5729 11437 5763
rect 11437 5729 11471 5763
rect 11471 5729 11480 5763
rect 11428 5720 11480 5729
rect 11520 5720 11572 5772
rect 11336 5584 11388 5636
rect 3976 5516 4028 5568
rect 4252 5516 4304 5568
rect 4988 5516 5040 5568
rect 6460 5516 6512 5568
rect 7012 5516 7064 5568
rect 9588 5516 9640 5568
rect 10232 5559 10284 5568
rect 10232 5525 10241 5559
rect 10241 5525 10275 5559
rect 10275 5525 10284 5559
rect 10232 5516 10284 5525
rect 10324 5516 10376 5568
rect 11612 5695 11664 5704
rect 11612 5661 11621 5695
rect 11621 5661 11655 5695
rect 11655 5661 11664 5695
rect 11612 5652 11664 5661
rect 12440 5720 12492 5772
rect 13728 5720 13780 5772
rect 14464 5720 14516 5772
rect 13820 5695 13872 5704
rect 13820 5661 13829 5695
rect 13829 5661 13863 5695
rect 13863 5661 13872 5695
rect 13820 5652 13872 5661
rect 14004 5652 14056 5704
rect 16212 5695 16264 5704
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16212 5652 16264 5661
rect 16580 5695 16632 5704
rect 16580 5661 16582 5695
rect 16582 5661 16632 5695
rect 16580 5652 16632 5661
rect 16856 5720 16908 5772
rect 18788 5695 18840 5704
rect 18788 5661 18790 5695
rect 18790 5661 18840 5695
rect 18788 5652 18840 5661
rect 20628 5788 20680 5840
rect 21180 5720 21232 5772
rect 21824 5720 21876 5772
rect 22192 5652 22244 5704
rect 24216 5695 24268 5704
rect 24216 5661 24225 5695
rect 24225 5661 24259 5695
rect 24259 5661 24268 5695
rect 24216 5652 24268 5661
rect 26056 5720 26108 5772
rect 26332 5720 26384 5772
rect 29092 5720 29144 5772
rect 26792 5652 26844 5704
rect 27160 5695 27212 5704
rect 27160 5661 27169 5695
rect 27169 5661 27203 5695
rect 27203 5661 27212 5695
rect 27160 5652 27212 5661
rect 27252 5652 27304 5704
rect 20628 5627 20680 5636
rect 20628 5593 20637 5627
rect 20637 5593 20671 5627
rect 20671 5593 20680 5627
rect 20628 5584 20680 5593
rect 28356 5584 28408 5636
rect 11796 5516 11848 5568
rect 14280 5516 14332 5568
rect 15476 5516 15528 5568
rect 16396 5516 16448 5568
rect 18328 5516 18380 5568
rect 18604 5516 18656 5568
rect 20812 5516 20864 5568
rect 21456 5516 21508 5568
rect 23112 5516 23164 5568
rect 24216 5516 24268 5568
rect 24952 5516 25004 5568
rect 25964 5559 26016 5568
rect 25964 5525 25973 5559
rect 25973 5525 26007 5559
rect 26007 5525 26016 5559
rect 25964 5516 26016 5525
rect 26056 5516 26108 5568
rect 27160 5516 27212 5568
rect 28264 5559 28316 5568
rect 28264 5525 28273 5559
rect 28273 5525 28307 5559
rect 28307 5525 28316 5559
rect 28264 5516 28316 5525
rect 28448 5516 28500 5568
rect 29276 5559 29328 5568
rect 29276 5525 29285 5559
rect 29285 5525 29319 5559
rect 29319 5525 29328 5559
rect 29276 5516 29328 5525
rect 4193 5414 4245 5466
rect 4257 5414 4309 5466
rect 4321 5414 4373 5466
rect 4385 5414 4437 5466
rect 4449 5414 4501 5466
rect 11783 5414 11835 5466
rect 11847 5414 11899 5466
rect 11911 5414 11963 5466
rect 11975 5414 12027 5466
rect 12039 5414 12091 5466
rect 19373 5414 19425 5466
rect 19437 5414 19489 5466
rect 19501 5414 19553 5466
rect 19565 5414 19617 5466
rect 19629 5414 19681 5466
rect 26963 5414 27015 5466
rect 27027 5414 27079 5466
rect 27091 5414 27143 5466
rect 27155 5414 27207 5466
rect 27219 5414 27271 5466
rect 664 5176 716 5228
rect 2872 5312 2924 5364
rect 4068 5312 4120 5364
rect 6276 5312 6328 5364
rect 3424 5244 3476 5296
rect 6092 5244 6144 5296
rect 4252 5176 4304 5228
rect 5080 5176 5132 5228
rect 6276 5176 6328 5228
rect 7012 5176 7064 5228
rect 1676 5151 1728 5160
rect 1676 5117 1685 5151
rect 1685 5117 1719 5151
rect 1719 5117 1728 5151
rect 1676 5108 1728 5117
rect 3516 5108 3568 5160
rect 2872 5040 2924 5092
rect 3700 5040 3752 5092
rect 3792 5040 3844 5092
rect 5356 5108 5408 5160
rect 6736 5108 6788 5160
rect 10232 5312 10284 5364
rect 7564 5176 7616 5228
rect 8852 5176 8904 5228
rect 9404 5219 9456 5228
rect 9404 5185 9406 5219
rect 9406 5185 9456 5219
rect 9404 5176 9456 5185
rect 9588 5176 9640 5228
rect 7840 5108 7892 5160
rect 8944 5108 8996 5160
rect 9036 5151 9088 5160
rect 9036 5117 9045 5151
rect 9045 5117 9079 5151
rect 9079 5117 9088 5151
rect 9036 5108 9088 5117
rect 11060 5176 11112 5228
rect 1768 4972 1820 5024
rect 2136 4972 2188 5024
rect 3884 4972 3936 5024
rect 6368 4972 6420 5024
rect 6552 5015 6604 5024
rect 6552 4981 6567 5015
rect 6567 4981 6601 5015
rect 6601 4981 6604 5015
rect 6552 4972 6604 4981
rect 9772 5151 9824 5160
rect 9772 5117 9781 5151
rect 9781 5117 9815 5151
rect 9815 5117 9824 5151
rect 9772 5108 9824 5117
rect 13728 5312 13780 5364
rect 21732 5312 21784 5364
rect 23020 5312 23072 5364
rect 23112 5287 23164 5296
rect 23112 5253 23121 5287
rect 23121 5253 23155 5287
rect 23155 5253 23164 5287
rect 23112 5244 23164 5253
rect 11428 5176 11480 5228
rect 11612 5176 11664 5228
rect 11704 5219 11756 5228
rect 11704 5185 11716 5219
rect 11716 5185 11750 5219
rect 11750 5185 11756 5219
rect 11704 5176 11756 5185
rect 12808 5176 12860 5228
rect 13636 5176 13688 5228
rect 9496 4972 9548 5024
rect 11888 5108 11940 5160
rect 13820 5108 13872 5160
rect 13912 5151 13964 5160
rect 13912 5117 13921 5151
rect 13921 5117 13955 5151
rect 13955 5117 13964 5151
rect 13912 5108 13964 5117
rect 11152 5083 11204 5092
rect 11152 5049 11161 5083
rect 11161 5049 11195 5083
rect 11195 5049 11204 5083
rect 11152 5040 11204 5049
rect 14556 5176 14608 5228
rect 16948 5219 17000 5228
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 20260 5176 20312 5228
rect 21456 5176 21508 5228
rect 16304 5108 16356 5160
rect 18328 5040 18380 5092
rect 11520 4972 11572 5024
rect 13636 4972 13688 5024
rect 13728 5015 13780 5024
rect 13728 4981 13737 5015
rect 13737 4981 13771 5015
rect 13771 4981 13780 5015
rect 13728 4972 13780 4981
rect 14004 4972 14056 5024
rect 16580 4972 16632 5024
rect 16856 4972 16908 5024
rect 17316 4972 17368 5024
rect 18788 4972 18840 5024
rect 20720 5108 20772 5160
rect 21180 5108 21232 5160
rect 22744 5108 22796 5160
rect 29368 5312 29420 5364
rect 25504 5244 25556 5296
rect 24952 5176 25004 5228
rect 25964 5176 26016 5228
rect 26608 5176 26660 5228
rect 23848 5108 23900 5160
rect 21272 4972 21324 5024
rect 21548 4972 21600 5024
rect 21640 4972 21692 5024
rect 23664 5040 23716 5092
rect 26332 5040 26384 5092
rect 26700 5151 26752 5160
rect 26700 5117 26709 5151
rect 26709 5117 26743 5151
rect 26743 5117 26752 5151
rect 26700 5108 26752 5117
rect 27528 5176 27580 5228
rect 27804 5176 27856 5228
rect 29092 5176 29144 5228
rect 26516 5040 26568 5092
rect 22744 5015 22796 5024
rect 22744 4981 22753 5015
rect 22753 4981 22787 5015
rect 22787 4981 22796 5015
rect 22744 4972 22796 4981
rect 24400 4972 24452 5024
rect 25228 4972 25280 5024
rect 29000 4972 29052 5024
rect 29460 5015 29512 5024
rect 29460 4981 29469 5015
rect 29469 4981 29503 5015
rect 29503 4981 29512 5015
rect 29460 4972 29512 4981
rect 7988 4870 8040 4922
rect 8052 4870 8104 4922
rect 8116 4870 8168 4922
rect 8180 4870 8232 4922
rect 8244 4870 8296 4922
rect 15578 4870 15630 4922
rect 15642 4870 15694 4922
rect 15706 4870 15758 4922
rect 15770 4870 15822 4922
rect 15834 4870 15886 4922
rect 23168 4870 23220 4922
rect 23232 4870 23284 4922
rect 23296 4870 23348 4922
rect 23360 4870 23412 4922
rect 23424 4870 23476 4922
rect 30758 4870 30810 4922
rect 30822 4870 30874 4922
rect 30886 4870 30938 4922
rect 30950 4870 31002 4922
rect 31014 4870 31066 4922
rect 848 4768 900 4820
rect 1952 4768 2004 4820
rect 3884 4768 3936 4820
rect 6276 4811 6328 4820
rect 6276 4777 6291 4811
rect 6291 4777 6325 4811
rect 6325 4777 6328 4811
rect 6276 4768 6328 4777
rect 8668 4768 8720 4820
rect 8852 4768 8904 4820
rect 9772 4768 9824 4820
rect 10876 4768 10928 4820
rect 10968 4768 11020 4820
rect 848 4564 900 4616
rect 1492 4564 1544 4616
rect 2780 4632 2832 4684
rect 2044 4607 2096 4616
rect 2044 4573 2053 4607
rect 2053 4573 2087 4607
rect 2087 4573 2096 4607
rect 2044 4564 2096 4573
rect 940 4428 992 4480
rect 3148 4564 3200 4616
rect 3424 4564 3476 4616
rect 3976 4607 4028 4616
rect 3976 4573 3988 4607
rect 3988 4573 4022 4607
rect 4022 4573 4028 4607
rect 3976 4564 4028 4573
rect 5264 4564 5316 4616
rect 5816 4607 5868 4616
rect 5816 4573 5825 4607
rect 5825 4573 5859 4607
rect 5859 4573 5868 4607
rect 5816 4564 5868 4573
rect 6368 4564 6420 4616
rect 6736 4564 6788 4616
rect 7748 4564 7800 4616
rect 8576 4632 8628 4684
rect 8852 4632 8904 4684
rect 11060 4632 11112 4684
rect 11336 4768 11388 4820
rect 11520 4768 11572 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 13728 4768 13780 4820
rect 16856 4768 16908 4820
rect 17776 4768 17828 4820
rect 21640 4768 21692 4820
rect 21732 4811 21784 4820
rect 21732 4777 21741 4811
rect 21741 4777 21775 4811
rect 21775 4777 21784 4811
rect 21732 4768 21784 4777
rect 21824 4768 21876 4820
rect 22468 4768 22520 4820
rect 26056 4768 26108 4820
rect 11888 4632 11940 4684
rect 13084 4632 13136 4684
rect 20536 4743 20588 4752
rect 20536 4709 20545 4743
rect 20545 4709 20579 4743
rect 20579 4709 20588 4743
rect 20536 4700 20588 4709
rect 21272 4700 21324 4752
rect 11428 4564 11480 4616
rect 12072 4609 12124 4616
rect 12072 4575 12084 4609
rect 12084 4575 12118 4609
rect 12118 4575 12124 4609
rect 12072 4564 12124 4575
rect 13820 4607 13872 4616
rect 13820 4573 13829 4607
rect 13829 4573 13863 4607
rect 13863 4573 13872 4607
rect 13820 4564 13872 4573
rect 14004 4564 14056 4616
rect 14280 4607 14332 4616
rect 14280 4573 14292 4607
rect 14292 4573 14326 4607
rect 14326 4573 14332 4607
rect 14280 4564 14332 4573
rect 16396 4564 16448 4616
rect 17224 4632 17276 4684
rect 9496 4496 9548 4548
rect 11520 4496 11572 4548
rect 18788 4607 18840 4616
rect 18788 4573 18790 4607
rect 18790 4573 18840 4607
rect 18788 4564 18840 4573
rect 18972 4632 19024 4684
rect 20812 4675 20864 4684
rect 20812 4641 20821 4675
rect 20821 4641 20855 4675
rect 20855 4641 20864 4675
rect 20812 4632 20864 4641
rect 21180 4632 21232 4684
rect 21364 4632 21416 4684
rect 24308 4700 24360 4752
rect 28448 4768 28500 4820
rect 29644 4768 29696 4820
rect 22192 4632 22244 4684
rect 22744 4632 22796 4684
rect 22836 4675 22888 4684
rect 22836 4641 22845 4675
rect 22845 4641 22879 4675
rect 22879 4641 22888 4675
rect 22836 4632 22888 4641
rect 23664 4632 23716 4684
rect 26148 4632 26200 4684
rect 27160 4700 27212 4752
rect 27804 4632 27856 4684
rect 27896 4675 27948 4684
rect 27896 4641 27905 4675
rect 27905 4641 27939 4675
rect 27939 4641 27948 4675
rect 27896 4632 27948 4641
rect 19248 4564 19300 4616
rect 3148 4471 3200 4480
rect 3148 4437 3157 4471
rect 3157 4437 3191 4471
rect 3191 4437 3200 4471
rect 3148 4428 3200 4437
rect 3516 4428 3568 4480
rect 8852 4428 8904 4480
rect 10048 4471 10100 4480
rect 10048 4437 10057 4471
rect 10057 4437 10091 4471
rect 10091 4437 10100 4471
rect 10048 4428 10100 4437
rect 12164 4428 12216 4480
rect 12256 4428 12308 4480
rect 16672 4428 16724 4480
rect 18328 4428 18380 4480
rect 19064 4428 19116 4480
rect 20996 4428 21048 4480
rect 21456 4428 21508 4480
rect 26516 4564 26568 4616
rect 28172 4564 28224 4616
rect 28540 4632 28592 4684
rect 26792 4496 26844 4548
rect 27896 4496 27948 4548
rect 24768 4428 24820 4480
rect 26608 4428 26660 4480
rect 26700 4471 26752 4480
rect 26700 4437 26709 4471
rect 26709 4437 26743 4471
rect 26743 4437 26752 4471
rect 26700 4428 26752 4437
rect 26884 4428 26936 4480
rect 4193 4326 4245 4378
rect 4257 4326 4309 4378
rect 4321 4326 4373 4378
rect 4385 4326 4437 4378
rect 4449 4326 4501 4378
rect 11783 4326 11835 4378
rect 11847 4326 11899 4378
rect 11911 4326 11963 4378
rect 11975 4326 12027 4378
rect 12039 4326 12091 4378
rect 19373 4326 19425 4378
rect 19437 4326 19489 4378
rect 19501 4326 19553 4378
rect 19565 4326 19617 4378
rect 19629 4326 19681 4378
rect 26963 4326 27015 4378
rect 27027 4326 27079 4378
rect 27091 4326 27143 4378
rect 27155 4326 27207 4378
rect 27219 4326 27271 4378
rect 3056 4224 3108 4276
rect 848 4131 900 4140
rect 848 4097 857 4131
rect 857 4097 891 4131
rect 891 4097 900 4131
rect 848 4088 900 4097
rect 1308 4113 1360 4140
rect 1308 4088 1353 4113
rect 1353 4088 1360 4113
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 1676 4088 1728 4140
rect 3976 4088 4028 4140
rect 4344 4088 4396 4140
rect 4528 4131 4580 4140
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 4528 4088 4580 4097
rect 5908 4131 5960 4140
rect 5908 4097 5917 4131
rect 5917 4097 5951 4131
rect 5951 4097 5960 4131
rect 5908 4088 5960 4097
rect 7564 4224 7616 4276
rect 9036 4156 9088 4208
rect 11704 4224 11756 4276
rect 2964 4063 3016 4072
rect 2964 4029 2973 4063
rect 2973 4029 3007 4063
rect 3007 4029 3016 4063
rect 2964 4020 3016 4029
rect 5448 4020 5500 4072
rect 5632 4020 5684 4072
rect 6184 4088 6236 4140
rect 9680 4088 9732 4140
rect 1492 3884 1544 3936
rect 1584 3884 1636 3936
rect 3056 3884 3108 3936
rect 3700 3884 3752 3936
rect 5632 3884 5684 3936
rect 8944 4020 8996 4072
rect 7840 3927 7892 3936
rect 7840 3893 7849 3927
rect 7849 3893 7883 3927
rect 7883 3893 7892 3927
rect 7840 3884 7892 3893
rect 8668 3995 8720 4004
rect 8668 3961 8677 3995
rect 8677 3961 8711 3995
rect 8711 3961 8720 3995
rect 8668 3952 8720 3961
rect 8852 3952 8904 4004
rect 12256 4156 12308 4208
rect 10048 4088 10100 4140
rect 10692 4088 10744 4140
rect 13820 4088 13872 4140
rect 14648 4088 14700 4140
rect 26884 4224 26936 4276
rect 10508 4020 10560 4072
rect 12808 4020 12860 4072
rect 14832 4020 14884 4072
rect 15200 4020 15252 4072
rect 17868 4088 17920 4140
rect 19248 4156 19300 4208
rect 18788 4088 18840 4140
rect 20720 4088 20772 4140
rect 20812 4131 20864 4140
rect 20812 4097 20824 4131
rect 20824 4097 20858 4131
rect 20858 4097 20864 4131
rect 20812 4088 20864 4097
rect 20996 4088 21048 4140
rect 22468 4088 22520 4140
rect 16212 4020 16264 4072
rect 16488 4020 16540 4072
rect 17776 4020 17828 4072
rect 18696 4063 18748 4072
rect 18696 4029 18705 4063
rect 18705 4029 18739 4063
rect 18739 4029 18748 4063
rect 18696 4020 18748 4029
rect 9404 3952 9456 4004
rect 9772 3884 9824 3936
rect 12900 3952 12952 4004
rect 11244 3884 11296 3936
rect 11336 3884 11388 3936
rect 16304 3995 16356 4004
rect 16304 3961 16313 3995
rect 16313 3961 16347 3995
rect 16347 3961 16356 3995
rect 16304 3952 16356 3961
rect 16396 3884 16448 3936
rect 18880 3952 18932 4004
rect 16672 3884 16724 3936
rect 16764 3884 16816 3936
rect 19248 3952 19300 4004
rect 19892 4020 19944 4072
rect 21180 4020 21232 4072
rect 23756 4088 23808 4140
rect 23572 4020 23624 4072
rect 24768 4020 24820 4072
rect 25872 4088 25924 4140
rect 26424 4088 26476 4140
rect 26516 4088 26568 4140
rect 27252 4088 27304 4140
rect 30380 4088 30432 4140
rect 25136 4020 25188 4072
rect 26792 4020 26844 4072
rect 29184 4020 29236 4072
rect 19800 3884 19852 3936
rect 21548 3884 21600 3936
rect 22468 3884 22520 3936
rect 23020 3884 23072 3936
rect 24400 3952 24452 4004
rect 29092 3952 29144 4004
rect 23664 3884 23716 3936
rect 26056 3884 26108 3936
rect 26516 3927 26568 3936
rect 26516 3893 26525 3927
rect 26525 3893 26559 3927
rect 26559 3893 26568 3927
rect 26516 3884 26568 3893
rect 28080 3884 28132 3936
rect 29460 3884 29512 3936
rect 7988 3782 8040 3834
rect 8052 3782 8104 3834
rect 8116 3782 8168 3834
rect 8180 3782 8232 3834
rect 8244 3782 8296 3834
rect 15578 3782 15630 3834
rect 15642 3782 15694 3834
rect 15706 3782 15758 3834
rect 15770 3782 15822 3834
rect 15834 3782 15886 3834
rect 23168 3782 23220 3834
rect 23232 3782 23284 3834
rect 23296 3782 23348 3834
rect 23360 3782 23412 3834
rect 23424 3782 23476 3834
rect 30758 3782 30810 3834
rect 30822 3782 30874 3834
rect 30886 3782 30938 3834
rect 30950 3782 31002 3834
rect 31014 3782 31066 3834
rect 3792 3680 3844 3732
rect 3884 3680 3936 3732
rect 4344 3680 4396 3732
rect 5816 3680 5868 3732
rect 6736 3680 6788 3732
rect 7840 3680 7892 3732
rect 8576 3680 8628 3732
rect 9404 3680 9456 3732
rect 11612 3680 11664 3732
rect 16212 3680 16264 3732
rect 16488 3680 16540 3732
rect 16856 3680 16908 3732
rect 5724 3612 5776 3664
rect 1676 3587 1728 3596
rect 1676 3553 1678 3587
rect 1678 3553 1728 3587
rect 1032 3476 1084 3528
rect 1676 3544 1728 3553
rect 8484 3612 8536 3664
rect 2412 3476 2464 3528
rect 3516 3519 3568 3528
rect 3516 3485 3525 3519
rect 3525 3485 3559 3519
rect 3559 3485 3568 3519
rect 3516 3476 3568 3485
rect 3976 3519 4028 3528
rect 3976 3485 3988 3519
rect 3988 3485 4022 3519
rect 4022 3485 4028 3519
rect 3976 3476 4028 3485
rect 4896 3476 4948 3528
rect 5264 3476 5316 3528
rect 6368 3519 6420 3528
rect 6368 3485 6370 3519
rect 6370 3485 6420 3519
rect 6368 3476 6420 3485
rect 6460 3519 6512 3528
rect 6460 3485 6472 3519
rect 6472 3485 6506 3519
rect 6506 3485 6512 3519
rect 6460 3476 6512 3485
rect 6736 3519 6788 3528
rect 6736 3485 6745 3519
rect 6745 3485 6779 3519
rect 6779 3485 6788 3519
rect 6736 3476 6788 3485
rect 6920 3476 6972 3528
rect 8944 3544 8996 3596
rect 9036 3476 9088 3528
rect 9220 3476 9272 3528
rect 9496 3544 9548 3596
rect 11244 3544 11296 3596
rect 11428 3544 11480 3596
rect 12164 3544 12216 3596
rect 5816 3408 5868 3460
rect 6460 3340 6512 3392
rect 13820 3519 13872 3528
rect 13820 3485 13829 3519
rect 13829 3485 13863 3519
rect 13863 3485 13872 3519
rect 13820 3476 13872 3485
rect 14004 3476 14056 3528
rect 14372 3476 14424 3528
rect 16396 3476 16448 3528
rect 16672 3544 16724 3596
rect 20812 3680 20864 3732
rect 21088 3680 21140 3732
rect 22560 3680 22612 3732
rect 24216 3680 24268 3732
rect 24860 3680 24912 3732
rect 26148 3680 26200 3732
rect 21548 3655 21600 3664
rect 21548 3621 21557 3655
rect 21557 3621 21591 3655
rect 21591 3621 21600 3655
rect 21548 3612 21600 3621
rect 24308 3612 24360 3664
rect 17960 3476 18012 3528
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 18328 3476 18380 3485
rect 18696 3519 18748 3528
rect 18696 3485 18698 3519
rect 18698 3485 18748 3519
rect 18696 3476 18748 3485
rect 19064 3587 19116 3596
rect 19064 3553 19073 3587
rect 19073 3553 19107 3587
rect 19107 3553 19116 3587
rect 19064 3544 19116 3553
rect 19892 3544 19944 3596
rect 20720 3544 20772 3596
rect 21364 3476 21416 3528
rect 21732 3476 21784 3528
rect 22192 3544 22244 3596
rect 23020 3587 23072 3596
rect 23020 3553 23029 3587
rect 23029 3553 23063 3587
rect 23063 3553 23072 3587
rect 23020 3544 23072 3553
rect 23756 3544 23808 3596
rect 22468 3476 22520 3528
rect 23480 3476 23532 3528
rect 25688 3544 25740 3596
rect 26884 3612 26936 3664
rect 29184 3680 29236 3732
rect 29828 3723 29880 3732
rect 29828 3689 29837 3723
rect 29837 3689 29871 3723
rect 29871 3689 29880 3723
rect 29828 3680 29880 3689
rect 27896 3544 27948 3596
rect 28816 3544 28868 3596
rect 27620 3519 27672 3528
rect 27620 3485 27629 3519
rect 27629 3485 27663 3519
rect 27663 3485 27672 3519
rect 27620 3476 27672 3485
rect 28172 3476 28224 3528
rect 28448 3519 28500 3528
rect 28448 3485 28460 3519
rect 28460 3485 28494 3519
rect 28494 3485 28500 3519
rect 28448 3476 28500 3485
rect 28540 3476 28592 3528
rect 30104 3544 30156 3596
rect 29092 3476 29144 3528
rect 14004 3340 14056 3392
rect 14464 3340 14516 3392
rect 15936 3340 15988 3392
rect 18052 3340 18104 3392
rect 19892 3408 19944 3460
rect 19248 3340 19300 3392
rect 21824 3383 21876 3392
rect 21824 3349 21833 3383
rect 21833 3349 21867 3383
rect 21867 3349 21876 3383
rect 21824 3340 21876 3349
rect 24584 3340 24636 3392
rect 25320 3383 25372 3392
rect 25320 3349 25329 3383
rect 25329 3349 25363 3383
rect 25363 3349 25372 3383
rect 25320 3340 25372 3349
rect 25596 3383 25648 3392
rect 25596 3349 25605 3383
rect 25605 3349 25639 3383
rect 25639 3349 25648 3383
rect 25596 3340 25648 3349
rect 25688 3340 25740 3392
rect 29552 3340 29604 3392
rect 4193 3238 4245 3290
rect 4257 3238 4309 3290
rect 4321 3238 4373 3290
rect 4385 3238 4437 3290
rect 4449 3238 4501 3290
rect 11783 3238 11835 3290
rect 11847 3238 11899 3290
rect 11911 3238 11963 3290
rect 11975 3238 12027 3290
rect 12039 3238 12091 3290
rect 19373 3238 19425 3290
rect 19437 3238 19489 3290
rect 19501 3238 19553 3290
rect 19565 3238 19617 3290
rect 19629 3238 19681 3290
rect 26963 3238 27015 3290
rect 27027 3238 27079 3290
rect 27091 3238 27143 3290
rect 27155 3238 27207 3290
rect 27219 3238 27271 3290
rect 3240 3179 3292 3188
rect 3240 3145 3249 3179
rect 3249 3145 3283 3179
rect 3283 3145 3292 3179
rect 3240 3136 3292 3145
rect 5632 3136 5684 3188
rect 5724 3179 5776 3188
rect 5724 3145 5733 3179
rect 5733 3145 5767 3179
rect 5767 3145 5776 3179
rect 5724 3136 5776 3145
rect 9220 3136 9272 3188
rect 9680 3136 9732 3188
rect 15936 3136 15988 3188
rect 5816 3068 5868 3120
rect 6000 3068 6052 3120
rect 13176 3068 13228 3120
rect 4252 3000 4304 3052
rect 5540 3000 5592 3052
rect 7656 3000 7708 3052
rect 7840 3000 7892 3052
rect 9404 3043 9456 3052
rect 1584 2932 1636 2984
rect 2136 2932 2188 2984
rect 3700 2932 3752 2984
rect 3056 2907 3108 2916
rect 3056 2873 3065 2907
rect 3065 2873 3099 2907
rect 3099 2873 3108 2907
rect 3056 2864 3108 2873
rect 3516 2864 3568 2916
rect 3884 2975 3936 2984
rect 3884 2941 3893 2975
rect 3893 2941 3927 2975
rect 3927 2941 3936 2975
rect 3884 2932 3936 2941
rect 4620 2975 4672 2984
rect 4620 2941 4629 2975
rect 4629 2941 4663 2975
rect 4663 2941 4672 2975
rect 4620 2932 4672 2941
rect 6092 2975 6144 2984
rect 6092 2941 6101 2975
rect 6101 2941 6135 2975
rect 6135 2941 6144 2975
rect 6092 2932 6144 2941
rect 6184 2932 6236 2984
rect 3884 2796 3936 2848
rect 4160 2796 4212 2848
rect 6552 2839 6604 2848
rect 6552 2805 6567 2839
rect 6567 2805 6601 2839
rect 6601 2805 6604 2839
rect 8484 2932 8536 2984
rect 8668 2932 8720 2984
rect 9036 2975 9088 2984
rect 9036 2941 9045 2975
rect 9045 2941 9079 2975
rect 9079 2941 9088 2975
rect 9036 2932 9088 2941
rect 9404 3009 9406 3043
rect 9406 3009 9456 3043
rect 9404 3000 9456 3009
rect 9588 3000 9640 3052
rect 11336 2932 11388 2984
rect 11520 2932 11572 2984
rect 16396 3136 16448 3188
rect 19800 3136 19852 3188
rect 19248 3000 19300 3052
rect 19340 3000 19392 3052
rect 21824 3136 21876 3188
rect 22284 3136 22336 3188
rect 20720 3000 20772 3052
rect 21456 3000 21508 3052
rect 23572 3136 23624 3188
rect 23848 3136 23900 3188
rect 25780 3136 25832 3188
rect 28540 3136 28592 3188
rect 30196 3179 30248 3188
rect 30196 3145 30205 3179
rect 30205 3145 30239 3179
rect 30239 3145 30248 3179
rect 30196 3136 30248 3145
rect 23848 3043 23900 3052
rect 23848 3009 23857 3043
rect 23857 3009 23891 3043
rect 23891 3009 23900 3043
rect 23848 3000 23900 3009
rect 24032 3000 24084 3052
rect 25228 3000 25280 3052
rect 26332 3000 26384 3052
rect 26608 3000 26660 3052
rect 27712 3000 27764 3052
rect 29920 3000 29972 3052
rect 13912 2932 13964 2984
rect 13176 2864 13228 2916
rect 16028 2932 16080 2984
rect 6552 2796 6604 2805
rect 7748 2796 7800 2848
rect 8944 2796 8996 2848
rect 11336 2796 11388 2848
rect 11612 2796 11664 2848
rect 14372 2796 14424 2848
rect 14464 2839 14516 2848
rect 14464 2805 14479 2839
rect 14479 2805 14513 2839
rect 14513 2805 14516 2839
rect 14464 2796 14516 2805
rect 15108 2796 15160 2848
rect 18512 2932 18564 2984
rect 18788 2864 18840 2916
rect 16856 2796 16908 2848
rect 21548 2932 21600 2984
rect 23664 2932 23716 2984
rect 24492 2932 24544 2984
rect 26424 2932 26476 2984
rect 28172 2932 28224 2984
rect 23572 2864 23624 2916
rect 29920 2864 29972 2916
rect 30380 2864 30432 2916
rect 23940 2796 23992 2848
rect 24216 2796 24268 2848
rect 24676 2796 24728 2848
rect 26056 2796 26108 2848
rect 26884 2796 26936 2848
rect 28080 2839 28132 2848
rect 28080 2805 28089 2839
rect 28089 2805 28123 2839
rect 28123 2805 28132 2839
rect 28080 2796 28132 2805
rect 7988 2694 8040 2746
rect 8052 2694 8104 2746
rect 8116 2694 8168 2746
rect 8180 2694 8232 2746
rect 8244 2694 8296 2746
rect 15578 2694 15630 2746
rect 15642 2694 15694 2746
rect 15706 2694 15758 2746
rect 15770 2694 15822 2746
rect 15834 2694 15886 2746
rect 23168 2694 23220 2746
rect 23232 2694 23284 2746
rect 23296 2694 23348 2746
rect 23360 2694 23412 2746
rect 23424 2694 23476 2746
rect 30758 2694 30810 2746
rect 30822 2694 30874 2746
rect 30886 2694 30938 2746
rect 30950 2694 31002 2746
rect 31014 2694 31066 2746
rect 940 2635 992 2644
rect 940 2601 949 2635
rect 949 2601 983 2635
rect 983 2601 992 2635
rect 940 2592 992 2601
rect 1768 2635 1820 2644
rect 1768 2601 1783 2635
rect 1783 2601 1817 2635
rect 1817 2601 1820 2635
rect 1768 2592 1820 2601
rect 3516 2592 3568 2644
rect 4160 2592 4212 2644
rect 5540 2635 5592 2644
rect 5540 2601 5549 2635
rect 5549 2601 5583 2635
rect 5583 2601 5592 2635
rect 5540 2592 5592 2601
rect 6368 2635 6420 2644
rect 6368 2601 6383 2635
rect 6383 2601 6417 2635
rect 6417 2601 6420 2635
rect 6368 2592 6420 2601
rect 756 2456 808 2508
rect 1676 2388 1728 2440
rect 3148 2456 3200 2508
rect 4252 2499 4304 2508
rect 4252 2465 4261 2499
rect 4261 2465 4295 2499
rect 4295 2465 4304 2499
rect 4252 2456 4304 2465
rect 5724 2456 5776 2508
rect 1676 2252 1728 2304
rect 2136 2252 2188 2304
rect 3792 2388 3844 2440
rect 5264 2320 5316 2372
rect 5448 2320 5500 2372
rect 6276 2388 6328 2440
rect 6460 2388 6512 2440
rect 6644 2499 6696 2508
rect 6644 2465 6653 2499
rect 6653 2465 6687 2499
rect 6687 2465 6696 2499
rect 6644 2456 6696 2465
rect 9588 2592 9640 2644
rect 10048 2592 10100 2644
rect 8484 2499 8536 2508
rect 7380 2388 7432 2440
rect 7748 2388 7800 2440
rect 8484 2465 8486 2499
rect 8486 2465 8536 2499
rect 8484 2456 8536 2465
rect 10324 2456 10376 2508
rect 7564 2320 7616 2372
rect 12992 2592 13044 2644
rect 14280 2635 14332 2644
rect 14280 2601 14295 2635
rect 14295 2601 14329 2635
rect 14329 2601 14332 2635
rect 14280 2592 14332 2601
rect 14464 2592 14516 2644
rect 16856 2592 16908 2644
rect 18788 2635 18840 2644
rect 18788 2601 18803 2635
rect 18803 2601 18837 2635
rect 18837 2601 18840 2635
rect 18788 2592 18840 2601
rect 20720 2592 20772 2644
rect 21548 2592 21600 2644
rect 24032 2592 24084 2644
rect 11612 2524 11664 2576
rect 25688 2592 25740 2644
rect 25780 2592 25832 2644
rect 27344 2592 27396 2644
rect 27712 2592 27764 2644
rect 27988 2592 28040 2644
rect 11428 2456 11480 2508
rect 10508 2388 10560 2440
rect 11244 2388 11296 2440
rect 11796 2388 11848 2440
rect 12348 2431 12400 2440
rect 12348 2397 12357 2431
rect 12357 2397 12391 2431
rect 12391 2397 12400 2431
rect 12348 2388 12400 2397
rect 13820 2431 13872 2440
rect 13820 2397 13829 2431
rect 13829 2397 13863 2431
rect 13863 2397 13872 2431
rect 13820 2388 13872 2397
rect 14464 2456 14516 2508
rect 16028 2388 16080 2440
rect 8116 2252 8168 2304
rect 10968 2252 11020 2304
rect 11152 2252 11204 2304
rect 18328 2431 18380 2440
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18328 2388 18380 2397
rect 22284 2456 22336 2508
rect 23756 2456 23808 2508
rect 25320 2456 25372 2508
rect 25504 2456 25556 2508
rect 26424 2456 26476 2508
rect 27528 2456 27580 2508
rect 20352 2363 20404 2372
rect 20352 2329 20361 2363
rect 20361 2329 20395 2363
rect 20395 2329 20404 2363
rect 20352 2320 20404 2329
rect 20536 2252 20588 2304
rect 20720 2320 20772 2372
rect 21640 2388 21692 2440
rect 23480 2388 23532 2440
rect 23572 2388 23624 2440
rect 24124 2431 24176 2440
rect 24124 2397 24133 2431
rect 24133 2397 24167 2431
rect 24167 2397 24176 2431
rect 24124 2388 24176 2397
rect 24308 2388 24360 2440
rect 24584 2431 24636 2440
rect 24584 2397 24596 2431
rect 24596 2397 24630 2431
rect 24630 2397 24636 2431
rect 24584 2388 24636 2397
rect 24768 2388 24820 2440
rect 27896 2456 27948 2508
rect 30012 2635 30064 2644
rect 30012 2601 30021 2635
rect 30021 2601 30055 2635
rect 30055 2601 30064 2635
rect 30012 2592 30064 2601
rect 29736 2456 29788 2508
rect 21916 2252 21968 2304
rect 22192 2252 22244 2304
rect 24492 2252 24544 2304
rect 25964 2295 26016 2304
rect 25964 2261 25973 2295
rect 25973 2261 26007 2295
rect 26007 2261 26016 2295
rect 25964 2252 26016 2261
rect 26424 2252 26476 2304
rect 28172 2388 28224 2440
rect 28540 2388 28592 2440
rect 4193 2150 4245 2202
rect 4257 2150 4309 2202
rect 4321 2150 4373 2202
rect 4385 2150 4437 2202
rect 4449 2150 4501 2202
rect 11783 2150 11835 2202
rect 11847 2150 11899 2202
rect 11911 2150 11963 2202
rect 11975 2150 12027 2202
rect 12039 2150 12091 2202
rect 19373 2150 19425 2202
rect 19437 2150 19489 2202
rect 19501 2150 19553 2202
rect 19565 2150 19617 2202
rect 19629 2150 19681 2202
rect 26963 2150 27015 2202
rect 27027 2150 27079 2202
rect 27091 2150 27143 2202
rect 27155 2150 27207 2202
rect 27219 2150 27271 2202
rect 1124 2048 1176 2100
rect 2780 1912 2832 1964
rect 1308 1844 1360 1896
rect 2504 1844 2556 1896
rect 3608 2048 3660 2100
rect 4528 2048 4580 2100
rect 5632 2048 5684 2100
rect 3792 1912 3844 1964
rect 3976 1955 4028 1964
rect 3976 1921 3978 1955
rect 3978 1921 4028 1955
rect 3976 1912 4028 1921
rect 4068 1912 4120 1964
rect 4344 1955 4396 1964
rect 4344 1921 4353 1955
rect 4353 1921 4387 1955
rect 4387 1921 4396 1955
rect 4344 1912 4396 1921
rect 6000 1912 6052 1964
rect 6368 1912 6420 1964
rect 7656 2091 7708 2100
rect 7656 2057 7665 2091
rect 7665 2057 7699 2091
rect 7699 2057 7708 2091
rect 7656 2048 7708 2057
rect 7840 2048 7892 2100
rect 8852 2048 8904 2100
rect 7748 1980 7800 2032
rect 12348 2048 12400 2100
rect 15108 2048 15160 2100
rect 3056 1819 3108 1828
rect 3056 1785 3065 1819
rect 3065 1785 3099 1819
rect 3099 1785 3108 1819
rect 3056 1776 3108 1785
rect 1768 1708 1820 1760
rect 4436 1844 4488 1896
rect 5448 1844 5500 1896
rect 5632 1776 5684 1828
rect 8116 1844 8168 1896
rect 8852 1912 8904 1964
rect 9036 1887 9088 1896
rect 9036 1853 9045 1887
rect 9045 1853 9079 1887
rect 9079 1853 9088 1887
rect 9036 1844 9088 1853
rect 11244 1887 11296 1896
rect 11244 1853 11253 1887
rect 11253 1853 11287 1887
rect 11287 1853 11296 1887
rect 11244 1844 11296 1853
rect 11612 1887 11664 1896
rect 11612 1853 11614 1887
rect 11614 1853 11664 1887
rect 11612 1844 11664 1853
rect 11980 1887 12032 1896
rect 11980 1853 11989 1887
rect 11989 1853 12023 1887
rect 12023 1853 12032 1887
rect 11980 1844 12032 1853
rect 5356 1708 5408 1760
rect 5724 1708 5776 1760
rect 9036 1708 9088 1760
rect 9404 1708 9456 1760
rect 9680 1708 9732 1760
rect 11980 1708 12032 1760
rect 13912 1887 13964 1896
rect 13912 1853 13921 1887
rect 13921 1853 13955 1887
rect 13955 1853 13964 1887
rect 13912 1844 13964 1853
rect 14280 1887 14332 1896
rect 14280 1853 14282 1887
rect 14282 1853 14332 1887
rect 14280 1844 14332 1853
rect 14648 1887 14700 1896
rect 14648 1853 14657 1887
rect 14657 1853 14691 1887
rect 14691 1853 14700 1887
rect 14648 1844 14700 1853
rect 17960 2048 18012 2100
rect 21732 2048 21784 2100
rect 24032 2048 24084 2100
rect 24768 2048 24820 2100
rect 27804 2048 27856 2100
rect 16028 1912 16080 1964
rect 20720 1912 20772 1964
rect 21272 1955 21324 1964
rect 21272 1921 21274 1955
rect 21274 1921 21324 1955
rect 21272 1912 21324 1921
rect 16672 1844 16724 1896
rect 18328 1844 18380 1896
rect 18512 1887 18564 1896
rect 18512 1853 18521 1887
rect 18521 1853 18555 1887
rect 18555 1853 18564 1887
rect 18512 1844 18564 1853
rect 18788 1844 18840 1896
rect 19432 1887 19484 1896
rect 19432 1853 19441 1887
rect 19441 1853 19475 1887
rect 19475 1853 19484 1887
rect 19432 1844 19484 1853
rect 20904 1887 20956 1896
rect 20904 1853 20913 1887
rect 20913 1853 20947 1887
rect 20947 1853 20956 1887
rect 20904 1844 20956 1853
rect 21732 1844 21784 1896
rect 23756 1980 23808 2032
rect 23388 1912 23440 1964
rect 23848 1955 23900 1964
rect 23848 1921 23857 1955
rect 23857 1921 23891 1955
rect 23891 1921 23900 1955
rect 23848 1912 23900 1921
rect 24216 1955 24268 1964
rect 24216 1921 24218 1955
rect 24218 1921 24268 1955
rect 24216 1912 24268 1921
rect 24492 1912 24544 1964
rect 24952 1912 25004 1964
rect 26424 1912 26476 1964
rect 26884 1912 26936 1964
rect 27436 1912 27488 1964
rect 29368 2048 29420 2100
rect 29460 2048 29512 2100
rect 28264 1912 28316 1964
rect 20996 1776 21048 1828
rect 22468 1776 22520 1828
rect 16856 1708 16908 1760
rect 17132 1708 17184 1760
rect 19248 1708 19300 1760
rect 20076 1708 20128 1760
rect 22928 1776 22980 1828
rect 26056 1844 26108 1896
rect 27712 1776 27764 1828
rect 28724 1776 28776 1828
rect 22744 1708 22796 1760
rect 23480 1708 23532 1760
rect 23664 1708 23716 1760
rect 24492 1708 24544 1760
rect 24860 1708 24912 1760
rect 24952 1708 25004 1760
rect 26608 1708 26660 1760
rect 28632 1708 28684 1760
rect 28816 1751 28868 1760
rect 28816 1717 28825 1751
rect 28825 1717 28859 1751
rect 28859 1717 28868 1751
rect 28816 1708 28868 1717
rect 29092 1708 29144 1760
rect 7988 1606 8040 1658
rect 8052 1606 8104 1658
rect 8116 1606 8168 1658
rect 8180 1606 8232 1658
rect 8244 1606 8296 1658
rect 15578 1606 15630 1658
rect 15642 1606 15694 1658
rect 15706 1606 15758 1658
rect 15770 1606 15822 1658
rect 15834 1606 15886 1658
rect 23168 1606 23220 1658
rect 23232 1606 23284 1658
rect 23296 1606 23348 1658
rect 23360 1606 23412 1658
rect 23424 1606 23476 1658
rect 30758 1606 30810 1658
rect 30822 1606 30874 1658
rect 30886 1606 30938 1658
rect 30950 1606 31002 1658
rect 31014 1606 31066 1658
rect 1216 1504 1268 1556
rect 1768 1547 1820 1556
rect 1768 1513 1783 1547
rect 1783 1513 1817 1547
rect 1817 1513 1820 1547
rect 1768 1504 1820 1513
rect 3056 1504 3108 1556
rect 5540 1547 5592 1556
rect 5540 1513 5549 1547
rect 5549 1513 5583 1547
rect 5583 1513 5592 1547
rect 5540 1504 5592 1513
rect 5908 1547 5960 1556
rect 5908 1513 5917 1547
rect 5917 1513 5951 1547
rect 5951 1513 5960 1547
rect 5908 1504 5960 1513
rect 1032 1368 1084 1420
rect 1308 1411 1360 1420
rect 1308 1377 1317 1411
rect 1317 1377 1351 1411
rect 1351 1377 1360 1411
rect 1308 1368 1360 1377
rect 2136 1368 2188 1420
rect 5816 1368 5868 1420
rect 6000 1368 6052 1420
rect 6184 1368 6236 1420
rect 2044 1343 2096 1352
rect 2044 1309 2053 1343
rect 2053 1309 2087 1343
rect 2087 1309 2096 1343
rect 2044 1300 2096 1309
rect 3516 1343 3568 1352
rect 3516 1309 3525 1343
rect 3525 1309 3559 1343
rect 3559 1309 3568 1343
rect 3516 1300 3568 1309
rect 3884 1343 3936 1352
rect 3884 1309 3886 1343
rect 3886 1309 3936 1343
rect 3884 1300 3936 1309
rect 4068 1300 4120 1352
rect 4252 1343 4304 1352
rect 4252 1309 4261 1343
rect 4261 1309 4295 1343
rect 4295 1309 4304 1343
rect 4252 1300 4304 1309
rect 4344 1300 4396 1352
rect 5632 1232 5684 1284
rect 1676 1164 1728 1216
rect 4436 1164 4488 1216
rect 4620 1164 4672 1216
rect 11244 1436 11296 1488
rect 11612 1504 11664 1556
rect 14280 1547 14332 1556
rect 14280 1513 14295 1547
rect 14295 1513 14329 1547
rect 14329 1513 14332 1547
rect 14280 1504 14332 1513
rect 16856 1504 16908 1556
rect 18788 1547 18840 1556
rect 18788 1513 18803 1547
rect 18803 1513 18837 1547
rect 18837 1513 18840 1547
rect 18788 1504 18840 1513
rect 19432 1504 19484 1556
rect 20904 1504 20956 1556
rect 11704 1436 11756 1488
rect 20076 1436 20128 1488
rect 7196 1343 7248 1352
rect 7196 1309 7205 1343
rect 7205 1309 7239 1343
rect 7239 1309 7248 1343
rect 7196 1300 7248 1309
rect 9036 1343 9088 1352
rect 9036 1309 9038 1343
rect 9038 1309 9088 1343
rect 9036 1300 9088 1309
rect 9128 1343 9180 1352
rect 9128 1309 9140 1343
rect 9140 1309 9174 1343
rect 9174 1309 9180 1343
rect 9128 1300 9180 1309
rect 10140 1300 10192 1352
rect 8944 1164 8996 1216
rect 11244 1232 11296 1284
rect 12164 1300 12216 1352
rect 13820 1343 13872 1352
rect 13820 1309 13829 1343
rect 13829 1309 13863 1343
rect 13863 1309 13872 1343
rect 13820 1300 13872 1309
rect 14372 1300 14424 1352
rect 16028 1300 16080 1352
rect 16856 1343 16908 1352
rect 16856 1309 16865 1343
rect 16865 1309 16899 1343
rect 16899 1309 16908 1343
rect 16856 1300 16908 1309
rect 18328 1343 18380 1352
rect 18328 1309 18337 1343
rect 18337 1309 18371 1343
rect 18371 1309 18380 1343
rect 18328 1300 18380 1309
rect 20904 1300 20956 1352
rect 13360 1232 13412 1284
rect 20536 1275 20588 1284
rect 20536 1241 20545 1275
rect 20545 1241 20579 1275
rect 20579 1241 20588 1275
rect 20536 1232 20588 1241
rect 21548 1504 21600 1556
rect 21916 1504 21968 1556
rect 21364 1368 21416 1420
rect 22468 1368 22520 1420
rect 22928 1504 22980 1556
rect 23112 1436 23164 1488
rect 23664 1504 23716 1556
rect 24860 1504 24912 1556
rect 24216 1436 24268 1488
rect 26332 1436 26384 1488
rect 27528 1547 27580 1556
rect 27528 1513 27537 1547
rect 27537 1513 27571 1547
rect 27571 1513 27580 1547
rect 27528 1504 27580 1513
rect 28172 1504 28224 1556
rect 29000 1504 29052 1556
rect 22744 1300 22796 1352
rect 11152 1164 11204 1216
rect 13820 1164 13872 1216
rect 14648 1164 14700 1216
rect 16304 1164 16356 1216
rect 17776 1164 17828 1216
rect 21272 1232 21324 1284
rect 23756 1368 23808 1420
rect 23940 1411 23992 1420
rect 23940 1377 23949 1411
rect 23949 1377 23983 1411
rect 23983 1377 23992 1411
rect 23940 1368 23992 1377
rect 25320 1368 25372 1420
rect 24032 1300 24084 1352
rect 23112 1232 23164 1284
rect 24308 1300 24360 1352
rect 24676 1300 24728 1352
rect 25596 1300 25648 1352
rect 26608 1411 26660 1420
rect 26608 1377 26617 1411
rect 26617 1377 26651 1411
rect 26651 1377 26660 1411
rect 26608 1368 26660 1377
rect 27436 1368 27488 1420
rect 27712 1368 27764 1420
rect 29460 1368 29512 1420
rect 27804 1300 27856 1352
rect 28080 1343 28132 1352
rect 28080 1309 28092 1343
rect 28092 1309 28126 1343
rect 28126 1309 28132 1343
rect 28080 1300 28132 1309
rect 28356 1343 28408 1352
rect 28356 1309 28365 1343
rect 28365 1309 28399 1343
rect 28399 1309 28408 1343
rect 28356 1300 28408 1309
rect 29920 1300 29972 1352
rect 21088 1164 21140 1216
rect 26424 1207 26476 1216
rect 26424 1173 26433 1207
rect 26433 1173 26467 1207
rect 26467 1173 26476 1207
rect 26424 1164 26476 1173
rect 4193 1062 4245 1114
rect 4257 1062 4309 1114
rect 4321 1062 4373 1114
rect 4385 1062 4437 1114
rect 4449 1062 4501 1114
rect 11783 1062 11835 1114
rect 11847 1062 11899 1114
rect 11911 1062 11963 1114
rect 11975 1062 12027 1114
rect 12039 1062 12091 1114
rect 19373 1062 19425 1114
rect 19437 1062 19489 1114
rect 19501 1062 19553 1114
rect 19565 1062 19617 1114
rect 19629 1062 19681 1114
rect 26963 1062 27015 1114
rect 27027 1062 27079 1114
rect 27091 1062 27143 1114
rect 27155 1062 27207 1114
rect 27219 1062 27271 1114
rect 2596 960 2648 1012
rect 2780 1003 2832 1012
rect 2780 969 2789 1003
rect 2789 969 2823 1003
rect 2823 969 2832 1003
rect 2780 960 2832 969
rect 3332 960 3384 1012
rect 4620 960 4672 1012
rect 4988 960 5040 1012
rect 5080 1003 5132 1012
rect 5080 969 5089 1003
rect 5089 969 5123 1003
rect 5123 969 5132 1003
rect 5080 960 5132 969
rect 5172 1003 5224 1012
rect 5172 969 5181 1003
rect 5181 969 5215 1003
rect 5215 969 5224 1003
rect 5172 960 5224 969
rect 4804 892 4856 944
rect 5816 935 5868 944
rect 5816 901 5825 935
rect 5825 901 5859 935
rect 5859 901 5868 935
rect 5816 892 5868 901
rect 940 867 992 876
rect 940 833 949 867
rect 949 833 983 867
rect 983 833 992 867
rect 940 824 992 833
rect 1676 867 1728 876
rect 1676 833 1685 867
rect 1685 833 1719 867
rect 1719 833 1728 867
rect 1676 824 1728 833
rect 1768 824 1820 876
rect 5448 824 5500 876
rect 3056 620 3108 672
rect 3608 756 3660 808
rect 3700 688 3752 740
rect 4252 756 4304 808
rect 4436 756 4488 808
rect 5540 756 5592 808
rect 7288 960 7340 1012
rect 8668 960 8720 1012
rect 10508 1003 10560 1012
rect 10508 969 10517 1003
rect 10517 969 10551 1003
rect 10551 969 10560 1003
rect 10508 960 10560 969
rect 11336 960 11388 1012
rect 12256 960 12308 1012
rect 13176 1003 13228 1012
rect 13176 969 13185 1003
rect 13185 969 13219 1003
rect 13219 969 13228 1003
rect 13176 960 13228 969
rect 14188 960 14240 1012
rect 16672 960 16724 1012
rect 16856 960 16908 1012
rect 20812 1003 20864 1012
rect 20812 969 20821 1003
rect 20821 969 20855 1003
rect 20855 969 20864 1003
rect 20812 960 20864 969
rect 20904 960 20956 1012
rect 21548 960 21600 1012
rect 23020 960 23072 1012
rect 23480 960 23532 1012
rect 10784 892 10836 944
rect 12716 892 12768 944
rect 13728 892 13780 944
rect 16396 892 16448 944
rect 18972 892 19024 944
rect 26424 960 26476 1012
rect 26608 1003 26660 1012
rect 26608 969 26617 1003
rect 26617 969 26651 1003
rect 26651 969 26660 1003
rect 26608 960 26660 969
rect 28540 1003 28592 1012
rect 28540 969 28549 1003
rect 28549 969 28583 1003
rect 28583 969 28592 1003
rect 28540 960 28592 969
rect 29460 1003 29512 1012
rect 29460 969 29469 1003
rect 29469 969 29503 1003
rect 29503 969 29512 1003
rect 29460 960 29512 969
rect 6276 824 6328 876
rect 6644 824 6696 876
rect 6736 824 6788 876
rect 8852 824 8904 876
rect 9220 824 9272 876
rect 6092 799 6144 808
rect 6092 765 6101 799
rect 6101 765 6135 799
rect 6135 765 6144 799
rect 6092 756 6144 765
rect 8300 756 8352 808
rect 9036 799 9088 808
rect 9036 765 9038 799
rect 9038 765 9088 799
rect 11152 824 11204 876
rect 11520 824 11572 876
rect 5908 688 5960 740
rect 8392 688 8444 740
rect 9036 756 9088 765
rect 10784 756 10836 808
rect 11428 756 11480 808
rect 12256 799 12308 808
rect 12256 765 12265 799
rect 12265 765 12299 799
rect 12299 765 12308 799
rect 12256 756 12308 765
rect 12440 756 12492 808
rect 13360 799 13412 808
rect 13360 765 13369 799
rect 13369 765 13403 799
rect 13403 765 13412 799
rect 13360 756 13412 765
rect 13544 756 13596 808
rect 14280 824 14332 876
rect 17132 867 17184 876
rect 17132 833 17141 867
rect 17141 833 17175 867
rect 17175 833 17184 867
rect 17132 824 17184 833
rect 17868 824 17920 876
rect 19340 867 19392 876
rect 19340 833 19342 867
rect 19342 833 19392 867
rect 19340 824 19392 833
rect 14464 756 14516 808
rect 14556 799 14608 808
rect 14556 765 14565 799
rect 14565 765 14599 799
rect 14599 765 14608 799
rect 14556 756 14608 765
rect 16304 799 16356 808
rect 16304 765 16313 799
rect 16313 765 16347 799
rect 16347 765 16356 799
rect 16304 756 16356 765
rect 16396 799 16448 808
rect 16396 765 16405 799
rect 16405 765 16439 799
rect 16439 765 16448 799
rect 16396 756 16448 765
rect 10968 688 11020 740
rect 12164 688 12216 740
rect 19708 867 19760 876
rect 19708 833 19717 867
rect 19717 833 19751 867
rect 19751 833 19760 867
rect 19708 824 19760 833
rect 21364 824 21416 876
rect 4712 620 4764 672
rect 10784 620 10836 672
rect 11152 620 11204 672
rect 12808 663 12860 672
rect 12808 629 12817 663
rect 12817 629 12851 663
rect 12851 629 12860 663
rect 12808 620 12860 629
rect 15292 620 15344 672
rect 16764 620 16816 672
rect 17868 620 17920 672
rect 19064 688 19116 740
rect 21548 688 21600 740
rect 22192 824 22244 876
rect 26700 892 26752 944
rect 23848 867 23900 876
rect 23848 833 23857 867
rect 23857 833 23891 867
rect 23891 833 23900 867
rect 23848 824 23900 833
rect 24308 867 24360 876
rect 24308 833 24320 867
rect 24320 833 24354 867
rect 24354 833 24360 867
rect 24308 824 24360 833
rect 23848 688 23900 740
rect 24400 756 24452 808
rect 25228 824 25280 876
rect 27344 824 27396 876
rect 29276 824 29328 876
rect 26516 756 26568 808
rect 28632 756 28684 808
rect 24124 620 24176 672
rect 25688 663 25740 672
rect 25688 629 25697 663
rect 25697 629 25731 663
rect 25731 629 25740 663
rect 25688 620 25740 629
rect 26056 663 26108 672
rect 26056 629 26065 663
rect 26065 629 26099 663
rect 26099 629 26108 663
rect 26056 620 26108 629
rect 26240 620 26292 672
rect 27804 620 27856 672
rect 29184 663 29236 672
rect 29184 629 29193 663
rect 29193 629 29227 663
rect 29227 629 29236 663
rect 29184 620 29236 629
rect 7988 518 8040 570
rect 8052 518 8104 570
rect 8116 518 8168 570
rect 8180 518 8232 570
rect 8244 518 8296 570
rect 15578 518 15630 570
rect 15642 518 15694 570
rect 15706 518 15758 570
rect 15770 518 15822 570
rect 15834 518 15886 570
rect 23168 518 23220 570
rect 23232 518 23284 570
rect 23296 518 23348 570
rect 23360 518 23412 570
rect 23424 518 23476 570
rect 30758 518 30810 570
rect 30822 518 30874 570
rect 30886 518 30938 570
rect 30950 518 31002 570
rect 31014 518 31066 570
rect 3056 416 3108 468
rect 5724 416 5776 468
rect 5816 416 5868 468
rect 14372 416 14424 468
rect 14556 416 14608 468
rect 26056 416 26108 468
rect 3516 348 3568 400
rect 8392 348 8444 400
rect 3884 280 3936 332
rect 9036 280 9088 332
rect 12808 348 12860 400
rect 19064 348 19116 400
rect 24492 348 24544 400
rect 25688 348 25740 400
rect 11520 280 11572 332
rect 14280 280 14332 332
rect 11336 212 11388 264
rect 12716 212 12768 264
rect 15568 212 15620 264
rect 1308 144 1360 196
rect 6092 144 6144 196
rect 12256 144 12308 196
rect 14464 144 14516 196
rect 24032 212 24084 264
rect 17868 144 17920 196
rect 26240 144 26292 196
rect 5540 8 5592 60
rect 12440 8 12492 60
rect 15476 76 15528 128
rect 16396 8 16448 60
<< metal2 >>
rect 7656 22296 7708 22302
rect 7656 22238 7708 22244
rect 7748 22296 7800 22302
rect 14924 22296 14976 22302
rect 7748 22238 7800 22244
rect 9126 22264 9182 22273
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 1768 22160 1820 22166
rect 1768 22102 1820 22108
rect 1676 21888 1728 21894
rect 1676 21830 1728 21836
rect 1688 21486 1716 21830
rect 1216 21480 1268 21486
rect 1216 21422 1268 21428
rect 1676 21480 1728 21486
rect 1676 21422 1728 21428
rect 756 20936 808 20942
rect 756 20878 808 20884
rect 664 19236 716 19242
rect 664 19178 716 19184
rect 676 11286 704 19178
rect 768 13938 796 20878
rect 848 20800 900 20806
rect 848 20742 900 20748
rect 860 19310 888 20742
rect 1228 19514 1256 21422
rect 1780 21146 1808 22102
rect 3608 22092 3660 22098
rect 3608 22034 3660 22040
rect 1952 22024 2004 22030
rect 1952 21966 2004 21972
rect 2502 21992 2558 22001
rect 1768 21140 1820 21146
rect 1768 21082 1820 21088
rect 1492 20936 1544 20942
rect 1492 20878 1544 20884
rect 1308 20392 1360 20398
rect 1308 20334 1360 20340
rect 1320 19922 1348 20334
rect 1308 19916 1360 19922
rect 1308 19858 1360 19864
rect 1216 19508 1268 19514
rect 1216 19450 1268 19456
rect 1320 19378 1348 19858
rect 1308 19372 1360 19378
rect 1308 19314 1360 19320
rect 848 19304 900 19310
rect 848 19246 900 19252
rect 860 18329 888 19246
rect 1216 18828 1268 18834
rect 1216 18770 1268 18776
rect 1228 18426 1256 18770
rect 1308 18760 1360 18766
rect 1308 18702 1360 18708
rect 1216 18420 1268 18426
rect 1216 18362 1268 18368
rect 846 18320 902 18329
rect 846 18255 902 18264
rect 1320 18170 1348 18702
rect 1228 18142 1348 18170
rect 1228 18086 1256 18142
rect 1216 18080 1268 18086
rect 1216 18022 1268 18028
rect 1228 17542 1256 18022
rect 1308 17876 1360 17882
rect 1308 17818 1360 17824
rect 1216 17536 1268 17542
rect 1216 17478 1268 17484
rect 1228 17202 1256 17478
rect 1216 17196 1268 17202
rect 1216 17138 1268 17144
rect 1216 16788 1268 16794
rect 1216 16730 1268 16736
rect 1032 16584 1084 16590
rect 1032 16526 1084 16532
rect 940 16448 992 16454
rect 940 16390 992 16396
rect 848 15360 900 15366
rect 848 15302 900 15308
rect 756 13932 808 13938
rect 756 13874 808 13880
rect 664 11280 716 11286
rect 664 11222 716 11228
rect 768 8514 796 13874
rect 860 13394 888 15302
rect 952 14618 980 16390
rect 1044 16046 1072 16526
rect 1032 16040 1084 16046
rect 1032 15982 1084 15988
rect 1044 15722 1072 15982
rect 1044 15694 1164 15722
rect 1136 15366 1164 15694
rect 1124 15360 1176 15366
rect 1124 15302 1176 15308
rect 1136 15026 1164 15302
rect 1124 15020 1176 15026
rect 1124 14962 1176 14968
rect 940 14612 992 14618
rect 940 14554 992 14560
rect 1228 14550 1256 16730
rect 1320 15026 1348 17818
rect 1400 15156 1452 15162
rect 1400 15098 1452 15104
rect 1308 15020 1360 15026
rect 1308 14962 1360 14968
rect 1412 14550 1440 15098
rect 1216 14544 1268 14550
rect 1216 14486 1268 14492
rect 1400 14544 1452 14550
rect 1400 14486 1452 14492
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 13410 1440 14350
rect 1320 13394 1440 13410
rect 848 13388 900 13394
rect 848 13330 900 13336
rect 1216 13388 1268 13394
rect 1216 13330 1268 13336
rect 1308 13388 1440 13394
rect 1360 13382 1440 13388
rect 1308 13330 1360 13336
rect 1228 12986 1256 13330
rect 1216 12980 1268 12986
rect 1216 12922 1268 12928
rect 1320 12850 1348 13330
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 1320 12306 1348 12786
rect 1504 12481 1532 20878
rect 1676 20392 1728 20398
rect 1676 20334 1728 20340
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 20058 1624 20198
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1596 19378 1624 19790
rect 1584 19372 1636 19378
rect 1584 19314 1636 19320
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1596 18086 1624 18906
rect 1688 18306 1716 20334
rect 1780 18442 1808 21082
rect 1964 19854 1992 21966
rect 2502 21927 2558 21936
rect 2320 21344 2372 21350
rect 2320 21286 2372 21292
rect 1952 19848 2004 19854
rect 1952 19790 2004 19796
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 1780 18414 1992 18442
rect 1688 18278 1900 18306
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 1584 18080 1636 18086
rect 1688 18057 1716 18158
rect 1768 18080 1820 18086
rect 1584 18022 1636 18028
rect 1674 18048 1730 18057
rect 1768 18022 1820 18028
rect 1674 17983 1730 17992
rect 1780 17882 1808 18022
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1676 17672 1728 17678
rect 1674 17640 1676 17649
rect 1728 17640 1730 17649
rect 1674 17575 1730 17584
rect 1780 16998 1808 17818
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1768 16584 1820 16590
rect 1768 16526 1820 16532
rect 1596 16266 1624 16526
rect 1596 16238 1716 16266
rect 1688 15910 1716 16238
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15502 1716 15846
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1688 14822 1716 15438
rect 1780 14929 1808 16526
rect 1766 14920 1822 14929
rect 1766 14855 1822 14864
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1688 13530 1716 14350
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 12850 1624 13126
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1688 12646 1716 13466
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1490 12472 1546 12481
rect 1490 12407 1546 12416
rect 1688 12306 1716 12582
rect 1308 12300 1360 12306
rect 1308 12242 1360 12248
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 940 11688 992 11694
rect 940 11630 992 11636
rect 848 10600 900 10606
rect 848 10542 900 10548
rect 676 8486 796 8514
rect 676 5778 704 8486
rect 756 8424 808 8430
rect 756 8366 808 8372
rect 768 7342 796 8366
rect 756 7336 808 7342
rect 756 7278 808 7284
rect 768 6934 796 7278
rect 756 6928 808 6934
rect 756 6870 808 6876
rect 768 6254 796 6870
rect 756 6248 808 6254
rect 756 6190 808 6196
rect 664 5772 716 5778
rect 664 5714 716 5720
rect 676 5234 704 5714
rect 664 5228 716 5234
rect 664 5170 716 5176
rect 676 2774 704 5170
rect 768 4604 796 6190
rect 860 4826 888 10542
rect 952 8634 980 11630
rect 1320 11218 1348 12242
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 1412 11354 1440 11834
rect 1688 11778 1716 12242
rect 1780 12238 1808 14214
rect 1872 13977 1900 18278
rect 1964 14634 1992 18414
rect 2056 16561 2084 19790
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2042 16552 2098 16561
rect 2042 16487 2098 16496
rect 2042 15600 2098 15609
rect 2042 15535 2098 15544
rect 2056 15502 2084 15535
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 2148 15065 2176 17138
rect 2134 15056 2190 15065
rect 2134 14991 2190 15000
rect 1964 14606 2084 14634
rect 2240 14618 2268 19314
rect 2332 19145 2360 21286
rect 2412 20936 2464 20942
rect 2412 20878 2464 20884
rect 2318 19136 2374 19145
rect 2318 19071 2374 19080
rect 2332 16794 2360 19071
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 1950 14512 2006 14521
rect 1950 14447 2006 14456
rect 1964 14414 1992 14447
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 2056 14226 2084 14606
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2424 14498 2452 20878
rect 2516 19310 2544 21927
rect 3148 21548 3200 21554
rect 3148 21490 3200 21496
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2688 20800 2740 20806
rect 2688 20742 2740 20748
rect 2504 19304 2556 19310
rect 2504 19246 2556 19252
rect 2504 18760 2556 18766
rect 2504 18702 2556 18708
rect 2516 15473 2544 18702
rect 2700 17354 2728 20742
rect 2792 17649 2820 21422
rect 3056 21412 3108 21418
rect 3056 21354 3108 21360
rect 2964 19236 3016 19242
rect 2964 19178 3016 19184
rect 2976 18834 3004 19178
rect 3068 18970 3096 21354
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 2872 18828 2924 18834
rect 2872 18770 2924 18776
rect 2964 18828 3016 18834
rect 2964 18770 3016 18776
rect 2778 17640 2834 17649
rect 2778 17575 2834 17584
rect 2700 17326 2820 17354
rect 2792 17082 2820 17326
rect 2608 17054 2820 17082
rect 2502 15464 2558 15473
rect 2502 15399 2558 15408
rect 2424 14470 2544 14498
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 1964 14198 2084 14226
rect 1858 13968 1914 13977
rect 1858 13903 1914 13912
rect 1964 13734 1992 14198
rect 2148 14090 2176 14350
rect 2056 14062 2176 14090
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 12434 1992 13670
rect 1872 12406 1992 12434
rect 1768 12232 1820 12238
rect 1768 12174 1820 12180
rect 1688 11750 1808 11778
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1308 11212 1360 11218
rect 1308 11154 1360 11160
rect 1320 10674 1348 11154
rect 1688 11014 1716 11630
rect 1780 11354 1808 11750
rect 1872 11506 1900 12406
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1964 12102 1992 12174
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 2056 11762 2084 14062
rect 2228 13320 2280 13326
rect 2226 13288 2228 13297
rect 2280 13288 2282 13297
rect 2226 13223 2282 13232
rect 2320 12776 2372 12782
rect 2240 12736 2320 12764
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 1872 11478 2084 11506
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 1320 10062 1348 10610
rect 1780 10470 1808 11290
rect 1950 11248 2006 11257
rect 1950 11183 2006 11192
rect 1964 11150 1992 11183
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 2056 10554 2084 11478
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2148 11218 2176 11290
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 1872 10526 2084 10554
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1780 10266 1808 10406
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1308 10056 1360 10062
rect 1308 9998 1360 10004
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1320 9586 1348 9998
rect 1412 9722 1440 9998
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1308 9580 1360 9586
rect 1308 9522 1360 9528
rect 1032 9512 1084 9518
rect 1032 9454 1084 9460
rect 940 8628 992 8634
rect 940 8570 992 8576
rect 940 6656 992 6662
rect 940 6598 992 6604
rect 848 4820 900 4826
rect 848 4762 900 4768
rect 848 4616 900 4622
rect 768 4576 848 4604
rect 848 4558 900 4564
rect 860 4146 888 4558
rect 952 4486 980 6598
rect 1044 5914 1072 9454
rect 1320 9178 1348 9522
rect 1308 9172 1360 9178
rect 1308 9114 1360 9120
rect 1308 7812 1360 7818
rect 1308 7754 1360 7760
rect 1124 7744 1176 7750
rect 1124 7686 1176 7692
rect 1136 7410 1164 7686
rect 1124 7404 1176 7410
rect 1124 7346 1176 7352
rect 1216 6656 1268 6662
rect 1216 6598 1268 6604
rect 1228 6458 1256 6598
rect 1216 6452 1268 6458
rect 1216 6394 1268 6400
rect 1032 5908 1084 5914
rect 1032 5850 1084 5856
rect 1320 5352 1348 7754
rect 1412 6866 1440 9658
rect 1780 9382 1808 10202
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1780 9042 1808 9318
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 1768 8900 1820 8906
rect 1768 8842 1820 8848
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1688 8430 1716 8774
rect 1584 8424 1636 8430
rect 1504 8384 1584 8412
rect 1504 7886 1532 8384
rect 1584 8366 1636 8372
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1780 7954 1808 8842
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1768 7948 1820 7954
rect 1768 7890 1820 7896
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1504 7206 1532 7822
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1398 6760 1454 6769
rect 1398 6695 1454 6704
rect 1412 5778 1440 6695
rect 1504 6236 1532 7142
rect 1596 7041 1624 7890
rect 1780 7206 1808 7890
rect 1768 7200 1820 7206
rect 1688 7160 1768 7188
rect 1582 7032 1638 7041
rect 1582 6967 1638 6976
rect 1688 6798 1716 7160
rect 1768 7142 1820 7148
rect 1768 6928 1820 6934
rect 1872 6916 1900 10526
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 2056 9722 2084 10406
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1964 9110 1992 9318
rect 1952 9104 2004 9110
rect 1952 9046 2004 9052
rect 1952 8900 2004 8906
rect 1952 8842 2004 8848
rect 1820 6888 1900 6916
rect 1768 6870 1820 6876
rect 1780 6854 1814 6870
rect 1676 6792 1728 6798
rect 1786 6780 1814 6854
rect 1676 6734 1728 6740
rect 1780 6752 1814 6780
rect 1584 6248 1636 6254
rect 1504 6208 1584 6236
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1136 5324 1348 5352
rect 940 4480 992 4486
rect 940 4422 992 4428
rect 848 4140 900 4146
rect 848 4082 900 4088
rect 938 3904 994 3913
rect 938 3839 994 3848
rect 676 2746 796 2774
rect 768 2514 796 2746
rect 952 2650 980 3839
rect 1032 3528 1084 3534
rect 1032 3470 1084 3476
rect 940 2644 992 2650
rect 940 2586 992 2592
rect 756 2508 808 2514
rect 756 2450 808 2456
rect 1044 2088 1072 3470
rect 1136 2774 1164 5324
rect 1504 4622 1532 6208
rect 1584 6190 1636 6196
rect 1780 5914 1808 6752
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1582 5808 1638 5817
rect 1582 5743 1638 5752
rect 1492 4616 1544 4622
rect 1492 4558 1544 4564
rect 1308 4140 1360 4146
rect 1308 4082 1360 4088
rect 1320 4049 1348 4082
rect 1306 4040 1362 4049
rect 1306 3975 1362 3984
rect 1504 3942 1532 4558
rect 1596 4146 1624 5743
rect 1674 5672 1730 5681
rect 1674 5607 1730 5616
rect 1688 5166 1716 5607
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1596 2990 1624 3878
rect 1688 3602 1716 4082
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 1136 2746 1256 2774
rect 1124 2100 1176 2106
rect 1044 2060 1124 2088
rect 938 1728 994 1737
rect 938 1663 994 1672
rect 952 882 980 1663
rect 1044 1426 1072 2060
rect 1124 2042 1176 2048
rect 1228 1562 1256 2746
rect 1780 2650 1808 4966
rect 1872 4468 1900 6666
rect 1964 4826 1992 8842
rect 2240 8090 2268 12736
rect 2320 12718 2372 12724
rect 2318 10024 2374 10033
rect 2318 9959 2374 9968
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2044 8016 2096 8022
rect 2044 7958 2096 7964
rect 2056 7342 2084 7958
rect 2226 7848 2282 7857
rect 2226 7783 2282 7792
rect 2044 7336 2096 7342
rect 2044 7278 2096 7284
rect 2056 6934 2084 7278
rect 2044 6928 2096 6934
rect 2044 6870 2096 6876
rect 2134 6352 2190 6361
rect 2134 6287 2136 6296
rect 2188 6287 2190 6296
rect 2136 6258 2188 6264
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 2148 5914 2176 6054
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2042 5128 2098 5137
rect 2042 5063 2098 5072
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 2056 4622 2084 5063
rect 2148 5030 2176 5850
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 1872 4440 2084 4468
rect 2056 2774 2084 4440
rect 2134 4176 2190 4185
rect 2134 4111 2190 4120
rect 2148 2990 2176 4111
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 2056 2746 2176 2774
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1688 2310 1716 2382
rect 2148 2310 2176 2746
rect 1676 2304 1728 2310
rect 1676 2246 1728 2252
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 1308 1896 1360 1902
rect 1308 1838 1360 1844
rect 1216 1556 1268 1562
rect 1216 1498 1268 1504
rect 1320 1426 1348 1838
rect 1688 1442 1716 2246
rect 2240 2122 2268 7783
rect 2056 2094 2268 2122
rect 1766 1864 1822 1873
rect 1766 1799 1822 1808
rect 1780 1766 1808 1799
rect 1768 1760 1820 1766
rect 1768 1702 1820 1708
rect 1780 1562 1808 1702
rect 1768 1556 1820 1562
rect 1768 1498 1820 1504
rect 1032 1420 1084 1426
rect 1032 1362 1084 1368
rect 1308 1420 1360 1426
rect 1688 1414 1808 1442
rect 1308 1362 1360 1368
rect 940 876 992 882
rect 940 818 992 824
rect 1320 202 1348 1362
rect 1676 1216 1728 1222
rect 1676 1158 1728 1164
rect 1688 882 1716 1158
rect 1780 882 1808 1414
rect 2056 1358 2084 2094
rect 2136 1420 2188 1426
rect 2332 1408 2360 9959
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2424 8566 2452 8978
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2516 8514 2544 14470
rect 2608 14414 2636 17054
rect 2778 16824 2834 16833
rect 2778 16759 2834 16768
rect 2792 15042 2820 16759
rect 2884 15162 2912 18770
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2976 16250 3004 17070
rect 3068 16794 3096 18226
rect 3160 17882 3188 21490
rect 3514 21040 3570 21049
rect 3514 20975 3570 20984
rect 3528 20534 3556 20975
rect 3516 20528 3568 20534
rect 3516 20470 3568 20476
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 3344 20058 3372 20198
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 3620 19990 3648 22034
rect 3976 21956 4028 21962
rect 3976 21898 4028 21904
rect 3988 20942 4016 21898
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 4193 21788 4501 21797
rect 4193 21786 4199 21788
rect 4255 21786 4279 21788
rect 4335 21786 4359 21788
rect 4415 21786 4439 21788
rect 4495 21786 4501 21788
rect 4255 21734 4257 21786
rect 4437 21734 4439 21786
rect 4193 21732 4199 21734
rect 4255 21732 4279 21734
rect 4335 21732 4359 21734
rect 4415 21732 4439 21734
rect 4495 21732 4501 21734
rect 4193 21723 4501 21732
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 4080 21185 4108 21490
rect 4066 21176 4122 21185
rect 4066 21111 4122 21120
rect 3700 20936 3752 20942
rect 3700 20878 3752 20884
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 4252 20936 4304 20942
rect 4304 20896 4844 20924
rect 4252 20878 4304 20884
rect 3712 20534 3740 20878
rect 4712 20800 4764 20806
rect 4618 20768 4674 20777
rect 4712 20742 4764 20748
rect 4193 20700 4501 20709
rect 4618 20703 4674 20712
rect 4193 20698 4199 20700
rect 4255 20698 4279 20700
rect 4335 20698 4359 20700
rect 4415 20698 4439 20700
rect 4495 20698 4501 20700
rect 4255 20646 4257 20698
rect 4437 20646 4439 20698
rect 4193 20644 4199 20646
rect 4255 20644 4279 20646
rect 4335 20644 4359 20646
rect 4415 20644 4439 20646
rect 4495 20644 4501 20646
rect 4193 20635 4501 20644
rect 3700 20528 3752 20534
rect 3700 20470 3752 20476
rect 4526 20496 4582 20505
rect 4526 20431 4582 20440
rect 3792 20392 3844 20398
rect 3792 20334 3844 20340
rect 3608 19984 3660 19990
rect 3422 19952 3478 19961
rect 3608 19926 3660 19932
rect 3422 19887 3478 19896
rect 3700 19916 3752 19922
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3252 18970 3280 19110
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3148 17740 3200 17746
rect 3148 17682 3200 17688
rect 3056 16788 3108 16794
rect 3056 16730 3108 16736
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 3054 16144 3110 16153
rect 2976 16102 3054 16130
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2792 15014 2912 15042
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2608 9722 2636 13806
rect 2596 9716 2648 9722
rect 2596 9658 2648 9664
rect 2792 8634 2820 13874
rect 2884 11898 2912 15014
rect 2976 12782 3004 16102
rect 3054 16079 3110 16088
rect 3054 15872 3110 15881
rect 3054 15807 3110 15816
rect 3068 15026 3096 15807
rect 3160 15706 3188 17682
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2884 9178 2912 11494
rect 2962 10704 3018 10713
rect 2962 10639 3018 10648
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2780 8628 2832 8634
rect 2884 8616 2912 9114
rect 2976 8974 3004 10639
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2884 8588 3004 8616
rect 2780 8570 2832 8576
rect 2516 8486 2912 8514
rect 2976 8498 3004 8588
rect 3068 8498 3096 13806
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 12442 3188 13126
rect 3252 12442 3280 17614
rect 3344 17320 3372 19790
rect 3436 18902 3464 19887
rect 3700 19858 3752 19864
rect 3606 19816 3662 19825
rect 3606 19751 3662 19760
rect 3424 18896 3476 18902
rect 3424 18838 3476 18844
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3436 17882 3464 18566
rect 3620 18426 3648 19751
rect 3712 18766 3740 19858
rect 3804 19514 3832 20334
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 3896 19922 3924 20198
rect 3884 19916 3936 19922
rect 3884 19858 3936 19864
rect 4448 19802 4476 20198
rect 4540 19990 4568 20431
rect 4528 19984 4580 19990
rect 4528 19926 4580 19932
rect 4448 19774 4568 19802
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 3792 19508 3844 19514
rect 3792 19450 3844 19456
rect 3792 19372 3844 19378
rect 3792 19314 3844 19320
rect 3700 18760 3752 18766
rect 3700 18702 3752 18708
rect 3712 18426 3740 18702
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3608 18216 3660 18222
rect 3608 18158 3660 18164
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3620 17762 3648 18158
rect 3700 18080 3752 18086
rect 3700 18022 3752 18028
rect 3712 17785 3740 18022
rect 3528 17746 3648 17762
rect 3516 17740 3648 17746
rect 3568 17734 3648 17740
rect 3698 17776 3754 17785
rect 3698 17711 3754 17720
rect 3516 17682 3568 17688
rect 3344 17292 3464 17320
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3344 16794 3372 17138
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3344 15978 3372 16730
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 3332 14272 3384 14278
rect 3436 14260 3464 17292
rect 3528 17202 3556 17682
rect 3804 17241 3832 19314
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3988 18193 4016 19246
rect 4080 18873 4108 19654
rect 4193 19612 4501 19621
rect 4193 19610 4199 19612
rect 4255 19610 4279 19612
rect 4335 19610 4359 19612
rect 4415 19610 4439 19612
rect 4495 19610 4501 19612
rect 4255 19558 4257 19610
rect 4437 19558 4439 19610
rect 4193 19556 4199 19558
rect 4255 19556 4279 19558
rect 4335 19556 4359 19558
rect 4415 19556 4439 19558
rect 4495 19556 4501 19558
rect 4193 19547 4501 19556
rect 4066 18864 4122 18873
rect 4066 18799 4122 18808
rect 4193 18524 4501 18533
rect 4193 18522 4199 18524
rect 4255 18522 4279 18524
rect 4335 18522 4359 18524
rect 4415 18522 4439 18524
rect 4495 18522 4501 18524
rect 4255 18470 4257 18522
rect 4437 18470 4439 18522
rect 4193 18468 4199 18470
rect 4255 18468 4279 18470
rect 4335 18468 4359 18470
rect 4415 18468 4439 18470
rect 4495 18468 4501 18470
rect 4193 18459 4501 18468
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 3974 18184 4030 18193
rect 4264 18170 4292 18226
rect 4540 18222 4568 19774
rect 4528 18216 4580 18222
rect 4264 18142 4476 18170
rect 4528 18158 4580 18164
rect 3974 18119 4030 18128
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 4448 18034 4476 18142
rect 4632 18034 4660 20703
rect 4724 19990 4752 20742
rect 4712 19984 4764 19990
rect 4712 19926 4764 19932
rect 4816 19334 4844 20896
rect 4896 20392 4948 20398
rect 4894 20360 4896 20369
rect 4948 20360 4950 20369
rect 4894 20295 4950 20304
rect 5000 19802 5028 21830
rect 5368 21554 5396 22170
rect 5356 21548 5408 21554
rect 5356 21490 5408 21496
rect 5264 21480 5316 21486
rect 5264 21422 5316 21428
rect 5276 21078 5304 21422
rect 5356 21412 5408 21418
rect 5356 21354 5408 21360
rect 5264 21072 5316 21078
rect 5184 21032 5264 21060
rect 5078 20632 5134 20641
rect 5078 20567 5134 20576
rect 5092 19990 5120 20567
rect 5080 19984 5132 19990
rect 5080 19926 5132 19932
rect 5000 19774 5120 19802
rect 4816 19306 4936 19334
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 3896 17678 3924 18022
rect 4448 18006 4660 18034
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3790 17232 3846 17241
rect 3516 17196 3568 17202
rect 3790 17167 3846 17176
rect 3516 17138 3568 17144
rect 3896 17116 3924 17614
rect 4193 17436 4501 17445
rect 4193 17434 4199 17436
rect 4255 17434 4279 17436
rect 4335 17434 4359 17436
rect 4415 17434 4439 17436
rect 4495 17434 4501 17436
rect 4255 17382 4257 17434
rect 4437 17382 4439 17434
rect 4193 17380 4199 17382
rect 4255 17380 4279 17382
rect 4335 17380 4359 17382
rect 4415 17380 4439 17382
rect 4495 17380 4501 17382
rect 4193 17371 4501 17380
rect 3976 17128 4028 17134
rect 3896 17088 3976 17116
rect 3896 16998 3924 17088
rect 3976 17070 4028 17076
rect 4528 17128 4580 17134
rect 4528 17070 4580 17076
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 4540 16776 4568 17070
rect 4724 16946 4752 18158
rect 4724 16918 4844 16946
rect 4540 16748 4752 16776
rect 3608 16652 3660 16658
rect 3608 16594 3660 16600
rect 4528 16652 4580 16658
rect 4528 16594 4580 16600
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3528 15502 3556 15846
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 3620 14550 3648 16594
rect 3700 16584 3752 16590
rect 3700 16526 3752 16532
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 3712 16046 3740 16526
rect 3700 16040 3752 16046
rect 3700 15982 3752 15988
rect 3712 15910 3740 15982
rect 3896 15910 3924 16526
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 15502 3924 15846
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 15026 3832 15302
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3896 14958 3924 15438
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 3988 14634 4016 15438
rect 4080 14822 4108 16526
rect 4193 16348 4501 16357
rect 4193 16346 4199 16348
rect 4255 16346 4279 16348
rect 4335 16346 4359 16348
rect 4415 16346 4439 16348
rect 4495 16346 4501 16348
rect 4255 16294 4257 16346
rect 4437 16294 4439 16346
rect 4193 16292 4199 16294
rect 4255 16292 4279 16294
rect 4335 16292 4359 16294
rect 4415 16292 4439 16294
rect 4495 16292 4501 16294
rect 4193 16283 4501 16292
rect 4436 16040 4488 16046
rect 4436 15982 4488 15988
rect 4448 15910 4476 15982
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 4193 15260 4501 15269
rect 4193 15258 4199 15260
rect 4255 15258 4279 15260
rect 4335 15258 4359 15260
rect 4415 15258 4439 15260
rect 4495 15258 4501 15260
rect 4255 15206 4257 15258
rect 4437 15206 4439 15258
rect 4193 15204 4199 15206
rect 4255 15204 4279 15206
rect 4335 15204 4359 15206
rect 4415 15204 4439 15206
rect 4495 15204 4501 15206
rect 4193 15195 4501 15204
rect 4540 15042 4568 16594
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4448 15014 4568 15042
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 3792 14612 3844 14618
rect 3988 14606 4108 14634
rect 4448 14618 4476 15014
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4540 14618 4568 14894
rect 3792 14554 3844 14560
rect 3608 14544 3660 14550
rect 3608 14486 3660 14492
rect 3384 14232 3464 14260
rect 3516 14272 3568 14278
rect 3332 14214 3384 14220
rect 3516 14214 3568 14220
rect 3528 14074 3556 14214
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3698 13968 3754 13977
rect 3620 13926 3698 13954
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3252 11694 3280 12174
rect 3344 12170 3372 13670
rect 3436 13530 3464 13806
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3436 13002 3464 13466
rect 3528 13190 3556 13806
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3436 12974 3556 13002
rect 3424 12912 3476 12918
rect 3422 12880 3424 12889
rect 3476 12880 3478 12889
rect 3422 12815 3478 12824
rect 3424 12776 3476 12782
rect 3422 12744 3424 12753
rect 3476 12744 3478 12753
rect 3422 12679 3478 12688
rect 3528 12646 3556 12974
rect 3620 12782 3648 13926
rect 3698 13903 3754 13912
rect 3804 13734 3832 14554
rect 3700 13728 3752 13734
rect 3700 13670 3752 13676
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3528 12238 3556 12582
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3332 12164 3384 12170
rect 3332 12106 3384 12112
rect 3514 11792 3570 11801
rect 3514 11727 3516 11736
rect 3568 11727 3570 11736
rect 3516 11698 3568 11704
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3252 10606 3280 11630
rect 3620 11354 3648 11630
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3712 11098 3740 13670
rect 3988 13530 4016 13670
rect 4080 13546 4108 14606
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4632 14278 4660 15438
rect 4724 14618 4752 16748
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4816 14346 4844 16918
rect 4908 16153 4936 19306
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 5000 19009 5028 19110
rect 4986 19000 5042 19009
rect 4986 18935 5042 18944
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 5000 16402 5028 18702
rect 5092 18086 5120 19774
rect 5184 19446 5212 21032
rect 5264 21014 5316 21020
rect 5264 20528 5316 20534
rect 5264 20470 5316 20476
rect 5276 20398 5304 20470
rect 5264 20392 5316 20398
rect 5368 20380 5396 21354
rect 5316 20352 5396 20380
rect 5264 20334 5316 20340
rect 5276 19990 5304 20334
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5264 19984 5316 19990
rect 5264 19926 5316 19932
rect 5264 19780 5316 19786
rect 5264 19722 5316 19728
rect 5172 19440 5224 19446
rect 5172 19382 5224 19388
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5184 18630 5212 19246
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 5276 17202 5304 19722
rect 5368 18737 5396 20198
rect 5460 19174 5488 22170
rect 7668 22166 7696 22238
rect 7288 22160 7340 22166
rect 7288 22102 7340 22108
rect 7656 22160 7708 22166
rect 7656 22102 7708 22108
rect 6828 21888 6880 21894
rect 6550 21856 6606 21865
rect 6828 21830 6880 21836
rect 6550 21791 6606 21800
rect 5814 21720 5870 21729
rect 5814 21655 5870 21664
rect 5540 21480 5592 21486
rect 5540 21422 5592 21428
rect 5552 21010 5580 21422
rect 5828 21146 5856 21655
rect 6000 21548 6052 21554
rect 6000 21490 6052 21496
rect 5908 21412 5960 21418
rect 5908 21354 5960 21360
rect 5920 21146 5948 21354
rect 5816 21140 5868 21146
rect 5816 21082 5868 21088
rect 5908 21140 5960 21146
rect 5908 21082 5960 21088
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5552 20262 5580 20946
rect 5828 20913 5856 20946
rect 5814 20904 5870 20913
rect 5814 20839 5870 20848
rect 6012 20602 6040 21490
rect 6564 21486 6592 21791
rect 6552 21480 6604 21486
rect 6552 21422 6604 21428
rect 6460 20936 6512 20942
rect 6458 20904 6460 20913
rect 6736 20936 6788 20942
rect 6512 20904 6514 20913
rect 6458 20839 6514 20848
rect 6642 20904 6698 20913
rect 6736 20878 6788 20884
rect 6642 20839 6698 20848
rect 6000 20596 6052 20602
rect 6000 20538 6052 20544
rect 6000 20392 6052 20398
rect 6460 20392 6512 20398
rect 6000 20334 6052 20340
rect 6090 20360 6146 20369
rect 5540 20256 5592 20262
rect 5908 20256 5960 20262
rect 5592 20216 5764 20244
rect 5540 20198 5592 20204
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 5540 19712 5592 19718
rect 5644 19689 5672 19858
rect 5736 19786 5764 20216
rect 5908 20198 5960 20204
rect 5920 19990 5948 20198
rect 5908 19984 5960 19990
rect 5908 19926 5960 19932
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 5540 19654 5592 19660
rect 5630 19680 5686 19689
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5354 18728 5410 18737
rect 5552 18698 5580 19654
rect 5630 19615 5686 19624
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5644 18902 5672 19314
rect 5736 19174 5764 19722
rect 5828 19553 5856 19858
rect 5814 19544 5870 19553
rect 5814 19479 5870 19488
rect 5816 19440 5868 19446
rect 5920 19428 5948 19926
rect 5868 19400 5948 19428
rect 5816 19382 5868 19388
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5814 19136 5870 19145
rect 5814 19071 5870 19080
rect 5828 18902 5856 19071
rect 5632 18896 5684 18902
rect 5632 18838 5684 18844
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 5540 18692 5592 18698
rect 5354 18663 5410 18672
rect 5460 18652 5540 18680
rect 5460 18222 5488 18652
rect 5540 18634 5592 18640
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5354 18048 5410 18057
rect 5354 17983 5410 17992
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5080 16992 5132 16998
rect 5080 16934 5132 16940
rect 5092 16726 5120 16934
rect 5080 16720 5132 16726
rect 5080 16662 5132 16668
rect 5264 16448 5316 16454
rect 5000 16374 5120 16402
rect 5264 16390 5316 16396
rect 4894 16144 4950 16153
rect 4894 16079 4950 16088
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4908 14346 4936 15982
rect 4988 15700 5040 15706
rect 4988 15642 5040 15648
rect 5000 14482 5028 15642
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4896 14340 4948 14346
rect 4896 14282 4948 14288
rect 5000 14278 5028 14418
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 4193 14172 4501 14181
rect 4193 14170 4199 14172
rect 4255 14170 4279 14172
rect 4335 14170 4359 14172
rect 4415 14170 4439 14172
rect 4495 14170 4501 14172
rect 4255 14118 4257 14170
rect 4437 14118 4439 14170
rect 4193 14116 4199 14118
rect 4255 14116 4279 14118
rect 4335 14116 4359 14118
rect 4415 14116 4439 14118
rect 4495 14116 4501 14118
rect 4193 14107 4501 14116
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4172 13938 4200 14010
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4158 13560 4214 13569
rect 3976 13524 4028 13530
rect 4080 13518 4158 13546
rect 4158 13495 4214 13504
rect 3976 13466 4028 13472
rect 3792 13320 3844 13326
rect 3976 13320 4028 13326
rect 3844 13280 3976 13308
rect 3792 13262 3844 13268
rect 3976 13262 4028 13268
rect 4193 13084 4501 13093
rect 4193 13082 4199 13084
rect 4255 13082 4279 13084
rect 4335 13082 4359 13084
rect 4415 13082 4439 13084
rect 4495 13082 4501 13084
rect 4255 13030 4257 13082
rect 4437 13030 4439 13082
rect 4193 13028 4199 13030
rect 4255 13028 4279 13030
rect 4335 13028 4359 13030
rect 4415 13028 4439 13030
rect 4495 13028 4501 13030
rect 4193 13019 4501 13028
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4264 12850 4292 12922
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4540 12646 4568 13670
rect 5092 13410 5120 16374
rect 5276 14385 5304 16390
rect 5262 14376 5318 14385
rect 5262 14311 5318 14320
rect 5000 13382 5120 13410
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 4540 12442 4568 12582
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 3804 11150 3832 12378
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3896 11354 3924 12174
rect 3988 11558 4016 12378
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4080 12102 4108 12174
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4193 11996 4501 12005
rect 4193 11994 4199 11996
rect 4255 11994 4279 11996
rect 4335 11994 4359 11996
rect 4415 11994 4439 11996
rect 4495 11994 4501 11996
rect 4255 11942 4257 11994
rect 4437 11942 4439 11994
rect 4193 11940 4199 11942
rect 4255 11940 4279 11942
rect 4335 11940 4359 11942
rect 4415 11940 4439 11942
rect 4495 11940 4501 11942
rect 4193 11931 4501 11940
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3988 11286 4016 11494
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 3620 11082 3740 11098
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3608 11076 3740 11082
rect 3660 11070 3740 11076
rect 3608 11018 3660 11024
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3252 10044 3280 10542
rect 3988 10470 4016 11222
rect 4080 11082 4108 11494
rect 4724 11218 4752 11630
rect 5000 11354 5028 13382
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5092 12238 5120 13262
rect 5368 13258 5396 17983
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5460 16153 5488 17614
rect 5552 16794 5580 18226
rect 5644 17814 5672 18226
rect 5736 17814 5764 18362
rect 5908 18080 5960 18086
rect 5908 18022 5960 18028
rect 5632 17808 5684 17814
rect 5632 17750 5684 17756
rect 5724 17808 5776 17814
rect 5724 17750 5776 17756
rect 5814 17776 5870 17785
rect 5814 17711 5816 17720
rect 5868 17711 5870 17720
rect 5816 17682 5868 17688
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5552 16250 5580 16390
rect 5644 16250 5672 17614
rect 5816 17536 5868 17542
rect 5722 17504 5778 17513
rect 5816 17478 5868 17484
rect 5722 17439 5778 17448
rect 5736 17338 5764 17439
rect 5828 17338 5856 17478
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5816 17332 5868 17338
rect 5816 17274 5868 17280
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5632 16244 5684 16250
rect 5632 16186 5684 16192
rect 5446 16144 5502 16153
rect 5446 16079 5502 16088
rect 5736 15502 5764 16934
rect 5920 16776 5948 18022
rect 5828 16748 5948 16776
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5446 15328 5502 15337
rect 5446 15263 5502 15272
rect 5460 14618 5488 15263
rect 5722 15192 5778 15201
rect 5722 15127 5724 15136
rect 5776 15127 5778 15136
rect 5724 15098 5776 15104
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5552 13802 5580 14486
rect 5644 13938 5672 14894
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5644 12442 5672 12786
rect 5736 12442 5764 14214
rect 5828 13954 5856 16748
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 5920 15162 5948 16594
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5920 14113 5948 14418
rect 5906 14104 5962 14113
rect 5906 14039 5962 14048
rect 5828 13926 5948 13954
rect 5816 13864 5868 13870
rect 5816 13806 5868 13812
rect 5828 13530 5856 13806
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5170 12200 5226 12209
rect 5170 12135 5226 12144
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4632 11098 4660 11154
rect 4068 11076 4120 11082
rect 4632 11070 4752 11098
rect 4068 11018 4120 11024
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4193 10908 4501 10917
rect 4193 10906 4199 10908
rect 4255 10906 4279 10908
rect 4335 10906 4359 10908
rect 4415 10906 4439 10908
rect 4495 10906 4501 10908
rect 4255 10854 4257 10906
rect 4437 10854 4439 10906
rect 4193 10852 4199 10854
rect 4255 10852 4279 10854
rect 4335 10852 4359 10854
rect 4415 10852 4439 10854
rect 4495 10852 4501 10854
rect 4193 10843 4501 10852
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4448 10470 4476 10610
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 3988 10266 4016 10406
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3332 10056 3384 10062
rect 3252 10016 3332 10044
rect 3332 9998 3384 10004
rect 3344 9500 3372 9998
rect 3988 9518 4016 10202
rect 4540 10130 4568 10950
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4193 9820 4501 9829
rect 4193 9818 4199 9820
rect 4255 9818 4279 9820
rect 4335 9818 4359 9820
rect 4415 9818 4439 9820
rect 4495 9818 4501 9820
rect 4255 9766 4257 9818
rect 4437 9766 4439 9818
rect 4193 9764 4199 9766
rect 4255 9764 4279 9766
rect 4335 9764 4359 9766
rect 4415 9764 4439 9766
rect 4495 9764 4501 9766
rect 4193 9755 4501 9764
rect 3424 9512 3476 9518
rect 3344 9472 3424 9500
rect 3424 9454 3476 9460
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3436 9382 3464 9454
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 4632 9178 4660 10542
rect 4724 10470 4752 11070
rect 5078 10840 5134 10849
rect 5078 10775 5080 10784
rect 5132 10775 5134 10784
rect 5080 10746 5132 10752
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4724 9586 4752 10406
rect 5184 9602 5212 12135
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5368 10577 5396 11018
rect 5354 10568 5410 10577
rect 5354 10503 5410 10512
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 5092 9574 5212 9602
rect 5092 9450 5120 9574
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 3332 8968 3384 8974
rect 3330 8936 3332 8945
rect 3384 8936 3386 8945
rect 3330 8871 3386 8880
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 4193 8732 4501 8741
rect 4193 8730 4199 8732
rect 4255 8730 4279 8732
rect 4335 8730 4359 8732
rect 4415 8730 4439 8732
rect 4495 8730 4501 8732
rect 4255 8678 4257 8730
rect 4437 8678 4439 8730
rect 4193 8676 4199 8678
rect 4255 8676 4279 8678
rect 4335 8676 4359 8678
rect 4415 8676 4439 8678
rect 4495 8676 4501 8678
rect 4193 8667 4501 8676
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2410 8256 2466 8265
rect 2410 8191 2466 8200
rect 2424 3534 2452 8191
rect 2700 8129 2728 8298
rect 2686 8120 2742 8129
rect 2686 8055 2742 8064
rect 2884 7313 2912 8486
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 3252 8430 3280 8502
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3252 8072 3280 8366
rect 3252 8044 3556 8072
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3252 7750 3280 7890
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7342 3280 7686
rect 3240 7336 3292 7342
rect 2870 7304 2926 7313
rect 3240 7278 3292 7284
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 2870 7239 2926 7248
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 2778 6896 2834 6905
rect 2778 6831 2834 6840
rect 2792 6458 2820 6831
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2502 5944 2558 5953
rect 2502 5879 2558 5888
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2516 1902 2544 5879
rect 2504 1896 2556 1902
rect 2504 1838 2556 1844
rect 2188 1380 2360 1408
rect 2136 1362 2188 1368
rect 2044 1352 2096 1358
rect 2044 1294 2096 1300
rect 2608 1018 2636 6190
rect 2884 5370 2912 6190
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2778 5264 2834 5273
rect 2778 5199 2834 5208
rect 2792 4690 2820 5199
rect 2884 5098 2912 5306
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 3068 4282 3096 7210
rect 3146 7032 3202 7041
rect 3252 7002 3280 7278
rect 3146 6967 3202 6976
rect 3240 6996 3292 7002
rect 3160 4622 3188 6967
rect 3240 6938 3292 6944
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2964 4072 3016 4078
rect 2778 4040 2834 4049
rect 2778 3975 2834 3984
rect 2962 4040 2964 4049
rect 3016 4040 3018 4049
rect 2962 3975 3018 3984
rect 2792 3777 2820 3975
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 3068 3777 3096 3878
rect 2778 3768 2834 3777
rect 2778 3703 2834 3712
rect 3054 3768 3110 3777
rect 3054 3703 3110 3712
rect 3054 2952 3110 2961
rect 3054 2887 3056 2896
rect 3108 2887 3110 2896
rect 3056 2858 3108 2864
rect 3160 2514 3188 4422
rect 3252 3194 3280 6734
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 2780 1964 2832 1970
rect 2780 1906 2832 1912
rect 2792 1018 2820 1906
rect 3056 1828 3108 1834
rect 3056 1770 3108 1776
rect 3068 1562 3096 1770
rect 3056 1556 3108 1562
rect 3056 1498 3108 1504
rect 3344 1018 3372 7278
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3436 5302 3464 6938
rect 3528 5710 3556 8044
rect 3620 6934 3648 8366
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 3608 6928 3660 6934
rect 3976 6928 4028 6934
rect 3608 6870 3660 6876
rect 3882 6896 3938 6905
rect 3976 6870 4028 6876
rect 3882 6831 3938 6840
rect 3896 6798 3924 6831
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 3528 5166 3556 5646
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3424 4616 3476 4622
rect 3422 4584 3424 4593
rect 3476 4584 3478 4593
rect 3422 4519 3478 4528
rect 3436 1442 3464 4519
rect 3528 4486 3556 5102
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3528 3534 3556 4422
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3528 2825 3556 2858
rect 3514 2816 3570 2825
rect 3514 2751 3570 2760
rect 3514 2680 3570 2689
rect 3514 2615 3516 2624
rect 3568 2615 3570 2624
rect 3516 2586 3568 2592
rect 3620 2106 3648 6190
rect 3896 5914 3924 6598
rect 3988 5914 4016 6870
rect 4080 6322 4108 7686
rect 4193 7644 4501 7653
rect 4193 7642 4199 7644
rect 4255 7642 4279 7644
rect 4335 7642 4359 7644
rect 4415 7642 4439 7644
rect 4495 7642 4501 7644
rect 4255 7590 4257 7642
rect 4437 7590 4439 7642
rect 4193 7588 4199 7590
rect 4255 7588 4279 7590
rect 4335 7588 4359 7590
rect 4415 7588 4439 7590
rect 4495 7588 4501 7590
rect 4193 7579 4501 7588
rect 4436 7200 4488 7206
rect 4434 7168 4436 7177
rect 4620 7200 4672 7206
rect 4488 7168 4490 7177
rect 4434 7103 4490 7112
rect 4540 7160 4620 7188
rect 4344 6860 4396 6866
rect 4448 6848 4476 7103
rect 4396 6820 4476 6848
rect 4344 6802 4396 6808
rect 4193 6556 4501 6565
rect 4193 6554 4199 6556
rect 4255 6554 4279 6556
rect 4335 6554 4359 6556
rect 4415 6554 4439 6556
rect 4495 6554 4501 6556
rect 4255 6502 4257 6554
rect 4437 6502 4439 6554
rect 4193 6500 4199 6502
rect 4255 6500 4279 6502
rect 4335 6500 4359 6502
rect 4415 6500 4439 6502
rect 4495 6500 4501 6502
rect 4193 6491 4501 6500
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3988 5658 4016 5850
rect 3896 5630 4016 5658
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3700 5092 3752 5098
rect 3700 5034 3752 5040
rect 3792 5092 3844 5098
rect 3792 5034 3844 5040
rect 3712 4049 3740 5034
rect 3698 4040 3754 4049
rect 3698 3975 3754 3984
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3712 2990 3740 3878
rect 3804 3738 3832 5034
rect 3896 5030 3924 5630
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 4826 3924 4966
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3896 4128 3924 4762
rect 3988 4622 4016 5510
rect 4080 5370 4108 5646
rect 4264 5574 4292 6054
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4193 5468 4501 5477
rect 4193 5466 4199 5468
rect 4255 5466 4279 5468
rect 4335 5466 4359 5468
rect 4415 5466 4439 5468
rect 4495 5466 4501 5468
rect 4255 5414 4257 5466
rect 4437 5414 4439 5466
rect 4193 5412 4199 5414
rect 4255 5412 4279 5414
rect 4335 5412 4359 5414
rect 4415 5412 4439 5414
rect 4495 5412 4501 5414
rect 4193 5403 4501 5412
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4540 5250 4568 7160
rect 4620 7142 4672 7148
rect 4618 7032 4674 7041
rect 4618 6967 4674 6976
rect 4632 6934 4660 6967
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4264 5234 4568 5250
rect 4252 5228 4568 5234
rect 4304 5222 4568 5228
rect 4252 5170 4304 5176
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 4193 4380 4501 4389
rect 4193 4378 4199 4380
rect 4255 4378 4279 4380
rect 4335 4378 4359 4380
rect 4415 4378 4439 4380
rect 4495 4378 4501 4380
rect 4255 4326 4257 4378
rect 4437 4326 4439 4378
rect 4193 4324 4199 4326
rect 4255 4324 4279 4326
rect 4335 4324 4359 4326
rect 4415 4324 4439 4326
rect 4495 4324 4501 4326
rect 4193 4315 4501 4324
rect 3976 4140 4028 4146
rect 3896 4100 3976 4128
rect 3896 3738 3924 4100
rect 3976 4082 4028 4088
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4356 3738 4384 4082
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 3976 3528 4028 3534
rect 4540 3505 4568 4082
rect 4632 3913 4660 5646
rect 4618 3904 4674 3913
rect 4618 3839 4674 3848
rect 3976 3470 4028 3476
rect 4526 3496 4582 3505
rect 3700 2984 3752 2990
rect 3884 2984 3936 2990
rect 3700 2926 3752 2932
rect 3804 2932 3884 2938
rect 3804 2926 3936 2932
rect 3804 2910 3924 2926
rect 3804 2446 3832 2910
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3792 2440 3844 2446
rect 3790 2408 3792 2417
rect 3844 2408 3846 2417
rect 3790 2343 3846 2352
rect 3608 2100 3660 2106
rect 3608 2042 3660 2048
rect 3804 1970 3832 2343
rect 3792 1964 3844 1970
rect 3792 1906 3844 1912
rect 3896 1850 3924 2790
rect 3988 2689 4016 3470
rect 4526 3431 4582 3440
rect 4193 3292 4501 3301
rect 4193 3290 4199 3292
rect 4255 3290 4279 3292
rect 4335 3290 4359 3292
rect 4415 3290 4439 3292
rect 4495 3290 4501 3292
rect 4255 3238 4257 3290
rect 4437 3238 4439 3290
rect 4193 3236 4199 3238
rect 4255 3236 4279 3238
rect 4335 3236 4359 3238
rect 4415 3236 4439 3238
rect 4495 3236 4501 3238
rect 4193 3227 4501 3236
rect 4158 3088 4214 3097
rect 4158 3023 4214 3032
rect 4252 3052 4304 3058
rect 4172 2854 4200 3023
rect 4252 2994 4304 3000
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 3974 2680 4030 2689
rect 4172 2666 4200 2790
rect 4264 2774 4292 2994
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4264 2746 4568 2774
rect 3974 2615 4030 2624
rect 4080 2650 4200 2666
rect 4080 2644 4212 2650
rect 4080 2638 4160 2644
rect 4080 2530 4108 2638
rect 4160 2586 4212 2592
rect 3988 2502 4108 2530
rect 4250 2544 4306 2553
rect 3988 1970 4016 2502
rect 4250 2479 4252 2488
rect 4304 2479 4306 2488
rect 4252 2450 4304 2456
rect 4193 2204 4501 2213
rect 4193 2202 4199 2204
rect 4255 2202 4279 2204
rect 4335 2202 4359 2204
rect 4415 2202 4439 2204
rect 4495 2202 4501 2204
rect 4255 2150 4257 2202
rect 4437 2150 4439 2202
rect 4193 2148 4199 2150
rect 4255 2148 4279 2150
rect 4335 2148 4359 2150
rect 4415 2148 4439 2150
rect 4495 2148 4501 2150
rect 4193 2139 4501 2148
rect 4540 2106 4568 2746
rect 4528 2100 4580 2106
rect 4528 2042 4580 2048
rect 4342 2000 4398 2009
rect 3976 1964 4028 1970
rect 3976 1906 4028 1912
rect 4068 1964 4120 1970
rect 4342 1935 4344 1944
rect 4068 1906 4120 1912
rect 4396 1935 4398 1944
rect 4344 1906 4396 1912
rect 3804 1822 3924 1850
rect 3606 1456 3662 1465
rect 3436 1414 3606 1442
rect 3606 1391 3662 1400
rect 3516 1352 3568 1358
rect 3516 1294 3568 1300
rect 2596 1012 2648 1018
rect 2596 954 2648 960
rect 2780 1012 2832 1018
rect 2780 954 2832 960
rect 3332 1012 3384 1018
rect 3332 954 3384 960
rect 1676 876 1728 882
rect 1676 818 1728 824
rect 1768 876 1820 882
rect 1768 818 1820 824
rect 3056 672 3108 678
rect 3056 614 3108 620
rect 3068 474 3096 614
rect 3056 468 3108 474
rect 3056 410 3108 416
rect 3528 406 3556 1294
rect 3620 814 3648 1391
rect 3608 808 3660 814
rect 3608 750 3660 756
rect 3700 740 3752 746
rect 3804 728 3832 1822
rect 4080 1442 4108 1906
rect 4436 1896 4488 1902
rect 4436 1838 4488 1844
rect 4448 1737 4476 1838
rect 4434 1728 4490 1737
rect 4632 1714 4660 2926
rect 4434 1663 4490 1672
rect 4540 1686 4660 1714
rect 3988 1414 4108 1442
rect 4250 1456 4306 1465
rect 3884 1352 3936 1358
rect 3884 1294 3936 1300
rect 3752 700 3832 728
rect 3700 682 3752 688
rect 3516 400 3568 406
rect 3516 342 3568 348
rect 3896 338 3924 1294
rect 3884 332 3936 338
rect 3884 274 3936 280
rect 1308 196 1360 202
rect 1308 138 1360 144
rect 3988 105 4016 1414
rect 4434 1456 4490 1465
rect 4306 1414 4384 1442
rect 4250 1391 4306 1400
rect 4356 1358 4384 1414
rect 4434 1391 4490 1400
rect 4068 1352 4120 1358
rect 4252 1352 4304 1358
rect 4068 1294 4120 1300
rect 4250 1320 4252 1329
rect 4344 1352 4396 1358
rect 4304 1320 4306 1329
rect 4080 921 4108 1294
rect 4344 1294 4396 1300
rect 4250 1255 4306 1264
rect 4448 1222 4476 1391
rect 4436 1216 4488 1222
rect 4436 1158 4488 1164
rect 4193 1116 4501 1125
rect 4193 1114 4199 1116
rect 4255 1114 4279 1116
rect 4335 1114 4359 1116
rect 4415 1114 4439 1116
rect 4495 1114 4501 1116
rect 4255 1062 4257 1114
rect 4437 1062 4439 1114
rect 4193 1060 4199 1062
rect 4255 1060 4279 1062
rect 4335 1060 4359 1062
rect 4415 1060 4439 1062
rect 4495 1060 4501 1062
rect 4193 1051 4501 1060
rect 4066 912 4122 921
rect 4066 847 4122 856
rect 4252 808 4304 814
rect 4436 808 4488 814
rect 4304 768 4436 796
rect 4252 750 4304 756
rect 4436 750 4488 756
rect 4540 762 4568 1686
rect 4620 1216 4672 1222
rect 4620 1158 4672 1164
rect 4632 1018 4660 1158
rect 4620 1012 4672 1018
rect 4620 954 4672 960
rect 4618 776 4674 785
rect 4540 734 4618 762
rect 4618 711 4674 720
rect 4724 678 4752 8502
rect 4816 950 4844 8774
rect 4908 3534 4936 8774
rect 5000 5710 5028 8774
rect 5092 7936 5120 8842
rect 5184 8090 5212 9454
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5368 8906 5396 9318
rect 5460 8906 5488 11154
rect 5552 10606 5580 11630
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5722 11520 5778 11529
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5552 10266 5580 10542
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5172 7948 5224 7954
rect 5092 7908 5172 7936
rect 5172 7890 5224 7896
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 5092 7002 5120 7278
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5092 6644 5120 6802
rect 5184 6769 5212 7890
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5276 7410 5304 7754
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5170 6760 5226 6769
rect 5170 6695 5226 6704
rect 5092 6616 5212 6644
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 5000 4457 5028 5510
rect 5092 5234 5120 6054
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4986 4448 5042 4457
rect 4986 4383 5042 4392
rect 4986 3904 5042 3913
rect 4986 3839 5042 3848
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 5000 1018 5028 3839
rect 5078 2816 5134 2825
rect 5184 2802 5212 6616
rect 5276 6254 5304 7346
rect 5368 6780 5396 8842
rect 5552 8498 5580 10202
rect 5644 10130 5672 11494
rect 5722 11455 5778 11464
rect 5736 11218 5764 11455
rect 5828 11218 5856 13330
rect 5920 12442 5948 13926
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 6012 11354 6040 20334
rect 6460 20334 6512 20340
rect 6090 20295 6146 20304
rect 6104 18766 6132 20295
rect 6472 19718 6500 20334
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6472 19334 6500 19654
rect 6288 19306 6500 19334
rect 6184 18828 6236 18834
rect 6184 18770 6236 18776
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 6104 18222 6132 18702
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 6104 17678 6132 18158
rect 6196 18086 6224 18770
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 6104 17134 6132 17614
rect 6196 17134 6224 18022
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 6104 13530 6132 15846
rect 6196 15366 6224 15982
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 6196 14958 6224 15302
rect 6184 14952 6236 14958
rect 6184 14894 6236 14900
rect 6182 14784 6238 14793
rect 6182 14719 6238 14728
rect 6196 14618 6224 14719
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6288 14482 6316 19306
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6380 18426 6408 18702
rect 6458 18456 6514 18465
rect 6368 18420 6420 18426
rect 6458 18391 6514 18400
rect 6368 18362 6420 18368
rect 6472 18170 6500 18391
rect 6380 18142 6500 18170
rect 6279 14476 6331 14482
rect 6196 14436 6279 14464
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6196 13394 6224 14436
rect 6279 14418 6331 14424
rect 6276 14340 6328 14346
rect 6276 14282 6328 14288
rect 6288 13938 6316 14282
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6104 13025 6132 13126
rect 6090 13016 6146 13025
rect 6090 12951 6146 12960
rect 6196 12170 6224 13330
rect 6380 13258 6408 18142
rect 6458 18048 6514 18057
rect 6458 17983 6514 17992
rect 6472 15994 6500 17983
rect 6564 16776 6592 19246
rect 6656 18766 6684 20839
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6748 18465 6776 20878
rect 6840 19922 6868 21830
rect 7300 21622 7328 22102
rect 7760 22030 7788 22238
rect 9126 22199 9182 22208
rect 14370 22264 14426 22273
rect 22284 22296 22336 22302
rect 14924 22238 14976 22244
rect 22282 22264 22284 22273
rect 22376 22296 22428 22302
rect 22336 22264 22338 22273
rect 14370 22199 14372 22208
rect 9034 22128 9090 22137
rect 9034 22063 9090 22072
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 8392 21888 8444 21894
rect 8312 21848 8392 21876
rect 7288 21616 7340 21622
rect 7288 21558 7340 21564
rect 8312 21486 8340 21848
rect 8392 21830 8444 21836
rect 8666 21720 8722 21729
rect 8576 21684 8628 21690
rect 8666 21655 8722 21664
rect 8576 21626 8628 21632
rect 7196 21480 7248 21486
rect 7010 21448 7066 21457
rect 7196 21422 7248 21428
rect 8300 21480 8352 21486
rect 8300 21422 8352 21428
rect 7010 21383 7066 21392
rect 7024 19922 7052 21383
rect 7102 21176 7158 21185
rect 7102 21111 7158 21120
rect 7116 20602 7144 21111
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 7012 19916 7064 19922
rect 7012 19858 7064 19864
rect 7208 19825 7236 21422
rect 8392 21412 8444 21418
rect 8392 21354 8444 21360
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7840 21344 7892 21350
rect 8404 21321 8432 21354
rect 7840 21286 7892 21292
rect 8390 21312 8446 21321
rect 7194 19816 7250 19825
rect 7194 19751 7250 19760
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 6918 19000 6974 19009
rect 6918 18935 6974 18944
rect 6734 18456 6790 18465
rect 6932 18426 6960 18935
rect 6734 18391 6790 18400
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6748 17746 6776 18022
rect 6736 17740 6788 17746
rect 6736 17682 6788 17688
rect 6644 17672 6696 17678
rect 6840 17626 6868 18022
rect 6696 17620 6868 17626
rect 6644 17614 6868 17620
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 6656 17598 6868 17614
rect 6826 17368 6882 17377
rect 6826 17303 6882 17312
rect 6840 17202 6868 17303
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6840 17105 6868 17138
rect 6826 17096 6882 17105
rect 6826 17031 6882 17040
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6564 16748 6684 16776
rect 6550 16688 6606 16697
rect 6550 16623 6552 16632
rect 6604 16623 6606 16632
rect 6552 16594 6604 16600
rect 6472 15966 6592 15994
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6472 15638 6500 15846
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 6472 14958 6500 15574
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6472 13938 6500 14894
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 6472 13394 6500 13670
rect 6564 13433 6592 15966
rect 6656 14550 6684 16748
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6840 15337 6868 15982
rect 6826 15328 6882 15337
rect 6826 15263 6882 15272
rect 6932 14958 6960 16934
rect 7024 16794 7052 17614
rect 7104 17128 7156 17134
rect 7102 17096 7104 17105
rect 7156 17096 7158 17105
rect 7102 17031 7158 17040
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 7104 16040 7156 16046
rect 7010 16008 7066 16017
rect 7104 15982 7156 15988
rect 7010 15943 7066 15952
rect 7024 15337 7052 15943
rect 7116 15881 7144 15982
rect 7102 15872 7158 15881
rect 7102 15807 7158 15816
rect 7208 15586 7236 19246
rect 7300 16726 7328 21286
rect 7852 21128 7880 21286
rect 7988 21244 8296 21253
rect 8390 21247 8446 21256
rect 7988 21242 7994 21244
rect 8050 21242 8074 21244
rect 8130 21242 8154 21244
rect 8210 21242 8234 21244
rect 8290 21242 8296 21244
rect 8050 21190 8052 21242
rect 8232 21190 8234 21242
rect 7988 21188 7994 21190
rect 8050 21188 8074 21190
rect 8130 21188 8154 21190
rect 8210 21188 8234 21190
rect 8290 21188 8296 21190
rect 7988 21179 8296 21188
rect 8482 21176 8538 21185
rect 7852 21100 8432 21128
rect 8482 21111 8538 21120
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7484 18902 7512 20946
rect 8404 20942 8432 21100
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7564 20324 7616 20330
rect 7564 20266 7616 20272
rect 7472 18896 7524 18902
rect 7472 18838 7524 18844
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7392 17785 7420 18770
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7378 17776 7434 17785
rect 7378 17711 7434 17720
rect 7288 16720 7340 16726
rect 7288 16662 7340 16668
rect 7116 15558 7236 15586
rect 7010 15328 7066 15337
rect 7010 15263 7066 15272
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6644 14544 6696 14550
rect 6644 14486 6696 14492
rect 6748 14498 6776 14894
rect 6840 14618 6868 14894
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6748 14470 6960 14498
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6656 14113 6684 14214
rect 6642 14104 6698 14113
rect 6642 14039 6698 14048
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 6656 13569 6684 13670
rect 6642 13560 6698 13569
rect 6642 13495 6698 13504
rect 6550 13424 6606 13433
rect 6460 13388 6512 13394
rect 6840 13394 6868 14350
rect 6932 13870 6960 14470
rect 7012 14272 7064 14278
rect 7116 14260 7144 15558
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7208 14793 7236 15438
rect 7392 15201 7420 17711
rect 7378 15192 7434 15201
rect 7378 15127 7434 15136
rect 7194 14784 7250 14793
rect 7194 14719 7250 14728
rect 7392 14618 7420 15127
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7064 14232 7144 14260
rect 7012 14214 7064 14220
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 7208 13530 7236 14350
rect 7300 14074 7328 14350
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 6550 13359 6606 13368
rect 6828 13388 6880 13394
rect 6460 13330 6512 13336
rect 6828 13330 6880 13336
rect 6276 13252 6328 13258
rect 6276 13194 6328 13200
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6288 12442 6316 13194
rect 6472 12832 6500 13330
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6748 12850 6776 13194
rect 6380 12804 6500 12832
rect 6736 12844 6788 12850
rect 6380 12753 6408 12804
rect 6736 12786 6788 12792
rect 6644 12776 6696 12782
rect 6366 12744 6422 12753
rect 6366 12679 6422 12688
rect 6472 12724 6644 12730
rect 6840 12730 6868 13330
rect 6696 12724 6868 12730
rect 6472 12702 6868 12724
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6380 12306 6408 12679
rect 6472 12424 6500 12702
rect 6932 12646 6960 13466
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6472 12396 6592 12424
rect 6472 12306 6500 12396
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6104 11898 6132 12038
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5816 11212 5868 11218
rect 5868 11172 5948 11200
rect 5816 11154 5868 11160
rect 5920 10606 5948 11172
rect 6104 10810 6132 11698
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6288 11354 6316 11630
rect 6564 11506 6592 12396
rect 6932 12322 6960 12582
rect 6840 12294 6960 12322
rect 7116 12306 7144 13126
rect 7104 12300 7156 12306
rect 6840 12238 6868 12294
rect 7104 12242 7156 12248
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6656 11694 6684 12174
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6736 11552 6788 11558
rect 6564 11478 6684 11506
rect 6840 11540 6868 12174
rect 6932 11898 6960 12174
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6788 11512 6868 11540
rect 6736 11494 6788 11500
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6656 11150 6684 11478
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6460 11008 6512 11014
rect 6460 10950 6512 10956
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 5828 10198 5856 10542
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 10198 6224 10406
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5460 7002 5488 7346
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5448 6792 5500 6798
rect 5368 6752 5448 6780
rect 5448 6734 5500 6740
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5368 5166 5396 6598
rect 5460 5914 5488 6598
rect 5552 6118 5580 7822
rect 5644 7177 5672 10066
rect 5724 9988 5776 9994
rect 5724 9930 5776 9936
rect 5736 9722 5764 9930
rect 5724 9716 5776 9722
rect 6196 9674 6224 10134
rect 6288 9722 6316 10542
rect 6472 10452 6500 10950
rect 6656 10452 6684 11086
rect 6472 10424 6684 10452
rect 6472 10266 6500 10424
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 6748 10130 6776 11222
rect 6840 11200 6868 11512
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6920 11212 6972 11218
rect 6840 11172 6920 11200
rect 6840 10266 6868 11172
rect 6920 11154 6972 11160
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 5724 9658 5776 9664
rect 6012 9646 6224 9674
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5814 9072 5870 9081
rect 5736 9030 5814 9058
rect 5736 8242 5764 9030
rect 5814 9007 5870 9016
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8498 5856 8774
rect 5920 8498 5948 9386
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 6012 8294 6040 9646
rect 6366 9616 6422 9625
rect 6472 9586 6500 9658
rect 6366 9551 6422 9560
rect 6460 9580 6512 9586
rect 6380 9382 6408 9551
rect 6460 9522 6512 9528
rect 6748 9518 6776 10066
rect 7024 9586 7052 11494
rect 7208 11132 7236 13262
rect 7300 12986 7328 13262
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7484 12306 7512 18158
rect 7576 15201 7604 20266
rect 7668 19446 7696 20742
rect 7748 20528 7800 20534
rect 7748 20470 7800 20476
rect 7656 19440 7708 19446
rect 7656 19382 7708 19388
rect 7654 19000 7710 19009
rect 7654 18935 7710 18944
rect 7668 18680 7696 18935
rect 7760 18834 7788 20470
rect 7852 19922 7880 20878
rect 8496 20777 8524 21111
rect 8588 21010 8616 21626
rect 8680 21486 8708 21655
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 8760 21412 8812 21418
rect 8760 21354 8812 21360
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8576 21004 8628 21010
rect 8576 20946 8628 20952
rect 8482 20768 8538 20777
rect 8482 20703 8538 20712
rect 8680 20618 8708 21082
rect 8772 20924 8800 21354
rect 8944 21344 8996 21350
rect 8864 21321 8944 21332
rect 8850 21312 8944 21321
rect 8906 21304 8944 21312
rect 8944 21286 8996 21292
rect 8850 21247 8906 21256
rect 8852 20936 8904 20942
rect 8772 20896 8852 20924
rect 8852 20878 8904 20884
rect 9048 20618 9076 22063
rect 9140 21554 9168 22199
rect 14424 22199 14426 22208
rect 14372 22170 14424 22176
rect 9956 22160 10008 22166
rect 9956 22102 10008 22108
rect 13176 22160 13228 22166
rect 13176 22102 13228 22108
rect 9494 21856 9550 21865
rect 9494 21791 9550 21800
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 9220 21480 9272 21486
rect 9220 21422 9272 21428
rect 9232 21321 9260 21422
rect 9218 21312 9274 21321
rect 9218 21247 9274 21256
rect 9508 21146 9536 21791
rect 9496 21140 9548 21146
rect 9496 21082 9548 21088
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 9496 20936 9548 20942
rect 9496 20878 9548 20884
rect 8312 20590 8708 20618
rect 8772 20590 9076 20618
rect 8312 20398 8340 20590
rect 8484 20528 8536 20534
rect 8536 20488 8616 20516
rect 8484 20470 8536 20476
rect 8588 20398 8616 20488
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 7988 20156 8296 20165
rect 7988 20154 7994 20156
rect 8050 20154 8074 20156
rect 8130 20154 8154 20156
rect 8210 20154 8234 20156
rect 8290 20154 8296 20156
rect 8050 20102 8052 20154
rect 8232 20102 8234 20154
rect 7988 20100 7994 20102
rect 8050 20100 8074 20102
rect 8130 20100 8154 20102
rect 8210 20100 8234 20102
rect 8290 20100 8296 20102
rect 7988 20091 8296 20100
rect 8404 19972 8432 20334
rect 8128 19944 8432 19972
rect 8576 19984 8628 19990
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 8128 19258 8156 19944
rect 8772 19972 8800 20590
rect 8852 20460 8904 20466
rect 8852 20402 8904 20408
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 9404 20460 9456 20466
rect 9404 20402 9456 20408
rect 8628 19944 8800 19972
rect 8576 19926 8628 19932
rect 8392 19848 8444 19854
rect 8206 19816 8262 19825
rect 8392 19790 8444 19796
rect 8206 19751 8262 19760
rect 8220 19514 8248 19751
rect 8404 19700 8432 19790
rect 8312 19672 8432 19700
rect 8312 19514 8340 19672
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8404 19468 8800 19496
rect 8404 19378 8432 19468
rect 8666 19408 8722 19417
rect 8392 19372 8444 19378
rect 8576 19372 8628 19378
rect 8392 19314 8444 19320
rect 8496 19332 8576 19360
rect 8128 19230 8432 19258
rect 7988 19068 8296 19077
rect 7988 19066 7994 19068
rect 8050 19066 8074 19068
rect 8130 19066 8154 19068
rect 8210 19066 8234 19068
rect 8290 19066 8296 19068
rect 8050 19014 8052 19066
rect 8232 19014 8234 19066
rect 7988 19012 7994 19014
rect 8050 19012 8074 19014
rect 8130 19012 8154 19014
rect 8210 19012 8234 19014
rect 8290 19012 8296 19014
rect 7988 19003 8296 19012
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 8404 18748 8432 19230
rect 8496 19122 8524 19332
rect 8666 19343 8722 19352
rect 8576 19314 8628 19320
rect 8680 19310 8708 19343
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8772 19224 8800 19468
rect 8864 19292 8892 20402
rect 8956 19938 8984 20402
rect 9416 20369 9444 20402
rect 9402 20360 9458 20369
rect 9402 20295 9458 20304
rect 8956 19910 9168 19938
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8956 19417 8984 19790
rect 9140 19718 9168 19910
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9404 19848 9456 19854
rect 9404 19790 9456 19796
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 9048 19530 9076 19654
rect 9048 19502 9168 19530
rect 8942 19408 8998 19417
rect 8942 19343 8998 19352
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 8864 19281 8984 19292
rect 8864 19272 8998 19281
rect 8864 19264 8942 19272
rect 8772 19196 8892 19224
rect 8942 19207 8998 19216
rect 8668 19168 8720 19174
rect 8496 19094 8527 19122
rect 8864 19156 8892 19196
rect 8864 19128 8984 19156
rect 8668 19110 8720 19116
rect 8499 18986 8527 19094
rect 8496 18970 8527 18986
rect 8484 18964 8536 18970
rect 8680 18952 8708 19110
rect 8680 18924 8892 18952
rect 8484 18906 8536 18912
rect 8864 18873 8892 18924
rect 8666 18864 8722 18873
rect 8666 18799 8722 18808
rect 8850 18864 8906 18873
rect 8956 18850 8984 19128
rect 9048 18970 9076 19314
rect 9140 18970 9168 19502
rect 9324 19378 9352 19790
rect 9416 19718 9444 19790
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9312 19372 9364 19378
rect 9312 19314 9364 19320
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 8956 18822 9168 18850
rect 8850 18799 8906 18808
rect 8484 18760 8536 18766
rect 8404 18720 8484 18748
rect 8484 18702 8536 18708
rect 7668 18652 7880 18680
rect 7654 18456 7710 18465
rect 7654 18391 7710 18400
rect 7668 15502 7696 18391
rect 7746 18048 7802 18057
rect 7746 17983 7802 17992
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7562 15192 7618 15201
rect 7562 15127 7618 15136
rect 7562 15056 7618 15065
rect 7562 14991 7618 15000
rect 7576 14890 7604 14991
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7576 11898 7604 14350
rect 7654 13696 7710 13705
rect 7654 13631 7710 13640
rect 7668 13190 7696 13631
rect 7760 13546 7788 17983
rect 7852 15688 7880 18652
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 7988 17980 8296 17989
rect 7988 17978 7994 17980
rect 8050 17978 8074 17980
rect 8130 17978 8154 17980
rect 8210 17978 8234 17980
rect 8290 17978 8296 17980
rect 8050 17926 8052 17978
rect 8232 17926 8234 17978
rect 7988 17924 7994 17926
rect 8050 17924 8074 17926
rect 8130 17924 8154 17926
rect 8210 17924 8234 17926
rect 8290 17924 8296 17926
rect 7988 17915 8296 17924
rect 8206 17776 8262 17785
rect 8206 17711 8262 17720
rect 8220 17678 8248 17711
rect 8208 17672 8260 17678
rect 8208 17614 8260 17620
rect 8404 17610 8432 18226
rect 8496 18222 8524 18702
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8496 17660 8524 18022
rect 8574 17912 8630 17921
rect 8574 17847 8630 17856
rect 8588 17814 8616 17847
rect 8680 17814 8708 18799
rect 8944 18760 8996 18766
rect 8864 18720 8944 18748
rect 8758 18456 8814 18465
rect 8758 18391 8814 18400
rect 8772 17882 8800 18391
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 8576 17808 8628 17814
rect 8576 17750 8628 17756
rect 8668 17808 8720 17814
rect 8668 17750 8720 17756
rect 8864 17762 8892 18720
rect 8944 18702 8996 18708
rect 8942 18592 8998 18601
rect 9140 18578 9168 18822
rect 8998 18550 9168 18578
rect 8942 18527 8998 18536
rect 8956 18290 8984 18527
rect 9232 18408 9260 19110
rect 9508 18884 9536 20878
rect 9600 20602 9628 20946
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 9588 20460 9640 20466
rect 9588 20402 9640 20408
rect 9600 19854 9628 20402
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9586 19680 9642 19689
rect 9586 19615 9642 19624
rect 9600 19292 9628 19615
rect 9600 19264 9720 19292
rect 9692 19009 9720 19264
rect 9678 19000 9734 19009
rect 9678 18935 9734 18944
rect 9310 18864 9366 18873
rect 9508 18856 9628 18884
rect 9310 18799 9366 18808
rect 9048 18380 9260 18408
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 9048 18086 9076 18380
rect 9324 18290 9352 18799
rect 9402 18456 9458 18465
rect 9458 18414 9536 18442
rect 9402 18391 9458 18400
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9036 18080 9088 18086
rect 8956 18040 9036 18068
rect 8956 17882 8984 18040
rect 9140 18068 9168 18226
rect 9140 18040 9444 18068
rect 9036 18022 9088 18028
rect 9416 17921 9444 18040
rect 9402 17912 9458 17921
rect 8944 17876 8996 17882
rect 9402 17847 9458 17856
rect 8944 17818 8996 17824
rect 8864 17734 8984 17762
rect 9508 17746 9536 18414
rect 8852 17672 8904 17678
rect 8496 17632 8852 17660
rect 8852 17614 8904 17620
rect 8392 17604 8444 17610
rect 8444 17564 8524 17592
rect 8392 17546 8444 17552
rect 8496 17270 8524 17564
rect 8484 17264 8536 17270
rect 8484 17206 8536 17212
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8576 17128 8628 17134
rect 8956 17116 8984 17734
rect 9220 17740 9272 17746
rect 9140 17700 9220 17728
rect 9036 17128 9088 17134
rect 8956 17088 9036 17116
rect 8576 17070 8628 17076
rect 9036 17070 9088 17076
rect 7988 16892 8296 16901
rect 7988 16890 7994 16892
rect 8050 16890 8074 16892
rect 8130 16890 8154 16892
rect 8210 16890 8234 16892
rect 8290 16890 8296 16892
rect 8050 16838 8052 16890
rect 8232 16838 8234 16890
rect 7988 16836 7994 16838
rect 8050 16836 8074 16838
rect 8130 16836 8154 16838
rect 8210 16836 8234 16838
rect 8290 16836 8296 16838
rect 7988 16827 8296 16836
rect 8404 16114 8432 17070
rect 8588 16833 8616 17070
rect 8666 16960 8722 16969
rect 8666 16895 8722 16904
rect 8574 16824 8630 16833
rect 8680 16794 8708 16895
rect 8574 16759 8630 16768
rect 8668 16788 8720 16794
rect 8482 16688 8538 16697
rect 8482 16623 8538 16632
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8312 16017 8340 16050
rect 8496 16046 8524 16623
rect 8484 16040 8536 16046
rect 8298 16008 8354 16017
rect 8484 15982 8536 15988
rect 8298 15943 8354 15952
rect 8588 15910 8616 16759
rect 8668 16730 8720 16736
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8680 16046 8708 16526
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 7988 15804 8296 15813
rect 7988 15802 7994 15804
rect 8050 15802 8074 15804
rect 8130 15802 8154 15804
rect 8210 15802 8234 15804
rect 8290 15802 8296 15804
rect 8050 15750 8052 15802
rect 8232 15750 8234 15802
rect 7988 15748 7994 15750
rect 8050 15748 8074 15750
rect 8130 15748 8154 15750
rect 8210 15748 8234 15750
rect 8290 15748 8296 15750
rect 7988 15739 8296 15748
rect 7852 15660 7972 15688
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7852 13802 7880 15438
rect 7944 15065 7972 15660
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8312 15162 8340 15302
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 7930 15056 7986 15065
rect 7930 14991 7986 15000
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 7988 14716 8296 14725
rect 7988 14714 7994 14716
rect 8050 14714 8074 14716
rect 8130 14714 8154 14716
rect 8210 14714 8234 14716
rect 8290 14714 8296 14716
rect 8050 14662 8052 14714
rect 8232 14662 8234 14714
rect 7988 14660 7994 14662
rect 8050 14660 8074 14662
rect 8130 14660 8154 14662
rect 8210 14660 8234 14662
rect 8290 14660 8296 14662
rect 7988 14651 8296 14660
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8220 13870 8248 14214
rect 8208 13864 8260 13870
rect 8312 13852 8340 14554
rect 8404 14006 8432 14894
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 8392 13864 8444 13870
rect 8312 13824 8392 13852
rect 8208 13806 8260 13812
rect 8392 13806 8444 13812
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 7988 13628 8296 13637
rect 7988 13626 7994 13628
rect 8050 13626 8074 13628
rect 8130 13626 8154 13628
rect 8210 13626 8234 13628
rect 8290 13626 8296 13628
rect 8050 13574 8052 13626
rect 8232 13574 8234 13626
rect 7988 13572 7994 13574
rect 8050 13572 8074 13574
rect 8130 13572 8154 13574
rect 8210 13572 8234 13574
rect 8290 13572 8296 13574
rect 7988 13563 8296 13572
rect 7760 13530 7880 13546
rect 7760 13524 7892 13530
rect 7760 13518 7840 13524
rect 7840 13466 7892 13472
rect 8404 13310 8432 13806
rect 8496 13462 8524 14826
rect 8588 14600 8616 15846
rect 8680 15502 8708 15982
rect 8956 15910 8984 16730
rect 9034 16416 9090 16425
rect 9034 16351 9090 16360
rect 8944 15904 8996 15910
rect 8864 15864 8944 15892
rect 8864 15502 8892 15864
rect 8944 15846 8996 15852
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 8680 14958 8708 15438
rect 8864 15026 8892 15438
rect 8852 15020 8904 15026
rect 8772 14980 8852 15008
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8680 14793 8708 14894
rect 8666 14784 8722 14793
rect 8666 14719 8722 14728
rect 8588 14572 8708 14600
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8484 13456 8536 13462
rect 8484 13398 8536 13404
rect 8404 13282 8524 13310
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 8390 13016 8446 13025
rect 8390 12951 8446 12960
rect 8404 12918 8432 12951
rect 8392 12912 8444 12918
rect 8392 12854 8444 12860
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7852 11762 7880 12718
rect 7988 12540 8296 12549
rect 7988 12538 7994 12540
rect 8050 12538 8074 12540
rect 8130 12538 8154 12540
rect 8210 12538 8234 12540
rect 8290 12538 8296 12540
rect 8050 12486 8052 12538
rect 8232 12486 8234 12538
rect 7988 12484 7994 12486
rect 8050 12484 8074 12486
rect 8130 12484 8154 12486
rect 8210 12484 8234 12486
rect 8290 12484 8296 12486
rect 7988 12475 8296 12484
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7564 11552 7616 11558
rect 7852 11529 7880 11698
rect 8036 11694 8064 12038
rect 8312 11694 8340 12378
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 7564 11494 7616 11500
rect 7838 11520 7894 11529
rect 7576 11218 7604 11494
rect 7838 11455 7894 11464
rect 7988 11452 8296 11461
rect 7988 11450 7994 11452
rect 8050 11450 8074 11452
rect 8130 11450 8154 11452
rect 8210 11450 8234 11452
rect 8290 11450 8296 11452
rect 8050 11398 8052 11450
rect 8232 11398 8234 11450
rect 7988 11396 7994 11398
rect 8050 11396 8074 11398
rect 8130 11396 8154 11398
rect 8210 11396 8234 11398
rect 8290 11396 8296 11398
rect 7988 11387 8296 11396
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7288 11144 7340 11150
rect 7208 11104 7288 11132
rect 7288 11086 7340 11092
rect 7668 10690 7696 11154
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7576 10662 7696 10690
rect 7470 10160 7526 10169
rect 7392 10118 7470 10146
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6090 9208 6146 9217
rect 6090 9143 6146 9152
rect 6104 9042 6132 9143
rect 6380 9042 6408 9318
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6288 8906 6592 8922
rect 6276 8900 6592 8906
rect 6328 8894 6592 8900
rect 6276 8842 6328 8848
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6000 8288 6052 8294
rect 5736 8214 5856 8242
rect 6000 8230 6052 8236
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5630 7168 5686 7177
rect 5630 7103 5686 7112
rect 5632 6860 5684 6866
rect 5736 6848 5764 8026
rect 5828 8022 5856 8214
rect 5816 8016 5868 8022
rect 5868 7976 6132 8004
rect 5816 7958 5868 7964
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5828 7002 5856 7822
rect 6012 7750 6040 7822
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 5908 7404 5960 7410
rect 6012 7392 6040 7686
rect 5960 7364 6040 7392
rect 5908 7346 5960 7352
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5684 6820 5764 6848
rect 5814 6896 5870 6905
rect 5920 6866 5948 7346
rect 5814 6831 5870 6840
rect 5908 6860 5960 6866
rect 5632 6802 5684 6808
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5644 5545 5672 6802
rect 5828 6662 5856 6831
rect 5908 6802 5960 6808
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5920 6322 5948 6802
rect 6104 6610 6132 7976
rect 6380 7857 6408 8774
rect 6366 7848 6422 7857
rect 6366 7783 6422 7792
rect 6366 6896 6422 6905
rect 6366 6831 6422 6840
rect 6380 6798 6408 6831
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6012 6582 6132 6610
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5630 5536 5686 5545
rect 5630 5471 5686 5480
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5644 4706 5672 5471
rect 5368 4678 5672 4706
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5276 3534 5304 4558
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5134 2774 5212 2802
rect 5078 2751 5134 2760
rect 5276 2378 5304 3470
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 5368 1766 5396 4678
rect 5736 4298 5764 6258
rect 5814 6080 5870 6089
rect 5814 6015 5870 6024
rect 5828 5710 5856 6015
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5828 4622 5856 5646
rect 5906 4720 5962 4729
rect 5906 4655 5962 4664
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5736 4270 5856 4298
rect 5448 4072 5500 4078
rect 5632 4072 5684 4078
rect 5448 4014 5500 4020
rect 5630 4040 5632 4049
rect 5684 4040 5686 4049
rect 5460 3369 5488 4014
rect 5630 3975 5686 3984
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5644 3641 5672 3878
rect 5828 3738 5856 4270
rect 5920 4146 5948 4655
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5724 3664 5776 3670
rect 5630 3632 5686 3641
rect 5724 3606 5776 3612
rect 5630 3567 5686 3576
rect 5446 3360 5502 3369
rect 5446 3295 5502 3304
rect 5736 3194 5764 3606
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 5552 2774 5580 2994
rect 5460 2746 5580 2774
rect 5460 2530 5488 2746
rect 5538 2680 5594 2689
rect 5538 2615 5540 2624
rect 5592 2615 5594 2624
rect 5540 2586 5592 2592
rect 5460 2502 5580 2530
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 5460 1902 5488 2314
rect 5448 1896 5500 1902
rect 5448 1838 5500 1844
rect 5356 1760 5408 1766
rect 5078 1728 5134 1737
rect 5356 1702 5408 1708
rect 5078 1663 5134 1672
rect 5092 1018 5120 1663
rect 5552 1562 5580 2502
rect 5644 2106 5672 3130
rect 5828 3126 5856 3402
rect 6012 3210 6040 6582
rect 6090 6488 6146 6497
rect 6090 6423 6146 6432
rect 6104 6322 6132 6423
rect 6472 6322 6500 8774
rect 6564 6798 6592 8894
rect 6656 8090 6684 8978
rect 6748 8956 6776 9454
rect 7012 8968 7064 8974
rect 6748 8928 7012 8956
rect 7012 8910 7064 8916
rect 7012 8832 7064 8838
rect 7012 8774 7064 8780
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6748 7562 6776 8434
rect 6656 7534 6776 7562
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6104 5302 6132 5850
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6288 5370 6316 5646
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6288 4826 6316 5170
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 6182 4448 6238 4457
rect 6182 4383 6238 4392
rect 6196 4146 6224 4383
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6288 3516 6316 4762
rect 6380 4622 6408 4966
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6472 3534 6500 5510
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6368 3528 6420 3534
rect 6288 3488 6368 3516
rect 6368 3470 6420 3476
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 5920 3182 6040 3210
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 5632 2100 5684 2106
rect 5632 2042 5684 2048
rect 5632 1828 5684 1834
rect 5632 1770 5684 1776
rect 5540 1556 5592 1562
rect 5540 1498 5592 1504
rect 5644 1290 5672 1770
rect 5736 1766 5764 2450
rect 5724 1760 5776 1766
rect 5724 1702 5776 1708
rect 5814 1728 5870 1737
rect 5632 1284 5684 1290
rect 5632 1226 5684 1232
rect 5170 1184 5226 1193
rect 5170 1119 5226 1128
rect 5184 1018 5212 1119
rect 5446 1048 5502 1057
rect 4988 1012 5040 1018
rect 4988 954 5040 960
rect 5080 1012 5132 1018
rect 5080 954 5132 960
rect 5172 1012 5224 1018
rect 5446 983 5502 992
rect 5172 954 5224 960
rect 4804 944 4856 950
rect 4804 886 4856 892
rect 5460 882 5488 983
rect 5448 876 5500 882
rect 5448 818 5500 824
rect 5540 808 5592 814
rect 5540 750 5592 756
rect 4712 672 4764 678
rect 4712 614 4764 620
rect 3974 96 4030 105
rect 5552 66 5580 750
rect 5736 474 5764 1702
rect 5920 1714 5948 3182
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 6012 1970 6040 3062
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 6104 2281 6132 2926
rect 6090 2272 6146 2281
rect 6090 2207 6146 2216
rect 6000 1964 6052 1970
rect 6000 1906 6052 1912
rect 5920 1686 6040 1714
rect 5814 1663 5870 1672
rect 5828 1426 5856 1663
rect 5906 1592 5962 1601
rect 5906 1527 5908 1536
rect 5960 1527 5962 1536
rect 5908 1498 5960 1504
rect 6012 1426 6040 1686
rect 5816 1420 5868 1426
rect 5816 1362 5868 1368
rect 6000 1420 6052 1426
rect 6000 1362 6052 1368
rect 5816 944 5868 950
rect 5816 886 5868 892
rect 5828 474 5856 886
rect 5908 740 5960 746
rect 6012 728 6040 1362
rect 6104 814 6132 2207
rect 6196 1426 6224 2926
rect 6380 2650 6408 3470
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 6472 2446 6500 3334
rect 6564 2854 6592 4966
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6276 2440 6328 2446
rect 6460 2440 6512 2446
rect 6328 2400 6408 2428
rect 6276 2382 6328 2388
rect 6380 1970 6408 2400
rect 6460 2382 6512 2388
rect 6368 1964 6420 1970
rect 6368 1906 6420 1912
rect 6274 1864 6330 1873
rect 6564 1850 6592 2790
rect 6656 2774 6684 7534
rect 6734 7440 6790 7449
rect 6734 7375 6736 7384
rect 6788 7375 6790 7384
rect 6736 7346 6788 7352
rect 7024 5953 7052 8774
rect 7116 8634 7144 9998
rect 7208 9178 7236 9998
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7194 9072 7250 9081
rect 7194 9007 7196 9016
rect 7248 9007 7250 9016
rect 7196 8978 7248 8984
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7300 6497 7328 9998
rect 7286 6488 7342 6497
rect 7286 6423 7342 6432
rect 7392 6338 7420 10118
rect 7470 10095 7526 10104
rect 7470 9208 7526 9217
rect 7576 9178 7604 10662
rect 7656 10532 7708 10538
rect 7656 10474 7708 10480
rect 7668 9178 7696 10474
rect 7470 9143 7526 9152
rect 7564 9172 7616 9178
rect 7484 9058 7512 9143
rect 7564 9114 7616 9120
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7760 9058 7788 10746
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7852 10266 7880 10474
rect 7988 10364 8296 10373
rect 7988 10362 7994 10364
rect 8050 10362 8074 10364
rect 8130 10362 8154 10364
rect 8210 10362 8234 10364
rect 8290 10362 8296 10364
rect 8050 10310 8052 10362
rect 8232 10310 8234 10362
rect 7988 10308 7994 10310
rect 8050 10308 8074 10310
rect 8130 10308 8154 10310
rect 8210 10308 8234 10310
rect 8290 10308 8296 10310
rect 7988 10299 8296 10308
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 7852 9450 7880 10202
rect 8404 9625 8432 12854
rect 8496 12442 8524 13282
rect 8588 12782 8616 14418
rect 8680 14090 8708 14572
rect 8772 14278 8800 14980
rect 8852 14962 8904 14968
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8680 14062 8800 14090
rect 8666 13968 8722 13977
rect 8666 13903 8722 13912
rect 8680 13734 8708 13903
rect 8668 13728 8720 13734
rect 8772 13716 8800 14062
rect 8864 13841 8892 14214
rect 8850 13832 8906 13841
rect 8850 13767 8906 13776
rect 8772 13688 8892 13716
rect 8668 13670 8720 13676
rect 8680 12866 8708 13670
rect 8864 13394 8892 13688
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8772 12986 8800 13262
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8680 12838 8800 12866
rect 8772 12782 8800 12838
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11762 8524 12038
rect 8588 11898 8616 12174
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8482 10976 8538 10985
rect 8538 10934 8616 10962
rect 8482 10911 8538 10920
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8390 9616 8446 9625
rect 8496 9586 8524 9998
rect 8588 9994 8616 10934
rect 8668 10600 8720 10606
rect 8772 10588 8800 11630
rect 8864 11558 8892 12174
rect 9048 11898 9076 16351
rect 9140 15502 9168 17700
rect 9220 17682 9272 17688
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9232 17202 9260 17274
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9324 17134 9352 17274
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9508 16697 9536 17070
rect 9494 16688 9550 16697
rect 9404 16652 9456 16658
rect 9494 16623 9550 16632
rect 9404 16594 9456 16600
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9126 15328 9182 15337
rect 9182 15286 9260 15314
rect 9126 15263 9182 15272
rect 9126 14376 9182 14385
rect 9126 14311 9182 14320
rect 9140 14006 9168 14311
rect 9128 14000 9180 14006
rect 9128 13942 9180 13948
rect 9232 13530 9260 15286
rect 9324 14618 9352 15438
rect 9416 14618 9444 16594
rect 9600 15337 9628 18856
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9692 16998 9720 17818
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9678 16144 9734 16153
rect 9678 16079 9734 16088
rect 9692 16046 9720 16079
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9586 15328 9642 15337
rect 9586 15263 9642 15272
rect 9784 14822 9812 21082
rect 9862 20088 9918 20097
rect 9862 20023 9918 20032
rect 9876 19310 9904 20023
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 9312 13864 9364 13870
rect 9404 13864 9456 13870
rect 9312 13806 9364 13812
rect 9402 13832 9404 13841
rect 9496 13864 9548 13870
rect 9456 13832 9458 13841
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9128 13456 9180 13462
rect 9128 13398 9180 13404
rect 9140 13326 9168 13398
rect 9324 13394 9352 13806
rect 9496 13806 9548 13812
rect 9402 13767 9458 13776
rect 9312 13388 9364 13394
rect 9508 13376 9536 13806
rect 9588 13456 9640 13462
rect 9312 13330 9364 13336
rect 9416 13348 9536 13376
rect 9586 13424 9588 13433
rect 9640 13424 9642 13433
rect 9586 13359 9642 13368
rect 9784 13376 9812 14486
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 14074 9904 14214
rect 9968 14074 9996 22102
rect 12716 22024 12768 22030
rect 10966 21992 11022 22001
rect 10966 21927 11022 21936
rect 11426 21992 11482 22001
rect 12716 21966 12768 21972
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 11426 21927 11482 21936
rect 10980 21894 11008 21927
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10140 21684 10192 21690
rect 10140 21626 10192 21632
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 10060 15178 10088 21422
rect 10152 19310 10180 21626
rect 10244 21078 10272 21626
rect 10600 21412 10652 21418
rect 10600 21354 10652 21360
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 10508 21344 10560 21350
rect 10508 21286 10560 21292
rect 10232 21072 10284 21078
rect 10232 21014 10284 21020
rect 10336 20466 10364 21286
rect 10416 21072 10468 21078
rect 10416 21014 10468 21020
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10244 19514 10272 20402
rect 10428 20097 10456 21014
rect 10520 20777 10548 21286
rect 10506 20768 10562 20777
rect 10506 20703 10562 20712
rect 10506 20496 10562 20505
rect 10506 20431 10562 20440
rect 10414 20088 10470 20097
rect 10414 20023 10470 20032
rect 10520 19961 10548 20431
rect 10506 19952 10562 19961
rect 10506 19887 10562 19896
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 10140 19304 10192 19310
rect 10140 19246 10192 19252
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10244 18873 10272 19178
rect 10230 18864 10286 18873
rect 10230 18799 10286 18808
rect 10138 17640 10194 17649
rect 10138 17575 10194 17584
rect 10152 16998 10180 17575
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10152 16182 10180 16390
rect 10140 16176 10192 16182
rect 10140 16118 10192 16124
rect 10060 15150 10180 15178
rect 10046 14784 10102 14793
rect 10046 14719 10102 14728
rect 10060 14550 10088 14719
rect 10048 14544 10100 14550
rect 10048 14486 10100 14492
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 9864 13388 9916 13394
rect 9784 13348 9864 13376
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9324 13190 9352 13330
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9232 12986 9260 13126
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 9140 11354 9168 12174
rect 9324 11694 9352 13126
rect 9416 12918 9444 13348
rect 9864 13330 9916 13336
rect 9508 13258 9812 13274
rect 9496 13252 9812 13258
rect 9548 13246 9812 13252
rect 9784 13240 9812 13246
rect 9784 13212 9996 13240
rect 9496 13194 9548 13200
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 9416 12102 9444 12854
rect 9968 12850 9996 13212
rect 10060 12866 10088 13806
rect 10152 13433 10180 15150
rect 10138 13424 10194 13433
rect 10138 13359 10194 13368
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 10152 13025 10180 13194
rect 10138 13016 10194 13025
rect 10138 12951 10194 12960
rect 9956 12844 10008 12850
rect 10060 12838 10183 12866
rect 9956 12786 10008 12792
rect 10155 12764 10183 12838
rect 10060 12736 10183 12764
rect 10060 12730 10088 12736
rect 9968 12702 10088 12730
rect 9968 12646 9996 12702
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9692 12345 9720 12582
rect 9678 12336 9734 12345
rect 9678 12271 9734 12280
rect 9864 12300 9916 12306
rect 9968 12288 9996 12582
rect 9916 12260 10180 12288
rect 9864 12242 9916 12248
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9678 12064 9734 12073
rect 9416 11694 9444 12038
rect 9678 11999 9734 12008
rect 9682 11914 9710 11999
rect 9682 11886 9720 11914
rect 9692 11830 9720 11886
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9324 11218 9352 11630
rect 9416 11354 9444 11630
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 10048 11552 10100 11558
rect 10152 11540 10180 12260
rect 10100 11512 10180 11540
rect 10048 11494 10100 11500
rect 9968 11393 9996 11494
rect 9954 11384 10010 11393
rect 9404 11348 9456 11354
rect 9954 11319 10010 11328
rect 9404 11290 9456 11296
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8720 10560 8800 10588
rect 8668 10542 8720 10548
rect 8680 10441 8708 10542
rect 8760 10464 8812 10470
rect 8666 10432 8722 10441
rect 8760 10406 8812 10412
rect 8666 10367 8722 10376
rect 8576 9988 8628 9994
rect 8576 9930 8628 9936
rect 8772 9722 8800 10406
rect 8864 9722 8892 10746
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8390 9551 8446 9560
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 7852 9178 7880 9386
rect 7988 9276 8296 9285
rect 7988 9274 7994 9276
rect 8050 9274 8074 9276
rect 8130 9274 8154 9276
rect 8210 9274 8234 9276
rect 8290 9274 8296 9276
rect 8050 9222 8052 9274
rect 8232 9222 8234 9274
rect 7988 9220 7994 9222
rect 8050 9220 8074 9222
rect 8130 9220 8154 9222
rect 8210 9220 8234 9222
rect 8290 9220 8296 9222
rect 7988 9211 8296 9220
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7484 9042 7788 9058
rect 7472 9036 7788 9042
rect 7524 9030 7788 9036
rect 8208 9036 8260 9042
rect 7472 8978 7524 8984
rect 8208 8978 8260 8984
rect 7470 8528 7526 8537
rect 7470 8463 7526 8472
rect 7208 6310 7420 6338
rect 7010 5944 7066 5953
rect 7010 5879 7066 5888
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6748 5545 6776 5646
rect 7012 5568 7064 5574
rect 6734 5536 6790 5545
rect 7012 5510 7064 5516
rect 6734 5471 6790 5480
rect 7024 5234 7052 5510
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6748 4622 6776 5102
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6748 3534 6776 3674
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6932 2825 6960 3470
rect 6918 2816 6974 2825
rect 6656 2746 6776 2774
rect 6918 2751 6974 2760
rect 6642 2680 6698 2689
rect 6642 2615 6698 2624
rect 6656 2514 6684 2615
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 6330 1822 6592 1850
rect 6274 1799 6330 1808
rect 6184 1420 6236 1426
rect 6184 1362 6236 1368
rect 6288 882 6316 1799
rect 6748 882 6776 2746
rect 7208 1358 7236 6310
rect 7484 6236 7512 8463
rect 7840 8288 7892 8294
rect 8220 8276 8248 8978
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8312 8634 8340 8910
rect 8404 8634 8432 9454
rect 8484 8968 8536 8974
rect 8482 8936 8484 8945
rect 8536 8936 8538 8945
rect 8482 8871 8538 8880
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8496 8634 8524 8774
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8496 8498 8524 8570
rect 8680 8498 8708 8774
rect 8772 8566 8800 9658
rect 9048 9382 9076 9998
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 8760 8560 8812 8566
rect 8760 8502 8812 8508
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8668 8492 8720 8498
rect 8956 8480 8984 9318
rect 9140 8634 9168 11018
rect 9324 10606 9352 11018
rect 9416 10674 9444 11290
rect 10060 11218 10088 11494
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9416 10130 9444 10406
rect 9508 10266 9536 11154
rect 9862 10976 9918 10985
rect 9862 10911 9918 10920
rect 9586 10840 9642 10849
rect 9586 10775 9642 10784
rect 9600 10452 9628 10775
rect 9876 10674 9904 10911
rect 10060 10674 10088 11154
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9600 10424 9720 10452
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9232 9178 9260 9454
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9312 8560 9364 8566
rect 9218 8528 9274 8537
rect 9128 8492 9180 8498
rect 8956 8452 9128 8480
rect 8668 8434 8720 8440
rect 9312 8502 9364 8508
rect 9218 8463 9274 8472
rect 9128 8434 9180 8440
rect 9232 8430 9260 8463
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9036 8288 9088 8294
rect 8220 8248 8432 8276
rect 7840 8230 7892 8236
rect 7654 8120 7710 8129
rect 7654 8055 7656 8064
rect 7708 8055 7710 8064
rect 7656 8026 7708 8032
rect 7852 7818 7880 8230
rect 7988 8188 8296 8197
rect 7988 8186 7994 8188
rect 8050 8186 8074 8188
rect 8130 8186 8154 8188
rect 8210 8186 8234 8188
rect 8290 8186 8296 8188
rect 8050 8134 8052 8186
rect 8232 8134 8234 8186
rect 7988 8132 7994 8134
rect 8050 8132 8074 8134
rect 8130 8132 8154 8134
rect 8210 8132 8234 8134
rect 8290 8132 8296 8134
rect 7988 8123 8296 8132
rect 8404 7954 8432 8248
rect 9036 8230 9088 8236
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7576 7478 7604 7686
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7668 7206 7696 7482
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7656 7200 7708 7206
rect 7852 7177 7880 7278
rect 8312 7188 8340 7754
rect 8404 7342 8432 7890
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8588 7410 8616 7822
rect 9048 7800 9076 8230
rect 9140 7954 9168 8230
rect 9324 7954 9352 8502
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9048 7772 9168 7800
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8576 7404 8628 7410
rect 8576 7346 8628 7352
rect 8392 7336 8444 7342
rect 8444 7296 8524 7324
rect 8392 7278 8444 7284
rect 7656 7142 7708 7148
rect 7838 7168 7894 7177
rect 8312 7160 8432 7188
rect 7838 7103 7894 7112
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7760 6361 7788 6598
rect 7746 6352 7802 6361
rect 7746 6287 7802 6296
rect 7300 6208 7512 6236
rect 7196 1352 7248 1358
rect 7196 1294 7248 1300
rect 7300 1018 7328 6208
rect 7748 6180 7800 6186
rect 7748 6122 7800 6128
rect 7656 6112 7708 6118
rect 7654 6080 7656 6089
rect 7708 6080 7710 6089
rect 7654 6015 7710 6024
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7576 5234 7604 5850
rect 7760 5710 7788 6122
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7760 4622 7788 5646
rect 7852 5166 7880 7103
rect 7988 7100 8296 7109
rect 7988 7098 7994 7100
rect 8050 7098 8074 7100
rect 8130 7098 8154 7100
rect 8210 7098 8234 7100
rect 8290 7098 8296 7100
rect 8050 7046 8052 7098
rect 8232 7046 8234 7098
rect 7988 7044 7994 7046
rect 8050 7044 8074 7046
rect 8130 7044 8154 7046
rect 8210 7044 8234 7046
rect 8290 7044 8296 7046
rect 7988 7035 8296 7044
rect 8404 6225 8432 7160
rect 8496 6866 8524 7296
rect 8588 7002 8616 7346
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8496 6254 8524 6802
rect 8588 6322 8616 6938
rect 8956 6798 8984 7686
rect 9140 7410 9168 7772
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8484 6248 8536 6254
rect 8390 6216 8446 6225
rect 8484 6190 8536 6196
rect 8390 6151 8446 6160
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 7988 6012 8296 6021
rect 7988 6010 7994 6012
rect 8050 6010 8074 6012
rect 8130 6010 8154 6012
rect 8210 6010 8234 6012
rect 8290 6010 8296 6012
rect 8050 5958 8052 6010
rect 8232 5958 8234 6010
rect 7988 5956 7994 5958
rect 8050 5956 8074 5958
rect 8130 5956 8154 5958
rect 8210 5956 8234 5958
rect 8290 5956 8296 5958
rect 7988 5947 8296 5956
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7988 4924 8296 4933
rect 7988 4922 7994 4924
rect 8050 4922 8074 4924
rect 8130 4922 8154 4924
rect 8210 4922 8234 4924
rect 8290 4922 8296 4924
rect 8050 4870 8052 4922
rect 8232 4870 8234 4922
rect 7988 4868 7994 4870
rect 8050 4868 8074 4870
rect 8130 4868 8154 4870
rect 8210 4868 8234 4870
rect 8290 4868 8296 4870
rect 7988 4859 8296 4868
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7392 2281 7420 2382
rect 7576 2378 7604 4218
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7378 2272 7434 2281
rect 7378 2207 7434 2216
rect 7668 2106 7696 2994
rect 7760 2854 7788 4558
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7852 3738 7880 3878
rect 7988 3836 8296 3845
rect 7988 3834 7994 3836
rect 8050 3834 8074 3836
rect 8130 3834 8154 3836
rect 8210 3834 8234 3836
rect 8290 3834 8296 3836
rect 8050 3782 8052 3834
rect 8232 3782 8234 3834
rect 7988 3780 7994 3782
rect 8050 3780 8074 3782
rect 8130 3780 8154 3782
rect 8210 3780 8234 3782
rect 8290 3780 8296 3782
rect 7988 3771 8296 3780
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 8496 3670 8524 5646
rect 8680 4826 8708 5850
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8588 3738 8616 4626
rect 8680 4010 8708 4762
rect 8668 4004 8720 4010
rect 8668 3946 8720 3952
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7760 2446 7788 2790
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7852 2106 7880 2994
rect 8680 2990 8708 3946
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 7988 2748 8296 2757
rect 7988 2746 7994 2748
rect 8050 2746 8074 2748
rect 8130 2746 8154 2748
rect 8210 2746 8234 2748
rect 8290 2746 8296 2748
rect 8050 2694 8052 2746
rect 8232 2694 8234 2746
rect 7988 2692 7994 2694
rect 8050 2692 8074 2694
rect 8130 2692 8154 2694
rect 8210 2692 8234 2694
rect 8290 2692 8296 2694
rect 7988 2683 8296 2692
rect 8496 2514 8524 2926
rect 8772 2774 8800 5646
rect 8956 5273 8984 6054
rect 9416 5386 9444 8842
rect 9508 8430 9536 10202
rect 9692 10130 9720 10424
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9862 9616 9918 9625
rect 9862 9551 9918 9560
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 8430 9628 9318
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9692 7857 9720 8026
rect 9678 7848 9734 7857
rect 9678 7783 9734 7792
rect 9876 6458 9904 9551
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9416 5358 9536 5386
rect 8942 5264 8998 5273
rect 8852 5228 8904 5234
rect 8942 5199 8998 5208
rect 9404 5228 9456 5234
rect 8852 5170 8904 5176
rect 9404 5170 9456 5176
rect 8864 4826 8892 5170
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8864 4593 8892 4626
rect 8850 4584 8906 4593
rect 8850 4519 8906 4528
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8864 4010 8892 4422
rect 8956 4078 8984 5102
rect 9048 4214 9076 5102
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 8680 2746 8800 2774
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7840 2100 7892 2106
rect 7840 2042 7892 2048
rect 7748 2032 7800 2038
rect 7748 1974 7800 1980
rect 7760 1601 7788 1974
rect 8128 1902 8156 2246
rect 8116 1896 8168 1902
rect 8116 1838 8168 1844
rect 7988 1660 8296 1669
rect 7988 1658 7994 1660
rect 8050 1658 8074 1660
rect 8130 1658 8154 1660
rect 8210 1658 8234 1660
rect 8290 1658 8296 1660
rect 8050 1606 8052 1658
rect 8232 1606 8234 1658
rect 7988 1604 7994 1606
rect 8050 1604 8074 1606
rect 8130 1604 8154 1606
rect 8210 1604 8234 1606
rect 8290 1604 8296 1606
rect 7746 1592 7802 1601
rect 7988 1595 8296 1604
rect 7746 1527 7802 1536
rect 8298 1048 8354 1057
rect 7288 1012 7340 1018
rect 8680 1018 8708 2746
rect 8864 2106 8892 3946
rect 8956 3602 8984 4014
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 9048 3534 9076 4150
rect 9416 4010 9444 5170
rect 9508 5030 9536 5358
rect 9600 5234 9628 5510
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9784 4826 9812 5102
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9416 3738 9444 3946
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9310 3496 9366 3505
rect 8942 3360 8998 3369
rect 8942 3295 8998 3304
rect 8956 2854 8984 3295
rect 9048 2990 9076 3470
rect 9232 3194 9260 3470
rect 9310 3431 9366 3440
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 8852 2100 8904 2106
rect 8852 2042 8904 2048
rect 8852 1964 8904 1970
rect 8852 1906 8904 1912
rect 8298 983 8354 992
rect 8668 1012 8720 1018
rect 7288 954 7340 960
rect 6276 876 6328 882
rect 6276 818 6328 824
rect 6644 876 6696 882
rect 6644 818 6696 824
rect 6736 876 6788 882
rect 6736 818 6788 824
rect 6092 808 6144 814
rect 6092 750 6144 756
rect 5960 700 6040 728
rect 5908 682 5960 688
rect 5724 468 5776 474
rect 5724 410 5776 416
rect 5816 468 5868 474
rect 5816 410 5868 416
rect 6104 202 6132 750
rect 6656 241 6684 818
rect 8312 814 8340 983
rect 8668 954 8720 960
rect 8864 882 8892 1906
rect 9048 1902 9076 2926
rect 9036 1896 9088 1902
rect 8956 1856 9036 1884
rect 8956 1222 8984 1856
rect 9324 1873 9352 3431
rect 9416 3058 9444 3674
rect 9508 3602 9536 4490
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10060 4146 10088 4422
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9692 3194 9720 4082
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9036 1838 9088 1844
rect 9126 1864 9182 1873
rect 9126 1799 9182 1808
rect 9310 1864 9366 1873
rect 9310 1799 9366 1808
rect 9036 1760 9088 1766
rect 9036 1702 9088 1708
rect 9048 1358 9076 1702
rect 9140 1358 9168 1799
rect 9416 1766 9444 2994
rect 9600 2650 9628 2994
rect 9588 2644 9640 2650
rect 9784 2632 9812 3878
rect 10048 2644 10100 2650
rect 9784 2604 10048 2632
rect 9588 2586 9640 2592
rect 10048 2586 10100 2592
rect 9404 1760 9456 1766
rect 9404 1702 9456 1708
rect 9680 1760 9732 1766
rect 9680 1702 9732 1708
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 9128 1352 9180 1358
rect 9128 1294 9180 1300
rect 8944 1216 8996 1222
rect 9692 1193 9720 1702
rect 10152 1358 10180 11086
rect 10244 10130 10272 18799
rect 10416 17536 10468 17542
rect 10612 17513 10640 21354
rect 10704 21010 10732 21830
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 10692 21004 10744 21010
rect 10692 20946 10744 20952
rect 10692 20528 10744 20534
rect 10692 20470 10744 20476
rect 10704 18154 10732 20470
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10416 17478 10468 17484
rect 10598 17504 10654 17513
rect 10428 16833 10456 17478
rect 10598 17439 10654 17448
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10414 16824 10470 16833
rect 10520 16794 10548 17070
rect 10414 16759 10470 16768
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 10324 16584 10376 16590
rect 10324 16526 10376 16532
rect 10336 16250 10364 16526
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10322 15736 10378 15745
rect 10322 15671 10378 15680
rect 10336 12209 10364 15671
rect 10506 14920 10562 14929
rect 10506 14855 10562 14864
rect 10520 14822 10548 14855
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10428 14618 10456 14758
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10508 13864 10560 13870
rect 10612 13852 10640 17206
rect 10704 14929 10732 17818
rect 10796 17814 10824 21490
rect 10968 21480 11020 21486
rect 11020 21440 11100 21468
rect 10968 21422 11020 21428
rect 10968 21344 11020 21350
rect 10874 21312 10930 21321
rect 10968 21286 11020 21292
rect 10874 21247 10930 21256
rect 10888 21078 10916 21247
rect 10876 21072 10928 21078
rect 10876 21014 10928 21020
rect 10874 20768 10930 20777
rect 10874 20703 10930 20712
rect 10888 20602 10916 20703
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 10980 20398 11008 21286
rect 11072 20534 11100 21440
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 10968 20392 11020 20398
rect 11020 20352 11100 20380
rect 10968 20334 11020 20340
rect 10874 19544 10930 19553
rect 10874 19479 10930 19488
rect 10784 17808 10836 17814
rect 10784 17750 10836 17756
rect 10888 17270 10916 19479
rect 11072 18970 11100 20352
rect 11164 20330 11192 20878
rect 11256 20398 11284 20878
rect 11440 20466 11468 21927
rect 11783 21788 12091 21797
rect 11783 21786 11789 21788
rect 11845 21786 11869 21788
rect 11925 21786 11949 21788
rect 12005 21786 12029 21788
rect 12085 21786 12091 21788
rect 11845 21734 11847 21786
rect 12027 21734 12029 21786
rect 11783 21732 11789 21734
rect 11845 21732 11869 21734
rect 11925 21732 11949 21734
rect 12005 21732 12029 21734
rect 12085 21732 12091 21734
rect 11783 21723 12091 21732
rect 12162 21720 12218 21729
rect 12162 21655 12218 21664
rect 11704 21480 11756 21486
rect 11532 21440 11704 21468
rect 11532 21146 11560 21440
rect 11704 21422 11756 21428
rect 11520 21140 11572 21146
rect 11520 21082 11572 21088
rect 11612 21140 11664 21146
rect 11612 21082 11664 21088
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 11532 20777 11560 20878
rect 11518 20768 11574 20777
rect 11518 20703 11574 20712
rect 11624 20584 11652 21082
rect 12176 21049 12204 21655
rect 12162 21040 12218 21049
rect 12162 20975 12218 20984
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11808 20806 11836 20878
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11783 20700 12091 20709
rect 11783 20698 11789 20700
rect 11845 20698 11869 20700
rect 11925 20698 11949 20700
rect 12005 20698 12029 20700
rect 12085 20698 12091 20700
rect 11845 20646 11847 20698
rect 12027 20646 12029 20698
rect 11783 20644 11789 20646
rect 11845 20644 11869 20646
rect 11925 20644 11949 20646
rect 12005 20644 12029 20646
rect 12085 20644 12091 20646
rect 11783 20635 12091 20644
rect 11532 20556 11652 20584
rect 11428 20460 11480 20466
rect 11428 20402 11480 20408
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 11152 20324 11204 20330
rect 11152 20266 11204 20272
rect 11256 19514 11284 20334
rect 11336 20324 11388 20330
rect 11388 20284 11468 20312
rect 11336 20266 11388 20272
rect 11440 19786 11468 20284
rect 11532 20262 11560 20556
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11520 20256 11572 20262
rect 11520 20198 11572 20204
rect 11336 19780 11388 19786
rect 11336 19722 11388 19728
rect 11428 19780 11480 19786
rect 11428 19722 11480 19728
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11152 19440 11204 19446
rect 11152 19382 11204 19388
rect 11060 18964 11112 18970
rect 11060 18906 11112 18912
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 10980 18601 11008 18702
rect 10966 18592 11022 18601
rect 10966 18527 11022 18536
rect 11072 18086 11100 18906
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11164 17882 11192 19382
rect 11256 19310 11284 19450
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11256 18766 11284 19110
rect 11250 18760 11302 18766
rect 11250 18702 11302 18708
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11348 17814 11376 19722
rect 11428 19372 11480 19378
rect 11532 19360 11560 20198
rect 11624 19990 11652 20402
rect 12072 20392 12124 20398
rect 11900 20352 12072 20380
rect 11612 19984 11664 19990
rect 11612 19926 11664 19932
rect 11900 19922 11928 20352
rect 12072 20334 12124 20340
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 12440 19916 12492 19922
rect 12492 19876 12572 19904
rect 12440 19858 12492 19864
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 11480 19332 11560 19360
rect 11428 19314 11480 19320
rect 11440 18970 11468 19314
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11428 18964 11480 18970
rect 11428 18906 11480 18912
rect 11532 18766 11560 19110
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11336 17808 11388 17814
rect 11336 17750 11388 17756
rect 11624 17746 11652 19790
rect 11704 19780 11756 19786
rect 11704 19722 11756 19728
rect 11716 19145 11744 19722
rect 11783 19612 12091 19621
rect 11783 19610 11789 19612
rect 11845 19610 11869 19612
rect 11925 19610 11949 19612
rect 12005 19610 12029 19612
rect 12085 19610 12091 19612
rect 11845 19558 11847 19610
rect 12027 19558 12029 19610
rect 11783 19556 11789 19558
rect 11845 19556 11869 19558
rect 11925 19556 11949 19558
rect 12005 19556 12029 19558
rect 12085 19556 12091 19558
rect 11783 19547 12091 19556
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11702 19136 11758 19145
rect 11702 19071 11758 19080
rect 11808 18766 11836 19450
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 10876 17264 10928 17270
rect 10876 17206 10928 17212
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10796 15026 10824 16458
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10690 14920 10746 14929
rect 10690 14855 10746 14864
rect 10560 13824 10640 13852
rect 10508 13806 10560 13812
rect 10322 12200 10378 12209
rect 10322 12135 10378 12144
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10336 11393 10364 11494
rect 10322 11384 10378 11393
rect 10428 11354 10456 13806
rect 10520 11506 10548 13806
rect 10704 13326 10732 14855
rect 10782 14240 10838 14249
rect 10888 14226 10916 17070
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10980 15094 11008 17002
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 11072 16153 11100 16594
rect 11058 16144 11114 16153
rect 11058 16079 11114 16088
rect 11072 15473 11100 16079
rect 11164 15745 11192 17682
rect 11256 17134 11284 17682
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 11256 16590 11284 17070
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11256 16114 11284 16526
rect 11348 16522 11376 16934
rect 11716 16697 11744 18702
rect 11783 18524 12091 18533
rect 11783 18522 11789 18524
rect 11845 18522 11869 18524
rect 11925 18522 11949 18524
rect 12005 18522 12029 18524
rect 12085 18522 12091 18524
rect 11845 18470 11847 18522
rect 12027 18470 12029 18522
rect 11783 18468 11789 18470
rect 11845 18468 11869 18470
rect 11925 18468 11949 18470
rect 12005 18468 12029 18470
rect 12085 18468 12091 18470
rect 11783 18459 12091 18468
rect 12176 17882 12204 19790
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12268 18290 12296 19654
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 11783 17436 12091 17445
rect 11783 17434 11789 17436
rect 11845 17434 11869 17436
rect 11925 17434 11949 17436
rect 12005 17434 12029 17436
rect 12085 17434 12091 17436
rect 11845 17382 11847 17434
rect 12027 17382 12029 17434
rect 11783 17380 11789 17382
rect 11845 17380 11869 17382
rect 11925 17380 11949 17382
rect 12005 17380 12029 17382
rect 12085 17380 12091 17382
rect 11783 17371 12091 17380
rect 12176 17338 12204 17818
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12268 17542 12296 17614
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 16794 11928 16934
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11702 16688 11758 16697
rect 11702 16623 11758 16632
rect 11796 16584 11848 16590
rect 11716 16544 11796 16572
rect 11336 16516 11388 16522
rect 11336 16458 11388 16464
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11150 15736 11206 15745
rect 11150 15671 11206 15680
rect 11256 15570 11284 16050
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11058 15464 11114 15473
rect 11058 15399 11114 15408
rect 11150 15328 11206 15337
rect 11150 15263 11206 15272
rect 11058 15192 11114 15201
rect 11058 15127 11114 15136
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10980 14482 11008 14758
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10838 14198 10916 14226
rect 10782 14175 10838 14184
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10600 13184 10652 13190
rect 10598 13152 10600 13161
rect 10652 13152 10654 13161
rect 10598 13087 10654 13096
rect 10704 12646 10732 13262
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 11762 10640 12038
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10598 11520 10654 11529
rect 10520 11478 10598 11506
rect 10598 11455 10654 11464
rect 10322 11319 10378 11328
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10612 11218 10640 11455
rect 10704 11354 10732 12106
rect 10796 11694 10824 14175
rect 10980 13394 11008 14418
rect 11072 13870 11100 15127
rect 11164 14657 11192 15263
rect 11256 15026 11284 15506
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11150 14648 11206 14657
rect 11150 14583 11206 14592
rect 11164 14550 11192 14583
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 11256 14346 11284 14962
rect 11348 14958 11376 16458
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 11164 14006 11192 14282
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 11348 13938 11376 14350
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11440 13802 11468 16050
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11624 14550 11652 15982
rect 11716 15910 11744 16544
rect 11796 16526 11848 16532
rect 11980 16584 12032 16590
rect 12176 16572 12204 17274
rect 12254 17232 12310 17241
rect 12254 17167 12310 17176
rect 12268 17134 12296 17167
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 12032 16544 12204 16572
rect 11980 16526 12032 16532
rect 11783 16348 12091 16357
rect 11783 16346 11789 16348
rect 11845 16346 11869 16348
rect 11925 16346 11949 16348
rect 12005 16346 12029 16348
rect 12085 16346 12091 16348
rect 11845 16294 11847 16346
rect 12027 16294 12029 16346
rect 11783 16292 11789 16294
rect 11845 16292 11869 16294
rect 11925 16292 11949 16294
rect 12005 16292 12029 16294
rect 12085 16292 12091 16294
rect 11783 16283 12091 16292
rect 12360 16153 12388 17274
rect 12346 16144 12402 16153
rect 12346 16079 12402 16088
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11716 15638 11744 15846
rect 11900 15706 11928 15846
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11716 15042 11744 15574
rect 11992 15366 12020 15642
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11783 15260 12091 15269
rect 11783 15258 11789 15260
rect 11845 15258 11869 15260
rect 11925 15258 11949 15260
rect 12005 15258 12029 15260
rect 12085 15258 12091 15260
rect 11845 15206 11847 15258
rect 12027 15206 12029 15258
rect 11783 15204 11789 15206
rect 11845 15204 11869 15206
rect 11925 15204 11949 15206
rect 12005 15204 12029 15206
rect 12085 15204 12091 15206
rect 11783 15195 12091 15204
rect 11716 15014 12112 15042
rect 11716 14822 11744 15014
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 11150 13696 11206 13705
rect 11150 13631 11206 13640
rect 11058 13560 11114 13569
rect 11164 13530 11192 13631
rect 11058 13495 11114 13504
rect 11152 13524 11204 13530
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 11072 13326 11100 13495
rect 11152 13466 11204 13472
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11164 12889 11192 13466
rect 11624 13394 11652 14010
rect 11716 13938 11744 14758
rect 11992 14618 12020 14894
rect 12084 14618 12112 15014
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 11783 14172 12091 14181
rect 11783 14170 11789 14172
rect 11845 14170 11869 14172
rect 11925 14170 11949 14172
rect 12005 14170 12029 14172
rect 12085 14170 12091 14172
rect 11845 14118 11847 14170
rect 12027 14118 12029 14170
rect 11783 14116 11789 14118
rect 11845 14116 11869 14118
rect 11925 14116 11949 14118
rect 12005 14116 12029 14118
rect 12085 14116 12091 14118
rect 11783 14107 12091 14116
rect 12360 14074 12388 14350
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 11886 13968 11942 13977
rect 11704 13932 11756 13938
rect 11886 13903 11942 13912
rect 11704 13874 11756 13880
rect 11900 13870 11928 13903
rect 11888 13864 11940 13870
rect 12452 13818 12480 19654
rect 12544 14074 12572 19876
rect 12636 19514 12664 20334
rect 12624 19508 12676 19514
rect 12624 19450 12676 19456
rect 12728 19394 12756 21966
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12820 20466 12848 21286
rect 12912 21078 12940 21966
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 12900 21072 12952 21078
rect 12900 21014 12952 21020
rect 13004 20874 13032 21490
rect 13096 21486 13124 21966
rect 13188 21690 13216 22102
rect 14004 22024 14056 22030
rect 14002 21992 14004 22001
rect 14056 21992 14058 22001
rect 14002 21927 14058 21936
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 13084 21480 13136 21486
rect 13544 21480 13596 21486
rect 13084 21422 13136 21428
rect 13372 21440 13544 21468
rect 13268 21412 13320 21418
rect 13268 21354 13320 21360
rect 12992 20868 13044 20874
rect 12992 20810 13044 20816
rect 12808 20460 12860 20466
rect 12808 20402 12860 20408
rect 12900 20392 12952 20398
rect 12900 20334 12952 20340
rect 12636 19366 12756 19394
rect 12912 19378 12940 20334
rect 13280 19718 13308 21354
rect 13372 20942 13400 21440
rect 13544 21422 13596 21428
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 14016 21010 14044 21286
rect 14094 21040 14150 21049
rect 14004 21004 14056 21010
rect 14200 21026 14228 21490
rect 14936 21146 14964 22238
rect 18972 22228 19024 22234
rect 18972 22170 19024 22176
rect 21732 22228 21784 22234
rect 22376 22238 22428 22244
rect 23664 22296 23716 22302
rect 23756 22296 23808 22302
rect 23664 22238 23716 22244
rect 23754 22264 23756 22273
rect 28540 22296 28592 22302
rect 23808 22264 23810 22273
rect 22282 22199 22338 22208
rect 21732 22170 21784 22176
rect 18512 22092 18564 22098
rect 18512 22034 18564 22040
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 15752 21684 15804 21690
rect 15752 21626 15804 21632
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15016 21480 15068 21486
rect 15016 21422 15068 21428
rect 14924 21140 14976 21146
rect 14924 21082 14976 21088
rect 14150 20998 14228 21026
rect 14646 21040 14702 21049
rect 14094 20975 14150 20984
rect 14702 20998 14780 21026
rect 14646 20975 14702 20984
rect 14004 20946 14056 20952
rect 13360 20936 13412 20942
rect 14096 20936 14148 20942
rect 13360 20878 13412 20884
rect 13740 20884 14096 20890
rect 13740 20878 14148 20884
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 13372 20602 13400 20878
rect 13740 20862 14136 20878
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13372 20233 13400 20538
rect 13358 20224 13414 20233
rect 13358 20159 13414 20168
rect 13740 19938 13768 20862
rect 13818 20768 13874 20777
rect 13818 20703 13874 20712
rect 13832 20466 13860 20703
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 13910 20088 13966 20097
rect 13910 20023 13966 20032
rect 13372 19910 13768 19938
rect 13268 19712 13320 19718
rect 13268 19654 13320 19660
rect 12900 19372 12952 19378
rect 12636 19334 12664 19366
rect 12636 19306 12756 19334
rect 12728 18698 12756 19306
rect 12820 19320 12900 19334
rect 12820 19314 12952 19320
rect 12820 19306 12940 19314
rect 12716 18692 12768 18698
rect 12716 18634 12768 18640
rect 12820 17626 12848 19306
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 13004 18086 13032 19178
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 12636 17598 12848 17626
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 11888 13806 11940 13812
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 12176 13790 12480 13818
rect 11808 13530 11836 13738
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11428 13388 11480 13394
rect 11428 13330 11480 13336
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11256 12986 11284 13262
rect 11348 13025 11376 13262
rect 11334 13016 11390 13025
rect 11244 12980 11296 12986
rect 11334 12951 11390 12960
rect 11244 12922 11296 12928
rect 11150 12880 11206 12889
rect 10876 12844 10928 12850
rect 11150 12815 11206 12824
rect 10876 12786 10928 12792
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10782 11520 10838 11529
rect 10782 11455 10838 11464
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10796 11286 10824 11455
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10336 9722 10364 10542
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10336 8022 10364 9658
rect 10428 9466 10456 10406
rect 10520 9586 10548 11018
rect 10612 10713 10640 11154
rect 10598 10704 10654 10713
rect 10598 10639 10654 10648
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10428 9438 10548 9466
rect 10520 9042 10548 9438
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10520 8129 10548 8978
rect 10612 8906 10640 10066
rect 10704 9353 10732 11154
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10796 9518 10824 9998
rect 10888 9761 10916 12786
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11256 12442 11284 12718
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11150 12336 11206 12345
rect 11150 12271 11152 12280
rect 11204 12271 11206 12280
rect 11152 12242 11204 12248
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10966 11656 11022 11665
rect 10966 11591 11022 11600
rect 10980 11286 11008 11591
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10874 9752 10930 9761
rect 10874 9687 10930 9696
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10690 9344 10746 9353
rect 10690 9279 10746 9288
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10704 8786 10732 9279
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10888 8786 10916 8910
rect 10704 8758 10916 8786
rect 10888 8378 10916 8758
rect 10980 8498 11008 11018
rect 11072 10674 11100 12038
rect 11348 11830 11376 12582
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11164 10810 11192 10950
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11440 10441 11468 13330
rect 11716 12850 11744 13330
rect 11783 13084 12091 13093
rect 11783 13082 11789 13084
rect 11845 13082 11869 13084
rect 11925 13082 11949 13084
rect 12005 13082 12029 13084
rect 12085 13082 12091 13084
rect 11845 13030 11847 13082
rect 12027 13030 12029 13082
rect 11783 13028 11789 13030
rect 11845 13028 11869 13030
rect 11925 13028 11949 13030
rect 12005 13028 12029 13030
rect 12085 13028 12091 13030
rect 11783 13019 12091 13028
rect 12072 12980 12124 12986
rect 12176 12968 12204 13790
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 12124 12940 12204 12968
rect 12072 12922 12124 12928
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11610 12472 11666 12481
rect 11610 12407 11666 12416
rect 11624 12220 11652 12407
rect 11532 12192 11652 12220
rect 11532 11898 11560 12192
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11612 11076 11664 11082
rect 11612 11018 11664 11024
rect 11426 10432 11482 10441
rect 11426 10367 11482 10376
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11164 9674 11192 9862
rect 11164 9646 11284 9674
rect 11256 9586 11284 9646
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11072 9466 11100 9522
rect 11348 9466 11376 9998
rect 11440 9586 11468 9998
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11072 9438 11376 9466
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11348 9382 11376 9438
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11164 8974 11192 9318
rect 11348 9042 11376 9318
rect 11532 9178 11560 9454
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11624 9042 11652 11018
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11612 9036 11664 9042
rect 11612 8978 11664 8984
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11164 8566 11192 8910
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 11348 8430 11376 8774
rect 11532 8634 11560 8910
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11426 8528 11482 8537
rect 11426 8463 11482 8472
rect 11336 8424 11388 8430
rect 10888 8350 11008 8378
rect 11336 8366 11388 8372
rect 10874 8256 10930 8265
rect 10874 8191 10930 8200
rect 10506 8120 10562 8129
rect 10506 8055 10562 8064
rect 10324 8016 10376 8022
rect 10324 7958 10376 7964
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10336 5658 10364 7686
rect 10520 7206 10548 8055
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10428 6254 10456 6598
rect 10520 6338 10548 7142
rect 10612 6458 10640 7822
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10520 6310 10640 6338
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10336 5630 10456 5658
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10244 5370 10272 5510
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10336 2514 10364 5510
rect 10428 4049 10456 5630
rect 10520 4078 10548 6190
rect 10612 6089 10640 6310
rect 10598 6080 10654 6089
rect 10598 6015 10654 6024
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10612 4162 10640 5850
rect 10704 5681 10732 7686
rect 10690 5672 10746 5681
rect 10690 5607 10746 5616
rect 10796 5137 10824 7686
rect 10782 5128 10838 5137
rect 10782 5063 10838 5072
rect 10888 4826 10916 8191
rect 10980 7342 11008 8350
rect 11348 8090 11376 8366
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10980 4826 11008 7278
rect 11164 6866 11192 7822
rect 11256 7478 11284 7890
rect 11348 7886 11376 8026
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11244 7336 11296 7342
rect 11348 7290 11376 7822
rect 11296 7284 11376 7290
rect 11244 7278 11376 7284
rect 11256 7262 11376 7278
rect 11256 6866 11284 7262
rect 11440 7188 11468 8463
rect 11716 8430 11744 12786
rect 11796 12708 11848 12714
rect 11796 12650 11848 12656
rect 11808 12306 11836 12650
rect 11980 12640 12032 12646
rect 12162 12608 12218 12617
rect 11980 12582 12032 12588
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11992 12209 12020 12582
rect 12084 12566 12162 12594
rect 12084 12306 12112 12566
rect 12162 12543 12218 12552
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 11978 12200 12034 12209
rect 11978 12135 12034 12144
rect 11783 11996 12091 12005
rect 11783 11994 11789 11996
rect 11845 11994 11869 11996
rect 11925 11994 11949 11996
rect 12005 11994 12029 11996
rect 12085 11994 12091 11996
rect 11845 11942 11847 11994
rect 12027 11942 12029 11994
rect 11783 11940 11789 11942
rect 11845 11940 11869 11942
rect 11925 11940 11949 11942
rect 12005 11940 12029 11942
rect 12085 11940 12091 11942
rect 11783 11931 12091 11940
rect 12176 11937 12204 12378
rect 12162 11928 12218 11937
rect 12162 11863 12218 11872
rect 12268 11694 12296 13670
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12360 12986 12388 13262
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12452 12306 12480 13262
rect 12636 12424 12664 17598
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12728 16454 12756 17478
rect 13096 17202 13124 18566
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 13188 17746 13216 18022
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 12808 17196 12860 17202
rect 12808 17138 12860 17144
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12820 16794 12848 17138
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 13174 16280 13230 16289
rect 13174 16215 13230 16224
rect 13084 15904 13136 15910
rect 12990 15872 13046 15881
rect 13084 15846 13136 15852
rect 12990 15807 13046 15816
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12728 14006 12756 15438
rect 12808 14952 12860 14958
rect 12806 14920 12808 14929
rect 12860 14920 12862 14929
rect 12806 14855 12862 14864
rect 13004 14618 13032 15807
rect 13096 15706 13124 15846
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13188 14657 13216 16215
rect 13280 15609 13308 18566
rect 13266 15600 13322 15609
rect 13266 15535 13322 15544
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13174 14648 13230 14657
rect 12992 14612 13044 14618
rect 13174 14583 13230 14592
rect 12992 14554 13044 14560
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 13096 13394 13124 13670
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12544 12396 12664 12424
rect 12714 12472 12770 12481
rect 12714 12407 12770 12416
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12346 12064 12402 12073
rect 12346 11999 12402 12008
rect 12360 11898 12388 11999
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 11794 11112 11850 11121
rect 11794 11047 11796 11056
rect 11848 11047 11850 11056
rect 11796 11018 11848 11024
rect 11783 10908 12091 10917
rect 11783 10906 11789 10908
rect 11845 10906 11869 10908
rect 11925 10906 11949 10908
rect 12005 10906 12029 10908
rect 12085 10906 12091 10908
rect 11845 10854 11847 10906
rect 12027 10854 12029 10906
rect 11783 10852 11789 10854
rect 11845 10852 11869 10854
rect 11925 10852 11949 10854
rect 12005 10852 12029 10854
rect 12085 10852 12091 10854
rect 11783 10843 12091 10852
rect 12176 10606 12204 11154
rect 12452 11150 12480 12242
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 12084 10266 12112 10406
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 11783 9820 12091 9829
rect 11783 9818 11789 9820
rect 11845 9818 11869 9820
rect 11925 9818 11949 9820
rect 12005 9818 12029 9820
rect 12085 9818 12091 9820
rect 11845 9766 11847 9818
rect 12027 9766 12029 9818
rect 11783 9764 11789 9766
rect 11845 9764 11869 9766
rect 11925 9764 11949 9766
rect 12005 9764 12029 9766
rect 12085 9764 12091 9766
rect 11783 9755 12091 9764
rect 11783 8732 12091 8741
rect 11783 8730 11789 8732
rect 11845 8730 11869 8732
rect 11925 8730 11949 8732
rect 12005 8730 12029 8732
rect 12085 8730 12091 8732
rect 11845 8678 11847 8730
rect 12027 8678 12029 8730
rect 11783 8676 11789 8678
rect 11845 8676 11869 8678
rect 11925 8676 11949 8678
rect 12005 8676 12029 8678
rect 12085 8676 12091 8678
rect 11783 8667 12091 8676
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 11348 7160 11468 7188
rect 11624 7177 11652 8230
rect 12084 8129 12112 8230
rect 12070 8120 12126 8129
rect 12070 8055 12126 8064
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11796 7880 11848 7886
rect 12176 7868 12204 9862
rect 12268 9024 12296 11018
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12360 10146 12388 10542
rect 12452 10470 12480 11086
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12360 10118 12480 10146
rect 12360 9217 12388 10118
rect 12346 9208 12402 9217
rect 12346 9143 12402 9152
rect 12348 9036 12400 9042
rect 12268 8996 12348 9024
rect 12268 8537 12296 8996
rect 12348 8978 12400 8984
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12254 8528 12310 8537
rect 12254 8463 12310 8472
rect 11848 7840 12204 7868
rect 11796 7822 11848 7828
rect 11716 7206 11744 7822
rect 11783 7644 12091 7653
rect 11783 7642 11789 7644
rect 11845 7642 11869 7644
rect 11925 7642 11949 7644
rect 12005 7642 12029 7644
rect 12085 7642 12091 7644
rect 11845 7590 11847 7642
rect 12027 7590 12029 7642
rect 11783 7588 11789 7590
rect 11845 7588 11869 7590
rect 11925 7588 11949 7590
rect 12005 7588 12029 7590
rect 12085 7588 12091 7590
rect 11783 7579 12091 7588
rect 11704 7200 11756 7206
rect 11610 7168 11666 7177
rect 11348 6866 11376 7160
rect 11704 7142 11756 7148
rect 11610 7103 11666 7112
rect 11716 7002 11744 7142
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 12360 6798 12388 8774
rect 12452 7342 12480 10118
rect 12544 9625 12572 12396
rect 12624 12232 12676 12238
rect 12728 12220 12756 12407
rect 12820 12306 12848 13262
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12912 12442 12940 12718
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12676 12192 12756 12220
rect 12624 12174 12676 12180
rect 12622 11928 12678 11937
rect 12622 11863 12678 11872
rect 12636 10606 12664 11863
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12636 10305 12664 10406
rect 12622 10296 12678 10305
rect 12622 10231 12678 10240
rect 12530 9616 12586 9625
rect 12530 9551 12586 9560
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12348 6792 12400 6798
rect 11058 6760 11114 6769
rect 12348 6734 12400 6740
rect 11058 6695 11114 6704
rect 11072 6662 11100 6695
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11783 6556 12091 6565
rect 11783 6554 11789 6556
rect 11845 6554 11869 6556
rect 11925 6554 11949 6556
rect 12005 6554 12029 6556
rect 12085 6554 12091 6556
rect 11845 6502 11847 6554
rect 12027 6502 12029 6554
rect 11783 6500 11789 6502
rect 11845 6500 11869 6502
rect 11925 6500 11949 6502
rect 12005 6500 12029 6502
rect 12085 6500 12091 6502
rect 11783 6491 12091 6500
rect 12544 6440 12572 8502
rect 12636 7410 12664 9318
rect 12728 9042 12756 11766
rect 12820 11150 12848 12242
rect 12912 11778 12940 12378
rect 13004 11898 13032 13262
rect 13188 12782 13216 14583
rect 13280 14074 13308 15098
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13372 13190 13400 19910
rect 13924 19786 13952 20023
rect 13912 19780 13964 19786
rect 13912 19722 13964 19728
rect 13636 19712 13688 19718
rect 13542 19680 13598 19689
rect 13636 19654 13688 19660
rect 13542 19615 13598 19624
rect 13556 19334 13584 19615
rect 13648 19417 13676 19654
rect 14016 19417 14044 20402
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14096 19780 14148 19786
rect 14096 19722 14148 19728
rect 14108 19514 14136 19722
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 13634 19408 13690 19417
rect 13634 19343 13690 19352
rect 14002 19408 14058 19417
rect 14002 19343 14058 19352
rect 13464 19306 13584 19334
rect 13464 19009 13492 19306
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 13450 19000 13506 19009
rect 13450 18935 13506 18944
rect 13464 18834 13492 18935
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13464 17082 13492 18770
rect 13542 18456 13598 18465
rect 13542 18391 13598 18400
rect 13636 18420 13688 18426
rect 13556 18222 13584 18391
rect 13636 18362 13688 18368
rect 13544 18216 13596 18222
rect 13544 18158 13596 18164
rect 13544 17808 13596 17814
rect 13544 17750 13596 17756
rect 13556 17270 13584 17750
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 13464 17054 13584 17082
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13464 16250 13492 16390
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13556 15978 13584 17054
rect 13648 16998 13676 18362
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13740 16250 13768 18158
rect 13832 17678 13860 18158
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13832 16590 13860 17614
rect 13924 16726 13952 18022
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 14016 16674 14044 19110
rect 14200 18714 14228 19858
rect 14292 19174 14320 20878
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14384 18766 14412 20198
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14372 18760 14424 18766
rect 14278 18728 14334 18737
rect 14108 18686 14278 18714
rect 14108 17338 14136 18686
rect 14372 18702 14424 18708
rect 14278 18663 14334 18672
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14200 17678 14228 18226
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 14016 16646 14136 16674
rect 14200 16658 14228 17614
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13464 15570 13492 15914
rect 13452 15564 13504 15570
rect 13452 15506 13504 15512
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13464 14414 13492 15302
rect 13542 15056 13598 15065
rect 13542 14991 13544 15000
rect 13596 14991 13598 15000
rect 13544 14962 13596 14968
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13740 13938 13768 16186
rect 13832 15570 13860 16526
rect 14004 15972 14056 15978
rect 14004 15914 14056 15920
rect 13820 15564 13872 15570
rect 13872 15524 13952 15552
rect 13820 15506 13872 15512
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13832 14385 13860 14758
rect 13924 14482 13952 15524
rect 14016 15094 14044 15914
rect 14004 15088 14056 15094
rect 14004 15030 14056 15036
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13818 14376 13874 14385
rect 13818 14311 13874 14320
rect 13924 13938 13952 14418
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 14016 14006 14044 14350
rect 14108 14278 14136 16646
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14200 15910 14228 16594
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14292 15978 14320 16390
rect 14280 15972 14332 15978
rect 14280 15914 14332 15920
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14200 15706 14228 15846
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14200 14414 14228 15642
rect 14188 14408 14240 14414
rect 14188 14350 14240 14356
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 13452 13932 13504 13938
rect 13728 13932 13780 13938
rect 13452 13874 13504 13880
rect 13648 13892 13728 13920
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 13096 11898 13124 12582
rect 13268 12436 13320 12442
rect 13268 12378 13320 12384
rect 13280 12238 13308 12378
rect 13372 12238 13400 12854
rect 13464 12782 13492 13874
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13464 12617 13492 12718
rect 13450 12608 13506 12617
rect 13450 12543 13506 12552
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13176 11824 13228 11830
rect 12912 11772 13176 11778
rect 12912 11766 13228 11772
rect 12912 11750 13216 11766
rect 13280 11762 13308 12174
rect 13464 11937 13492 12242
rect 13450 11928 13506 11937
rect 13450 11863 13506 11872
rect 13268 11756 13320 11762
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12820 9722 12848 11086
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12912 10130 12940 10542
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12360 6412 12572 6440
rect 11060 6316 11112 6322
rect 11060 6258 11112 6264
rect 11072 5234 11100 6258
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11164 4865 11192 5034
rect 11150 4856 11206 4865
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10968 4820 11020 4826
rect 11150 4791 11206 4800
rect 10968 4762 11020 4768
rect 11060 4684 11112 4690
rect 10980 4644 11060 4672
rect 10612 4146 10732 4162
rect 10612 4140 10744 4146
rect 10612 4134 10692 4140
rect 10692 4082 10744 4088
rect 10508 4072 10560 4078
rect 10414 4040 10470 4049
rect 10508 4014 10560 4020
rect 10414 3975 10470 3984
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10140 1352 10192 1358
rect 10140 1294 10192 1300
rect 8944 1158 8996 1164
rect 9678 1184 9734 1193
rect 9678 1119 9734 1128
rect 10520 1018 10548 2382
rect 10980 2310 11008 4644
rect 11060 4626 11112 4632
rect 11256 3942 11284 6054
rect 11348 5642 11376 6190
rect 11796 6112 11848 6118
rect 11426 6080 11482 6089
rect 11796 6054 11848 6060
rect 11426 6015 11482 6024
rect 11440 5778 11468 6015
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11440 5522 11468 5714
rect 11348 5494 11468 5522
rect 11348 4826 11376 5494
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11440 4622 11468 5170
rect 11532 5030 11560 5714
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11624 5234 11652 5646
rect 11808 5574 11836 6054
rect 12360 5817 12388 6412
rect 12820 6338 12848 8910
rect 12544 6310 12848 6338
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12346 5808 12402 5817
rect 12452 5778 12480 6054
rect 12346 5743 12402 5752
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11783 5468 12091 5477
rect 11783 5466 11789 5468
rect 11845 5466 11869 5468
rect 11925 5466 11949 5468
rect 12005 5466 12029 5468
rect 12085 5466 12091 5468
rect 11845 5414 11847 5466
rect 12027 5414 12029 5466
rect 11783 5412 11789 5414
rect 11845 5412 11869 5414
rect 11925 5412 11949 5414
rect 12005 5412 12029 5414
rect 12085 5412 12091 5414
rect 11783 5403 12091 5412
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4826 11560 4966
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11532 4706 11560 4762
rect 11532 4678 11652 4706
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11348 3754 11376 3878
rect 11256 3726 11376 3754
rect 11256 3602 11284 3726
rect 11440 3602 11468 4558
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11336 2984 11388 2990
rect 11440 2938 11468 3538
rect 11532 2990 11560 4490
rect 11624 3738 11652 4678
rect 11716 4282 11744 5170
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11900 4690 11928 5102
rect 11978 4856 12034 4865
rect 12034 4814 12112 4842
rect 11978 4791 12034 4800
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 12084 4622 12112 4814
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 11783 4380 12091 4389
rect 11783 4378 11789 4380
rect 11845 4378 11869 4380
rect 11925 4378 11949 4380
rect 12005 4378 12029 4380
rect 12085 4378 12091 4380
rect 11845 4326 11847 4378
rect 12027 4326 12029 4378
rect 11783 4324 11789 4326
rect 11845 4324 11869 4326
rect 11925 4324 11949 4326
rect 12005 4324 12029 4326
rect 12085 4324 12091 4326
rect 11783 4315 12091 4324
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11388 2932 11468 2938
rect 11336 2926 11468 2932
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11348 2910 11468 2926
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11164 1222 11192 2246
rect 11256 1902 11284 2382
rect 11244 1896 11296 1902
rect 11244 1838 11296 1844
rect 11256 1494 11284 1838
rect 11244 1488 11296 1494
rect 11244 1430 11296 1436
rect 11256 1290 11284 1430
rect 11244 1284 11296 1290
rect 11244 1226 11296 1232
rect 11152 1216 11204 1222
rect 11152 1158 11204 1164
rect 11348 1018 11376 2790
rect 11440 2514 11468 2910
rect 11624 2854 11652 3674
rect 12176 3602 12204 4422
rect 12268 4214 12296 4422
rect 12256 4208 12308 4214
rect 12256 4150 12308 4156
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 11783 3292 12091 3301
rect 11783 3290 11789 3292
rect 11845 3290 11869 3292
rect 11925 3290 11949 3292
rect 12005 3290 12029 3292
rect 12085 3290 12091 3292
rect 11845 3238 11847 3290
rect 12027 3238 12029 3290
rect 11783 3236 11789 3238
rect 11845 3236 11869 3238
rect 11925 3236 11949 3238
rect 12005 3236 12029 3238
rect 12085 3236 12091 3238
rect 11783 3227 12091 3236
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11624 2582 11652 2790
rect 12544 2774 12572 6310
rect 12716 6248 12768 6254
rect 12820 6225 12848 6310
rect 12716 6190 12768 6196
rect 12806 6216 12862 6225
rect 12728 5914 12756 6190
rect 12806 6151 12862 6160
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12820 5234 12848 6054
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12452 2746 12572 2774
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 11428 2508 11480 2514
rect 11428 2450 11480 2456
rect 11624 1902 11652 2518
rect 11796 2440 11848 2446
rect 11716 2388 11796 2394
rect 11716 2382 11848 2388
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 11716 2366 11836 2382
rect 11612 1896 11664 1902
rect 11612 1838 11664 1844
rect 11624 1562 11652 1838
rect 11612 1556 11664 1562
rect 11612 1498 11664 1504
rect 11716 1494 11744 2366
rect 11783 2204 12091 2213
rect 11783 2202 11789 2204
rect 11845 2202 11869 2204
rect 11925 2202 11949 2204
rect 12005 2202 12029 2204
rect 12085 2202 12091 2204
rect 11845 2150 11847 2202
rect 12027 2150 12029 2202
rect 11783 2148 11789 2150
rect 11845 2148 11869 2150
rect 11925 2148 11949 2150
rect 12005 2148 12029 2150
rect 12085 2148 12091 2150
rect 11783 2139 12091 2148
rect 12360 2106 12388 2382
rect 12348 2100 12400 2106
rect 12348 2042 12400 2048
rect 11980 1896 12032 1902
rect 11980 1838 12032 1844
rect 12254 1864 12310 1873
rect 11992 1766 12020 1838
rect 12254 1799 12310 1808
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 11704 1488 11756 1494
rect 11426 1456 11482 1465
rect 11704 1430 11756 1436
rect 11426 1391 11482 1400
rect 10508 1012 10560 1018
rect 10508 954 10560 960
rect 11336 1012 11388 1018
rect 11336 954 11388 960
rect 10784 944 10836 950
rect 10784 886 10836 892
rect 8852 876 8904 882
rect 8852 818 8904 824
rect 9220 876 9272 882
rect 9220 818 9272 824
rect 8300 808 8352 814
rect 8300 750 8352 756
rect 9036 808 9088 814
rect 9036 750 9088 756
rect 8392 740 8444 746
rect 8392 682 8444 688
rect 7988 572 8296 581
rect 7988 570 7994 572
rect 8050 570 8074 572
rect 8130 570 8154 572
rect 8210 570 8234 572
rect 8290 570 8296 572
rect 8050 518 8052 570
rect 8232 518 8234 570
rect 7988 516 7994 518
rect 8050 516 8074 518
rect 8130 516 8154 518
rect 8210 516 8234 518
rect 8290 516 8296 518
rect 7988 507 8296 516
rect 8404 406 8432 682
rect 8392 400 8444 406
rect 8392 342 8444 348
rect 9048 338 9076 750
rect 9232 377 9260 818
rect 10796 814 10824 886
rect 11152 876 11204 882
rect 11152 818 11204 824
rect 10784 808 10836 814
rect 10784 750 10836 756
rect 10968 740 11020 746
rect 10968 682 11020 688
rect 10784 672 10836 678
rect 10980 626 11008 682
rect 11164 678 11192 818
rect 10836 620 11008 626
rect 10784 614 11008 620
rect 11152 672 11204 678
rect 11152 614 11204 620
rect 10796 598 11008 614
rect 9218 368 9274 377
rect 9036 332 9088 338
rect 9218 303 9274 312
rect 9036 274 9088 280
rect 11348 270 11376 954
rect 11440 814 11468 1391
rect 12164 1352 12216 1358
rect 12164 1294 12216 1300
rect 11783 1116 12091 1125
rect 11783 1114 11789 1116
rect 11845 1114 11869 1116
rect 11925 1114 11949 1116
rect 12005 1114 12029 1116
rect 12085 1114 12091 1116
rect 11845 1062 11847 1114
rect 12027 1062 12029 1114
rect 11783 1060 11789 1062
rect 11845 1060 11869 1062
rect 11925 1060 11949 1062
rect 12005 1060 12029 1062
rect 12085 1060 12091 1062
rect 11783 1051 12091 1060
rect 11520 876 11572 882
rect 11520 818 11572 824
rect 11428 808 11480 814
rect 11428 750 11480 756
rect 11532 338 11560 818
rect 12176 746 12204 1294
rect 12268 1018 12296 1799
rect 12256 1012 12308 1018
rect 12256 954 12308 960
rect 12452 814 12480 2746
rect 12820 2417 12848 4014
rect 12912 4010 12940 10066
rect 13004 9722 13032 11750
rect 13268 11698 13320 11704
rect 13556 11694 13584 12718
rect 13648 11694 13676 13892
rect 13728 13874 13780 13880
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13726 13832 13782 13841
rect 13726 13767 13728 13776
rect 13780 13767 13782 13776
rect 13728 13738 13780 13744
rect 13740 13376 13768 13738
rect 14200 13734 14228 14350
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 13740 13348 13860 13376
rect 13726 13288 13782 13297
rect 13726 13223 13782 13232
rect 13740 12073 13768 13223
rect 13832 13190 13860 13348
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13726 12064 13782 12073
rect 13726 11999 13782 12008
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13096 11218 13124 11630
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 13556 11014 13584 11630
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13174 10432 13230 10441
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 13096 8974 13124 10406
rect 13174 10367 13230 10376
rect 13188 9586 13216 10367
rect 13372 10266 13400 10678
rect 13832 10674 13860 12786
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13464 10266 13492 10542
rect 13360 10260 13412 10266
rect 13280 10220 13360 10248
rect 13280 9586 13308 10220
rect 13360 10202 13412 10208
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13556 10130 13584 10542
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13188 9353 13216 9386
rect 13174 9344 13230 9353
rect 13174 9279 13230 9288
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 13096 8401 13124 8502
rect 13082 8392 13138 8401
rect 13082 8327 13138 8336
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13188 7546 13216 7686
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 12900 4004 12952 4010
rect 12900 3946 12952 3952
rect 13004 2650 13032 7278
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 13096 6322 13124 7142
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 13096 4690 13124 6054
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13188 3126 13216 7346
rect 13280 7342 13308 9522
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13280 6458 13308 6598
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13372 6322 13400 9386
rect 13464 6458 13492 9658
rect 13556 9586 13584 10066
rect 13924 10062 13952 10406
rect 14016 10062 14044 13126
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14200 12442 14228 12582
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14280 12232 14332 12238
rect 14094 12200 14150 12209
rect 14150 12158 14228 12186
rect 14280 12174 14332 12180
rect 14094 12135 14150 12144
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13556 9042 13584 9522
rect 13924 9382 13952 9998
rect 14108 9586 14136 12038
rect 14200 11762 14228 12158
rect 14292 11762 14320 12174
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14200 10674 14228 10950
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13924 9178 13952 9318
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13556 8498 13584 8978
rect 13924 8498 13952 9114
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13648 7970 13676 8230
rect 13726 7984 13782 7993
rect 13648 7942 13726 7970
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13556 5914 13584 6054
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13648 5234 13676 7942
rect 13726 7919 13728 7928
rect 13780 7919 13782 7928
rect 13728 7890 13780 7896
rect 13820 7744 13872 7750
rect 14200 7721 14228 8366
rect 14384 8265 14412 18702
rect 14476 16592 14504 19654
rect 14556 19236 14608 19242
rect 14556 19178 14608 19184
rect 14568 18873 14596 19178
rect 14554 18864 14610 18873
rect 14554 18799 14610 18808
rect 14660 17184 14688 20334
rect 14752 18630 14780 20998
rect 14936 19310 14964 21082
rect 15028 20942 15056 21422
rect 15396 21321 15424 21490
rect 15764 21486 15792 21626
rect 15752 21480 15804 21486
rect 15752 21422 15804 21428
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 15476 21344 15528 21350
rect 15382 21312 15438 21321
rect 16132 21321 16160 21422
rect 16212 21412 16264 21418
rect 16212 21354 16264 21360
rect 15476 21286 15528 21292
rect 16118 21312 16174 21321
rect 15382 21247 15438 21256
rect 15108 21004 15160 21010
rect 15108 20946 15160 20952
rect 15016 20936 15068 20942
rect 15016 20878 15068 20884
rect 15120 20330 15148 20946
rect 15198 20496 15254 20505
rect 15198 20431 15200 20440
rect 15252 20431 15254 20440
rect 15200 20402 15252 20408
rect 15108 20324 15160 20330
rect 15160 20284 15240 20312
rect 15108 20266 15160 20272
rect 15106 19408 15162 19417
rect 15106 19343 15162 19352
rect 15120 19310 15148 19343
rect 14924 19304 14976 19310
rect 15108 19304 15160 19310
rect 14924 19246 14976 19252
rect 15014 19272 15070 19281
rect 15108 19246 15160 19252
rect 15014 19207 15070 19216
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14924 19168 14976 19174
rect 14924 19110 14976 19116
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14568 17156 14688 17184
rect 14844 17218 14872 19110
rect 14936 18970 14964 19110
rect 15028 18970 15056 19207
rect 15108 19168 15160 19174
rect 15106 19136 15108 19145
rect 15160 19136 15162 19145
rect 15106 19071 15162 19080
rect 15106 19000 15162 19009
rect 14924 18964 14976 18970
rect 14924 18906 14976 18912
rect 15016 18964 15068 18970
rect 15106 18935 15162 18944
rect 15016 18906 15068 18912
rect 15120 17354 15148 18935
rect 15028 17338 15148 17354
rect 15016 17332 15148 17338
rect 15068 17326 15148 17332
rect 15016 17274 15068 17280
rect 14844 17190 15148 17218
rect 14568 16946 14596 17156
rect 14648 17060 14700 17066
rect 14844 17048 14872 17190
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14700 17020 14872 17048
rect 14648 17002 14700 17008
rect 14568 16918 14688 16946
rect 14554 16688 14610 16697
rect 14554 16623 14610 16632
rect 14464 16586 14516 16592
rect 14464 16528 14516 16534
rect 14462 16280 14518 16289
rect 14462 16215 14518 16224
rect 14476 16182 14504 16215
rect 14464 16176 14516 16182
rect 14464 16118 14516 16124
rect 14568 15586 14596 16623
rect 14476 15570 14596 15586
rect 14464 15564 14596 15570
rect 14516 15558 14596 15564
rect 14464 15506 14516 15512
rect 14462 15192 14518 15201
rect 14462 15127 14464 15136
rect 14516 15127 14518 15136
rect 14464 15098 14516 15104
rect 14554 14920 14610 14929
rect 14476 14890 14554 14906
rect 14464 14884 14554 14890
rect 14516 14878 14554 14884
rect 14554 14855 14610 14864
rect 14464 14826 14516 14832
rect 14660 14498 14688 16918
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14752 15502 14780 16050
rect 14936 16046 14964 17070
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14844 15706 14872 15982
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14752 14890 14780 15438
rect 15028 15026 15056 15846
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 15120 14521 15148 17190
rect 15212 16969 15240 20284
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15396 19961 15424 20198
rect 15382 19952 15438 19961
rect 15488 19922 15516 21286
rect 15578 21244 15886 21253
rect 16118 21247 16174 21256
rect 15578 21242 15584 21244
rect 15640 21242 15664 21244
rect 15720 21242 15744 21244
rect 15800 21242 15824 21244
rect 15880 21242 15886 21244
rect 15640 21190 15642 21242
rect 15822 21190 15824 21242
rect 15578 21188 15584 21190
rect 15640 21188 15664 21190
rect 15720 21188 15744 21190
rect 15800 21188 15824 21190
rect 15880 21188 15886 21190
rect 15578 21179 15886 21188
rect 15752 21004 15804 21010
rect 15752 20946 15804 20952
rect 16028 21004 16080 21010
rect 16224 20992 16252 21354
rect 16684 21146 16712 21966
rect 17316 21956 17368 21962
rect 17316 21898 17368 21904
rect 16762 21720 16818 21729
rect 16762 21655 16818 21664
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 16488 21004 16540 21010
rect 16224 20964 16488 20992
rect 16028 20946 16080 20952
rect 16488 20946 16540 20952
rect 15764 20505 15792 20946
rect 15750 20496 15806 20505
rect 15750 20431 15806 20440
rect 15578 20156 15886 20165
rect 15578 20154 15584 20156
rect 15640 20154 15664 20156
rect 15720 20154 15744 20156
rect 15800 20154 15824 20156
rect 15880 20154 15886 20156
rect 15640 20102 15642 20154
rect 15822 20102 15824 20154
rect 15578 20100 15584 20102
rect 15640 20100 15664 20102
rect 15720 20100 15744 20102
rect 15800 20100 15824 20102
rect 15880 20100 15886 20102
rect 15578 20091 15886 20100
rect 15752 19984 15804 19990
rect 15752 19926 15804 19932
rect 15382 19887 15438 19896
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 15304 17882 15332 19790
rect 15764 19553 15792 19926
rect 16040 19718 16068 20946
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 16132 20482 16160 20878
rect 16132 20454 16344 20482
rect 16120 20392 16172 20398
rect 16120 20334 16172 20340
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15750 19544 15806 19553
rect 15750 19479 15806 19488
rect 15936 19440 15988 19446
rect 15936 19382 15988 19388
rect 15384 19236 15436 19242
rect 15436 19196 15516 19224
rect 15384 19178 15436 19184
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15488 17649 15516 19196
rect 15578 19068 15886 19077
rect 15578 19066 15584 19068
rect 15640 19066 15664 19068
rect 15720 19066 15744 19068
rect 15800 19066 15824 19068
rect 15880 19066 15886 19068
rect 15640 19014 15642 19066
rect 15822 19014 15824 19066
rect 15578 19012 15584 19014
rect 15640 19012 15664 19014
rect 15720 19012 15744 19014
rect 15800 19012 15824 19014
rect 15880 19012 15886 19014
rect 15578 19003 15886 19012
rect 15948 18970 15976 19382
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 15948 18442 15976 18770
rect 15856 18414 15976 18442
rect 15856 18086 15884 18414
rect 15936 18352 15988 18358
rect 15936 18294 15988 18300
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15578 17980 15886 17989
rect 15578 17978 15584 17980
rect 15640 17978 15664 17980
rect 15720 17978 15744 17980
rect 15800 17978 15824 17980
rect 15880 17978 15886 17980
rect 15640 17926 15642 17978
rect 15822 17926 15824 17978
rect 15578 17924 15584 17926
rect 15640 17924 15664 17926
rect 15720 17924 15744 17926
rect 15800 17924 15824 17926
rect 15880 17924 15886 17926
rect 15578 17915 15886 17924
rect 15568 17808 15620 17814
rect 15568 17750 15620 17756
rect 15474 17640 15530 17649
rect 15474 17575 15530 17584
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15198 16960 15254 16969
rect 15198 16895 15254 16904
rect 15292 16040 15344 16046
rect 15212 16000 15292 16028
rect 15106 14512 15162 14521
rect 14660 14470 15056 14498
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14556 14408 14608 14414
rect 14556 14350 14608 14356
rect 14476 13530 14504 14350
rect 14568 14074 14596 14350
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14660 11354 14688 14214
rect 14752 13938 14780 14214
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14832 13864 14884 13870
rect 14832 13806 14884 13812
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14648 11348 14700 11354
rect 14648 11290 14700 11296
rect 14752 11200 14780 13194
rect 14844 12306 14872 13806
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14936 13462 14964 13670
rect 14924 13456 14976 13462
rect 14924 13398 14976 13404
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14832 11212 14884 11218
rect 14752 11172 14832 11200
rect 14832 11154 14884 11160
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14660 9586 14688 11018
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14936 9042 14964 11018
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 15028 8548 15056 14470
rect 15212 14482 15240 16000
rect 15292 15982 15344 15988
rect 15396 15366 15424 17478
rect 15488 16658 15516 17575
rect 15580 17202 15608 17750
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15578 16892 15886 16901
rect 15578 16890 15584 16892
rect 15640 16890 15664 16892
rect 15720 16890 15744 16892
rect 15800 16890 15824 16892
rect 15880 16890 15886 16892
rect 15640 16838 15642 16890
rect 15822 16838 15824 16890
rect 15578 16836 15584 16838
rect 15640 16836 15664 16838
rect 15720 16836 15744 16838
rect 15800 16836 15824 16838
rect 15880 16836 15886 16838
rect 15578 16827 15886 16836
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15948 16538 15976 18294
rect 16040 17814 16068 19654
rect 16132 18193 16160 20334
rect 16210 20224 16266 20233
rect 16210 20159 16266 20168
rect 16224 19689 16252 20159
rect 16316 19990 16344 20454
rect 16776 20262 16804 21655
rect 17328 21026 17356 21898
rect 17960 21616 18012 21622
rect 17960 21558 18012 21564
rect 17684 21480 17736 21486
rect 17684 21422 17736 21428
rect 17592 21344 17644 21350
rect 17592 21286 17644 21292
rect 17604 21049 17632 21286
rect 17144 20998 17356 21026
rect 17590 21040 17646 21049
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16304 19984 16356 19990
rect 16304 19926 16356 19932
rect 16210 19680 16266 19689
rect 16210 19615 16266 19624
rect 16316 19394 16344 19926
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16500 19514 16528 19790
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16316 19366 16620 19394
rect 16592 19334 16620 19366
rect 16316 19306 16620 19334
rect 16212 19236 16264 19242
rect 16212 19178 16264 19184
rect 16224 18358 16252 19178
rect 16212 18352 16264 18358
rect 16212 18294 16264 18300
rect 16118 18184 16174 18193
rect 16118 18119 16174 18128
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16028 17808 16080 17814
rect 16028 17750 16080 17756
rect 16224 17678 16252 17818
rect 16316 17746 16344 19306
rect 16776 19174 16804 19654
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16396 19168 16448 19174
rect 16764 19168 16816 19174
rect 16396 19110 16448 19116
rect 16486 19136 16542 19145
rect 16408 18329 16436 19110
rect 16764 19110 16816 19116
rect 16486 19071 16542 19080
rect 16500 18970 16528 19071
rect 16868 18986 16896 19450
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16592 18958 16896 18986
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 16394 18320 16450 18329
rect 16394 18255 16450 18264
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16224 17270 16252 17614
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16212 17264 16264 17270
rect 16212 17206 16264 17212
rect 16210 17096 16266 17105
rect 16210 17031 16266 17040
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16132 16561 16160 16730
rect 16224 16658 16252 17031
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16118 16552 16174 16561
rect 15476 16516 15528 16522
rect 15948 16510 16068 16538
rect 15476 16458 15528 16464
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15304 14550 15332 14894
rect 15292 14544 15344 14550
rect 15292 14486 15344 14492
rect 15106 14447 15162 14456
rect 15200 14476 15252 14482
rect 15120 14056 15148 14447
rect 15200 14418 15252 14424
rect 15120 14028 15240 14056
rect 15106 13968 15162 13977
rect 15106 13903 15162 13912
rect 15120 13394 15148 13903
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15120 12986 15148 13330
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15212 12442 15240 14028
rect 15396 13530 15424 14894
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15488 13394 15516 16458
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 15578 15804 15886 15813
rect 15578 15802 15584 15804
rect 15640 15802 15664 15804
rect 15720 15802 15744 15804
rect 15800 15802 15824 15804
rect 15880 15802 15886 15804
rect 15640 15750 15642 15802
rect 15822 15750 15824 15802
rect 15578 15748 15584 15750
rect 15640 15748 15664 15750
rect 15720 15748 15744 15750
rect 15800 15748 15824 15750
rect 15880 15748 15886 15750
rect 15578 15739 15886 15748
rect 15948 15570 15976 16390
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 16040 15450 16068 16510
rect 16118 16487 16174 16496
rect 16040 15422 16160 15450
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 15844 15156 15896 15162
rect 15896 15116 15976 15144
rect 15844 15098 15896 15104
rect 15578 14716 15886 14725
rect 15578 14714 15584 14716
rect 15640 14714 15664 14716
rect 15720 14714 15744 14716
rect 15800 14714 15824 14716
rect 15880 14714 15886 14716
rect 15640 14662 15642 14714
rect 15822 14662 15824 14714
rect 15578 14660 15584 14662
rect 15640 14660 15664 14662
rect 15720 14660 15744 14662
rect 15800 14660 15824 14662
rect 15880 14660 15886 14662
rect 15578 14651 15886 14660
rect 15578 13628 15886 13637
rect 15578 13626 15584 13628
rect 15640 13626 15664 13628
rect 15720 13626 15744 13628
rect 15800 13626 15824 13628
rect 15880 13626 15886 13628
rect 15640 13574 15642 13626
rect 15822 13574 15824 13626
rect 15578 13572 15584 13574
rect 15640 13572 15664 13574
rect 15720 13572 15744 13574
rect 15800 13572 15824 13574
rect 15880 13572 15886 13574
rect 15578 13563 15886 13572
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15200 12436 15252 12442
rect 15488 12434 15516 13330
rect 15578 12540 15886 12549
rect 15578 12538 15584 12540
rect 15640 12538 15664 12540
rect 15720 12538 15744 12540
rect 15800 12538 15824 12540
rect 15880 12538 15886 12540
rect 15640 12486 15642 12538
rect 15822 12486 15824 12538
rect 15578 12484 15584 12486
rect 15640 12484 15664 12486
rect 15720 12484 15744 12486
rect 15800 12484 15824 12486
rect 15880 12484 15886 12486
rect 15578 12475 15886 12484
rect 15948 12442 15976 15116
rect 16040 14006 16068 15302
rect 16132 14482 16160 15422
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16132 14385 16160 14418
rect 16118 14376 16174 14385
rect 16118 14311 16174 14320
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 15200 12378 15252 12384
rect 15396 12406 15516 12434
rect 15936 12436 15988 12442
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15212 8974 15240 11494
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15108 8560 15160 8566
rect 15028 8520 15108 8548
rect 15108 8502 15160 8508
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 15120 8401 15148 8502
rect 15106 8392 15162 8401
rect 15106 8327 15162 8336
rect 14556 8288 14608 8294
rect 14370 8256 14426 8265
rect 14556 8230 14608 8236
rect 14370 8191 14426 8200
rect 14568 7750 14596 8230
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14556 7744 14608 7750
rect 13820 7686 13872 7692
rect 14186 7712 14242 7721
rect 13726 6896 13782 6905
rect 13832 6866 13860 7686
rect 14556 7686 14608 7692
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14186 7647 14242 7656
rect 14464 7336 14516 7342
rect 14384 7296 14464 7324
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 13910 6896 13966 6905
rect 13726 6831 13782 6840
rect 13820 6860 13872 6866
rect 13740 6662 13768 6831
rect 14200 6866 14228 7142
rect 13910 6831 13912 6840
rect 13820 6802 13872 6808
rect 13964 6831 13966 6840
rect 14188 6860 14240 6866
rect 13912 6802 13964 6808
rect 14188 6802 14240 6808
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 14384 6322 14412 7296
rect 14568 7324 14596 7686
rect 14516 7296 14596 7324
rect 14464 7278 14516 7284
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14372 6316 14424 6322
rect 14372 6258 14424 6264
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13740 5370 13768 5714
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13636 5228 13688 5234
rect 13556 5188 13636 5216
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 13176 2916 13228 2922
rect 13176 2858 13228 2864
rect 12992 2644 13044 2650
rect 12992 2586 13044 2592
rect 12806 2408 12862 2417
rect 12806 2343 12862 2352
rect 12716 944 12768 950
rect 12716 886 12768 892
rect 12256 808 12308 814
rect 12256 750 12308 756
rect 12440 808 12492 814
rect 12440 750 12492 756
rect 12164 740 12216 746
rect 12164 682 12216 688
rect 11520 332 11572 338
rect 11520 274 11572 280
rect 11336 264 11388 270
rect 6642 232 6698 241
rect 6092 196 6144 202
rect 11336 206 11388 212
rect 12268 202 12296 750
rect 6642 167 6698 176
rect 12256 196 12308 202
rect 6092 138 6144 144
rect 12256 138 12308 144
rect 12452 66 12480 750
rect 12728 270 12756 886
rect 12820 678 12848 2343
rect 13188 1018 13216 2858
rect 13360 1284 13412 1290
rect 13360 1226 13412 1232
rect 13176 1012 13228 1018
rect 13176 954 13228 960
rect 13372 814 13400 1226
rect 13556 814 13584 5188
rect 13636 5170 13688 5176
rect 13832 5166 13860 5646
rect 13924 5166 13952 6122
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5778 14504 6054
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13648 4826 13676 4966
rect 13740 4826 13768 4966
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13832 4622 13860 5102
rect 14016 5030 14044 5646
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14016 4622 14044 4966
rect 14292 4622 14320 5510
rect 14568 5234 14596 6394
rect 14660 6225 14688 6394
rect 14752 6322 14780 7686
rect 14844 7206 14872 8026
rect 14832 7200 14884 7206
rect 15016 7200 15068 7206
rect 14832 7142 14884 7148
rect 14922 7168 14978 7177
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14646 6216 14702 6225
rect 14646 6151 14702 6160
rect 14844 6118 14872 7142
rect 14978 7148 15016 7154
rect 14978 7142 15068 7148
rect 14978 7126 15056 7142
rect 14922 7103 14978 7112
rect 15212 6322 15240 8502
rect 15304 7410 15332 10406
rect 15396 10248 15424 12406
rect 15936 12378 15988 12384
rect 15844 12232 15896 12238
rect 15842 12200 15844 12209
rect 15896 12200 15898 12209
rect 15842 12135 15898 12144
rect 15856 11694 15884 12135
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15578 11452 15886 11461
rect 15578 11450 15584 11452
rect 15640 11450 15664 11452
rect 15720 11450 15744 11452
rect 15800 11450 15824 11452
rect 15880 11450 15886 11452
rect 15640 11398 15642 11450
rect 15822 11398 15824 11450
rect 15578 11396 15584 11398
rect 15640 11396 15664 11398
rect 15720 11396 15744 11398
rect 15800 11396 15824 11398
rect 15880 11396 15886 11398
rect 15578 11387 15886 11396
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15488 11082 15516 11154
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15948 10713 15976 11494
rect 15934 10704 15990 10713
rect 15934 10639 15990 10648
rect 15578 10364 15886 10373
rect 15578 10362 15584 10364
rect 15640 10362 15664 10364
rect 15720 10362 15744 10364
rect 15800 10362 15824 10364
rect 15880 10362 15886 10364
rect 15640 10310 15642 10362
rect 15822 10310 15824 10362
rect 15578 10308 15584 10310
rect 15640 10308 15664 10310
rect 15720 10308 15744 10310
rect 15800 10308 15824 10310
rect 15880 10308 15886 10310
rect 15578 10299 15886 10308
rect 15476 10260 15528 10266
rect 15396 10220 15476 10248
rect 15476 10202 15528 10208
rect 15948 10130 15976 10639
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15396 7886 15424 9862
rect 15488 9722 15516 10066
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15488 9042 15516 9658
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 15578 9276 15886 9285
rect 15578 9274 15584 9276
rect 15640 9274 15664 9276
rect 15720 9274 15744 9276
rect 15800 9274 15824 9276
rect 15880 9274 15886 9276
rect 15640 9222 15642 9274
rect 15822 9222 15824 9274
rect 15578 9220 15584 9222
rect 15640 9220 15664 9222
rect 15720 9220 15744 9222
rect 15800 9220 15824 9222
rect 15880 9220 15886 9222
rect 15578 9211 15886 9220
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15476 8900 15528 8906
rect 15476 8842 15528 8848
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15488 6322 15516 8842
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15580 8566 15608 8774
rect 15568 8560 15620 8566
rect 15568 8502 15620 8508
rect 15672 8430 15700 9114
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15578 8188 15886 8197
rect 15578 8186 15584 8188
rect 15640 8186 15664 8188
rect 15720 8186 15744 8188
rect 15800 8186 15824 8188
rect 15880 8186 15886 8188
rect 15640 8134 15642 8186
rect 15822 8134 15824 8186
rect 15578 8132 15584 8134
rect 15640 8132 15664 8134
rect 15720 8132 15744 8134
rect 15800 8132 15824 8134
rect 15880 8132 15886 8134
rect 15578 8123 15886 8132
rect 15660 7744 15712 7750
rect 15566 7712 15622 7721
rect 15660 7686 15712 7692
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15566 7647 15622 7656
rect 15580 7410 15608 7647
rect 15672 7449 15700 7686
rect 15764 7546 15792 7686
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15658 7440 15714 7449
rect 15568 7404 15620 7410
rect 15658 7375 15714 7384
rect 15568 7346 15620 7352
rect 15578 7100 15886 7109
rect 15578 7098 15584 7100
rect 15640 7098 15664 7100
rect 15720 7098 15744 7100
rect 15800 7098 15824 7100
rect 15880 7098 15886 7100
rect 15640 7046 15642 7098
rect 15822 7046 15824 7098
rect 15578 7044 15584 7046
rect 15640 7044 15664 7046
rect 15720 7044 15744 7046
rect 15800 7044 15824 7046
rect 15880 7044 15886 7046
rect 15578 7035 15886 7044
rect 15948 6866 15976 9386
rect 16040 8634 16068 12650
rect 16132 11642 16160 14311
rect 16224 13190 16252 16594
rect 16316 16561 16344 17546
rect 16302 16552 16358 16561
rect 16302 16487 16358 16496
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16316 13394 16344 14214
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16408 12866 16436 18022
rect 16500 16250 16528 18566
rect 16592 17882 16620 18958
rect 16670 18864 16726 18873
rect 16670 18799 16726 18808
rect 16684 17882 16712 18799
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 16776 17921 16804 18702
rect 16854 18320 16910 18329
rect 17144 18290 17172 20998
rect 17590 20975 17646 20984
rect 17696 20874 17724 21422
rect 17972 21418 18000 21558
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 17960 21412 18012 21418
rect 17960 21354 18012 21360
rect 17972 21026 18000 21354
rect 18236 21344 18288 21350
rect 18340 21321 18368 21422
rect 18236 21286 18288 21292
rect 18326 21312 18382 21321
rect 17972 20998 18184 21026
rect 18050 20904 18106 20913
rect 17684 20868 17736 20874
rect 18050 20839 18106 20848
rect 17684 20810 17736 20816
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 16854 18255 16910 18264
rect 17040 18284 17092 18290
rect 16868 18222 16896 18255
rect 17040 18226 17092 18232
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 17052 18170 17080 18226
rect 17130 18184 17186 18193
rect 17052 18142 17130 18170
rect 17130 18119 17186 18128
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 16762 17912 16818 17921
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16672 17876 16724 17882
rect 16762 17847 16818 17856
rect 16672 17818 16724 17824
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16684 17134 16712 17614
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16684 16590 16712 17070
rect 16868 16998 16896 17614
rect 17144 17202 17172 18022
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 16868 16640 16896 16934
rect 17052 16794 17080 16934
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 17040 16652 17092 16658
rect 16868 16612 17040 16640
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16856 16040 16908 16046
rect 16856 15982 16908 15988
rect 16868 15609 16896 15982
rect 16960 15638 16988 16612
rect 17040 16594 17092 16600
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 17038 16144 17094 16153
rect 17038 16079 17094 16088
rect 16948 15632 17000 15638
rect 16854 15600 16910 15609
rect 16948 15574 17000 15580
rect 17052 15570 17080 16079
rect 17144 15910 17172 16526
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 16854 15535 16910 15544
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 17144 15502 17172 15846
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16578 14920 16634 14929
rect 16578 14855 16634 14864
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16500 14618 16528 14758
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16592 13394 16620 14855
rect 16684 14414 16712 15302
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16776 14618 16804 14758
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16684 13734 16712 14350
rect 16776 13938 16804 14418
rect 16868 14074 16896 15302
rect 17130 15056 17186 15065
rect 17130 14991 17132 15000
rect 17184 14991 17186 15000
rect 17132 14962 17184 14968
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16672 13728 16724 13734
rect 16672 13670 16724 13676
rect 16776 13462 16804 13874
rect 16960 13841 16988 14894
rect 16946 13832 17002 13841
rect 16946 13767 17002 13776
rect 16764 13456 16816 13462
rect 16764 13398 16816 13404
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16960 13308 16988 13767
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17144 13326 17172 13670
rect 16776 13280 16988 13308
rect 17132 13320 17184 13326
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16408 12838 16528 12866
rect 16396 12776 16448 12782
rect 16396 12718 16448 12724
rect 16132 11614 16252 11642
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16132 11354 16160 11494
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16224 11082 16252 11614
rect 16212 11076 16264 11082
rect 16264 11036 16344 11064
rect 16212 11018 16264 11024
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16132 9178 16160 9862
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 16040 8090 16068 8230
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 15658 6760 15714 6769
rect 15658 6695 15660 6704
rect 15712 6695 15714 6704
rect 15660 6666 15712 6672
rect 16040 6458 16068 6802
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 15578 6012 15886 6021
rect 15578 6010 15584 6012
rect 15640 6010 15664 6012
rect 15720 6010 15744 6012
rect 15800 6010 15824 6012
rect 15880 6010 15886 6012
rect 15640 5958 15642 6010
rect 15822 5958 15824 6010
rect 15578 5956 15584 5958
rect 15640 5956 15664 5958
rect 15720 5956 15744 5958
rect 15800 5956 15824 5958
rect 15880 5956 15886 5958
rect 15578 5947 15886 5956
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 13832 4146 13860 4558
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13832 3534 13860 4082
rect 14016 3534 14044 4558
rect 14660 4146 15240 4162
rect 14648 4140 15240 4146
rect 14700 4134 15240 4140
rect 14648 4082 14700 4088
rect 15212 4078 15240 4134
rect 14832 4072 14884 4078
rect 14752 4032 14832 4060
rect 14200 3590 14412 3618
rect 13820 3528 13872 3534
rect 14004 3528 14056 3534
rect 13872 3476 13952 3482
rect 13820 3470 13952 3476
rect 14004 3470 14056 3476
rect 13832 3454 13952 3470
rect 13924 2990 13952 3454
rect 14016 3398 14044 3470
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13820 2440 13872 2446
rect 13924 2428 13952 2926
rect 13872 2400 13952 2428
rect 13820 2382 13872 2388
rect 13924 1902 13952 2400
rect 13912 1896 13964 1902
rect 13912 1838 13964 1844
rect 13820 1352 13872 1358
rect 13924 1340 13952 1838
rect 13872 1312 13952 1340
rect 13820 1294 13872 1300
rect 13820 1216 13872 1222
rect 13820 1158 13872 1164
rect 13728 944 13780 950
rect 13832 898 13860 1158
rect 14200 1018 14228 3590
rect 14384 3534 14412 3590
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14476 2854 14504 3334
rect 14752 3097 14780 4032
rect 14832 4014 14884 4020
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 14738 3088 14794 3097
rect 14738 3023 14794 3032
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 14292 1902 14320 2586
rect 14384 2530 14412 2790
rect 14476 2650 14504 2790
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14384 2514 14504 2530
rect 14384 2508 14516 2514
rect 14384 2502 14464 2508
rect 14464 2450 14516 2456
rect 14280 1896 14332 1902
rect 14280 1838 14332 1844
rect 14648 1896 14700 1902
rect 14648 1838 14700 1844
rect 14292 1562 14320 1838
rect 14280 1556 14332 1562
rect 14280 1498 14332 1504
rect 14372 1352 14424 1358
rect 14372 1294 14424 1300
rect 14188 1012 14240 1018
rect 14188 954 14240 960
rect 13780 892 13860 898
rect 13728 886 13860 892
rect 13740 870 13860 886
rect 14280 876 14332 882
rect 14280 818 14332 824
rect 13360 808 13412 814
rect 13360 750 13412 756
rect 13544 808 13596 814
rect 13544 750 13596 756
rect 12808 672 12860 678
rect 12808 614 12860 620
rect 12820 406 12848 614
rect 12808 400 12860 406
rect 12808 342 12860 348
rect 14292 338 14320 818
rect 14384 474 14412 1294
rect 14660 1222 14688 1838
rect 14752 1465 14780 3023
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 15120 2106 15148 2790
rect 15108 2100 15160 2106
rect 15108 2042 15160 2048
rect 14738 1456 14794 1465
rect 14738 1391 14794 1400
rect 14648 1216 14700 1222
rect 14648 1158 14700 1164
rect 14464 808 14516 814
rect 14464 750 14516 756
rect 14556 808 14608 814
rect 14556 750 14608 756
rect 14372 468 14424 474
rect 14372 410 14424 416
rect 14280 332 14332 338
rect 14280 274 14332 280
rect 12716 264 12768 270
rect 12716 206 12768 212
rect 14476 202 14504 750
rect 14568 474 14596 750
rect 15292 672 15344 678
rect 15292 614 15344 620
rect 14556 468 14608 474
rect 14556 410 14608 416
rect 14464 196 14516 202
rect 14464 138 14516 144
rect 15304 105 15332 614
rect 15488 134 15516 5510
rect 15578 4924 15886 4933
rect 15578 4922 15584 4924
rect 15640 4922 15664 4924
rect 15720 4922 15744 4924
rect 15800 4922 15824 4924
rect 15880 4922 15886 4924
rect 15640 4870 15642 4922
rect 15822 4870 15824 4922
rect 15578 4868 15584 4870
rect 15640 4868 15664 4870
rect 15720 4868 15744 4870
rect 15800 4868 15824 4870
rect 15880 4868 15886 4870
rect 15578 4859 15886 4868
rect 16132 4060 16160 8978
rect 16224 8022 16252 10202
rect 16316 8022 16344 11036
rect 16408 10713 16436 12718
rect 16500 12434 16528 12838
rect 16684 12753 16712 13126
rect 16670 12744 16726 12753
rect 16670 12679 16726 12688
rect 16580 12436 16632 12442
rect 16500 12406 16580 12434
rect 16580 12378 16632 12384
rect 16592 12238 16620 12378
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16684 11150 16712 11630
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16394 10704 16450 10713
rect 16394 10639 16450 10648
rect 16408 10588 16436 10639
rect 16488 10600 16540 10606
rect 16408 10560 16488 10588
rect 16488 10542 16540 10548
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16212 8016 16264 8022
rect 16212 7958 16264 7964
rect 16304 8016 16356 8022
rect 16304 7958 16356 7964
rect 16408 7954 16436 9998
rect 16500 9042 16528 10542
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16210 7848 16266 7857
rect 16210 7783 16266 7792
rect 16224 7546 16252 7783
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16394 6896 16450 6905
rect 16394 6831 16396 6840
rect 16448 6831 16450 6840
rect 16396 6802 16448 6808
rect 16396 6724 16448 6730
rect 16396 6666 16448 6672
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16224 6458 16252 6598
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16224 5250 16252 5646
rect 16408 5574 16436 6666
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16224 5222 16344 5250
rect 16316 5166 16344 5222
rect 16304 5160 16356 5166
rect 16356 5108 16436 5114
rect 16304 5102 16436 5108
rect 16316 5086 16436 5102
rect 16408 4622 16436 5086
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16212 4072 16264 4078
rect 16132 4032 16212 4060
rect 16212 4014 16264 4020
rect 15578 3836 15886 3845
rect 15578 3834 15584 3836
rect 15640 3834 15664 3836
rect 15720 3834 15744 3836
rect 15800 3834 15824 3836
rect 15880 3834 15886 3836
rect 15640 3782 15642 3834
rect 15822 3782 15824 3834
rect 15578 3780 15584 3782
rect 15640 3780 15664 3782
rect 15720 3780 15744 3782
rect 15800 3780 15824 3782
rect 15880 3780 15886 3782
rect 15578 3771 15886 3780
rect 16224 3738 16252 4014
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15948 3194 15976 3334
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 15578 2748 15886 2757
rect 15578 2746 15584 2748
rect 15640 2746 15664 2748
rect 15720 2746 15744 2748
rect 15800 2746 15824 2748
rect 15880 2746 15886 2748
rect 15640 2694 15642 2746
rect 15822 2694 15824 2746
rect 15578 2692 15584 2694
rect 15640 2692 15664 2694
rect 15720 2692 15744 2694
rect 15800 2692 15824 2694
rect 15880 2692 15886 2694
rect 15578 2683 15886 2692
rect 16040 2446 16068 2926
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 16040 1970 16068 2382
rect 16028 1964 16080 1970
rect 16028 1906 16080 1912
rect 15578 1660 15886 1669
rect 15578 1658 15584 1660
rect 15640 1658 15664 1660
rect 15720 1658 15744 1660
rect 15800 1658 15824 1660
rect 15880 1658 15886 1660
rect 15640 1606 15642 1658
rect 15822 1606 15824 1658
rect 15578 1604 15584 1606
rect 15640 1604 15664 1606
rect 15720 1604 15744 1606
rect 15800 1604 15824 1606
rect 15880 1604 15886 1606
rect 15578 1595 15886 1604
rect 16040 1358 16068 1906
rect 16316 1850 16344 3946
rect 16408 3942 16436 4558
rect 16500 4078 16528 8774
rect 16592 7342 16620 11086
rect 16776 10810 16804 13280
rect 17132 13262 17184 13268
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16684 9908 16712 10406
rect 16776 10010 16804 10610
rect 16868 10470 16896 12582
rect 17236 12434 17264 20198
rect 17696 19990 17724 20810
rect 18064 20806 18092 20839
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17684 19984 17736 19990
rect 17684 19926 17736 19932
rect 17696 19514 17724 19926
rect 17972 19854 18000 20198
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17684 19508 17736 19514
rect 17684 19450 17736 19456
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17316 19304 17368 19310
rect 17314 19272 17316 19281
rect 17408 19304 17460 19310
rect 17368 19272 17370 19281
rect 17408 19246 17460 19252
rect 17314 19207 17370 19216
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 17328 17882 17356 18226
rect 17316 17876 17368 17882
rect 17316 17818 17368 17824
rect 17420 16289 17448 19246
rect 17774 19136 17830 19145
rect 17774 19071 17830 19080
rect 17788 18970 17816 19071
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17498 18592 17554 18601
rect 17498 18527 17554 18536
rect 17512 18057 17540 18527
rect 17498 18048 17554 18057
rect 17498 17983 17554 17992
rect 17406 16280 17462 16289
rect 17406 16215 17462 16224
rect 17406 16144 17462 16153
rect 17512 16130 17540 17983
rect 17512 16102 17632 16130
rect 17406 16079 17462 16088
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17328 15026 17356 15438
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17328 14482 17356 14962
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17420 13190 17448 16079
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17328 12628 17356 12922
rect 17408 12640 17460 12646
rect 17328 12600 17408 12628
rect 17408 12582 17460 12588
rect 17236 12406 17356 12434
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17052 11762 17080 12038
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17144 11150 17172 11494
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 16960 10810 16988 11086
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16960 10130 16988 10746
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 17052 10130 17080 10406
rect 17144 10266 17172 11086
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 16776 9982 17080 10010
rect 16948 9920 17000 9926
rect 16684 9880 16896 9908
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16776 9081 16804 9454
rect 16762 9072 16818 9081
rect 16672 9036 16724 9042
rect 16762 9007 16818 9016
rect 16672 8978 16724 8984
rect 16684 8634 16712 8978
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16684 7993 16712 8026
rect 16670 7984 16726 7993
rect 16670 7919 16726 7928
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16776 7342 16804 7686
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16776 6798 16804 7142
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16672 6656 16724 6662
rect 16868 6644 16896 9880
rect 16948 9862 17000 9868
rect 16960 9042 16988 9862
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16672 6598 16724 6604
rect 16776 6616 16896 6644
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16592 5030 16620 5646
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16684 4486 16712 6598
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 16776 3942 16804 6616
rect 17052 6390 17080 9982
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17144 9178 17172 9454
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17236 9178 17264 9318
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17130 9072 17186 9081
rect 17130 9007 17186 9016
rect 17144 8974 17172 9007
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17144 8498 17172 8910
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17222 7848 17278 7857
rect 17328 7834 17356 12406
rect 17420 12306 17448 12582
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17512 11801 17540 15982
rect 17604 14958 17632 16102
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17498 11792 17554 11801
rect 17498 11727 17554 11736
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17278 7806 17356 7834
rect 17222 7783 17278 7792
rect 17512 7750 17540 10610
rect 17590 9480 17646 9489
rect 17590 9415 17646 9424
rect 17604 8634 17632 9415
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17592 8424 17644 8430
rect 17592 8366 17644 8372
rect 17604 8090 17632 8366
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 17132 7336 17184 7342
rect 17132 7278 17184 7284
rect 17500 7336 17552 7342
rect 17500 7278 17552 7284
rect 17590 7304 17646 7313
rect 17144 6934 17172 7278
rect 17132 6928 17184 6934
rect 17132 6870 17184 6876
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17130 6488 17186 6497
rect 17130 6423 17186 6432
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 17144 6254 17172 6423
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 16868 5778 16896 6054
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16960 5234 16988 6054
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16868 4826 16896 4966
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16408 3534 16436 3878
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16408 3194 16436 3470
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16316 1822 16436 1850
rect 16028 1352 16080 1358
rect 16028 1294 16080 1300
rect 16304 1216 16356 1222
rect 16304 1158 16356 1164
rect 16316 814 16344 1158
rect 16408 950 16436 1822
rect 16396 944 16448 950
rect 16396 886 16448 892
rect 16304 808 16356 814
rect 16304 750 16356 756
rect 16396 808 16448 814
rect 16500 762 16528 3674
rect 16684 3602 16712 3878
rect 16776 3641 16804 3878
rect 16868 3777 16896 4762
rect 17236 4690 17264 6054
rect 17328 5030 17356 6734
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17420 6361 17448 6598
rect 17406 6352 17462 6361
rect 17406 6287 17462 6296
rect 17512 6254 17540 7278
rect 17590 7239 17646 7248
rect 17604 7206 17632 7239
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17696 6882 17724 18702
rect 17972 18442 18000 19450
rect 18156 19378 18184 20998
rect 18248 20777 18276 21286
rect 18326 21247 18382 21256
rect 18340 21078 18368 21247
rect 18328 21072 18380 21078
rect 18328 21014 18380 21020
rect 18234 20768 18290 20777
rect 18234 20703 18290 20712
rect 18418 20496 18474 20505
rect 18418 20431 18474 20440
rect 18234 19544 18290 19553
rect 18234 19479 18290 19488
rect 18248 19378 18276 19479
rect 18144 19372 18196 19378
rect 18144 19314 18196 19320
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18432 19310 18460 20431
rect 18524 19310 18552 22034
rect 18616 21622 18644 22034
rect 18604 21616 18656 21622
rect 18604 21558 18656 21564
rect 18984 21010 19012 22170
rect 21638 22128 21694 22137
rect 21638 22063 21694 22072
rect 20812 21956 20864 21962
rect 20812 21898 20864 21904
rect 21364 21956 21416 21962
rect 21364 21898 21416 21904
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 19373 21788 19681 21797
rect 19373 21786 19379 21788
rect 19435 21786 19459 21788
rect 19515 21786 19539 21788
rect 19595 21786 19619 21788
rect 19675 21786 19681 21788
rect 19435 21734 19437 21786
rect 19617 21734 19619 21786
rect 19373 21732 19379 21734
rect 19435 21732 19459 21734
rect 19515 21732 19539 21734
rect 19595 21732 19619 21734
rect 19675 21732 19681 21734
rect 19373 21723 19681 21732
rect 20732 21622 20760 21830
rect 20824 21622 20852 21898
rect 20720 21616 20772 21622
rect 20720 21558 20772 21564
rect 20812 21616 20864 21622
rect 20812 21558 20864 21564
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 20444 21480 20496 21486
rect 20444 21422 20496 21428
rect 19076 21146 19104 21422
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 19352 21078 19380 21422
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 19340 21072 19392 21078
rect 19340 21014 19392 21020
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 18972 21004 19024 21010
rect 18972 20946 19024 20952
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 18512 19304 18564 19310
rect 18512 19246 18564 19252
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 17880 18426 18000 18442
rect 17868 18420 18000 18426
rect 17920 18414 18000 18420
rect 18052 18420 18104 18426
rect 17868 18362 17920 18368
rect 18052 18362 18104 18368
rect 17960 18080 18012 18086
rect 17960 18022 18012 18028
rect 17972 16794 18000 18022
rect 18064 17338 18092 18362
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 18156 12434 18184 18566
rect 18340 18290 18368 19110
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18340 17542 18368 18226
rect 18432 17898 18460 19246
rect 18510 17912 18566 17921
rect 18432 17870 18510 17898
rect 18510 17847 18566 17856
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18616 17338 18644 20334
rect 18708 20330 18736 20742
rect 18696 20324 18748 20330
rect 18696 20266 18748 20272
rect 18708 19310 18736 20266
rect 18696 19304 18748 19310
rect 18696 19246 18748 19252
rect 18708 18766 18736 19246
rect 18800 18766 18828 20946
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19260 20466 19288 20878
rect 19373 20700 19681 20709
rect 19373 20698 19379 20700
rect 19435 20698 19459 20700
rect 19515 20698 19539 20700
rect 19595 20698 19619 20700
rect 19675 20698 19681 20700
rect 19435 20646 19437 20698
rect 19617 20646 19619 20698
rect 19373 20644 19379 20646
rect 19435 20644 19459 20646
rect 19515 20644 19539 20646
rect 19595 20644 19619 20646
rect 19675 20644 19681 20646
rect 19373 20635 19681 20644
rect 19982 20632 20038 20641
rect 19812 20590 19982 20618
rect 19064 20460 19116 20466
rect 19064 20402 19116 20408
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 19076 20058 19104 20402
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 18892 19961 18920 19994
rect 18878 19952 18934 19961
rect 18878 19887 18934 19896
rect 18972 19712 19024 19718
rect 18972 19654 19024 19660
rect 18984 18834 19012 19654
rect 19168 19514 19196 20266
rect 19812 19990 19840 20590
rect 19982 20567 20038 20576
rect 19982 20496 20038 20505
rect 19982 20431 20038 20440
rect 19800 19984 19852 19990
rect 19800 19926 19852 19932
rect 19373 19612 19681 19621
rect 19373 19610 19379 19612
rect 19435 19610 19459 19612
rect 19515 19610 19539 19612
rect 19595 19610 19619 19612
rect 19675 19610 19681 19612
rect 19435 19558 19437 19610
rect 19617 19558 19619 19610
rect 19373 19556 19379 19558
rect 19435 19556 19459 19558
rect 19515 19556 19539 19558
rect 19595 19556 19619 19558
rect 19675 19556 19681 19558
rect 19373 19547 19681 19556
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19706 19408 19762 19417
rect 19340 19372 19392 19378
rect 19706 19343 19762 19352
rect 19340 19314 19392 19320
rect 19352 19281 19380 19314
rect 19338 19272 19394 19281
rect 19338 19207 19394 19216
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18800 17746 18828 18702
rect 19373 18524 19681 18533
rect 19373 18522 19379 18524
rect 19435 18522 19459 18524
rect 19515 18522 19539 18524
rect 19595 18522 19619 18524
rect 19675 18522 19681 18524
rect 19435 18470 19437 18522
rect 19617 18470 19619 18522
rect 19373 18468 19379 18470
rect 19435 18468 19459 18470
rect 19515 18468 19539 18470
rect 19595 18468 19619 18470
rect 19675 18468 19681 18470
rect 19246 18456 19302 18465
rect 19373 18459 19681 18468
rect 19246 18391 19302 18400
rect 19260 18358 19288 18391
rect 19248 18352 19300 18358
rect 19720 18306 19748 19343
rect 19812 18902 19840 19926
rect 19892 19304 19944 19310
rect 19892 19246 19944 19252
rect 19800 18896 19852 18902
rect 19800 18838 19852 18844
rect 19248 18294 19300 18300
rect 19536 18278 19748 18306
rect 18788 17740 18840 17746
rect 18788 17682 18840 17688
rect 18800 17626 18828 17682
rect 19536 17678 19564 18278
rect 19812 18154 19840 18838
rect 19904 18358 19932 19246
rect 19892 18352 19944 18358
rect 19892 18294 19944 18300
rect 19616 18148 19668 18154
rect 19616 18090 19668 18096
rect 19800 18148 19852 18154
rect 19800 18090 19852 18096
rect 18708 17598 18828 17626
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19628 17626 19656 18090
rect 19996 18086 20024 20431
rect 20088 19922 20116 21286
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 20180 21049 20208 21082
rect 20260 21072 20312 21078
rect 20166 21040 20222 21049
rect 20260 21014 20312 21020
rect 20166 20975 20222 20984
rect 20180 19922 20208 20975
rect 20272 20330 20300 21014
rect 20260 20324 20312 20330
rect 20260 20266 20312 20272
rect 20272 19922 20300 20266
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20180 19802 20208 19858
rect 20180 19774 20300 19802
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 20088 17746 20116 19246
rect 20180 19242 20208 19654
rect 20168 19236 20220 19242
rect 20168 19178 20220 19184
rect 20180 18222 20208 19178
rect 20272 19174 20300 19774
rect 20456 19310 20484 21422
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20824 21146 20852 21286
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 21180 20936 21232 20942
rect 21180 20878 21232 20884
rect 21192 20466 21220 20878
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 20626 20360 20682 20369
rect 20626 20295 20682 20304
rect 20640 19990 20668 20295
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20628 19712 20680 19718
rect 20732 19689 20760 19994
rect 21088 19916 21140 19922
rect 21088 19858 21140 19864
rect 21100 19825 21128 19858
rect 21086 19816 21142 19825
rect 21086 19751 21142 19760
rect 20628 19654 20680 19660
rect 20718 19680 20774 19689
rect 20534 19408 20590 19417
rect 20534 19343 20590 19352
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20456 18834 20484 19110
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20168 18216 20220 18222
rect 20168 18158 20220 18164
rect 20076 17740 20128 17746
rect 20076 17682 20128 17688
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 19628 17598 19932 17626
rect 18604 17332 18656 17338
rect 18604 17274 18656 17280
rect 18708 17134 18736 17598
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 19156 17536 19208 17542
rect 19156 17478 19208 17484
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18432 16590 18460 16934
rect 18800 16697 18828 17478
rect 19168 16794 19196 17478
rect 19373 17436 19681 17445
rect 19373 17434 19379 17436
rect 19435 17434 19459 17436
rect 19515 17434 19539 17436
rect 19595 17434 19619 17436
rect 19675 17434 19681 17436
rect 19435 17382 19437 17434
rect 19617 17382 19619 17434
rect 19373 17380 19379 17382
rect 19435 17380 19459 17382
rect 19515 17380 19539 17382
rect 19595 17380 19619 17382
rect 19675 17380 19681 17382
rect 19373 17371 19681 17380
rect 19430 16960 19486 16969
rect 19430 16895 19486 16904
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 18786 16688 18842 16697
rect 18786 16623 18842 16632
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 19444 16522 19472 16895
rect 19432 16516 19484 16522
rect 19432 16458 19484 16464
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 19156 16448 19208 16454
rect 19156 16390 19208 16396
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 18432 16250 18460 16390
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18248 14074 18276 15642
rect 18604 15428 18656 15434
rect 18604 15370 18656 15376
rect 18328 14544 18380 14550
rect 18326 14512 18328 14521
rect 18380 14512 18382 14521
rect 18326 14447 18382 14456
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18156 12406 18276 12434
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17880 11830 17908 12174
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 17972 11762 18000 12174
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17788 9722 17816 9998
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17880 9178 17908 11630
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17960 8560 18012 8566
rect 17960 8502 18012 8508
rect 17774 7712 17830 7721
rect 17774 7647 17830 7656
rect 17788 7546 17816 7647
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17788 7002 17816 7142
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17604 6866 17724 6882
rect 17592 6860 17724 6866
rect 17644 6854 17724 6860
rect 17776 6860 17828 6866
rect 17592 6802 17644 6808
rect 17776 6802 17828 6808
rect 17788 6390 17816 6802
rect 17776 6384 17828 6390
rect 17776 6326 17828 6332
rect 17972 6254 18000 8502
rect 18064 6662 18092 9862
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18156 6254 18184 7890
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 17972 5522 18000 6190
rect 18052 6112 18104 6118
rect 18052 6054 18104 6060
rect 17696 5494 18000 5522
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 16854 3768 16910 3777
rect 16854 3703 16856 3712
rect 16908 3703 16910 3712
rect 16856 3674 16908 3680
rect 16762 3632 16818 3641
rect 16672 3596 16724 3602
rect 16762 3567 16818 3576
rect 16672 3538 16724 3544
rect 16672 1896 16724 1902
rect 16672 1838 16724 1844
rect 16684 1018 16712 1838
rect 16672 1012 16724 1018
rect 16672 954 16724 960
rect 16448 756 16528 762
rect 16396 750 16528 756
rect 16408 734 16528 750
rect 15578 572 15886 581
rect 15578 570 15584 572
rect 15640 570 15664 572
rect 15720 570 15744 572
rect 15800 570 15824 572
rect 15880 570 15886 572
rect 15640 518 15642 570
rect 15822 518 15824 570
rect 15578 516 15584 518
rect 15640 516 15664 518
rect 15720 516 15744 518
rect 15800 516 15824 518
rect 15880 516 15886 518
rect 15578 507 15886 516
rect 15568 264 15620 270
rect 15568 206 15620 212
rect 15476 128 15528 134
rect 15290 96 15346 105
rect 3974 31 4030 40
rect 5540 60 5592 66
rect 5540 2 5592 8
rect 12440 60 12492 66
rect 15580 105 15608 206
rect 15476 70 15528 76
rect 15566 96 15622 105
rect 15290 31 15346 40
rect 16408 66 16436 734
rect 16776 678 16804 3567
rect 16868 2854 16896 3674
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16868 2650 16896 2790
rect 17696 2774 17724 5494
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 17788 4078 17816 4762
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17880 3641 17908 4082
rect 17866 3632 17922 3641
rect 17866 3567 17922 3576
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17696 2746 17816 2774
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 16868 1766 16896 2586
rect 16856 1760 16908 1766
rect 16856 1702 16908 1708
rect 17132 1760 17184 1766
rect 17132 1702 17184 1708
rect 16868 1562 16896 1702
rect 16856 1556 16908 1562
rect 16856 1498 16908 1504
rect 16856 1352 16908 1358
rect 16856 1294 16908 1300
rect 16868 1018 16896 1294
rect 16856 1012 16908 1018
rect 16856 954 16908 960
rect 17144 882 17172 1702
rect 17788 1222 17816 2746
rect 17972 2106 18000 3470
rect 18064 3398 18092 6054
rect 18156 3913 18184 6190
rect 18142 3904 18198 3913
rect 18142 3839 18198 3848
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18064 3097 18092 3334
rect 18050 3088 18106 3097
rect 18050 3023 18106 3032
rect 17960 2100 18012 2106
rect 17960 2042 18012 2048
rect 17866 1456 17922 1465
rect 17866 1391 17922 1400
rect 17776 1216 17828 1222
rect 17776 1158 17828 1164
rect 17880 882 17908 1391
rect 17132 876 17184 882
rect 17132 818 17184 824
rect 17868 876 17920 882
rect 17868 818 17920 824
rect 16764 672 16816 678
rect 16764 614 16816 620
rect 17868 672 17920 678
rect 17868 614 17920 620
rect 17880 202 17908 614
rect 18248 241 18276 12406
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18340 11898 18368 12038
rect 18432 11898 18460 12174
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18616 11354 18644 15370
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18800 14521 18828 14894
rect 18786 14512 18842 14521
rect 18786 14447 18842 14456
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18708 13394 18736 13942
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18800 12646 18828 14447
rect 18984 14346 19012 15302
rect 19076 15026 19104 15846
rect 19168 15570 19196 16390
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19260 15434 19288 16390
rect 19373 16348 19681 16357
rect 19373 16346 19379 16348
rect 19435 16346 19459 16348
rect 19515 16346 19539 16348
rect 19595 16346 19619 16348
rect 19675 16346 19681 16348
rect 19435 16294 19437 16346
rect 19617 16294 19619 16346
rect 19373 16292 19379 16294
rect 19435 16292 19459 16294
rect 19515 16292 19539 16294
rect 19595 16292 19619 16294
rect 19675 16292 19681 16294
rect 19373 16283 19681 16292
rect 19800 15496 19852 15502
rect 19720 15444 19800 15450
rect 19720 15438 19852 15444
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19720 15422 19840 15438
rect 19373 15260 19681 15269
rect 19373 15258 19379 15260
rect 19435 15258 19459 15260
rect 19515 15258 19539 15260
rect 19595 15258 19619 15260
rect 19675 15258 19681 15260
rect 19435 15206 19437 15258
rect 19617 15206 19619 15258
rect 19373 15204 19379 15206
rect 19435 15204 19459 15206
rect 19515 15204 19539 15206
rect 19595 15204 19619 15206
rect 19675 15204 19681 15206
rect 19373 15195 19681 15204
rect 19720 15026 19748 15422
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 18972 14340 19024 14346
rect 18972 14282 19024 14288
rect 19076 14074 19104 14758
rect 19260 14618 19288 14758
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19156 14544 19208 14550
rect 19156 14486 19208 14492
rect 19168 14346 19196 14486
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 19373 14172 19681 14181
rect 19373 14170 19379 14172
rect 19435 14170 19459 14172
rect 19515 14170 19539 14172
rect 19595 14170 19619 14172
rect 19675 14170 19681 14172
rect 19435 14118 19437 14170
rect 19617 14118 19619 14170
rect 19373 14116 19379 14118
rect 19435 14116 19459 14118
rect 19515 14116 19539 14118
rect 19595 14116 19619 14118
rect 19675 14116 19681 14118
rect 19373 14107 19681 14116
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19720 13841 19748 14350
rect 19338 13832 19394 13841
rect 19706 13832 19762 13841
rect 19394 13790 19472 13818
rect 19338 13767 19394 13776
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 18970 13424 19026 13433
rect 18970 13359 19026 13368
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18892 12434 18920 12582
rect 18708 12406 18920 12434
rect 18708 12306 18736 12406
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18696 11756 18748 11762
rect 18696 11698 18748 11704
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18708 11082 18736 11698
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 11354 18828 11494
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18696 11076 18748 11082
rect 18748 11036 18828 11064
rect 18696 11018 18748 11024
rect 18800 10538 18828 11036
rect 18984 11014 19012 13359
rect 19352 13172 19380 13670
rect 19444 13326 19472 13790
rect 19706 13767 19762 13776
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19260 13144 19380 13172
rect 19708 13184 19760 13190
rect 19260 12900 19288 13144
rect 19708 13126 19760 13132
rect 19373 13084 19681 13093
rect 19373 13082 19379 13084
rect 19435 13082 19459 13084
rect 19515 13082 19539 13084
rect 19595 13082 19619 13084
rect 19675 13082 19681 13084
rect 19435 13030 19437 13082
rect 19617 13030 19619 13082
rect 19373 13028 19379 13030
rect 19435 13028 19459 13030
rect 19515 13028 19539 13030
rect 19595 13028 19619 13030
rect 19675 13028 19681 13030
rect 19373 13019 19681 13028
rect 19720 12918 19748 13126
rect 19340 12912 19392 12918
rect 19260 12872 19340 12900
rect 19340 12854 19392 12860
rect 19708 12912 19760 12918
rect 19708 12854 19760 12860
rect 19064 12776 19116 12782
rect 19064 12718 19116 12724
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19076 12442 19104 12718
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 19064 12232 19116 12238
rect 19352 12186 19380 12582
rect 19064 12174 19116 12180
rect 19076 11558 19104 12174
rect 19260 12158 19380 12186
rect 19260 11778 19288 12158
rect 19444 12102 19472 12718
rect 19812 12646 19840 15302
rect 19904 13326 19932 17598
rect 20272 17338 20300 17682
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19996 16833 20024 17138
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 19982 16824 20038 16833
rect 19982 16759 20038 16768
rect 20088 16658 20116 16934
rect 20076 16652 20128 16658
rect 20076 16594 20128 16600
rect 20168 15972 20220 15978
rect 20168 15914 20220 15920
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19892 12912 19944 12918
rect 19996 12900 20024 13806
rect 19944 12872 20024 12900
rect 19892 12854 19944 12860
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19904 12238 19932 12854
rect 20088 12782 20116 14758
rect 20180 13190 20208 15914
rect 20350 15464 20406 15473
rect 20272 15422 20350 15450
rect 20272 13410 20300 15422
rect 20350 15399 20406 15408
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20364 13530 20392 13670
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20272 13382 20392 13410
rect 20168 13184 20220 13190
rect 20168 13126 20220 13132
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20076 12776 20128 12782
rect 20074 12744 20076 12753
rect 20128 12744 20130 12753
rect 20074 12679 20130 12688
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19996 12186 20024 12582
rect 20180 12442 20208 12786
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20272 12442 20300 12718
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 19996 12158 20208 12186
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19373 11996 19681 12005
rect 19373 11994 19379 11996
rect 19435 11994 19459 11996
rect 19515 11994 19539 11996
rect 19595 11994 19619 11996
rect 19675 11994 19681 11996
rect 19435 11942 19437 11994
rect 19617 11942 19619 11994
rect 19373 11940 19379 11942
rect 19435 11940 19459 11942
rect 19515 11940 19539 11942
rect 19595 11940 19619 11942
rect 19675 11940 19681 11942
rect 19373 11931 19681 11940
rect 19260 11762 19380 11778
rect 19260 11756 19392 11762
rect 19260 11750 19340 11756
rect 19340 11698 19392 11704
rect 19892 11688 19944 11694
rect 19892 11630 19944 11636
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 19076 11286 19104 11494
rect 19064 11280 19116 11286
rect 19064 11222 19116 11228
rect 19524 11212 19576 11218
rect 19260 11172 19524 11200
rect 19156 11144 19208 11150
rect 19076 11104 19156 11132
rect 18972 11008 19024 11014
rect 18972 10950 19024 10956
rect 18696 10532 18748 10538
rect 18696 10474 18748 10480
rect 18788 10532 18840 10538
rect 18788 10474 18840 10480
rect 18708 10198 18736 10474
rect 18696 10192 18748 10198
rect 18696 10134 18748 10140
rect 18800 10062 18828 10474
rect 19076 10266 19104 11104
rect 19156 11086 19208 11092
rect 19260 10810 19288 11172
rect 19524 11154 19576 11160
rect 19373 10908 19681 10917
rect 19373 10906 19379 10908
rect 19435 10906 19459 10908
rect 19515 10906 19539 10908
rect 19595 10906 19619 10908
rect 19675 10906 19681 10908
rect 19435 10854 19437 10906
rect 19617 10854 19619 10906
rect 19373 10852 19379 10854
rect 19435 10852 19459 10854
rect 19515 10852 19539 10854
rect 19595 10852 19619 10854
rect 19675 10852 19681 10854
rect 19373 10843 19681 10852
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19904 10674 19932 11630
rect 19892 10668 19944 10674
rect 19892 10610 19944 10616
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 19168 9722 19196 10542
rect 19616 10464 19668 10470
rect 19616 10406 19668 10412
rect 19628 10198 19656 10406
rect 19616 10192 19668 10198
rect 19616 10134 19668 10140
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19536 9926 19564 10066
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19373 9820 19681 9829
rect 19373 9818 19379 9820
rect 19435 9818 19459 9820
rect 19515 9818 19539 9820
rect 19595 9818 19619 9820
rect 19675 9818 19681 9820
rect 19435 9766 19437 9818
rect 19617 9766 19619 9818
rect 19373 9764 19379 9766
rect 19435 9764 19459 9766
rect 19515 9764 19539 9766
rect 19595 9764 19619 9766
rect 19675 9764 19681 9766
rect 19373 9755 19681 9764
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 18616 8634 18644 9386
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18708 8498 18736 9454
rect 19352 9382 19380 9454
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19076 9058 19104 9318
rect 19444 9178 19472 9454
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19156 9104 19208 9110
rect 19076 9052 19156 9058
rect 19076 9046 19208 9052
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 19076 9030 19196 9046
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18420 8424 18472 8430
rect 18420 8366 18472 8372
rect 18432 7886 18460 8366
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18432 7342 18460 7822
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 18432 6798 18460 7278
rect 18524 7002 18552 7346
rect 18604 7268 18656 7274
rect 18604 7210 18656 7216
rect 18616 7154 18644 7210
rect 18800 7154 18828 8978
rect 19076 8498 19104 9030
rect 19720 8906 19748 10066
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19248 8832 19300 8838
rect 19248 8774 19300 8780
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 19156 8492 19208 8498
rect 19260 8480 19288 8774
rect 19373 8732 19681 8741
rect 19373 8730 19379 8732
rect 19435 8730 19459 8732
rect 19515 8730 19539 8732
rect 19595 8730 19619 8732
rect 19675 8730 19681 8732
rect 19435 8678 19437 8730
rect 19617 8678 19619 8730
rect 19373 8676 19379 8678
rect 19435 8676 19459 8678
rect 19515 8676 19539 8678
rect 19595 8676 19619 8678
rect 19675 8676 19681 8678
rect 19373 8667 19681 8676
rect 19340 8492 19392 8498
rect 19260 8452 19340 8480
rect 19156 8434 19208 8440
rect 19340 8434 19392 8440
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 19076 8090 19104 8230
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18892 7721 18920 7822
rect 18878 7712 18934 7721
rect 18878 7647 18934 7656
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18616 7126 18828 7154
rect 18708 7002 18736 7126
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18602 6896 18658 6905
rect 18602 6831 18658 6840
rect 18616 6798 18644 6831
rect 18420 6792 18472 6798
rect 18604 6792 18656 6798
rect 18472 6752 18552 6780
rect 18420 6734 18472 6740
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18432 5658 18460 6598
rect 18524 6338 18552 6752
rect 18604 6734 18656 6740
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18708 6390 18736 6734
rect 18696 6384 18748 6390
rect 18524 6310 18644 6338
rect 18696 6326 18748 6332
rect 18616 6254 18644 6310
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18892 5794 18920 7482
rect 19076 7410 19104 8026
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18984 6497 19012 6734
rect 18970 6488 19026 6497
rect 18970 6423 19026 6432
rect 19076 6118 19104 7346
rect 19168 6662 19196 8434
rect 19373 7644 19681 7653
rect 19373 7642 19379 7644
rect 19435 7642 19459 7644
rect 19515 7642 19539 7644
rect 19595 7642 19619 7644
rect 19675 7642 19681 7644
rect 19435 7590 19437 7642
rect 19617 7590 19619 7642
rect 19373 7588 19379 7590
rect 19435 7588 19459 7590
rect 19515 7588 19539 7590
rect 19595 7588 19619 7590
rect 19675 7588 19681 7590
rect 19373 7579 19681 7588
rect 19720 6866 19748 8842
rect 19904 8090 19932 9454
rect 19996 9042 20024 9862
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19996 7562 20024 8978
rect 19904 7546 20024 7562
rect 19892 7540 20024 7546
rect 19944 7534 20024 7540
rect 19892 7482 19944 7488
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 19708 6860 19760 6866
rect 19708 6802 19760 6808
rect 19246 6760 19302 6769
rect 19246 6695 19302 6704
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 19260 6322 19288 6695
rect 19373 6556 19681 6565
rect 19373 6554 19379 6556
rect 19435 6554 19459 6556
rect 19515 6554 19539 6556
rect 19595 6554 19619 6556
rect 19675 6554 19681 6556
rect 19435 6502 19437 6554
rect 19617 6502 19619 6554
rect 19373 6500 19379 6502
rect 19435 6500 19459 6502
rect 19515 6500 19539 6502
rect 19595 6500 19619 6502
rect 19675 6500 19681 6502
rect 19373 6491 19681 6500
rect 19248 6316 19300 6322
rect 19248 6258 19300 6264
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 19064 6112 19116 6118
rect 19064 6054 19116 6060
rect 18708 5766 18920 5794
rect 18432 5630 18644 5658
rect 18616 5574 18644 5630
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 18340 5098 18368 5510
rect 18328 5092 18380 5098
rect 18328 5034 18380 5040
rect 18340 4486 18368 5034
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18340 3534 18368 4422
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18512 2984 18564 2990
rect 18340 2932 18512 2938
rect 18340 2926 18564 2932
rect 18340 2910 18552 2926
rect 18340 2446 18368 2910
rect 18616 2774 18644 5510
rect 18708 4078 18736 5766
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18800 5030 18828 5646
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18800 4622 18828 4966
rect 18984 4690 19012 6054
rect 19373 5468 19681 5477
rect 19373 5466 19379 5468
rect 19435 5466 19459 5468
rect 19515 5466 19539 5468
rect 19595 5466 19619 5468
rect 19675 5466 19681 5468
rect 19435 5414 19437 5466
rect 19617 5414 19619 5466
rect 19373 5412 19379 5414
rect 19435 5412 19459 5414
rect 19515 5412 19539 5414
rect 19595 5412 19619 5414
rect 19675 5412 19681 5414
rect 19373 5403 19681 5412
rect 19246 5128 19302 5137
rect 19168 5086 19246 5114
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18788 4616 18840 4622
rect 18788 4558 18840 4564
rect 18800 4146 18828 4558
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18696 3528 18748 3534
rect 18800 3516 18828 4082
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 18892 3777 18920 3946
rect 18878 3768 18934 3777
rect 18878 3703 18934 3712
rect 19076 3602 19104 4422
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 18748 3488 18828 3516
rect 18696 3470 18748 3476
rect 18800 2922 18828 3488
rect 18970 3496 19026 3505
rect 18970 3431 19026 3440
rect 18788 2916 18840 2922
rect 18788 2858 18840 2864
rect 18524 2746 18644 2774
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 18340 1902 18368 2382
rect 18524 1902 18552 2746
rect 18800 2650 18828 2858
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 18800 1902 18828 2586
rect 18328 1896 18380 1902
rect 18328 1838 18380 1844
rect 18512 1896 18564 1902
rect 18512 1838 18564 1844
rect 18788 1896 18840 1902
rect 18788 1838 18840 1844
rect 18340 1358 18368 1838
rect 18800 1562 18828 1838
rect 18788 1556 18840 1562
rect 18788 1498 18840 1504
rect 18328 1352 18380 1358
rect 18328 1294 18380 1300
rect 18984 950 19012 3431
rect 19168 2774 19196 5086
rect 19246 5063 19302 5072
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19260 4214 19288 4558
rect 19373 4380 19681 4389
rect 19373 4378 19379 4380
rect 19435 4378 19459 4380
rect 19515 4378 19539 4380
rect 19595 4378 19619 4380
rect 19675 4378 19681 4380
rect 19435 4326 19437 4378
rect 19617 4326 19619 4378
rect 19373 4324 19379 4326
rect 19435 4324 19459 4326
rect 19515 4324 19539 4326
rect 19595 4324 19619 4326
rect 19675 4324 19681 4326
rect 19373 4315 19681 4324
rect 19248 4208 19300 4214
rect 19248 4150 19300 4156
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 19248 4004 19300 4010
rect 19248 3946 19300 3952
rect 19260 3398 19288 3946
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19260 3058 19288 3334
rect 19373 3292 19681 3301
rect 19373 3290 19379 3292
rect 19435 3290 19459 3292
rect 19515 3290 19539 3292
rect 19595 3290 19619 3292
rect 19675 3290 19681 3292
rect 19435 3238 19437 3290
rect 19617 3238 19619 3290
rect 19373 3236 19379 3238
rect 19435 3236 19459 3238
rect 19515 3236 19539 3238
rect 19595 3236 19619 3238
rect 19675 3236 19681 3238
rect 19373 3227 19681 3236
rect 19812 3194 19840 3878
rect 19904 3602 19932 4014
rect 19892 3596 19944 3602
rect 19892 3538 19944 3544
rect 19892 3460 19944 3466
rect 19892 3402 19944 3408
rect 19800 3188 19852 3194
rect 19800 3130 19852 3136
rect 19338 3088 19394 3097
rect 19248 3052 19300 3058
rect 19904 3074 19932 3402
rect 19338 3023 19340 3032
rect 19248 2994 19300 3000
rect 19392 3023 19394 3032
rect 19720 3046 19932 3074
rect 19340 2994 19392 3000
rect 19168 2746 19288 2774
rect 19260 1766 19288 2746
rect 19373 2204 19681 2213
rect 19373 2202 19379 2204
rect 19435 2202 19459 2204
rect 19515 2202 19539 2204
rect 19595 2202 19619 2204
rect 19675 2202 19681 2204
rect 19435 2150 19437 2202
rect 19617 2150 19619 2202
rect 19373 2148 19379 2150
rect 19435 2148 19459 2150
rect 19515 2148 19539 2150
rect 19595 2148 19619 2150
rect 19675 2148 19681 2150
rect 19373 2139 19681 2148
rect 19432 1896 19484 1902
rect 19432 1838 19484 1844
rect 19248 1760 19300 1766
rect 19248 1702 19300 1708
rect 19338 1592 19394 1601
rect 19444 1562 19472 1838
rect 19338 1527 19394 1536
rect 19432 1556 19484 1562
rect 19352 1306 19380 1527
rect 19432 1498 19484 1504
rect 19260 1278 19380 1306
rect 19260 1000 19288 1278
rect 19373 1116 19681 1125
rect 19373 1114 19379 1116
rect 19435 1114 19459 1116
rect 19515 1114 19539 1116
rect 19595 1114 19619 1116
rect 19675 1114 19681 1116
rect 19435 1062 19437 1114
rect 19617 1062 19619 1114
rect 19373 1060 19379 1062
rect 19435 1060 19459 1062
rect 19515 1060 19539 1062
rect 19595 1060 19619 1062
rect 19675 1060 19681 1062
rect 19373 1051 19681 1060
rect 19260 972 19380 1000
rect 18972 944 19024 950
rect 18972 886 19024 892
rect 19352 882 19380 972
rect 19720 882 19748 3046
rect 20088 1766 20116 6938
rect 20180 5273 20208 12158
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20272 10266 20300 10542
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20258 10160 20314 10169
rect 20258 10095 20260 10104
rect 20312 10095 20314 10104
rect 20260 10066 20312 10072
rect 20364 8906 20392 13382
rect 20456 9178 20484 18770
rect 20548 18442 20576 19343
rect 20640 18970 20668 19654
rect 20718 19615 20774 19624
rect 20812 19304 20864 19310
rect 20812 19246 20864 19252
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20824 18766 20852 19246
rect 21272 18896 21324 18902
rect 21272 18838 21324 18844
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20548 18414 20668 18442
rect 21284 18426 21312 18838
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20548 17134 20576 18226
rect 20640 17241 20668 18414
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 20718 18320 20774 18329
rect 20718 18255 20774 18264
rect 20732 17785 20760 18255
rect 20812 18080 20864 18086
rect 20996 18080 21048 18086
rect 20812 18022 20864 18028
rect 20902 18048 20958 18057
rect 20718 17776 20774 17785
rect 20718 17711 20774 17720
rect 20626 17232 20682 17241
rect 20626 17167 20682 17176
rect 20824 17134 20852 18022
rect 20958 18028 20996 18034
rect 20958 18022 21048 18028
rect 20958 18006 21036 18022
rect 20902 17983 20958 17992
rect 21086 17776 21142 17785
rect 21086 17711 21142 17720
rect 21100 17202 21128 17711
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 21192 17513 21220 17546
rect 21178 17504 21234 17513
rect 21178 17439 21234 17448
rect 21178 17232 21234 17241
rect 21088 17196 21140 17202
rect 21178 17167 21180 17176
rect 21088 17138 21140 17144
rect 21232 17167 21234 17176
rect 21180 17138 21232 17144
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20812 17128 20864 17134
rect 20812 17070 20864 17076
rect 20548 16590 20576 17070
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21086 16688 21142 16697
rect 21086 16623 21088 16632
rect 21140 16623 21142 16632
rect 21088 16594 21140 16600
rect 20536 16584 20588 16590
rect 20904 16584 20956 16590
rect 20536 16526 20588 16532
rect 20718 16552 20774 16561
rect 20904 16526 20956 16532
rect 20718 16487 20774 16496
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20548 16153 20576 16186
rect 20732 16182 20760 16487
rect 20720 16176 20772 16182
rect 20534 16144 20590 16153
rect 20720 16118 20772 16124
rect 20534 16079 20590 16088
rect 20916 16046 20944 16526
rect 21192 16454 21220 16730
rect 21284 16590 21312 17614
rect 21376 16658 21404 21898
rect 21456 21888 21508 21894
rect 21456 21830 21508 21836
rect 21468 21554 21496 21830
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21548 20392 21600 20398
rect 21548 20334 21600 20340
rect 21560 19990 21588 20334
rect 21548 19984 21600 19990
rect 21548 19926 21600 19932
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21468 18426 21496 18702
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21652 17762 21680 22063
rect 21744 18222 21772 22170
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 21836 20913 21864 21966
rect 22388 21894 22416 22238
rect 22468 22160 22520 22166
rect 22744 22160 22796 22166
rect 22468 22102 22520 22108
rect 22558 22128 22614 22137
rect 22376 21888 22428 21894
rect 21914 21856 21970 21865
rect 22376 21830 22428 21836
rect 21914 21791 21970 21800
rect 21928 21690 21956 21791
rect 22098 21720 22154 21729
rect 21916 21684 21968 21690
rect 22098 21655 22154 21664
rect 21916 21626 21968 21632
rect 22008 21548 22060 21554
rect 22112 21536 22140 21655
rect 22060 21508 22140 21536
rect 22008 21490 22060 21496
rect 22192 21480 22244 21486
rect 22309 21480 22361 21486
rect 22192 21422 22244 21428
rect 22296 21428 22309 21468
rect 22296 21422 22361 21428
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 22020 21162 22048 21286
rect 22020 21134 22140 21162
rect 22204 21146 22232 21422
rect 21822 20904 21878 20913
rect 21822 20839 21878 20848
rect 21822 20632 21878 20641
rect 21822 20567 21878 20576
rect 21916 20596 21968 20602
rect 21836 20330 21864 20567
rect 21916 20538 21968 20544
rect 22008 20596 22060 20602
rect 22008 20538 22060 20544
rect 21928 20369 21956 20538
rect 21914 20360 21970 20369
rect 21824 20324 21876 20330
rect 21914 20295 21970 20304
rect 21824 20266 21876 20272
rect 22020 20074 22048 20538
rect 21928 20046 22048 20074
rect 22112 20074 22140 21134
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22296 20448 22324 21422
rect 22204 20420 22324 20448
rect 22204 20262 22232 20420
rect 22282 20360 22338 20369
rect 22338 20318 22416 20346
rect 22282 20295 22338 20304
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22112 20046 22324 20074
rect 21928 19514 21956 20046
rect 22008 19916 22060 19922
rect 22008 19858 22060 19864
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 22020 18766 22048 19858
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22112 19514 22140 19654
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22204 19394 22232 19654
rect 22112 19366 22232 19394
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 21822 18456 21878 18465
rect 21822 18391 21878 18400
rect 21732 18216 21784 18222
rect 21732 18158 21784 18164
rect 21836 18034 21864 18391
rect 21560 17734 21680 17762
rect 21744 18006 21864 18034
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21468 17134 21496 17614
rect 21560 17542 21588 17734
rect 21548 17536 21600 17542
rect 21548 17478 21600 17484
rect 21638 17368 21694 17377
rect 21638 17303 21694 17312
rect 21456 17128 21508 17134
rect 21456 17070 21508 17076
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21468 16590 21496 17070
rect 21272 16584 21324 16590
rect 21272 16526 21324 16532
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 21180 16448 21232 16454
rect 21468 16436 21496 16526
rect 21180 16390 21232 16396
rect 21284 16408 21496 16436
rect 20812 16040 20864 16046
rect 20812 15982 20864 15988
rect 20904 16040 20956 16046
rect 20904 15982 20956 15988
rect 20824 14822 20852 15982
rect 20916 15502 20944 15982
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 20902 15192 20958 15201
rect 20902 15127 20958 15136
rect 20916 15026 20944 15127
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 20824 14618 20852 14758
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20548 11898 20576 13874
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20720 13864 20772 13870
rect 20720 13806 20772 13812
rect 20640 12850 20668 13806
rect 20732 13530 20760 13806
rect 20812 13728 20864 13734
rect 20812 13670 20864 13676
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20640 12442 20668 12786
rect 20824 12646 20852 13670
rect 20916 13394 20944 14758
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 21008 12102 21036 15302
rect 21100 13138 21128 16390
rect 21284 16114 21312 16408
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 21364 15564 21416 15570
rect 21468 15552 21496 16408
rect 21548 15564 21600 15570
rect 21468 15524 21548 15552
rect 21364 15506 21416 15512
rect 21548 15506 21600 15512
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21284 14482 21312 15438
rect 21376 15162 21404 15506
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 21272 14476 21324 14482
rect 21272 14418 21324 14424
rect 21468 14006 21496 14894
rect 21652 14550 21680 17303
rect 21640 14544 21692 14550
rect 21640 14486 21692 14492
rect 21548 14272 21600 14278
rect 21548 14214 21600 14220
rect 21456 14000 21508 14006
rect 21456 13942 21508 13948
rect 21560 13841 21588 14214
rect 21546 13832 21602 13841
rect 21546 13767 21602 13776
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21640 13388 21692 13394
rect 21640 13330 21692 13336
rect 21284 13138 21312 13330
rect 21652 13161 21680 13330
rect 21100 13110 21312 13138
rect 21180 12300 21232 12306
rect 21284 12288 21312 13110
rect 21638 13152 21694 13161
rect 21638 13087 21694 13096
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21232 12260 21312 12288
rect 21180 12242 21232 12248
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20548 9654 20576 11290
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 20640 10198 20668 11154
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20628 10192 20680 10198
rect 20628 10134 20680 10140
rect 20626 10024 20682 10033
rect 20626 9959 20682 9968
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20444 9172 20496 9178
rect 20444 9114 20496 9120
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 20548 7954 20576 8978
rect 20640 8974 20668 9959
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20732 8634 20760 10610
rect 21008 10538 21036 11766
rect 21192 11694 21220 12242
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21560 11898 21588 12174
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21180 11688 21232 11694
rect 21652 11665 21680 12922
rect 21180 11630 21232 11636
rect 21638 11656 21694 11665
rect 21638 11591 21694 11600
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 21100 10713 21128 11494
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21180 11008 21232 11014
rect 21180 10950 21232 10956
rect 21272 11008 21324 11014
rect 21272 10950 21324 10956
rect 21086 10704 21142 10713
rect 21086 10639 21142 10648
rect 20996 10532 21048 10538
rect 20996 10474 21048 10480
rect 21008 10266 21036 10474
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 21100 10169 21128 10639
rect 21086 10160 21142 10169
rect 21086 10095 21142 10104
rect 21192 9674 21220 10950
rect 21284 10742 21312 10950
rect 21560 10810 21588 11086
rect 21652 11014 21680 11494
rect 21640 11008 21692 11014
rect 21640 10950 21692 10956
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21272 10736 21324 10742
rect 21272 10678 21324 10684
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21468 10062 21496 10610
rect 21548 10532 21600 10538
rect 21548 10474 21600 10480
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21560 10010 21588 10474
rect 21652 10130 21680 10950
rect 21744 10674 21772 18006
rect 22112 17626 22140 19366
rect 22296 18834 22324 20046
rect 22284 18828 22336 18834
rect 22284 18770 22336 18776
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22020 17598 22140 17626
rect 22020 17270 22048 17598
rect 22008 17264 22060 17270
rect 22008 17206 22060 17212
rect 22204 16266 22232 18022
rect 22388 17338 22416 20318
rect 22480 19242 22508 22102
rect 22744 22102 22796 22108
rect 23294 22128 23350 22137
rect 22558 22063 22614 22072
rect 22572 21894 22600 22063
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22560 21004 22612 21010
rect 22560 20946 22612 20952
rect 22572 20330 22600 20946
rect 22652 20868 22704 20874
rect 22652 20810 22704 20816
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 22572 20058 22600 20266
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22664 19990 22692 20810
rect 22652 19984 22704 19990
rect 22652 19926 22704 19932
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 22468 19236 22520 19242
rect 22468 19178 22520 19184
rect 22664 18766 22692 19246
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22468 18148 22520 18154
rect 22468 18090 22520 18096
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 22112 16250 22232 16266
rect 22100 16244 22232 16250
rect 22152 16238 22232 16244
rect 22100 16186 22152 16192
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 21836 14822 21864 15438
rect 22020 15366 22048 15438
rect 22008 15360 22060 15366
rect 22008 15302 22060 15308
rect 22388 14958 22416 16594
rect 22480 16454 22508 18090
rect 22558 17912 22614 17921
rect 22558 17847 22614 17856
rect 22572 17134 22600 17847
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22664 16182 22692 18702
rect 22756 17082 22784 22102
rect 23294 22063 23350 22072
rect 22836 21956 22888 21962
rect 22836 21898 22888 21904
rect 22848 19514 22876 21898
rect 23308 21554 23336 22063
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 23112 21480 23164 21486
rect 22940 21428 23112 21434
rect 22940 21422 23164 21428
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 22940 21406 23152 21422
rect 22836 19508 22888 19514
rect 22836 19450 22888 19456
rect 22836 19372 22888 19378
rect 22836 19314 22888 19320
rect 22848 18154 22876 19314
rect 22940 18766 22968 21406
rect 23112 21344 23164 21350
rect 23032 21304 23112 21332
rect 23032 18970 23060 21304
rect 23112 21286 23164 21292
rect 23168 21244 23476 21253
rect 23168 21242 23174 21244
rect 23230 21242 23254 21244
rect 23310 21242 23334 21244
rect 23390 21242 23414 21244
rect 23470 21242 23476 21244
rect 23230 21190 23232 21242
rect 23412 21190 23414 21242
rect 23168 21188 23174 21190
rect 23230 21188 23254 21190
rect 23310 21188 23334 21190
rect 23390 21188 23414 21190
rect 23470 21188 23476 21190
rect 23168 21179 23476 21188
rect 23388 21140 23440 21146
rect 23388 21082 23440 21088
rect 23400 20398 23428 21082
rect 23584 20806 23612 21422
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23168 20156 23476 20165
rect 23168 20154 23174 20156
rect 23230 20154 23254 20156
rect 23310 20154 23334 20156
rect 23390 20154 23414 20156
rect 23470 20154 23476 20156
rect 23230 20102 23232 20154
rect 23412 20102 23414 20154
rect 23168 20100 23174 20102
rect 23230 20100 23254 20102
rect 23310 20100 23334 20102
rect 23390 20100 23414 20102
rect 23470 20100 23476 20102
rect 23168 20091 23476 20100
rect 23386 19952 23442 19961
rect 23386 19887 23442 19896
rect 23400 19786 23428 19887
rect 23570 19816 23626 19825
rect 23388 19780 23440 19786
rect 23676 19802 23704 22238
rect 28540 22238 28592 22244
rect 23754 22199 23810 22208
rect 25596 22160 25648 22166
rect 25042 22128 25098 22137
rect 23756 22092 23808 22098
rect 25596 22102 25648 22108
rect 25042 22063 25044 22072
rect 23756 22034 23808 22040
rect 25096 22063 25098 22072
rect 25044 22034 25096 22040
rect 23768 21865 23796 22034
rect 23754 21856 23810 21865
rect 23754 21791 23810 21800
rect 23768 21350 23796 21791
rect 24674 21720 24730 21729
rect 24674 21655 24730 21664
rect 24492 21548 24544 21554
rect 24688 21536 24716 21655
rect 24544 21508 24716 21536
rect 24492 21490 24544 21496
rect 25056 21486 25084 22034
rect 25608 21690 25636 22102
rect 27896 22024 27948 22030
rect 26330 21992 26386 22001
rect 25780 21956 25832 21962
rect 27896 21966 27948 21972
rect 26330 21927 26386 21936
rect 25780 21898 25832 21904
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25504 21616 25556 21622
rect 25504 21558 25556 21564
rect 23848 21480 23900 21486
rect 23848 21422 23900 21428
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 24768 21480 24820 21486
rect 24768 21422 24820 21428
rect 24952 21480 25004 21486
rect 24952 21422 25004 21428
rect 25044 21480 25096 21486
rect 25044 21422 25096 21428
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23860 20058 23888 21422
rect 23952 21350 23980 21422
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 23938 20904 23994 20913
rect 23938 20839 23994 20848
rect 23848 20052 23900 20058
rect 23848 19994 23900 20000
rect 23846 19952 23902 19961
rect 23846 19887 23902 19896
rect 23626 19774 23704 19802
rect 23570 19751 23626 19760
rect 23388 19722 23440 19728
rect 23584 19514 23612 19751
rect 23860 19689 23888 19887
rect 23846 19680 23902 19689
rect 23846 19615 23902 19624
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 23664 19236 23716 19242
rect 23664 19178 23716 19184
rect 23168 19068 23476 19077
rect 23168 19066 23174 19068
rect 23230 19066 23254 19068
rect 23310 19066 23334 19068
rect 23390 19066 23414 19068
rect 23470 19066 23476 19068
rect 23230 19014 23232 19066
rect 23412 19014 23414 19066
rect 23168 19012 23174 19014
rect 23230 19012 23254 19014
rect 23310 19012 23334 19014
rect 23390 19012 23414 19014
rect 23470 19012 23476 19014
rect 23168 19003 23476 19012
rect 23020 18964 23072 18970
rect 23020 18906 23072 18912
rect 23386 18864 23442 18873
rect 23386 18799 23442 18808
rect 22928 18760 22980 18766
rect 22928 18702 22980 18708
rect 23400 18193 23428 18799
rect 23676 18465 23704 19178
rect 23860 18834 23888 19615
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 23756 18624 23808 18630
rect 23756 18566 23808 18572
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23662 18456 23718 18465
rect 23768 18426 23796 18566
rect 23662 18391 23718 18400
rect 23756 18420 23808 18426
rect 23386 18184 23442 18193
rect 22836 18148 22888 18154
rect 23386 18119 23442 18128
rect 23570 18184 23626 18193
rect 23676 18170 23704 18391
rect 23756 18362 23808 18368
rect 23626 18142 23704 18170
rect 23756 18148 23808 18154
rect 23570 18119 23572 18128
rect 22836 18090 22888 18096
rect 23624 18119 23626 18128
rect 23572 18090 23624 18096
rect 23756 18090 23808 18096
rect 23168 17980 23476 17989
rect 23168 17978 23174 17980
rect 23230 17978 23254 17980
rect 23310 17978 23334 17980
rect 23390 17978 23414 17980
rect 23470 17978 23476 17980
rect 23230 17926 23232 17978
rect 23412 17926 23414 17978
rect 23168 17924 23174 17926
rect 23230 17924 23254 17926
rect 23310 17924 23334 17926
rect 23390 17924 23414 17926
rect 23470 17924 23476 17926
rect 23168 17915 23476 17924
rect 23020 17740 23072 17746
rect 23020 17682 23072 17688
rect 22756 17054 22968 17082
rect 22742 16824 22798 16833
rect 22742 16759 22798 16768
rect 22756 16522 22784 16759
rect 22744 16516 22796 16522
rect 22744 16458 22796 16464
rect 22836 16244 22888 16250
rect 22836 16186 22888 16192
rect 22652 16176 22704 16182
rect 22652 16118 22704 16124
rect 22744 15904 22796 15910
rect 22744 15846 22796 15852
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22296 14618 22324 14758
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 21928 13977 21956 14010
rect 21914 13968 21970 13977
rect 21914 13903 21970 13912
rect 21916 13728 21968 13734
rect 21916 13670 21968 13676
rect 21928 13530 21956 13670
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 21914 12744 21970 12753
rect 21914 12679 21970 12688
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21836 11354 21864 12174
rect 21824 11348 21876 11354
rect 21824 11290 21876 11296
rect 21928 10826 21956 12679
rect 22008 12640 22060 12646
rect 22008 12582 22060 12588
rect 22020 12442 22048 12582
rect 22008 12436 22060 12442
rect 22112 12434 22140 13262
rect 22296 13190 22324 14350
rect 22388 13433 22416 14894
rect 22664 13977 22692 15302
rect 22756 14278 22784 15846
rect 22848 14482 22876 16186
rect 22940 16046 22968 17054
rect 23032 16969 23060 17682
rect 23768 17626 23796 18090
rect 23860 17746 23888 18566
rect 23952 17882 23980 20839
rect 24124 20800 24176 20806
rect 24124 20742 24176 20748
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 24044 17882 24072 18226
rect 24136 18154 24164 20742
rect 24308 20596 24360 20602
rect 24308 20538 24360 20544
rect 24320 19854 24348 20538
rect 24780 20262 24808 21422
rect 24964 21298 24992 21422
rect 25320 21344 25372 21350
rect 24964 21270 25084 21298
rect 25320 21286 25372 21292
rect 25056 21146 25084 21270
rect 25332 21146 25360 21286
rect 25516 21146 25544 21558
rect 25792 21486 25820 21898
rect 25872 21888 25924 21894
rect 25872 21830 25924 21836
rect 25780 21480 25832 21486
rect 25780 21422 25832 21428
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25044 21140 25096 21146
rect 25044 21082 25096 21088
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 25504 21140 25556 21146
rect 25504 21082 25556 21088
rect 25228 21072 25280 21078
rect 25228 21014 25280 21020
rect 24858 20632 24914 20641
rect 25136 20596 25188 20602
rect 24858 20567 24914 20576
rect 24768 20256 24820 20262
rect 24768 20198 24820 20204
rect 24308 19848 24360 19854
rect 24308 19790 24360 19796
rect 24492 19304 24544 19310
rect 24412 19252 24492 19258
rect 24412 19246 24544 19252
rect 24412 19230 24532 19246
rect 24216 18896 24268 18902
rect 24214 18864 24216 18873
rect 24268 18864 24270 18873
rect 24214 18799 24270 18808
rect 24412 18630 24440 19230
rect 24492 19168 24544 19174
rect 24492 19110 24544 19116
rect 24504 18834 24532 19110
rect 24492 18828 24544 18834
rect 24492 18770 24544 18776
rect 24400 18624 24452 18630
rect 24400 18566 24452 18572
rect 24490 18456 24546 18465
rect 24490 18391 24546 18400
rect 24400 18352 24452 18358
rect 24398 18320 24400 18329
rect 24452 18320 24454 18329
rect 24216 18284 24268 18290
rect 24398 18255 24454 18264
rect 24216 18226 24268 18232
rect 24124 18148 24176 18154
rect 24124 18090 24176 18096
rect 23940 17876 23992 17882
rect 23940 17818 23992 17824
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24228 17746 24256 18226
rect 23848 17740 23900 17746
rect 23848 17682 23900 17688
rect 24216 17740 24268 17746
rect 24216 17682 24268 17688
rect 24400 17740 24452 17746
rect 24400 17682 24452 17688
rect 23768 17610 23980 17626
rect 23768 17604 23992 17610
rect 23768 17598 23940 17604
rect 23940 17546 23992 17552
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 23216 17134 23244 17274
rect 23204 17128 23256 17134
rect 23204 17070 23256 17076
rect 23018 16960 23074 16969
rect 23018 16895 23074 16904
rect 23168 16892 23476 16901
rect 23168 16890 23174 16892
rect 23230 16890 23254 16892
rect 23310 16890 23334 16892
rect 23390 16890 23414 16892
rect 23470 16890 23476 16892
rect 23230 16838 23232 16890
rect 23412 16838 23414 16890
rect 23168 16836 23174 16838
rect 23230 16836 23254 16838
rect 23310 16836 23334 16838
rect 23390 16836 23414 16838
rect 23470 16836 23476 16838
rect 23168 16827 23476 16836
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23860 16114 23888 16730
rect 23952 16658 23980 17546
rect 24228 17202 24256 17682
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24228 16794 24256 17138
rect 24412 16998 24440 17682
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24412 16794 24440 16934
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 24030 16552 24086 16561
rect 24030 16487 24086 16496
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 23168 15804 23476 15813
rect 23168 15802 23174 15804
rect 23230 15802 23254 15804
rect 23310 15802 23334 15804
rect 23390 15802 23414 15804
rect 23470 15802 23476 15804
rect 23230 15750 23232 15802
rect 23412 15750 23414 15802
rect 23168 15748 23174 15750
rect 23230 15748 23254 15750
rect 23310 15748 23334 15750
rect 23390 15748 23414 15750
rect 23470 15748 23476 15750
rect 23168 15739 23476 15748
rect 23756 15700 23808 15706
rect 23756 15642 23808 15648
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23676 15026 23704 15438
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23020 14884 23072 14890
rect 23020 14826 23072 14832
rect 22836 14476 22888 14482
rect 22836 14418 22888 14424
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22650 13968 22706 13977
rect 22650 13903 22706 13912
rect 22926 13968 22982 13977
rect 22926 13903 22982 13912
rect 22940 13870 22968 13903
rect 22928 13864 22980 13870
rect 22928 13806 22980 13812
rect 22560 13796 22612 13802
rect 22744 13796 22796 13802
rect 22612 13756 22744 13784
rect 22560 13738 22612 13744
rect 22744 13738 22796 13744
rect 22374 13424 22430 13433
rect 22374 13359 22430 13368
rect 22376 13320 22428 13326
rect 22376 13262 22428 13268
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22388 12918 22416 13262
rect 22572 12918 22600 13738
rect 23032 13734 23060 14826
rect 23168 14716 23476 14725
rect 23168 14714 23174 14716
rect 23230 14714 23254 14716
rect 23310 14714 23334 14716
rect 23390 14714 23414 14716
rect 23470 14714 23476 14716
rect 23230 14662 23232 14714
rect 23412 14662 23414 14714
rect 23168 14660 23174 14662
rect 23230 14660 23254 14662
rect 23310 14660 23334 14662
rect 23390 14660 23414 14662
rect 23470 14660 23476 14662
rect 23168 14651 23476 14660
rect 23676 14482 23704 14962
rect 23768 14550 23796 15642
rect 23860 15570 23888 16050
rect 23940 16040 23992 16046
rect 23940 15982 23992 15988
rect 23848 15564 23900 15570
rect 23848 15506 23900 15512
rect 23846 15192 23902 15201
rect 23846 15127 23848 15136
rect 23900 15127 23902 15136
rect 23848 15098 23900 15104
rect 23756 14544 23808 14550
rect 23756 14486 23808 14492
rect 23846 14512 23902 14521
rect 23664 14476 23716 14482
rect 23846 14447 23902 14456
rect 23664 14418 23716 14424
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23308 13870 23336 14214
rect 23860 13954 23888 14447
rect 23768 13926 23888 13954
rect 23768 13870 23796 13926
rect 23952 13870 23980 15982
rect 24044 15504 24072 16487
rect 24412 16266 24440 16730
rect 24228 16238 24440 16266
rect 24228 16114 24256 16238
rect 24216 16108 24268 16114
rect 24216 16050 24268 16056
rect 24124 15904 24176 15910
rect 24124 15846 24176 15852
rect 24032 15498 24084 15504
rect 24136 15502 24164 15846
rect 24228 15706 24256 16050
rect 24308 15904 24360 15910
rect 24308 15846 24360 15852
rect 24216 15700 24268 15706
rect 24216 15642 24268 15648
rect 24032 15440 24084 15446
rect 24124 15496 24176 15502
rect 24124 15438 24176 15444
rect 24032 15360 24084 15366
rect 24032 15302 24084 15308
rect 24044 15026 24072 15302
rect 24228 15026 24256 15642
rect 24032 15020 24084 15026
rect 24032 14962 24084 14968
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24228 14482 24256 14962
rect 24216 14476 24268 14482
rect 24216 14418 24268 14424
rect 24320 14414 24348 15846
rect 24504 15745 24532 18391
rect 24872 18290 24900 20567
rect 25056 20556 25136 20584
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24584 18216 24636 18222
rect 24584 18158 24636 18164
rect 24596 17105 24624 18158
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 24766 17912 24822 17921
rect 24766 17847 24822 17856
rect 24780 17678 24808 17847
rect 24964 17746 24992 18022
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24582 17096 24638 17105
rect 24582 17031 24638 17040
rect 25056 16590 25084 20556
rect 25136 20538 25188 20544
rect 25240 20398 25268 21014
rect 25228 20392 25280 20398
rect 25228 20334 25280 20340
rect 25240 20058 25268 20334
rect 25228 20052 25280 20058
rect 25228 19994 25280 20000
rect 25136 19304 25188 19310
rect 25134 19272 25136 19281
rect 25504 19304 25556 19310
rect 25188 19272 25190 19281
rect 25504 19246 25556 19252
rect 25134 19207 25190 19216
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 25332 17785 25360 18022
rect 25318 17776 25374 17785
rect 25228 17740 25280 17746
rect 25318 17711 25374 17720
rect 25228 17682 25280 17688
rect 25240 17377 25268 17682
rect 25226 17368 25282 17377
rect 25226 17303 25282 17312
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 25320 16176 25372 16182
rect 25318 16144 25320 16153
rect 25372 16144 25374 16153
rect 25318 16079 25374 16088
rect 24766 15872 24822 15881
rect 24766 15807 24822 15816
rect 24490 15736 24546 15745
rect 24490 15671 24546 15680
rect 24780 15026 24808 15807
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 25044 14952 25096 14958
rect 25044 14894 25096 14900
rect 24398 14648 24454 14657
rect 24398 14583 24454 14592
rect 24308 14408 24360 14414
rect 24308 14350 24360 14356
rect 24412 13977 24440 14583
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24504 14006 24532 14350
rect 24492 14000 24544 14006
rect 24398 13968 24454 13977
rect 24216 13932 24268 13938
rect 24492 13942 24544 13948
rect 24398 13903 24400 13912
rect 24216 13874 24268 13880
rect 24452 13903 24454 13912
rect 24400 13874 24452 13880
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 23388 13864 23440 13870
rect 23756 13864 23808 13870
rect 23440 13812 23612 13818
rect 23388 13806 23612 13812
rect 23756 13806 23808 13812
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 23400 13790 23612 13806
rect 23020 13728 23072 13734
rect 23584 13705 23612 13790
rect 23020 13670 23072 13676
rect 23570 13696 23626 13705
rect 23168 13628 23476 13637
rect 23570 13631 23626 13640
rect 23168 13626 23174 13628
rect 23230 13626 23254 13628
rect 23310 13626 23334 13628
rect 23390 13626 23414 13628
rect 23470 13626 23476 13628
rect 23230 13574 23232 13626
rect 23412 13574 23414 13626
rect 23168 13572 23174 13574
rect 23230 13572 23254 13574
rect 23310 13572 23334 13574
rect 23390 13572 23414 13574
rect 23470 13572 23476 13574
rect 23168 13563 23476 13572
rect 23938 13560 23994 13569
rect 23938 13495 23940 13504
rect 23992 13495 23994 13504
rect 23940 13466 23992 13472
rect 23848 13456 23900 13462
rect 23848 13398 23900 13404
rect 22652 13320 22704 13326
rect 22652 13262 22704 13268
rect 22664 12986 22692 13262
rect 23020 13184 23072 13190
rect 22940 13161 23020 13172
rect 22926 13152 23020 13161
rect 22982 13144 23020 13152
rect 23020 13126 23072 13132
rect 22926 13087 22982 13096
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22376 12912 22428 12918
rect 22376 12854 22428 12860
rect 22560 12912 22612 12918
rect 22560 12854 22612 12860
rect 22834 12880 22890 12889
rect 22834 12815 22890 12824
rect 22848 12646 22876 12815
rect 22940 12782 22968 13087
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 23768 12782 23796 12922
rect 23860 12782 23888 13398
rect 24044 13258 24072 13806
rect 24124 13728 24176 13734
rect 24124 13670 24176 13676
rect 24136 13530 24164 13670
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 24228 13462 24256 13874
rect 24584 13796 24636 13802
rect 24688 13784 24716 14418
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24768 13864 24820 13870
rect 24768 13806 24820 13812
rect 24636 13756 24716 13784
rect 24584 13738 24636 13744
rect 24216 13456 24268 13462
rect 24216 13398 24268 13404
rect 24398 13424 24454 13433
rect 24398 13359 24454 13368
rect 24308 13320 24360 13326
rect 24308 13262 24360 13268
rect 24032 13252 24084 13258
rect 24032 13194 24084 13200
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 22928 12776 22980 12782
rect 23756 12776 23808 12782
rect 23754 12744 23756 12753
rect 23848 12776 23900 12782
rect 23808 12744 23810 12753
rect 22928 12718 22980 12724
rect 23032 12714 23612 12730
rect 23032 12708 23624 12714
rect 23032 12702 23572 12708
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 23032 12434 23060 12702
rect 24044 12730 24072 12786
rect 23848 12718 23900 12724
rect 23754 12679 23810 12688
rect 23572 12650 23624 12656
rect 23168 12540 23476 12549
rect 23168 12538 23174 12540
rect 23230 12538 23254 12540
rect 23310 12538 23334 12540
rect 23390 12538 23414 12540
rect 23470 12538 23476 12540
rect 23230 12486 23232 12538
rect 23412 12486 23414 12538
rect 23168 12484 23174 12486
rect 23230 12484 23254 12486
rect 23310 12484 23334 12486
rect 23390 12484 23414 12486
rect 23470 12484 23476 12486
rect 23168 12475 23476 12484
rect 23860 12442 23888 12718
rect 23952 12714 24072 12730
rect 23940 12708 24072 12714
rect 23992 12702 24072 12708
rect 23940 12650 23992 12656
rect 24320 12646 24348 13262
rect 24124 12640 24176 12646
rect 24124 12582 24176 12588
rect 24308 12640 24360 12646
rect 24308 12582 24360 12588
rect 23112 12436 23164 12442
rect 22112 12406 22784 12434
rect 23032 12406 23112 12434
rect 22008 12378 22060 12384
rect 22020 11558 22048 12378
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 21836 10798 21956 10826
rect 22020 10826 22048 11086
rect 22112 11014 22140 11086
rect 22100 11008 22152 11014
rect 22100 10950 22152 10956
rect 22020 10798 22140 10826
rect 22296 10810 22324 11630
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 21732 10668 21784 10674
rect 21732 10610 21784 10616
rect 21836 10606 21864 10798
rect 21916 10736 21968 10742
rect 21916 10678 21968 10684
rect 21824 10600 21876 10606
rect 21824 10542 21876 10548
rect 21928 10418 21956 10678
rect 22112 10470 22140 10798
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22100 10464 22152 10470
rect 21928 10390 22048 10418
rect 22100 10406 22152 10412
rect 22020 10130 22048 10390
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 21916 10056 21968 10062
rect 21560 10004 21916 10010
rect 22190 10024 22246 10033
rect 21560 9998 21968 10004
rect 21560 9982 21956 9998
rect 22112 9982 22190 10010
rect 21192 9646 21312 9674
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20536 7948 20588 7954
rect 20536 7890 20588 7896
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20456 7342 20484 7686
rect 20444 7336 20496 7342
rect 20444 7278 20496 7284
rect 20548 6866 20576 7890
rect 20640 7313 20668 7890
rect 20626 7304 20682 7313
rect 20626 7239 20682 7248
rect 20536 6860 20588 6866
rect 20588 6820 20668 6848
rect 20536 6802 20588 6808
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20166 5264 20222 5273
rect 20272 5234 20300 6598
rect 20364 5914 20392 6598
rect 20640 6458 20668 6820
rect 20732 6458 20760 8434
rect 20824 7546 20852 8774
rect 21192 8673 21220 9522
rect 21178 8664 21234 8673
rect 21178 8599 21234 8608
rect 21284 8480 21312 9646
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 21376 9110 21404 9318
rect 21652 9178 21680 9522
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 21364 9104 21416 9110
rect 21364 9046 21416 9052
rect 22020 9042 22048 9114
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 21916 8900 21968 8906
rect 21916 8842 21968 8848
rect 21284 8452 21404 8480
rect 20994 8392 21050 8401
rect 20994 8327 21050 8336
rect 21270 8392 21326 8401
rect 21270 8327 21326 8336
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20166 5199 20222 5208
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20548 4758 20576 6190
rect 20640 5846 20668 6394
rect 20628 5840 20680 5846
rect 20626 5808 20628 5817
rect 20680 5808 20682 5817
rect 20626 5743 20682 5752
rect 20626 5672 20682 5681
rect 20626 5607 20628 5616
rect 20680 5607 20682 5616
rect 20628 5578 20680 5584
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 20536 4752 20588 4758
rect 20536 4694 20588 4700
rect 20732 4146 20760 5102
rect 20824 4690 20852 5510
rect 20812 4684 20864 4690
rect 20812 4626 20864 4632
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20732 3602 20760 4082
rect 20824 3738 20852 4082
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 20732 3058 20760 3538
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20732 2650 20760 2994
rect 20916 2774 20944 7278
rect 21008 6225 21036 8327
rect 21284 8022 21312 8327
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 21284 6916 21312 7958
rect 21376 7018 21404 8452
rect 21928 8430 21956 8842
rect 22006 8528 22062 8537
rect 22006 8463 22008 8472
rect 22060 8463 22062 8472
rect 22008 8434 22060 8440
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21916 8424 21968 8430
rect 21916 8366 21968 8372
rect 21468 7886 21496 8366
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21916 8288 21968 8294
rect 21916 8230 21968 8236
rect 21652 7886 21680 8230
rect 21928 8090 21956 8230
rect 21916 8084 21968 8090
rect 21916 8026 21968 8032
rect 21456 7880 21508 7886
rect 21640 7880 21692 7886
rect 21508 7840 21588 7868
rect 21456 7822 21508 7828
rect 21560 7342 21588 7840
rect 21640 7822 21692 7828
rect 21928 7410 21956 8026
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 22008 7404 22060 7410
rect 22008 7346 22060 7352
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21376 6990 21680 7018
rect 21284 6888 21404 6916
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 20994 6216 21050 6225
rect 20994 6151 21050 6160
rect 21100 5914 21128 6734
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 21192 5778 21220 6190
rect 21180 5772 21232 5778
rect 21180 5714 21232 5720
rect 21192 5166 21220 5714
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 21284 4758 21312 4966
rect 21272 4752 21324 4758
rect 21272 4694 21324 4700
rect 21376 4690 21404 6888
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21560 6254 21588 6598
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 21560 5914 21588 6054
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21468 5234 21496 5510
rect 21456 5228 21508 5234
rect 21456 5170 21508 5176
rect 21560 5030 21588 5850
rect 21652 5522 21680 6990
rect 21744 6254 21772 7346
rect 22020 6610 22048 7346
rect 22112 6934 22140 9982
rect 22190 9959 22246 9968
rect 22388 9654 22416 11086
rect 22652 11008 22704 11014
rect 22652 10950 22704 10956
rect 22664 10266 22692 10950
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22466 9888 22522 9897
rect 22466 9823 22522 9832
rect 22376 9648 22428 9654
rect 22376 9590 22428 9596
rect 22376 9444 22428 9450
rect 22376 9386 22428 9392
rect 22284 9036 22336 9042
rect 22284 8978 22336 8984
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22204 8498 22232 8774
rect 22296 8634 22324 8978
rect 22284 8628 22336 8634
rect 22284 8570 22336 8576
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22204 7410 22232 7686
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22388 7206 22416 9386
rect 22480 8276 22508 9823
rect 22560 9512 22612 9518
rect 22560 9454 22612 9460
rect 22572 9042 22600 9454
rect 22560 9036 22612 9042
rect 22560 8978 22612 8984
rect 22652 8900 22704 8906
rect 22652 8842 22704 8848
rect 22560 8288 22612 8294
rect 22480 8248 22560 8276
rect 22560 8230 22612 8236
rect 22664 7410 22692 8842
rect 22756 7698 22784 12406
rect 23112 12378 23164 12384
rect 23848 12436 23900 12442
rect 23848 12378 23900 12384
rect 24136 12306 24164 12582
rect 24124 12300 24176 12306
rect 24124 12242 24176 12248
rect 24320 12238 24348 12582
rect 23940 12232 23992 12238
rect 23940 12174 23992 12180
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 23952 11898 23980 12174
rect 23940 11892 23992 11898
rect 23940 11834 23992 11840
rect 24320 11762 24348 12174
rect 24308 11756 24360 11762
rect 24308 11698 24360 11704
rect 22928 11688 22980 11694
rect 22848 11636 22928 11642
rect 22848 11630 22980 11636
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 24214 11656 24270 11665
rect 22848 11614 22968 11630
rect 22848 10266 22876 11614
rect 23168 11452 23476 11461
rect 23168 11450 23174 11452
rect 23230 11450 23254 11452
rect 23310 11450 23334 11452
rect 23390 11450 23414 11452
rect 23470 11450 23476 11452
rect 23230 11398 23232 11450
rect 23412 11398 23414 11450
rect 23168 11396 23174 11398
rect 23230 11396 23254 11398
rect 23310 11396 23334 11398
rect 23390 11396 23414 11398
rect 23470 11396 23476 11398
rect 23168 11387 23476 11396
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 22940 10674 22968 11290
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 22940 10198 22968 10610
rect 23020 10600 23072 10606
rect 23492 10577 23520 10610
rect 23020 10542 23072 10548
rect 23478 10568 23534 10577
rect 22928 10192 22980 10198
rect 22928 10134 22980 10140
rect 23032 9738 23060 10542
rect 23478 10503 23534 10512
rect 23168 10364 23476 10373
rect 23168 10362 23174 10364
rect 23230 10362 23254 10364
rect 23310 10362 23334 10364
rect 23390 10362 23414 10364
rect 23470 10362 23476 10364
rect 23230 10310 23232 10362
rect 23412 10310 23414 10362
rect 23168 10308 23174 10310
rect 23230 10308 23254 10310
rect 23310 10308 23334 10310
rect 23390 10308 23414 10310
rect 23470 10308 23476 10310
rect 23168 10299 23476 10308
rect 23584 10266 23612 11086
rect 23848 11008 23900 11014
rect 23848 10950 23900 10956
rect 23860 10538 23888 10950
rect 23848 10532 23900 10538
rect 23848 10474 23900 10480
rect 23572 10260 23624 10266
rect 23572 10202 23624 10208
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23032 9710 23152 9738
rect 23124 9654 23152 9710
rect 23112 9648 23164 9654
rect 23112 9590 23164 9596
rect 23492 9518 23520 9998
rect 23572 9988 23624 9994
rect 23572 9930 23624 9936
rect 23480 9512 23532 9518
rect 23478 9480 23480 9489
rect 23532 9480 23534 9489
rect 23478 9415 23534 9424
rect 23584 9353 23612 9930
rect 23664 9920 23716 9926
rect 23664 9862 23716 9868
rect 23570 9344 23626 9353
rect 23168 9276 23476 9285
rect 23570 9279 23626 9288
rect 23168 9274 23174 9276
rect 23230 9274 23254 9276
rect 23310 9274 23334 9276
rect 23390 9274 23414 9276
rect 23470 9274 23476 9276
rect 23230 9222 23232 9274
rect 23412 9222 23414 9274
rect 23168 9220 23174 9222
rect 23230 9220 23254 9222
rect 23310 9220 23334 9222
rect 23390 9220 23414 9222
rect 23470 9220 23476 9222
rect 23168 9211 23476 9220
rect 23584 9178 23612 9279
rect 23676 9178 23704 9862
rect 23756 9716 23808 9722
rect 23756 9658 23808 9664
rect 23768 9625 23796 9658
rect 23754 9616 23810 9625
rect 23754 9551 23810 9560
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23572 9172 23624 9178
rect 23572 9114 23624 9120
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23768 9042 23796 9318
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 23572 8968 23624 8974
rect 23572 8910 23624 8916
rect 23018 8664 23074 8673
rect 23018 8599 23074 8608
rect 22928 8424 22980 8430
rect 22928 8366 22980 8372
rect 22940 7886 22968 8366
rect 23032 8090 23060 8599
rect 23168 8188 23476 8197
rect 23168 8186 23174 8188
rect 23230 8186 23254 8188
rect 23310 8186 23334 8188
rect 23390 8186 23414 8188
rect 23470 8186 23476 8188
rect 23230 8134 23232 8186
rect 23412 8134 23414 8186
rect 23168 8132 23174 8134
rect 23230 8132 23254 8134
rect 23310 8132 23334 8134
rect 23390 8132 23414 8134
rect 23470 8132 23476 8134
rect 23168 8123 23476 8132
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 22756 7670 22968 7698
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22376 7200 22428 7206
rect 22376 7142 22428 7148
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22100 6928 22152 6934
rect 22100 6870 22152 6876
rect 22100 6792 22152 6798
rect 22152 6752 22232 6780
rect 22100 6734 22152 6740
rect 22020 6582 22140 6610
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 22112 5794 22140 6582
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 22020 5766 22140 5794
rect 21836 5681 21864 5714
rect 22020 5681 22048 5766
rect 22204 5710 22232 6752
rect 22388 6662 22416 7142
rect 22468 6792 22520 6798
rect 22572 6769 22600 7142
rect 22940 6866 22968 7670
rect 23584 7546 23612 8910
rect 23768 8430 23796 8978
rect 23860 8430 23888 9522
rect 23756 8424 23808 8430
rect 23756 8366 23808 8372
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 23168 7100 23476 7109
rect 23168 7098 23174 7100
rect 23230 7098 23254 7100
rect 23310 7098 23334 7100
rect 23390 7098 23414 7100
rect 23470 7098 23476 7100
rect 23230 7046 23232 7098
rect 23412 7046 23414 7098
rect 23168 7044 23174 7046
rect 23230 7044 23254 7046
rect 23310 7044 23334 7046
rect 23390 7044 23414 7046
rect 23470 7044 23476 7046
rect 23168 7035 23476 7044
rect 23676 7002 23704 7822
rect 23952 7290 23980 11630
rect 24214 11591 24270 11600
rect 24124 11144 24176 11150
rect 24124 11086 24176 11092
rect 24136 10538 24164 11086
rect 24124 10532 24176 10538
rect 24124 10474 24176 10480
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 24044 9586 24072 10406
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 24030 8936 24086 8945
rect 24030 8871 24086 8880
rect 23768 7262 23980 7290
rect 24044 7290 24072 8871
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 24136 7546 24164 7822
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24122 7440 24178 7449
rect 24122 7375 24124 7384
rect 24176 7375 24178 7384
rect 24228 7392 24256 11591
rect 24308 10600 24360 10606
rect 24308 10542 24360 10548
rect 24320 9926 24348 10542
rect 24308 9920 24360 9926
rect 24308 9862 24360 9868
rect 24412 9602 24440 13359
rect 24780 13326 24808 13806
rect 24872 13394 24900 14010
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24964 12986 24992 14350
rect 25056 14278 25084 14894
rect 25516 14890 25544 19246
rect 25700 18970 25728 21286
rect 25884 21010 25912 21830
rect 25962 21720 26018 21729
rect 25962 21655 25964 21664
rect 26016 21655 26018 21664
rect 25964 21626 26016 21632
rect 26056 21480 26108 21486
rect 26056 21422 26108 21428
rect 25780 21004 25832 21010
rect 25780 20946 25832 20952
rect 25872 21004 25924 21010
rect 25872 20946 25924 20952
rect 25688 18964 25740 18970
rect 25688 18906 25740 18912
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25608 18290 25636 18566
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25596 17672 25648 17678
rect 25792 17626 25820 20946
rect 26068 20942 26096 21422
rect 26146 21176 26202 21185
rect 26146 21111 26202 21120
rect 26160 21078 26188 21111
rect 26148 21072 26200 21078
rect 26148 21014 26200 21020
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 26238 20904 26294 20913
rect 25964 20868 26016 20874
rect 26238 20839 26294 20848
rect 25964 20810 26016 20816
rect 25872 18828 25924 18834
rect 25872 18770 25924 18776
rect 25884 17746 25912 18770
rect 25872 17740 25924 17746
rect 25872 17682 25924 17688
rect 25596 17614 25648 17620
rect 25504 14884 25556 14890
rect 25504 14826 25556 14832
rect 25044 14272 25096 14278
rect 25044 14214 25096 14220
rect 25608 12986 25636 17614
rect 25700 17598 25820 17626
rect 25700 14521 25728 17598
rect 25780 17536 25832 17542
rect 25976 17490 26004 20810
rect 26252 20534 26280 20839
rect 26240 20528 26292 20534
rect 26240 20470 26292 20476
rect 26148 20256 26200 20262
rect 26148 20198 26200 20204
rect 26160 19718 26188 20198
rect 26240 20052 26292 20058
rect 26240 19994 26292 20000
rect 26056 19712 26108 19718
rect 26056 19654 26108 19660
rect 26148 19712 26200 19718
rect 26148 19654 26200 19660
rect 26068 19417 26096 19654
rect 26252 19553 26280 19994
rect 26344 19922 26372 21927
rect 26963 21788 27271 21797
rect 26963 21786 26969 21788
rect 27025 21786 27049 21788
rect 27105 21786 27129 21788
rect 27185 21786 27209 21788
rect 27265 21786 27271 21788
rect 27025 21734 27027 21786
rect 27207 21734 27209 21786
rect 26963 21732 26969 21734
rect 27025 21732 27049 21734
rect 27105 21732 27129 21734
rect 27185 21732 27209 21734
rect 27265 21732 27271 21734
rect 26963 21723 27271 21732
rect 26698 21584 26754 21593
rect 26698 21519 26754 21528
rect 26712 21486 26740 21519
rect 26700 21480 26752 21486
rect 26700 21422 26752 21428
rect 27802 21448 27858 21457
rect 27802 21383 27858 21392
rect 27816 21350 27844 21383
rect 27804 21344 27856 21350
rect 27804 21286 27856 21292
rect 27908 21146 27936 21966
rect 28448 21412 28500 21418
rect 28448 21354 28500 21360
rect 28356 21344 28408 21350
rect 28356 21286 28408 21292
rect 27896 21140 27948 21146
rect 27896 21082 27948 21088
rect 27344 21004 27396 21010
rect 27344 20946 27396 20952
rect 26424 20936 26476 20942
rect 26424 20878 26476 20884
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26436 20482 26464 20878
rect 26608 20800 26660 20806
rect 26608 20742 26660 20748
rect 26436 20454 26556 20482
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 26332 19916 26384 19922
rect 26332 19858 26384 19864
rect 26332 19780 26384 19786
rect 26332 19722 26384 19728
rect 26238 19544 26294 19553
rect 26238 19479 26294 19488
rect 26054 19408 26110 19417
rect 26054 19343 26110 19352
rect 26344 19258 26372 19722
rect 26252 19230 26372 19258
rect 26056 18760 26108 18766
rect 26056 18702 26108 18708
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 26068 18222 26096 18702
rect 26160 18358 26188 18702
rect 26148 18352 26200 18358
rect 26148 18294 26200 18300
rect 26056 18216 26108 18222
rect 26056 18158 26108 18164
rect 26252 18057 26280 19230
rect 26332 19168 26384 19174
rect 26332 19110 26384 19116
rect 26238 18048 26294 18057
rect 26238 17983 26294 17992
rect 26054 17776 26110 17785
rect 26054 17711 26110 17720
rect 26068 17513 26096 17711
rect 26148 17672 26200 17678
rect 26148 17614 26200 17620
rect 25780 17478 25832 17484
rect 25792 17338 25820 17478
rect 25884 17462 26004 17490
rect 26054 17504 26110 17513
rect 25780 17332 25832 17338
rect 25780 17274 25832 17280
rect 25884 17270 25912 17462
rect 26054 17439 26110 17448
rect 25964 17332 26016 17338
rect 25964 17274 26016 17280
rect 25872 17264 25924 17270
rect 25872 17206 25924 17212
rect 25884 16153 25912 17206
rect 25870 16144 25926 16153
rect 25976 16114 26004 17274
rect 26160 17134 26188 17614
rect 26344 17202 26372 19110
rect 26436 18630 26464 20334
rect 26528 19514 26556 20454
rect 26516 19508 26568 19514
rect 26516 19450 26568 19456
rect 26424 18624 26476 18630
rect 26424 18566 26476 18572
rect 26436 17678 26464 18566
rect 26528 18222 26556 19450
rect 26516 18216 26568 18222
rect 26516 18158 26568 18164
rect 26620 17921 26648 20742
rect 26804 20398 26832 20878
rect 26963 20700 27271 20709
rect 26963 20698 26969 20700
rect 27025 20698 27049 20700
rect 27105 20698 27129 20700
rect 27185 20698 27209 20700
rect 27265 20698 27271 20700
rect 27025 20646 27027 20698
rect 27207 20646 27209 20698
rect 26963 20644 26969 20646
rect 27025 20644 27049 20646
rect 27105 20644 27129 20646
rect 27185 20644 27209 20646
rect 27265 20644 27271 20646
rect 26963 20635 27271 20644
rect 26792 20392 26844 20398
rect 26792 20334 26844 20340
rect 27356 20262 27384 20946
rect 28170 20496 28226 20505
rect 28170 20431 28226 20440
rect 26792 20256 26844 20262
rect 26792 20198 26844 20204
rect 27344 20256 27396 20262
rect 27344 20198 27396 20204
rect 27804 20256 27856 20262
rect 27804 20198 27856 20204
rect 26700 19304 26752 19310
rect 26700 19246 26752 19252
rect 26712 18630 26740 19246
rect 26804 19174 26832 20198
rect 27618 19952 27674 19961
rect 27618 19887 27620 19896
rect 27672 19887 27674 19896
rect 27620 19858 27672 19864
rect 27816 19854 27844 20198
rect 27988 19916 28040 19922
rect 27988 19858 28040 19864
rect 27804 19848 27856 19854
rect 27804 19790 27856 19796
rect 26963 19612 27271 19621
rect 26963 19610 26969 19612
rect 27025 19610 27049 19612
rect 27105 19610 27129 19612
rect 27185 19610 27209 19612
rect 27265 19610 27271 19612
rect 27025 19558 27027 19610
rect 27207 19558 27209 19610
rect 26963 19556 26969 19558
rect 27025 19556 27049 19558
rect 27105 19556 27129 19558
rect 27185 19556 27209 19558
rect 27265 19556 27271 19558
rect 26963 19547 27271 19556
rect 27250 19408 27306 19417
rect 27250 19343 27252 19352
rect 27304 19343 27306 19352
rect 27344 19372 27396 19378
rect 27252 19314 27304 19320
rect 27396 19320 27476 19334
rect 27344 19314 27476 19320
rect 27356 19306 27476 19314
rect 26792 19168 26844 19174
rect 26792 19110 26844 19116
rect 26976 19168 27028 19174
rect 26976 19110 27028 19116
rect 26700 18624 26752 18630
rect 26700 18566 26752 18572
rect 26606 17912 26662 17921
rect 26606 17847 26662 17856
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 26332 17196 26384 17202
rect 26332 17138 26384 17144
rect 26148 17128 26200 17134
rect 26148 17070 26200 17076
rect 26516 17128 26568 17134
rect 26516 17070 26568 17076
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 25870 16079 25926 16088
rect 25964 16108 26016 16114
rect 25686 14512 25742 14521
rect 25686 14447 25742 14456
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 25700 12986 25728 13806
rect 24952 12980 25004 12986
rect 24952 12922 25004 12928
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25688 12980 25740 12986
rect 25688 12922 25740 12928
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24872 11694 24900 12718
rect 25608 12442 25636 12786
rect 25884 12782 25912 16079
rect 25964 16050 26016 16056
rect 26068 15162 26096 16594
rect 26160 16590 26188 17070
rect 26424 16992 26476 16998
rect 26424 16934 26476 16940
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 26160 16046 26188 16526
rect 26436 16114 26464 16934
rect 26424 16108 26476 16114
rect 26424 16050 26476 16056
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 26160 15502 26188 15982
rect 26436 15638 26464 16050
rect 26424 15632 26476 15638
rect 26424 15574 26476 15580
rect 26332 15564 26384 15570
rect 26332 15506 26384 15512
rect 26148 15496 26200 15502
rect 26344 15450 26372 15506
rect 26148 15438 26200 15444
rect 26252 15422 26372 15450
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 26252 15042 26280 15422
rect 26332 15360 26384 15366
rect 26332 15302 26384 15308
rect 26424 15360 26476 15366
rect 26424 15302 26476 15308
rect 25976 15014 26280 15042
rect 25872 12776 25924 12782
rect 25872 12718 25924 12724
rect 25596 12436 25648 12442
rect 25596 12378 25648 12384
rect 25780 12436 25832 12442
rect 25780 12378 25832 12384
rect 25792 12306 25820 12378
rect 25780 12300 25832 12306
rect 25700 12260 25780 12288
rect 25700 11898 25728 12260
rect 25780 12242 25832 12248
rect 25976 12209 26004 15014
rect 26344 14958 26372 15302
rect 26436 15026 26464 15302
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 26332 14952 26384 14958
rect 26330 14920 26332 14929
rect 26384 14920 26386 14929
rect 26148 14884 26200 14890
rect 26330 14855 26386 14864
rect 26148 14826 26200 14832
rect 26160 14618 26188 14826
rect 26240 14816 26292 14822
rect 26240 14758 26292 14764
rect 26148 14612 26200 14618
rect 26148 14554 26200 14560
rect 26252 14482 26280 14758
rect 26240 14476 26292 14482
rect 26240 14418 26292 14424
rect 26056 14272 26108 14278
rect 26056 14214 26108 14220
rect 26068 14074 26096 14214
rect 26344 14090 26372 14855
rect 26424 14816 26476 14822
rect 26424 14758 26476 14764
rect 26056 14068 26108 14074
rect 26056 14010 26108 14016
rect 26252 14062 26372 14090
rect 26148 12708 26200 12714
rect 26148 12650 26200 12656
rect 25962 12200 26018 12209
rect 25962 12135 26018 12144
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25688 11892 25740 11898
rect 25688 11834 25740 11840
rect 25410 11792 25466 11801
rect 25410 11727 25466 11736
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 25228 11688 25280 11694
rect 25228 11630 25280 11636
rect 24676 11144 24728 11150
rect 24676 11086 24728 11092
rect 24688 10266 24716 11086
rect 24952 10668 25004 10674
rect 24952 10610 25004 10616
rect 24964 10266 24992 10610
rect 25136 10464 25188 10470
rect 25136 10406 25188 10412
rect 24676 10260 24728 10266
rect 24952 10260 25004 10266
rect 24676 10202 24728 10208
rect 24780 10220 24952 10248
rect 24780 10146 24808 10220
rect 24952 10202 25004 10208
rect 24504 10130 24808 10146
rect 25148 10130 25176 10406
rect 24492 10124 24808 10130
rect 24544 10118 24808 10124
rect 25136 10124 25188 10130
rect 24492 10066 24544 10072
rect 25136 10066 25188 10072
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24674 9616 24730 9625
rect 24412 9574 24624 9602
rect 24492 9512 24544 9518
rect 24492 9454 24544 9460
rect 24504 9382 24532 9454
rect 24492 9376 24544 9382
rect 24492 9318 24544 9324
rect 24492 7948 24544 7954
rect 24492 7890 24544 7896
rect 24400 7404 24452 7410
rect 24228 7364 24400 7392
rect 24124 7346 24176 7352
rect 24400 7346 24452 7352
rect 24044 7262 24256 7290
rect 23664 6996 23716 7002
rect 23664 6938 23716 6944
rect 22928 6860 22980 6866
rect 22928 6802 22980 6808
rect 23664 6860 23716 6866
rect 23664 6802 23716 6808
rect 22744 6792 22796 6798
rect 22468 6734 22520 6740
rect 22558 6760 22614 6769
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 22480 5914 22508 6734
rect 22744 6734 22796 6740
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 22558 6695 22614 6704
rect 22756 6458 22784 6734
rect 22744 6452 22796 6458
rect 22744 6394 22796 6400
rect 22836 6112 22888 6118
rect 22836 6054 22888 6060
rect 22468 5908 22520 5914
rect 22468 5850 22520 5856
rect 22192 5704 22244 5710
rect 21822 5672 21878 5681
rect 21822 5607 21878 5616
rect 22006 5672 22062 5681
rect 22192 5646 22244 5652
rect 22006 5607 22062 5616
rect 21652 5494 21864 5522
rect 21732 5364 21784 5370
rect 21732 5306 21784 5312
rect 21548 5024 21600 5030
rect 21548 4966 21600 4972
rect 21640 5024 21692 5030
rect 21640 4966 21692 4972
rect 21180 4684 21232 4690
rect 21180 4626 21232 4632
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 21008 4146 21036 4422
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 21192 4078 21220 4626
rect 21180 4072 21232 4078
rect 21180 4014 21232 4020
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 20824 2746 20944 2774
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20350 2408 20406 2417
rect 20732 2378 20760 2586
rect 20350 2343 20352 2352
rect 20404 2343 20406 2352
rect 20720 2372 20772 2378
rect 20352 2314 20404 2320
rect 20720 2314 20772 2320
rect 20536 2304 20588 2310
rect 20536 2246 20588 2252
rect 20076 1760 20128 1766
rect 20076 1702 20128 1708
rect 20088 1494 20116 1702
rect 20076 1488 20128 1494
rect 20076 1430 20128 1436
rect 20548 1290 20576 2246
rect 20732 1970 20760 2314
rect 20720 1964 20772 1970
rect 20720 1906 20772 1912
rect 20536 1284 20588 1290
rect 20536 1226 20588 1232
rect 20824 1018 20852 2746
rect 20904 1896 20956 1902
rect 20904 1838 20956 1844
rect 20916 1562 20944 1838
rect 20996 1828 21048 1834
rect 20996 1770 21048 1776
rect 21008 1737 21036 1770
rect 20994 1728 21050 1737
rect 20994 1663 21050 1672
rect 20904 1556 20956 1562
rect 20904 1498 20956 1504
rect 20904 1352 20956 1358
rect 20904 1294 20956 1300
rect 20916 1018 20944 1294
rect 21100 1222 21128 3674
rect 21376 3534 21404 4626
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21468 3058 21496 4422
rect 21560 3942 21588 4966
rect 21652 4826 21680 4966
rect 21744 4826 21772 5306
rect 21836 4826 21864 5494
rect 21640 4820 21692 4826
rect 21640 4762 21692 4768
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 21824 4820 21876 4826
rect 21824 4762 21876 4768
rect 22204 4690 22232 5646
rect 22480 4826 22508 5850
rect 22742 5808 22798 5817
rect 22742 5743 22798 5752
rect 22756 5166 22784 5743
rect 22744 5160 22796 5166
rect 22744 5102 22796 5108
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22468 4820 22520 4826
rect 22468 4762 22520 4768
rect 22192 4684 22244 4690
rect 22192 4626 22244 4632
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21560 3670 21588 3878
rect 21548 3664 21600 3670
rect 21548 3606 21600 3612
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 21560 2990 21588 3606
rect 22204 3602 22232 4626
rect 22480 4146 22508 4762
rect 22756 4690 22784 4966
rect 22848 4690 22876 6054
rect 23032 5370 23060 6734
rect 23296 6656 23348 6662
rect 23296 6598 23348 6604
rect 23308 6390 23336 6598
rect 23296 6384 23348 6390
rect 23296 6326 23348 6332
rect 23168 6012 23476 6021
rect 23168 6010 23174 6012
rect 23230 6010 23254 6012
rect 23310 6010 23334 6012
rect 23390 6010 23414 6012
rect 23470 6010 23476 6012
rect 23230 5958 23232 6010
rect 23412 5958 23414 6010
rect 23168 5956 23174 5958
rect 23230 5956 23254 5958
rect 23310 5956 23334 5958
rect 23390 5956 23414 5958
rect 23470 5956 23476 5958
rect 23168 5947 23476 5956
rect 23112 5568 23164 5574
rect 23112 5510 23164 5516
rect 23020 5364 23072 5370
rect 23020 5306 23072 5312
rect 23124 5302 23152 5510
rect 23112 5296 23164 5302
rect 23112 5238 23164 5244
rect 23676 5098 23704 6802
rect 23664 5092 23716 5098
rect 23664 5034 23716 5040
rect 23168 4924 23476 4933
rect 23168 4922 23174 4924
rect 23230 4922 23254 4924
rect 23310 4922 23334 4924
rect 23390 4922 23414 4924
rect 23470 4922 23476 4924
rect 23230 4870 23232 4922
rect 23412 4870 23414 4922
rect 23168 4868 23174 4870
rect 23230 4868 23254 4870
rect 23310 4868 23334 4870
rect 23390 4868 23414 4870
rect 23470 4868 23476 4870
rect 23168 4859 23476 4868
rect 23676 4690 23704 5034
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 22836 4684 22888 4690
rect 22836 4626 22888 4632
rect 23664 4684 23716 4690
rect 23664 4626 23716 4632
rect 23768 4146 23796 7262
rect 24124 6656 24176 6662
rect 24124 6598 24176 6604
rect 23848 6248 23900 6254
rect 23848 6190 23900 6196
rect 23860 5166 23888 6190
rect 24136 5953 24164 6598
rect 24122 5944 24178 5953
rect 24122 5879 24178 5888
rect 24228 5794 24256 7262
rect 24504 7206 24532 7890
rect 24492 7200 24544 7206
rect 24492 7142 24544 7148
rect 24596 6866 24624 9574
rect 24730 9574 24808 9602
rect 24674 9551 24730 9560
rect 24780 7426 24808 9574
rect 24872 9178 24900 9998
rect 24964 9178 24992 9998
rect 25240 9722 25268 11630
rect 25424 10470 25452 11727
rect 25504 11688 25556 11694
rect 25504 11630 25556 11636
rect 25516 11354 25544 11630
rect 25504 11348 25556 11354
rect 25504 11290 25556 11296
rect 25792 10606 25820 12038
rect 25976 11801 26004 12135
rect 25962 11792 26018 11801
rect 25962 11727 26018 11736
rect 26160 11354 26188 12650
rect 26148 11348 26200 11354
rect 26148 11290 26200 11296
rect 25688 10600 25740 10606
rect 25688 10542 25740 10548
rect 25780 10600 25832 10606
rect 25780 10542 25832 10548
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 25700 9722 25728 10542
rect 26056 9920 26108 9926
rect 26056 9862 26108 9868
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25688 9716 25740 9722
rect 25688 9658 25740 9664
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24952 9172 25004 9178
rect 24952 9114 25004 9120
rect 25044 8288 25096 8294
rect 25044 8230 25096 8236
rect 25056 8022 25084 8230
rect 25332 8090 25360 9522
rect 26068 9518 26096 9862
rect 25688 9512 25740 9518
rect 25688 9454 25740 9460
rect 26056 9512 26108 9518
rect 26056 9454 26108 9460
rect 26146 9480 26202 9489
rect 25700 9178 25728 9454
rect 26146 9415 26202 9424
rect 25780 9376 25832 9382
rect 25780 9318 25832 9324
rect 25872 9376 25924 9382
rect 25872 9318 25924 9324
rect 25688 9172 25740 9178
rect 25688 9114 25740 9120
rect 25792 9042 25820 9318
rect 25596 9036 25648 9042
rect 25596 8978 25648 8984
rect 25780 9036 25832 9042
rect 25780 8978 25832 8984
rect 25504 8968 25556 8974
rect 25504 8910 25556 8916
rect 25412 8832 25464 8838
rect 25412 8774 25464 8780
rect 25424 8566 25452 8774
rect 25412 8560 25464 8566
rect 25412 8502 25464 8508
rect 25410 8392 25466 8401
rect 25516 8378 25544 8910
rect 25608 8634 25636 8978
rect 25884 8634 25912 9318
rect 26160 9160 26188 9415
rect 26068 9132 26188 9160
rect 25596 8628 25648 8634
rect 25596 8570 25648 8576
rect 25872 8628 25924 8634
rect 25872 8570 25924 8576
rect 25466 8350 25544 8378
rect 25410 8327 25466 8336
rect 25320 8084 25372 8090
rect 25320 8026 25372 8032
rect 25044 8016 25096 8022
rect 25044 7958 25096 7964
rect 25228 7744 25280 7750
rect 25228 7686 25280 7692
rect 24780 7398 24992 7426
rect 24860 7336 24912 7342
rect 24860 7278 24912 7284
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24584 6860 24636 6866
rect 24584 6802 24636 6808
rect 24308 6316 24360 6322
rect 24308 6258 24360 6264
rect 24136 5766 24256 5794
rect 23848 5160 23900 5166
rect 23848 5102 23900 5108
rect 22468 4140 22520 4146
rect 23756 4140 23808 4146
rect 22520 4100 22600 4128
rect 22468 4082 22520 4088
rect 22468 3936 22520 3942
rect 22468 3878 22520 3884
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 21732 3528 21784 3534
rect 21732 3470 21784 3476
rect 21548 2984 21600 2990
rect 21548 2926 21600 2932
rect 21560 2650 21588 2926
rect 21548 2644 21600 2650
rect 21548 2586 21600 2592
rect 21272 1964 21324 1970
rect 21560 1952 21588 2586
rect 21640 2440 21692 2446
rect 21638 2408 21640 2417
rect 21692 2408 21694 2417
rect 21638 2343 21694 2352
rect 21744 2106 21772 3470
rect 21824 3392 21876 3398
rect 21824 3334 21876 3340
rect 21836 3194 21864 3334
rect 21824 3188 21876 3194
rect 22204 3176 22232 3538
rect 22480 3534 22508 3878
rect 22572 3738 22600 4100
rect 23756 4082 23808 4088
rect 23572 4072 23624 4078
rect 23572 4014 23624 4020
rect 23020 3936 23072 3942
rect 22926 3904 22982 3913
rect 23020 3878 23072 3884
rect 22926 3839 22982 3848
rect 22560 3732 22612 3738
rect 22560 3674 22612 3680
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22284 3188 22336 3194
rect 22204 3148 22284 3176
rect 21824 3130 21876 3136
rect 22284 3130 22336 3136
rect 22296 2514 22324 3130
rect 22940 3097 22968 3839
rect 23032 3602 23060 3878
rect 23168 3836 23476 3845
rect 23168 3834 23174 3836
rect 23230 3834 23254 3836
rect 23310 3834 23334 3836
rect 23390 3834 23414 3836
rect 23470 3834 23476 3836
rect 23230 3782 23232 3834
rect 23412 3782 23414 3834
rect 23168 3780 23174 3782
rect 23230 3780 23254 3782
rect 23310 3780 23334 3782
rect 23390 3780 23414 3782
rect 23470 3780 23476 3782
rect 23168 3771 23476 3780
rect 23020 3596 23072 3602
rect 23020 3538 23072 3544
rect 23480 3528 23532 3534
rect 23584 3516 23612 4014
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 23532 3488 23612 3516
rect 23480 3470 23532 3476
rect 23572 3188 23624 3194
rect 23572 3130 23624 3136
rect 22926 3088 22982 3097
rect 22926 3023 22982 3032
rect 23584 2922 23612 3130
rect 23676 2990 23704 3878
rect 23768 3602 23796 4082
rect 23756 3596 23808 3602
rect 23756 3538 23808 3544
rect 23860 3194 23888 5102
rect 23848 3188 23900 3194
rect 23848 3130 23900 3136
rect 23848 3052 23900 3058
rect 24032 3052 24084 3058
rect 23848 2994 23900 3000
rect 23952 3012 24032 3040
rect 23664 2984 23716 2990
rect 23664 2926 23716 2932
rect 23572 2916 23624 2922
rect 23572 2858 23624 2864
rect 23168 2748 23476 2757
rect 23168 2746 23174 2748
rect 23230 2746 23254 2748
rect 23310 2746 23334 2748
rect 23390 2746 23414 2748
rect 23470 2746 23476 2748
rect 23230 2694 23232 2746
rect 23412 2694 23414 2746
rect 23168 2692 23174 2694
rect 23230 2692 23254 2694
rect 23310 2692 23334 2694
rect 23390 2692 23414 2694
rect 23470 2692 23476 2694
rect 23168 2683 23476 2692
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 23584 2446 23612 2858
rect 23756 2508 23808 2514
rect 23756 2450 23808 2456
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 21916 2304 21968 2310
rect 21916 2246 21968 2252
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 23386 2272 23442 2281
rect 21732 2100 21784 2106
rect 21732 2042 21784 2048
rect 21324 1924 21588 1952
rect 21272 1906 21324 1912
rect 21560 1562 21588 1924
rect 21732 1896 21784 1902
rect 21732 1838 21784 1844
rect 21638 1728 21694 1737
rect 21744 1714 21772 1838
rect 21694 1686 21772 1714
rect 21638 1663 21694 1672
rect 21928 1562 21956 2246
rect 21548 1556 21600 1562
rect 21548 1498 21600 1504
rect 21916 1556 21968 1562
rect 21916 1498 21968 1504
rect 21364 1420 21416 1426
rect 21364 1362 21416 1368
rect 21272 1284 21324 1290
rect 21376 1272 21404 1362
rect 21324 1244 21404 1272
rect 21272 1226 21324 1232
rect 21088 1216 21140 1222
rect 21088 1158 21140 1164
rect 21362 1184 21418 1193
rect 21362 1119 21418 1128
rect 20812 1012 20864 1018
rect 20812 954 20864 960
rect 20904 1012 20956 1018
rect 20904 954 20956 960
rect 21376 882 21404 1119
rect 21548 1012 21600 1018
rect 21548 954 21600 960
rect 19340 876 19392 882
rect 19340 818 19392 824
rect 19708 876 19760 882
rect 19708 818 19760 824
rect 21364 876 21416 882
rect 21364 818 21416 824
rect 21560 746 21588 954
rect 22204 882 22232 2246
rect 23386 2207 23442 2216
rect 22834 2136 22890 2145
rect 22834 2071 22890 2080
rect 22468 1828 22520 1834
rect 22468 1770 22520 1776
rect 22480 1426 22508 1770
rect 22744 1760 22796 1766
rect 22744 1702 22796 1708
rect 22468 1420 22520 1426
rect 22468 1362 22520 1368
rect 22756 1358 22784 1702
rect 22848 1601 22876 2071
rect 23400 1970 23428 2207
rect 23388 1964 23440 1970
rect 23388 1906 23440 1912
rect 23400 1850 23428 1906
rect 22928 1828 22980 1834
rect 22928 1770 22980 1776
rect 23032 1822 23428 1850
rect 22834 1592 22890 1601
rect 22940 1562 22968 1770
rect 22834 1527 22890 1536
rect 22928 1556 22980 1562
rect 22928 1498 22980 1504
rect 22744 1352 22796 1358
rect 22744 1294 22796 1300
rect 23032 1018 23060 1822
rect 23492 1766 23520 2382
rect 23768 2038 23796 2450
rect 23756 2032 23808 2038
rect 23756 1974 23808 1980
rect 23480 1760 23532 1766
rect 23480 1702 23532 1708
rect 23664 1760 23716 1766
rect 23768 1737 23796 1974
rect 23860 1970 23888 2994
rect 23952 2854 23980 3012
rect 24032 2994 24084 3000
rect 23940 2848 23992 2854
rect 23940 2790 23992 2796
rect 24030 2680 24086 2689
rect 24030 2615 24032 2624
rect 24084 2615 24086 2624
rect 24032 2586 24084 2592
rect 24136 2530 24164 5766
rect 24216 5704 24268 5710
rect 24216 5646 24268 5652
rect 24228 5574 24256 5646
rect 24216 5568 24268 5574
rect 24216 5510 24268 5516
rect 24320 4758 24348 6258
rect 24400 6112 24452 6118
rect 24400 6054 24452 6060
rect 24412 5030 24440 6054
rect 24400 5024 24452 5030
rect 24400 4966 24452 4972
rect 24308 4752 24360 4758
rect 24308 4694 24360 4700
rect 24412 4128 24440 4966
rect 24780 4486 24808 7142
rect 24872 6662 24900 7278
rect 24964 6798 24992 7398
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24858 6216 24914 6225
rect 24858 6151 24914 6160
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24320 4100 24440 4128
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 24228 2854 24256 3674
rect 24320 3670 24348 4100
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 24400 4004 24452 4010
rect 24400 3946 24452 3952
rect 24308 3664 24360 3670
rect 24308 3606 24360 3612
rect 24216 2848 24268 2854
rect 24216 2790 24268 2796
rect 24044 2502 24164 2530
rect 24044 2106 24072 2502
rect 24124 2440 24176 2446
rect 24124 2382 24176 2388
rect 24032 2100 24084 2106
rect 24032 2042 24084 2048
rect 24136 1986 24164 2382
rect 23848 1964 23900 1970
rect 23848 1906 23900 1912
rect 24044 1958 24164 1986
rect 24228 1970 24256 2790
rect 24320 2446 24348 3606
rect 24308 2440 24360 2446
rect 24308 2382 24360 2388
rect 24216 1964 24268 1970
rect 23664 1702 23716 1708
rect 23754 1728 23810 1737
rect 23168 1660 23476 1669
rect 23168 1658 23174 1660
rect 23230 1658 23254 1660
rect 23310 1658 23334 1660
rect 23390 1658 23414 1660
rect 23470 1658 23476 1660
rect 23230 1606 23232 1658
rect 23412 1606 23414 1658
rect 23168 1604 23174 1606
rect 23230 1604 23254 1606
rect 23310 1604 23334 1606
rect 23390 1604 23414 1606
rect 23470 1604 23476 1606
rect 23168 1595 23476 1604
rect 23676 1562 23704 1702
rect 23754 1663 23810 1672
rect 23664 1556 23716 1562
rect 23664 1498 23716 1504
rect 23112 1488 23164 1494
rect 23112 1430 23164 1436
rect 23754 1456 23810 1465
rect 23124 1290 23152 1430
rect 23754 1391 23756 1400
rect 23808 1391 23810 1400
rect 23756 1362 23808 1368
rect 23112 1284 23164 1290
rect 23112 1226 23164 1232
rect 23020 1012 23072 1018
rect 23020 954 23072 960
rect 23480 1012 23532 1018
rect 23480 954 23532 960
rect 23492 921 23520 954
rect 23478 912 23534 921
rect 22192 876 22244 882
rect 23860 882 23888 1906
rect 23938 1456 23994 1465
rect 23938 1391 23940 1400
rect 23992 1391 23994 1400
rect 23940 1362 23992 1368
rect 24044 1358 24072 1958
rect 24216 1906 24268 1912
rect 24228 1578 24256 1906
rect 24136 1550 24256 1578
rect 24032 1352 24084 1358
rect 24032 1294 24084 1300
rect 23478 847 23534 856
rect 23848 876 23900 882
rect 22192 818 22244 824
rect 23848 818 23900 824
rect 23860 746 23888 818
rect 19064 740 19116 746
rect 19064 682 19116 688
rect 21548 740 21600 746
rect 21548 682 21600 688
rect 23848 740 23900 746
rect 23848 682 23900 688
rect 19076 406 19104 682
rect 23168 572 23476 581
rect 23168 570 23174 572
rect 23230 570 23254 572
rect 23310 570 23334 572
rect 23390 570 23414 572
rect 23470 570 23476 572
rect 23230 518 23232 570
rect 23412 518 23414 570
rect 23168 516 23174 518
rect 23230 516 23254 518
rect 23310 516 23334 518
rect 23390 516 23414 518
rect 23470 516 23476 518
rect 23168 507 23476 516
rect 19064 400 19116 406
rect 19064 342 19116 348
rect 24044 270 24072 1294
rect 24136 678 24164 1550
rect 24216 1488 24268 1494
rect 24320 1476 24348 2382
rect 24268 1448 24348 1476
rect 24216 1430 24268 1436
rect 24308 1352 24360 1358
rect 24308 1294 24360 1300
rect 24320 882 24348 1294
rect 24308 876 24360 882
rect 24308 818 24360 824
rect 24412 814 24440 3946
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 24504 2689 24532 2926
rect 24490 2680 24546 2689
rect 24490 2615 24546 2624
rect 24596 2446 24624 3334
rect 24676 2848 24728 2854
rect 24676 2790 24728 2796
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 24504 1970 24532 2246
rect 24492 1964 24544 1970
rect 24492 1906 24544 1912
rect 24492 1760 24544 1766
rect 24492 1702 24544 1708
rect 24400 808 24452 814
rect 24400 750 24452 756
rect 24124 672 24176 678
rect 24124 614 24176 620
rect 24504 406 24532 1702
rect 24688 1358 24716 2790
rect 24780 2530 24808 4014
rect 24872 3738 24900 6151
rect 24952 5568 25004 5574
rect 24952 5510 25004 5516
rect 24964 5234 24992 5510
rect 24952 5228 25004 5234
rect 24952 5170 25004 5176
rect 25240 5030 25268 7686
rect 25688 7268 25740 7274
rect 25688 7210 25740 7216
rect 25504 6248 25556 6254
rect 25504 6190 25556 6196
rect 25516 5302 25544 6190
rect 25700 5914 25728 7210
rect 25780 6112 25832 6118
rect 25780 6054 25832 6060
rect 25872 6112 25924 6118
rect 25872 6054 25924 6060
rect 25792 5914 25820 6054
rect 25688 5908 25740 5914
rect 25688 5850 25740 5856
rect 25780 5908 25832 5914
rect 25780 5850 25832 5856
rect 25504 5296 25556 5302
rect 25504 5238 25556 5244
rect 25228 5024 25280 5030
rect 25228 4966 25280 4972
rect 25884 4146 25912 6054
rect 26068 5778 26096 9132
rect 26146 9072 26202 9081
rect 26146 9007 26148 9016
rect 26200 9007 26202 9016
rect 26148 8978 26200 8984
rect 26146 7440 26202 7449
rect 26146 7375 26202 7384
rect 26160 7342 26188 7375
rect 26148 7336 26200 7342
rect 26148 7278 26200 7284
rect 26160 6934 26188 7278
rect 26148 6928 26200 6934
rect 26148 6870 26200 6876
rect 26160 6322 26188 6870
rect 26252 6866 26280 14062
rect 26436 13938 26464 14758
rect 26528 14074 26556 17070
rect 26608 16040 26660 16046
rect 26608 15982 26660 15988
rect 26620 14074 26648 15982
rect 26712 14958 26740 18566
rect 26804 17882 26832 19110
rect 26988 18970 27016 19110
rect 26976 18964 27028 18970
rect 26976 18906 27028 18912
rect 26884 18828 26936 18834
rect 26884 18770 26936 18776
rect 26792 17876 26844 17882
rect 26896 17864 26924 18770
rect 26963 18524 27271 18533
rect 26963 18522 26969 18524
rect 27025 18522 27049 18524
rect 27105 18522 27129 18524
rect 27185 18522 27209 18524
rect 27265 18522 27271 18524
rect 27025 18470 27027 18522
rect 27207 18470 27209 18522
rect 26963 18468 26969 18470
rect 27025 18468 27049 18470
rect 27105 18468 27129 18470
rect 27185 18468 27209 18470
rect 27265 18468 27271 18470
rect 26963 18459 27271 18468
rect 27068 17876 27120 17882
rect 26896 17836 27068 17864
rect 26792 17818 26844 17824
rect 27068 17818 27120 17824
rect 26804 16998 26832 17818
rect 26884 17672 26936 17678
rect 26884 17614 26936 17620
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 26804 16590 26832 16934
rect 26792 16584 26844 16590
rect 26792 16526 26844 16532
rect 26792 16448 26844 16454
rect 26792 16390 26844 16396
rect 26804 15570 26832 16390
rect 26792 15564 26844 15570
rect 26792 15506 26844 15512
rect 26792 15360 26844 15366
rect 26792 15302 26844 15308
rect 26700 14952 26752 14958
rect 26700 14894 26752 14900
rect 26804 14550 26832 15302
rect 26792 14544 26844 14550
rect 26792 14486 26844 14492
rect 26700 14272 26752 14278
rect 26700 14214 26752 14220
rect 26792 14272 26844 14278
rect 26792 14214 26844 14220
rect 26516 14068 26568 14074
rect 26516 14010 26568 14016
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26424 13932 26476 13938
rect 26424 13874 26476 13880
rect 26436 13326 26464 13874
rect 26516 13728 26568 13734
rect 26516 13670 26568 13676
rect 26528 13546 26556 13670
rect 26528 13518 26648 13546
rect 26620 13326 26648 13518
rect 26424 13320 26476 13326
rect 26424 13262 26476 13268
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26436 12782 26464 13262
rect 26712 12850 26740 14214
rect 26804 13954 26832 14214
rect 26896 14056 26924 17614
rect 26963 17436 27271 17445
rect 26963 17434 26969 17436
rect 27025 17434 27049 17436
rect 27105 17434 27129 17436
rect 27185 17434 27209 17436
rect 27265 17434 27271 17436
rect 27025 17382 27027 17434
rect 27207 17382 27209 17434
rect 26963 17380 26969 17382
rect 27025 17380 27049 17382
rect 27105 17380 27129 17382
rect 27185 17380 27209 17382
rect 27265 17380 27271 17382
rect 26963 17371 27271 17380
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 27264 16538 27292 16594
rect 27264 16510 27384 16538
rect 26963 16348 27271 16357
rect 26963 16346 26969 16348
rect 27025 16346 27049 16348
rect 27105 16346 27129 16348
rect 27185 16346 27209 16348
rect 27265 16346 27271 16348
rect 27025 16294 27027 16346
rect 27207 16294 27209 16346
rect 26963 16292 26969 16294
rect 27025 16292 27049 16294
rect 27105 16292 27129 16294
rect 27185 16292 27209 16294
rect 27265 16292 27271 16294
rect 26963 16283 27271 16292
rect 27160 16244 27212 16250
rect 27160 16186 27212 16192
rect 26974 16144 27030 16153
rect 26974 16079 27030 16088
rect 26988 15570 27016 16079
rect 27172 16046 27200 16186
rect 27160 16040 27212 16046
rect 27160 15982 27212 15988
rect 26976 15564 27028 15570
rect 26976 15506 27028 15512
rect 26988 15366 27016 15506
rect 26976 15360 27028 15366
rect 26976 15302 27028 15308
rect 26963 15260 27271 15269
rect 26963 15258 26969 15260
rect 27025 15258 27049 15260
rect 27105 15258 27129 15260
rect 27185 15258 27209 15260
rect 27265 15258 27271 15260
rect 27025 15206 27027 15258
rect 27207 15206 27209 15258
rect 26963 15204 26969 15206
rect 27025 15204 27049 15206
rect 27105 15204 27129 15206
rect 27185 15204 27209 15206
rect 27265 15204 27271 15206
rect 26963 15195 27271 15204
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 27080 15026 27108 15098
rect 27068 15020 27120 15026
rect 27068 14962 27120 14968
rect 27252 15020 27304 15026
rect 27252 14962 27304 14968
rect 27080 14550 27108 14962
rect 27264 14634 27292 14962
rect 27172 14606 27292 14634
rect 27068 14544 27120 14550
rect 27068 14486 27120 14492
rect 27080 14278 27108 14486
rect 27172 14278 27200 14606
rect 27252 14544 27304 14550
rect 27252 14486 27304 14492
rect 27264 14385 27292 14486
rect 27250 14376 27306 14385
rect 27250 14311 27306 14320
rect 27068 14272 27120 14278
rect 27068 14214 27120 14220
rect 27160 14272 27212 14278
rect 27160 14214 27212 14220
rect 26963 14172 27271 14181
rect 26963 14170 26969 14172
rect 27025 14170 27049 14172
rect 27105 14170 27129 14172
rect 27185 14170 27209 14172
rect 27265 14170 27271 14172
rect 27025 14118 27027 14170
rect 27207 14118 27209 14170
rect 26963 14116 26969 14118
rect 27025 14116 27049 14118
rect 27105 14116 27129 14118
rect 27185 14116 27209 14118
rect 27265 14116 27271 14118
rect 26963 14107 27271 14116
rect 26896 14028 27292 14056
rect 26804 13926 27108 13954
rect 26804 13326 26832 13926
rect 26976 13864 27028 13870
rect 26896 13824 26976 13852
rect 26896 13569 26924 13824
rect 26976 13806 27028 13812
rect 27080 13818 27108 13926
rect 27264 13818 27292 14028
rect 27356 13938 27384 16510
rect 27448 16425 27476 19306
rect 27528 19304 27580 19310
rect 27528 19246 27580 19252
rect 27434 16416 27490 16425
rect 27434 16351 27490 16360
rect 27540 16130 27568 19246
rect 27618 18184 27674 18193
rect 27618 18119 27674 18128
rect 27632 16658 27660 18119
rect 27712 17264 27764 17270
rect 27712 17206 27764 17212
rect 27724 16969 27752 17206
rect 27710 16960 27766 16969
rect 27710 16895 27766 16904
rect 27620 16652 27672 16658
rect 27620 16594 27672 16600
rect 27448 16102 27568 16130
rect 27620 16176 27672 16182
rect 27620 16118 27672 16124
rect 27448 15162 27476 16102
rect 27528 15972 27580 15978
rect 27528 15914 27580 15920
rect 27540 15706 27568 15914
rect 27528 15700 27580 15706
rect 27528 15642 27580 15648
rect 27632 15570 27660 16118
rect 27710 15736 27766 15745
rect 27710 15671 27766 15680
rect 27620 15564 27672 15570
rect 27620 15506 27672 15512
rect 27632 15337 27660 15506
rect 27618 15328 27674 15337
rect 27618 15263 27674 15272
rect 27436 15156 27488 15162
rect 27436 15098 27488 15104
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27632 14362 27660 14962
rect 27540 14334 27660 14362
rect 27540 14074 27568 14334
rect 27620 14272 27672 14278
rect 27620 14214 27672 14220
rect 27436 14068 27488 14074
rect 27436 14010 27488 14016
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 27344 13932 27396 13938
rect 27344 13874 27396 13880
rect 27080 13790 27200 13818
rect 27264 13790 27384 13818
rect 27172 13734 27200 13790
rect 27160 13728 27212 13734
rect 27160 13670 27212 13676
rect 26882 13560 26938 13569
rect 26882 13495 26938 13504
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 26988 13394 27016 13466
rect 26976 13388 27028 13394
rect 26976 13330 27028 13336
rect 26792 13320 26844 13326
rect 26844 13268 26924 13274
rect 26792 13262 26924 13268
rect 26804 13246 26924 13262
rect 26792 13184 26844 13190
rect 26792 13126 26844 13132
rect 26700 12844 26752 12850
rect 26700 12786 26752 12792
rect 26424 12776 26476 12782
rect 26424 12718 26476 12724
rect 26804 12434 26832 13126
rect 26896 12646 26924 13246
rect 26963 13084 27271 13093
rect 26963 13082 26969 13084
rect 27025 13082 27049 13084
rect 27105 13082 27129 13084
rect 27185 13082 27209 13084
rect 27265 13082 27271 13084
rect 27025 13030 27027 13082
rect 27207 13030 27209 13082
rect 26963 13028 26969 13030
rect 27025 13028 27049 13030
rect 27105 13028 27129 13030
rect 27185 13028 27209 13030
rect 27265 13028 27271 13030
rect 26963 13019 27271 13028
rect 27160 12980 27212 12986
rect 27160 12922 27212 12928
rect 27172 12850 27200 12922
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 26884 12640 26936 12646
rect 27356 12628 27384 13790
rect 27448 13530 27476 14010
rect 27528 13864 27580 13870
rect 27528 13806 27580 13812
rect 27436 13524 27488 13530
rect 27436 13466 27488 13472
rect 27540 12889 27568 13806
rect 27526 12880 27582 12889
rect 27526 12815 27582 12824
rect 27528 12708 27580 12714
rect 27528 12650 27580 12656
rect 27436 12640 27488 12646
rect 27356 12600 27436 12628
rect 26884 12582 26936 12588
rect 27436 12582 27488 12588
rect 26712 12406 26832 12434
rect 27158 12472 27214 12481
rect 27540 12442 27568 12650
rect 27632 12442 27660 14214
rect 27724 12918 27752 15671
rect 27712 12912 27764 12918
rect 27712 12854 27764 12860
rect 27158 12407 27214 12416
rect 27528 12436 27580 12442
rect 26516 12300 26568 12306
rect 26516 12242 26568 12248
rect 26332 12096 26384 12102
rect 26384 12056 26464 12084
rect 26332 12038 26384 12044
rect 26436 11150 26464 12056
rect 26528 11762 26556 12242
rect 26516 11756 26568 11762
rect 26516 11698 26568 11704
rect 26424 11144 26476 11150
rect 26330 11112 26386 11121
rect 26424 11086 26476 11092
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26330 11047 26386 11056
rect 26344 10266 26372 11047
rect 26332 10260 26384 10266
rect 26332 10202 26384 10208
rect 26436 10062 26464 11086
rect 26516 10192 26568 10198
rect 26516 10134 26568 10140
rect 26424 10056 26476 10062
rect 26424 9998 26476 10004
rect 26436 9674 26464 9998
rect 26344 9646 26464 9674
rect 26344 9042 26372 9646
rect 26424 9512 26476 9518
rect 26424 9454 26476 9460
rect 26332 9036 26384 9042
rect 26332 8978 26384 8984
rect 26436 8634 26464 9454
rect 26528 9382 26556 10134
rect 26620 10062 26648 11086
rect 26608 10056 26660 10062
rect 26608 9998 26660 10004
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26620 8974 26648 9998
rect 26608 8968 26660 8974
rect 26514 8936 26570 8945
rect 26608 8910 26660 8916
rect 26514 8871 26570 8880
rect 26424 8628 26476 8634
rect 26424 8570 26476 8576
rect 26528 8430 26556 8871
rect 26516 8424 26568 8430
rect 26516 8366 26568 8372
rect 26424 7948 26476 7954
rect 26424 7890 26476 7896
rect 26240 6860 26292 6866
rect 26240 6802 26292 6808
rect 26148 6316 26200 6322
rect 26148 6258 26200 6264
rect 26436 6202 26464 7890
rect 26608 7880 26660 7886
rect 26608 7822 26660 7828
rect 26620 7206 26648 7822
rect 26608 7200 26660 7206
rect 26608 7142 26660 7148
rect 26252 6174 26464 6202
rect 26516 6248 26568 6254
rect 26516 6190 26568 6196
rect 26056 5772 26108 5778
rect 26108 5732 26188 5760
rect 26056 5714 26108 5720
rect 25964 5568 26016 5574
rect 25964 5510 26016 5516
rect 26056 5568 26108 5574
rect 26056 5510 26108 5516
rect 25976 5234 26004 5510
rect 25964 5228 26016 5234
rect 25964 5170 26016 5176
rect 26068 4826 26096 5510
rect 26056 4820 26108 4826
rect 26056 4762 26108 4768
rect 26160 4690 26188 5732
rect 26148 4684 26200 4690
rect 26148 4626 26200 4632
rect 25872 4140 25924 4146
rect 25872 4082 25924 4088
rect 25136 4072 25188 4078
rect 25188 4032 25268 4060
rect 25136 4014 25188 4020
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 25240 3058 25268 4032
rect 26252 4026 26280 6174
rect 26332 6112 26384 6118
rect 26332 6054 26384 6060
rect 26424 6112 26476 6118
rect 26424 6054 26476 6060
rect 26344 5778 26372 6054
rect 26332 5772 26384 5778
rect 26332 5714 26384 5720
rect 26332 5092 26384 5098
rect 26332 5034 26384 5040
rect 26160 3998 26280 4026
rect 26056 3936 26108 3942
rect 26056 3878 26108 3884
rect 25688 3596 25740 3602
rect 25688 3538 25740 3544
rect 25700 3398 25728 3538
rect 25320 3392 25372 3398
rect 25320 3334 25372 3340
rect 25596 3392 25648 3398
rect 25596 3334 25648 3340
rect 25688 3392 25740 3398
rect 25688 3334 25740 3340
rect 25228 3052 25280 3058
rect 25228 2994 25280 3000
rect 24780 2502 24900 2530
rect 24768 2440 24820 2446
rect 24768 2382 24820 2388
rect 24780 2106 24808 2382
rect 24768 2100 24820 2106
rect 24768 2042 24820 2048
rect 24872 1986 24900 2502
rect 24872 1970 24992 1986
rect 24872 1964 25004 1970
rect 24872 1958 24952 1964
rect 24872 1766 24900 1958
rect 24952 1906 25004 1912
rect 24860 1760 24912 1766
rect 24860 1702 24912 1708
rect 24952 1760 25004 1766
rect 24952 1702 25004 1708
rect 24860 1556 24912 1562
rect 24860 1498 24912 1504
rect 24676 1352 24728 1358
rect 24676 1294 24728 1300
rect 24492 400 24544 406
rect 24492 342 24544 348
rect 24032 264 24084 270
rect 18234 232 18290 241
rect 17868 196 17920 202
rect 24032 206 24084 212
rect 18234 167 18290 176
rect 17868 138 17920 144
rect 24872 105 24900 1498
rect 24964 377 24992 1702
rect 25240 882 25268 2994
rect 25332 2514 25360 3334
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 25504 2508 25556 2514
rect 25504 2450 25556 2456
rect 25516 2281 25544 2450
rect 25502 2272 25558 2281
rect 25502 2207 25558 2216
rect 25318 1728 25374 1737
rect 25318 1663 25374 1672
rect 25332 1426 25360 1663
rect 25320 1420 25372 1426
rect 25320 1362 25372 1368
rect 25608 1358 25636 3334
rect 25700 2650 25728 3334
rect 25780 3188 25832 3194
rect 25780 3130 25832 3136
rect 25792 2650 25820 3130
rect 26068 2854 26096 3878
rect 26160 3738 26188 3998
rect 26148 3732 26200 3738
rect 26148 3674 26200 3680
rect 26344 3058 26372 5034
rect 26436 4146 26464 6054
rect 26528 5098 26556 6190
rect 26620 6118 26648 7142
rect 26712 6866 26740 12406
rect 27172 12306 27200 12407
rect 27528 12378 27580 12384
rect 27620 12436 27672 12442
rect 27620 12378 27672 12384
rect 27160 12300 27212 12306
rect 27540 12288 27568 12378
rect 27160 12242 27212 12248
rect 27356 12260 27568 12288
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 26896 11898 26924 12174
rect 26963 11996 27271 12005
rect 26963 11994 26969 11996
rect 27025 11994 27049 11996
rect 27105 11994 27129 11996
rect 27185 11994 27209 11996
rect 27265 11994 27271 11996
rect 27025 11942 27027 11994
rect 27207 11942 27209 11994
rect 26963 11940 26969 11942
rect 27025 11940 27049 11942
rect 27105 11940 27129 11942
rect 27185 11940 27209 11942
rect 27265 11940 27271 11942
rect 26963 11931 27271 11940
rect 26884 11892 26936 11898
rect 26884 11834 26936 11840
rect 26976 11892 27028 11898
rect 26976 11834 27028 11840
rect 26988 11558 27016 11834
rect 26976 11552 27028 11558
rect 26976 11494 27028 11500
rect 26884 11144 26936 11150
rect 26804 11104 26884 11132
rect 26804 10810 26832 11104
rect 26884 11086 26936 11092
rect 26988 10996 27016 11494
rect 26896 10968 27016 10996
rect 26792 10804 26844 10810
rect 26792 10746 26844 10752
rect 26896 8922 26924 10968
rect 26963 10908 27271 10917
rect 26963 10906 26969 10908
rect 27025 10906 27049 10908
rect 27105 10906 27129 10908
rect 27185 10906 27209 10908
rect 27265 10906 27271 10908
rect 27025 10854 27027 10906
rect 27207 10854 27209 10906
rect 26963 10852 26969 10854
rect 27025 10852 27049 10854
rect 27105 10852 27129 10854
rect 27185 10852 27209 10854
rect 27265 10852 27271 10854
rect 26963 10843 27271 10852
rect 26963 9820 27271 9829
rect 26963 9818 26969 9820
rect 27025 9818 27049 9820
rect 27105 9818 27129 9820
rect 27185 9818 27209 9820
rect 27265 9818 27271 9820
rect 27025 9766 27027 9818
rect 27207 9766 27209 9818
rect 26963 9764 26969 9766
rect 27025 9764 27049 9766
rect 27105 9764 27129 9766
rect 27185 9764 27209 9766
rect 27265 9764 27271 9766
rect 26963 9755 27271 9764
rect 26976 9580 27028 9586
rect 26976 9522 27028 9528
rect 26988 9081 27016 9522
rect 26974 9072 27030 9081
rect 26974 9007 27030 9016
rect 26804 8894 26924 8922
rect 26804 8362 26832 8894
rect 26884 8832 26936 8838
rect 26884 8774 26936 8780
rect 26792 8356 26844 8362
rect 26792 8298 26844 8304
rect 26700 6860 26752 6866
rect 26700 6802 26752 6808
rect 26896 6322 26924 8774
rect 26963 8732 27271 8741
rect 26963 8730 26969 8732
rect 27025 8730 27049 8732
rect 27105 8730 27129 8732
rect 27185 8730 27209 8732
rect 27265 8730 27271 8732
rect 27025 8678 27027 8730
rect 27207 8678 27209 8730
rect 26963 8676 26969 8678
rect 27025 8676 27049 8678
rect 27105 8676 27129 8678
rect 27185 8676 27209 8678
rect 27265 8676 27271 8678
rect 26963 8667 27271 8676
rect 27356 8430 27384 12260
rect 27816 12238 27844 19790
rect 27896 18896 27948 18902
rect 27894 18864 27896 18873
rect 27948 18864 27950 18873
rect 27894 18799 27950 18808
rect 27908 18698 27936 18799
rect 27896 18692 27948 18698
rect 27896 18634 27948 18640
rect 27896 18148 27948 18154
rect 27896 18090 27948 18096
rect 27908 16794 27936 18090
rect 28000 16946 28028 19858
rect 28184 19242 28212 20431
rect 28264 19848 28316 19854
rect 28264 19790 28316 19796
rect 28172 19236 28224 19242
rect 28172 19178 28224 19184
rect 28184 18714 28212 19178
rect 28276 18834 28304 19790
rect 28264 18828 28316 18834
rect 28264 18770 28316 18776
rect 28092 18686 28212 18714
rect 28092 17134 28120 18686
rect 28172 18624 28224 18630
rect 28172 18566 28224 18572
rect 28080 17128 28132 17134
rect 28080 17070 28132 17076
rect 28000 16918 28120 16946
rect 27896 16788 27948 16794
rect 27896 16730 27948 16736
rect 27988 16720 28040 16726
rect 27986 16688 27988 16697
rect 28040 16688 28042 16697
rect 27986 16623 28042 16632
rect 27896 16584 27948 16590
rect 27896 16526 27948 16532
rect 27908 15745 27936 16526
rect 27894 15736 27950 15745
rect 27894 15671 27950 15680
rect 27908 15473 27936 15671
rect 27988 15496 28040 15502
rect 27894 15464 27950 15473
rect 27988 15438 28040 15444
rect 27894 15399 27950 15408
rect 27896 14952 27948 14958
rect 27896 14894 27948 14900
rect 27908 14550 27936 14894
rect 27896 14544 27948 14550
rect 27896 14486 27948 14492
rect 27908 14346 27936 14486
rect 28000 14482 28028 15438
rect 28092 15162 28120 16918
rect 28184 16590 28212 18566
rect 28368 18465 28396 21286
rect 28354 18456 28410 18465
rect 28354 18391 28410 18400
rect 28356 18080 28408 18086
rect 28356 18022 28408 18028
rect 28264 17808 28316 17814
rect 28264 17750 28316 17756
rect 28172 16584 28224 16590
rect 28276 16561 28304 17750
rect 28368 17241 28396 18022
rect 28460 17338 28488 21354
rect 28552 19922 28580 22238
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 30392 21690 30420 22170
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 29460 21684 29512 21690
rect 29460 21626 29512 21632
rect 30380 21684 30432 21690
rect 30380 21626 30432 21632
rect 29092 21480 29144 21486
rect 29092 21422 29144 21428
rect 29276 21480 29328 21486
rect 29276 21422 29328 21428
rect 28632 20936 28684 20942
rect 28632 20878 28684 20884
rect 28540 19916 28592 19922
rect 28540 19858 28592 19864
rect 28540 18624 28592 18630
rect 28540 18566 28592 18572
rect 28552 18222 28580 18566
rect 28540 18216 28592 18222
rect 28540 18158 28592 18164
rect 28540 17876 28592 17882
rect 28540 17818 28592 17824
rect 28552 17678 28580 17818
rect 28540 17672 28592 17678
rect 28540 17614 28592 17620
rect 28448 17332 28500 17338
rect 28448 17274 28500 17280
rect 28354 17232 28410 17241
rect 28354 17167 28410 17176
rect 28552 16998 28580 17614
rect 28540 16992 28592 16998
rect 28540 16934 28592 16940
rect 28356 16788 28408 16794
rect 28356 16730 28408 16736
rect 28172 16526 28224 16532
rect 28262 16552 28318 16561
rect 28262 16487 28318 16496
rect 28264 16448 28316 16454
rect 28264 16390 28316 16396
rect 28172 16040 28224 16046
rect 28172 15982 28224 15988
rect 28184 15502 28212 15982
rect 28276 15881 28304 16390
rect 28368 16250 28396 16730
rect 28448 16584 28500 16590
rect 28448 16526 28500 16532
rect 28538 16552 28594 16561
rect 28460 16250 28488 16526
rect 28538 16487 28594 16496
rect 28356 16244 28408 16250
rect 28356 16186 28408 16192
rect 28448 16244 28500 16250
rect 28448 16186 28500 16192
rect 28262 15872 28318 15881
rect 28262 15807 28318 15816
rect 28264 15700 28316 15706
rect 28264 15642 28316 15648
rect 28172 15496 28224 15502
rect 28172 15438 28224 15444
rect 28170 15328 28226 15337
rect 28170 15263 28226 15272
rect 28080 15156 28132 15162
rect 28080 15098 28132 15104
rect 27988 14476 28040 14482
rect 27988 14418 28040 14424
rect 27896 14340 27948 14346
rect 27896 14282 27948 14288
rect 28000 12782 28028 14418
rect 27988 12776 28040 12782
rect 27988 12718 28040 12724
rect 28000 12306 28028 12718
rect 27988 12300 28040 12306
rect 27988 12242 28040 12248
rect 27804 12232 27856 12238
rect 27804 12174 27856 12180
rect 27620 12096 27672 12102
rect 27620 12038 27672 12044
rect 27528 11552 27580 11558
rect 27632 11540 27660 12038
rect 27580 11512 27660 11540
rect 27712 11552 27764 11558
rect 27528 11494 27580 11500
rect 27712 11494 27764 11500
rect 27528 11144 27580 11150
rect 27528 11086 27580 11092
rect 27434 10160 27490 10169
rect 27434 10095 27490 10104
rect 27344 8424 27396 8430
rect 27264 8384 27344 8412
rect 27264 7886 27292 8384
rect 27344 8366 27396 8372
rect 27252 7880 27304 7886
rect 27448 7834 27476 10095
rect 27540 9654 27568 11086
rect 27528 9648 27580 9654
rect 27528 9590 27580 9596
rect 27528 9444 27580 9450
rect 27528 9386 27580 9392
rect 27540 9178 27568 9386
rect 27528 9172 27580 9178
rect 27528 9114 27580 9120
rect 27724 8922 27752 11494
rect 27816 10674 27844 12174
rect 28184 11218 28212 15263
rect 28276 14618 28304 15642
rect 28356 15360 28408 15366
rect 28356 15302 28408 15308
rect 28368 14958 28396 15302
rect 28356 14952 28408 14958
rect 28356 14894 28408 14900
rect 28460 14657 28488 16186
rect 28552 15609 28580 16487
rect 28538 15600 28594 15609
rect 28538 15535 28594 15544
rect 28540 15496 28592 15502
rect 28540 15438 28592 15444
rect 28446 14648 28502 14657
rect 28264 14612 28316 14618
rect 28446 14583 28502 14592
rect 28264 14554 28316 14560
rect 28276 12170 28304 14554
rect 28356 14408 28408 14414
rect 28356 14350 28408 14356
rect 28264 12164 28316 12170
rect 28264 12106 28316 12112
rect 28172 11212 28224 11218
rect 28172 11154 28224 11160
rect 28080 11076 28132 11082
rect 28080 11018 28132 11024
rect 27804 10668 27856 10674
rect 27804 10610 27856 10616
rect 27896 9376 27948 9382
rect 27896 9318 27948 9324
rect 27908 9178 27936 9318
rect 27896 9172 27948 9178
rect 27896 9114 27948 9120
rect 27540 8894 27752 8922
rect 27540 7954 27568 8894
rect 27804 8628 27856 8634
rect 27804 8570 27856 8576
rect 27816 8090 27844 8570
rect 28092 8498 28120 11018
rect 28184 10130 28212 11154
rect 28172 10124 28224 10130
rect 28172 10066 28224 10072
rect 28264 10056 28316 10062
rect 28264 9998 28316 10004
rect 28172 9920 28224 9926
rect 28172 9862 28224 9868
rect 28080 8492 28132 8498
rect 28080 8434 28132 8440
rect 28080 8288 28132 8294
rect 28080 8230 28132 8236
rect 27804 8084 27856 8090
rect 27804 8026 27856 8032
rect 27528 7948 27580 7954
rect 27528 7890 27580 7896
rect 27252 7822 27304 7828
rect 27356 7806 27476 7834
rect 27712 7880 27764 7886
rect 27712 7822 27764 7828
rect 26963 7644 27271 7653
rect 26963 7642 26969 7644
rect 27025 7642 27049 7644
rect 27105 7642 27129 7644
rect 27185 7642 27209 7644
rect 27265 7642 27271 7644
rect 27025 7590 27027 7642
rect 27207 7590 27209 7642
rect 26963 7588 26969 7590
rect 27025 7588 27049 7590
rect 27105 7588 27129 7590
rect 27185 7588 27209 7590
rect 27265 7588 27271 7590
rect 26963 7579 27271 7588
rect 26976 7200 27028 7206
rect 26976 7142 27028 7148
rect 26988 6905 27016 7142
rect 27356 6934 27384 7806
rect 27436 7744 27488 7750
rect 27436 7686 27488 7692
rect 27344 6928 27396 6934
rect 26974 6896 27030 6905
rect 27344 6870 27396 6876
rect 26974 6831 27030 6840
rect 27344 6724 27396 6730
rect 27344 6666 27396 6672
rect 26963 6556 27271 6565
rect 26963 6554 26969 6556
rect 27025 6554 27049 6556
rect 27105 6554 27129 6556
rect 27185 6554 27209 6556
rect 27265 6554 27271 6556
rect 27025 6502 27027 6554
rect 27207 6502 27209 6554
rect 26963 6500 26969 6502
rect 27025 6500 27049 6502
rect 27105 6500 27129 6502
rect 27185 6500 27209 6502
rect 27265 6500 27271 6502
rect 26963 6491 27271 6500
rect 26700 6316 26752 6322
rect 26700 6258 26752 6264
rect 26884 6316 26936 6322
rect 26884 6258 26936 6264
rect 26608 6112 26660 6118
rect 26608 6054 26660 6060
rect 26620 5234 26648 6054
rect 26608 5228 26660 5234
rect 26608 5170 26660 5176
rect 26516 5092 26568 5098
rect 26516 5034 26568 5040
rect 26516 4616 26568 4622
rect 26620 4570 26648 5170
rect 26712 5166 26740 6258
rect 26792 6180 26844 6186
rect 26792 6122 26844 6128
rect 26804 6066 26832 6122
rect 26804 6038 27292 6066
rect 26790 5944 26846 5953
rect 26790 5879 26846 5888
rect 26804 5710 26832 5879
rect 27264 5710 27292 6038
rect 26792 5704 26844 5710
rect 26792 5646 26844 5652
rect 27160 5704 27212 5710
rect 27160 5646 27212 5652
rect 27252 5704 27304 5710
rect 27252 5646 27304 5652
rect 27172 5574 27200 5646
rect 27160 5568 27212 5574
rect 27160 5510 27212 5516
rect 26963 5468 27271 5477
rect 26963 5466 26969 5468
rect 27025 5466 27049 5468
rect 27105 5466 27129 5468
rect 27185 5466 27209 5468
rect 27265 5466 27271 5468
rect 27025 5414 27027 5466
rect 27207 5414 27209 5466
rect 26963 5412 26969 5414
rect 27025 5412 27049 5414
rect 27105 5412 27129 5414
rect 27185 5412 27209 5414
rect 27265 5412 27271 5414
rect 26963 5403 27271 5412
rect 26700 5160 26752 5166
rect 26752 5120 26832 5148
rect 26700 5102 26752 5108
rect 26568 4564 26648 4570
rect 26516 4558 26648 4564
rect 26528 4542 26648 4558
rect 26804 4554 26832 5120
rect 27160 4752 27212 4758
rect 27158 4720 27160 4729
rect 27212 4720 27214 4729
rect 27158 4655 27214 4664
rect 26792 4548 26844 4554
rect 26528 4146 26556 4542
rect 26792 4490 26844 4496
rect 26608 4480 26660 4486
rect 26608 4422 26660 4428
rect 26700 4480 26752 4486
rect 26700 4422 26752 4428
rect 26424 4140 26476 4146
rect 26424 4082 26476 4088
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26516 3936 26568 3942
rect 26516 3878 26568 3884
rect 26332 3052 26384 3058
rect 26332 2994 26384 3000
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26528 2938 26556 3878
rect 26620 3058 26648 4422
rect 26712 3618 26740 4422
rect 26804 4078 26832 4490
rect 26884 4480 26936 4486
rect 26884 4422 26936 4428
rect 26896 4282 26924 4422
rect 26963 4380 27271 4389
rect 26963 4378 26969 4380
rect 27025 4378 27049 4380
rect 27105 4378 27129 4380
rect 27185 4378 27209 4380
rect 27265 4378 27271 4380
rect 27025 4326 27027 4378
rect 27207 4326 27209 4378
rect 26963 4324 26969 4326
rect 27025 4324 27049 4326
rect 27105 4324 27129 4326
rect 27185 4324 27209 4326
rect 27265 4324 27271 4326
rect 26963 4315 27271 4324
rect 26884 4276 26936 4282
rect 26884 4218 26936 4224
rect 27252 4140 27304 4146
rect 27252 4082 27304 4088
rect 26792 4072 26844 4078
rect 26792 4014 26844 4020
rect 26884 3664 26936 3670
rect 26712 3590 26832 3618
rect 26884 3606 26936 3612
rect 26608 3052 26660 3058
rect 26608 2994 26660 3000
rect 26056 2848 26108 2854
rect 26056 2790 26108 2796
rect 25688 2644 25740 2650
rect 25688 2586 25740 2592
rect 25780 2644 25832 2650
rect 25780 2586 25832 2592
rect 25964 2304 26016 2310
rect 25964 2246 26016 2252
rect 25596 1352 25648 1358
rect 25596 1294 25648 1300
rect 25976 1193 26004 2246
rect 26068 2145 26096 2790
rect 26330 2544 26386 2553
rect 26436 2514 26464 2926
rect 26528 2910 26740 2938
rect 26330 2479 26386 2488
rect 26424 2508 26476 2514
rect 26054 2136 26110 2145
rect 26054 2071 26110 2080
rect 26068 1902 26096 2071
rect 26056 1896 26108 1902
rect 26056 1838 26108 1844
rect 26344 1494 26372 2479
rect 26424 2450 26476 2456
rect 26436 2310 26464 2450
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 26436 1970 26464 2246
rect 26424 1964 26476 1970
rect 26424 1906 26476 1912
rect 26608 1760 26660 1766
rect 26608 1702 26660 1708
rect 26332 1488 26384 1494
rect 26332 1430 26384 1436
rect 26422 1456 26478 1465
rect 26620 1442 26648 1702
rect 26478 1426 26648 1442
rect 26478 1420 26660 1426
rect 26478 1414 26608 1420
rect 26422 1391 26478 1400
rect 26424 1216 26476 1222
rect 25962 1184 26018 1193
rect 26424 1158 26476 1164
rect 25962 1119 26018 1128
rect 26436 1018 26464 1158
rect 26424 1012 26476 1018
rect 26424 954 26476 960
rect 25228 876 25280 882
rect 25228 818 25280 824
rect 26528 814 26556 1414
rect 26608 1362 26660 1368
rect 26606 1320 26662 1329
rect 26606 1255 26662 1264
rect 26620 1018 26648 1255
rect 26608 1012 26660 1018
rect 26608 954 26660 960
rect 26712 950 26740 2910
rect 26804 1986 26832 3590
rect 26896 2854 26924 3606
rect 27264 3505 27292 4082
rect 27250 3496 27306 3505
rect 27250 3431 27306 3440
rect 26963 3292 27271 3301
rect 26963 3290 26969 3292
rect 27025 3290 27049 3292
rect 27105 3290 27129 3292
rect 27185 3290 27209 3292
rect 27265 3290 27271 3292
rect 27025 3238 27027 3290
rect 27207 3238 27209 3290
rect 26963 3236 26969 3238
rect 27025 3236 27049 3238
rect 27105 3236 27129 3238
rect 27185 3236 27209 3238
rect 27265 3236 27271 3238
rect 26963 3227 27271 3236
rect 26884 2848 26936 2854
rect 26884 2790 26936 2796
rect 27356 2650 27384 6666
rect 27448 6322 27476 7686
rect 27528 7540 27580 7546
rect 27528 7482 27580 7488
rect 27436 6316 27488 6322
rect 27436 6258 27488 6264
rect 27540 5234 27568 7482
rect 27620 6928 27672 6934
rect 27620 6870 27672 6876
rect 27528 5228 27580 5234
rect 27528 5170 27580 5176
rect 27632 3618 27660 6870
rect 27724 6866 27752 7822
rect 27816 6934 27844 8026
rect 28092 7954 28120 8230
rect 28080 7948 28132 7954
rect 28080 7890 28132 7896
rect 28184 7886 28212 9862
rect 28276 9722 28304 9998
rect 28264 9716 28316 9722
rect 28264 9658 28316 9664
rect 28264 8832 28316 8838
rect 28264 8774 28316 8780
rect 28172 7880 28224 7886
rect 28172 7822 28224 7828
rect 27894 7304 27950 7313
rect 27894 7239 27950 7248
rect 27804 6928 27856 6934
rect 27804 6870 27856 6876
rect 27712 6860 27764 6866
rect 27712 6802 27764 6808
rect 27908 6254 27936 7239
rect 28276 6798 28304 8774
rect 28368 8090 28396 14350
rect 28552 13977 28580 15438
rect 28644 15162 28672 20878
rect 29104 20330 29132 21422
rect 29288 20482 29316 21422
rect 29288 20454 29408 20482
rect 29380 20398 29408 20454
rect 29276 20392 29328 20398
rect 29276 20334 29328 20340
rect 29368 20392 29420 20398
rect 29368 20334 29420 20340
rect 29092 20324 29144 20330
rect 29092 20266 29144 20272
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 28828 19242 28856 19790
rect 28906 19408 28962 19417
rect 28906 19343 28962 19352
rect 28816 19236 28868 19242
rect 28816 19178 28868 19184
rect 28828 18970 28856 19178
rect 28816 18964 28868 18970
rect 28816 18906 28868 18912
rect 28920 18850 28948 19343
rect 29012 19145 29040 19790
rect 28998 19136 29054 19145
rect 28998 19071 29054 19080
rect 29104 18970 29132 20266
rect 29288 20058 29316 20334
rect 29276 20052 29328 20058
rect 29276 19994 29328 20000
rect 29380 19334 29408 20334
rect 29184 19304 29236 19310
rect 29288 19306 29408 19334
rect 29288 19292 29316 19306
rect 29236 19264 29316 19292
rect 29184 19246 29236 19252
rect 29092 18964 29144 18970
rect 29092 18906 29144 18912
rect 28998 18864 29054 18873
rect 28920 18822 28998 18850
rect 28998 18799 29054 18808
rect 29182 18864 29238 18873
rect 29182 18799 29238 18808
rect 28816 18760 28868 18766
rect 28816 18702 28868 18708
rect 29000 18760 29052 18766
rect 29000 18702 29052 18708
rect 29092 18760 29144 18766
rect 29092 18702 29144 18708
rect 28724 18352 28776 18358
rect 28724 18294 28776 18300
rect 28736 17882 28764 18294
rect 28828 18272 28856 18702
rect 28828 18244 28859 18272
rect 28831 18136 28859 18244
rect 28828 18108 28859 18136
rect 28908 18148 28960 18154
rect 28724 17876 28776 17882
rect 28724 17818 28776 17824
rect 28724 17332 28776 17338
rect 28724 17274 28776 17280
rect 28736 16046 28764 17274
rect 28724 16040 28776 16046
rect 28724 15982 28776 15988
rect 28724 15496 28776 15502
rect 28724 15438 28776 15444
rect 28632 15156 28684 15162
rect 28632 15098 28684 15104
rect 28630 14920 28686 14929
rect 28630 14855 28686 14864
rect 28538 13968 28594 13977
rect 28538 13903 28594 13912
rect 28538 13832 28594 13841
rect 28538 13767 28594 13776
rect 28448 12436 28500 12442
rect 28552 12434 28580 13767
rect 28644 13326 28672 14855
rect 28632 13320 28684 13326
rect 28632 13262 28684 13268
rect 28552 12406 28672 12434
rect 28448 12378 28500 12384
rect 28460 11830 28488 12378
rect 28448 11824 28500 11830
rect 28448 11766 28500 11772
rect 28540 11620 28592 11626
rect 28540 11562 28592 11568
rect 28448 11144 28500 11150
rect 28448 11086 28500 11092
rect 28356 8084 28408 8090
rect 28356 8026 28408 8032
rect 28460 7954 28488 11086
rect 28552 8634 28580 11562
rect 28644 9042 28672 12406
rect 28736 11762 28764 15438
rect 28828 11898 28856 18108
rect 28908 18090 28960 18096
rect 28920 17785 28948 18090
rect 28906 17776 28962 17785
rect 28906 17711 28962 17720
rect 28920 16250 28948 17711
rect 29012 17678 29040 18702
rect 29000 17672 29052 17678
rect 29000 17614 29052 17620
rect 28998 17096 29054 17105
rect 28998 17031 29054 17040
rect 28908 16244 28960 16250
rect 28908 16186 28960 16192
rect 29012 16182 29040 17031
rect 29000 16176 29052 16182
rect 29000 16118 29052 16124
rect 28908 16040 28960 16046
rect 28908 15982 28960 15988
rect 29000 16040 29052 16046
rect 29000 15982 29052 15988
rect 28920 14890 28948 15982
rect 29012 15706 29040 15982
rect 29000 15700 29052 15706
rect 29000 15642 29052 15648
rect 28908 14884 28960 14890
rect 28908 14826 28960 14832
rect 28920 13870 28948 14826
rect 29000 14816 29052 14822
rect 29000 14758 29052 14764
rect 28908 13864 28960 13870
rect 28908 13806 28960 13812
rect 28908 13184 28960 13190
rect 28908 13126 28960 13132
rect 28920 12306 28948 13126
rect 29012 12714 29040 14758
rect 29104 14074 29132 18702
rect 29196 14618 29224 18799
rect 29288 17882 29316 19264
rect 29368 19168 29420 19174
rect 29368 19110 29420 19116
rect 29380 18970 29408 19110
rect 29368 18964 29420 18970
rect 29368 18906 29420 18912
rect 29380 18834 29408 18906
rect 29368 18828 29420 18834
rect 29368 18770 29420 18776
rect 29276 17876 29328 17882
rect 29276 17818 29328 17824
rect 29276 17672 29328 17678
rect 29276 17614 29328 17620
rect 29288 17134 29316 17614
rect 29276 17128 29328 17134
rect 29472 17082 29500 21626
rect 29828 21548 29880 21554
rect 29828 21490 29880 21496
rect 31116 21548 31168 21554
rect 31116 21490 31168 21496
rect 29736 20868 29788 20874
rect 29736 20810 29788 20816
rect 29552 19848 29604 19854
rect 29552 19790 29604 19796
rect 29642 19816 29698 19825
rect 29276 17070 29328 17076
rect 29288 16590 29316 17070
rect 29380 17054 29500 17082
rect 29276 16584 29328 16590
rect 29276 16526 29328 16532
rect 29380 16454 29408 17054
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29368 16448 29420 16454
rect 29368 16390 29420 16396
rect 29472 16289 29500 16934
rect 29564 16697 29592 19790
rect 29642 19751 29698 19760
rect 29656 19310 29684 19751
rect 29644 19304 29696 19310
rect 29644 19246 29696 19252
rect 29642 19000 29698 19009
rect 29748 18986 29776 20810
rect 29840 20398 29868 21490
rect 30104 21344 30156 21350
rect 30104 21286 30156 21292
rect 29828 20392 29880 20398
rect 29828 20334 29880 20340
rect 29840 19378 29868 20334
rect 30116 20330 30144 21286
rect 30758 21244 31066 21253
rect 30758 21242 30764 21244
rect 30820 21242 30844 21244
rect 30900 21242 30924 21244
rect 30980 21242 31004 21244
rect 31060 21242 31066 21244
rect 30820 21190 30822 21242
rect 31002 21190 31004 21242
rect 30758 21188 30764 21190
rect 30820 21188 30844 21190
rect 30900 21188 30924 21190
rect 30980 21188 31004 21190
rect 31060 21188 31066 21190
rect 30758 21179 31066 21188
rect 30472 20936 30524 20942
rect 30472 20878 30524 20884
rect 30196 20392 30248 20398
rect 30196 20334 30248 20340
rect 30104 20324 30156 20330
rect 30104 20266 30156 20272
rect 29920 20256 29972 20262
rect 29920 20198 29972 20204
rect 29828 19372 29880 19378
rect 29828 19314 29880 19320
rect 29698 18958 29776 18986
rect 29642 18935 29698 18944
rect 29748 18358 29776 18958
rect 29736 18352 29788 18358
rect 29736 18294 29788 18300
rect 29736 18216 29788 18222
rect 29840 18204 29868 19314
rect 29788 18176 29868 18204
rect 29736 18158 29788 18164
rect 29840 18086 29868 18176
rect 29828 18080 29880 18086
rect 29828 18022 29880 18028
rect 29644 17876 29696 17882
rect 29644 17818 29696 17824
rect 29656 17134 29684 17818
rect 29828 17332 29880 17338
rect 29828 17274 29880 17280
rect 29644 17128 29696 17134
rect 29644 17070 29696 17076
rect 29656 16946 29684 17070
rect 29656 16918 29776 16946
rect 29642 16824 29698 16833
rect 29642 16759 29698 16768
rect 29550 16688 29606 16697
rect 29550 16623 29606 16632
rect 29656 16590 29684 16759
rect 29552 16584 29604 16590
rect 29552 16526 29604 16532
rect 29644 16584 29696 16590
rect 29644 16526 29696 16532
rect 29458 16280 29514 16289
rect 29458 16215 29514 16224
rect 29564 16182 29592 16526
rect 29552 16176 29604 16182
rect 29366 16144 29422 16153
rect 29276 16108 29328 16114
rect 29328 16088 29366 16096
rect 29552 16118 29604 16124
rect 29328 16079 29422 16088
rect 29328 16068 29408 16079
rect 29276 16050 29328 16056
rect 29276 15904 29328 15910
rect 29552 15904 29604 15910
rect 29276 15846 29328 15852
rect 29380 15864 29552 15892
rect 29184 14612 29236 14618
rect 29184 14554 29236 14560
rect 29092 14068 29144 14074
rect 29092 14010 29144 14016
rect 29184 14000 29236 14006
rect 29184 13942 29236 13948
rect 29092 13864 29144 13870
rect 29092 13806 29144 13812
rect 29000 12708 29052 12714
rect 29000 12650 29052 12656
rect 28908 12300 28960 12306
rect 28908 12242 28960 12248
rect 28908 12096 28960 12102
rect 28908 12038 28960 12044
rect 28816 11892 28868 11898
rect 28816 11834 28868 11840
rect 28814 11792 28870 11801
rect 28724 11756 28776 11762
rect 28814 11727 28870 11736
rect 28724 11698 28776 11704
rect 28632 9036 28684 9042
rect 28632 8978 28684 8984
rect 28540 8628 28592 8634
rect 28540 8570 28592 8576
rect 28632 8560 28684 8566
rect 28632 8502 28684 8508
rect 28448 7948 28500 7954
rect 28448 7890 28500 7896
rect 28644 7206 28672 8502
rect 28828 8362 28856 11727
rect 28920 10130 28948 12038
rect 29000 11620 29052 11626
rect 29000 11562 29052 11568
rect 29012 11354 29040 11562
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 29000 10464 29052 10470
rect 29000 10406 29052 10412
rect 28908 10124 28960 10130
rect 28908 10066 28960 10072
rect 29012 9602 29040 10406
rect 28920 9586 29040 9602
rect 29104 9586 29132 13806
rect 29196 12714 29224 13942
rect 29288 13870 29316 15846
rect 29276 13864 29328 13870
rect 29276 13806 29328 13812
rect 29276 13524 29328 13530
rect 29276 13466 29328 13472
rect 29184 12708 29236 12714
rect 29184 12650 29236 12656
rect 29184 10668 29236 10674
rect 29184 10610 29236 10616
rect 29196 10033 29224 10610
rect 29182 10024 29238 10033
rect 29182 9959 29238 9968
rect 28908 9580 29040 9586
rect 28960 9574 29040 9580
rect 29092 9580 29144 9586
rect 28908 9522 28960 9528
rect 29092 9522 29144 9528
rect 28920 8838 28948 9522
rect 29000 9376 29052 9382
rect 29000 9318 29052 9324
rect 29012 9178 29040 9318
rect 29000 9172 29052 9178
rect 29000 9114 29052 9120
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 28816 8356 28868 8362
rect 28816 8298 28868 8304
rect 28816 7744 28868 7750
rect 28816 7686 28868 7692
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 28632 7200 28684 7206
rect 28632 7142 28684 7148
rect 28264 6792 28316 6798
rect 28264 6734 28316 6740
rect 27896 6248 27948 6254
rect 27896 6190 27948 6196
rect 28078 5672 28134 5681
rect 28078 5607 28134 5616
rect 28356 5636 28408 5642
rect 27804 5228 27856 5234
rect 27804 5170 27856 5176
rect 27816 4690 27844 5170
rect 27804 4684 27856 4690
rect 27804 4626 27856 4632
rect 27896 4684 27948 4690
rect 27896 4626 27948 4632
rect 27908 4554 27936 4626
rect 27896 4548 27948 4554
rect 27896 4490 27948 4496
rect 27710 4176 27766 4185
rect 27710 4111 27766 4120
rect 27540 3590 27660 3618
rect 27344 2644 27396 2650
rect 27344 2586 27396 2592
rect 27540 2514 27568 3590
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27528 2508 27580 2514
rect 27448 2468 27528 2496
rect 26963 2204 27271 2213
rect 26963 2202 26969 2204
rect 27025 2202 27049 2204
rect 27105 2202 27129 2204
rect 27185 2202 27209 2204
rect 27265 2202 27271 2204
rect 27025 2150 27027 2202
rect 27207 2150 27209 2202
rect 26963 2148 26969 2150
rect 27025 2148 27049 2150
rect 27105 2148 27129 2150
rect 27185 2148 27209 2150
rect 27265 2148 27271 2150
rect 26963 2139 27271 2148
rect 26804 1970 26924 1986
rect 27448 1970 27476 2468
rect 27528 2450 27580 2456
rect 27526 2000 27582 2009
rect 26804 1964 26936 1970
rect 26804 1958 26884 1964
rect 26884 1906 26936 1912
rect 27436 1964 27488 1970
rect 27526 1935 27582 1944
rect 27436 1906 27488 1912
rect 27448 1426 27476 1906
rect 27540 1562 27568 1935
rect 27528 1556 27580 1562
rect 27528 1498 27580 1504
rect 27436 1420 27488 1426
rect 27356 1380 27436 1408
rect 26963 1116 27271 1125
rect 26963 1114 26969 1116
rect 27025 1114 27049 1116
rect 27105 1114 27129 1116
rect 27185 1114 27209 1116
rect 27265 1114 27271 1116
rect 27025 1062 27027 1114
rect 27207 1062 27209 1114
rect 26963 1060 26969 1062
rect 27025 1060 27049 1062
rect 27105 1060 27129 1062
rect 27185 1060 27209 1062
rect 27265 1060 27271 1062
rect 26963 1051 27271 1060
rect 26700 944 26752 950
rect 26700 886 26752 892
rect 27356 882 27384 1380
rect 27436 1362 27488 1368
rect 27632 1306 27660 3470
rect 27724 3058 27752 4111
rect 27802 3632 27858 3641
rect 27908 3602 27936 4490
rect 28092 3942 28120 5607
rect 28356 5578 28408 5584
rect 28264 5568 28316 5574
rect 28264 5510 28316 5516
rect 28172 4616 28224 4622
rect 28172 4558 28224 4564
rect 28080 3936 28132 3942
rect 28080 3878 28132 3884
rect 27802 3567 27858 3576
rect 27896 3596 27948 3602
rect 27712 3052 27764 3058
rect 27712 2994 27764 3000
rect 27712 2644 27764 2650
rect 27712 2586 27764 2592
rect 27724 1834 27752 2586
rect 27816 2106 27844 3567
rect 27896 3538 27948 3544
rect 27908 2514 27936 3538
rect 28184 3534 28212 4558
rect 28172 3528 28224 3534
rect 28000 3488 28172 3516
rect 28000 2650 28028 3488
rect 28172 3470 28224 3476
rect 28172 2984 28224 2990
rect 28172 2926 28224 2932
rect 28080 2848 28132 2854
rect 28080 2790 28132 2796
rect 27988 2644 28040 2650
rect 27988 2586 28040 2592
rect 27896 2508 27948 2514
rect 27896 2450 27948 2456
rect 27804 2100 27856 2106
rect 27804 2042 27856 2048
rect 27712 1828 27764 1834
rect 27712 1770 27764 1776
rect 27724 1426 27752 1770
rect 27712 1420 27764 1426
rect 27712 1362 27764 1368
rect 28092 1358 28120 2790
rect 28184 2446 28212 2926
rect 28172 2440 28224 2446
rect 28172 2382 28224 2388
rect 28184 1562 28212 2382
rect 28276 1970 28304 5510
rect 28264 1964 28316 1970
rect 28264 1906 28316 1912
rect 28172 1556 28224 1562
rect 28172 1498 28224 1504
rect 28368 1358 28396 5578
rect 28448 5568 28500 5574
rect 28448 5510 28500 5516
rect 28460 4826 28488 5510
rect 28448 4820 28500 4826
rect 28448 4762 28500 4768
rect 28552 4690 28580 7142
rect 28540 4684 28592 4690
rect 28540 4626 28592 4632
rect 28448 3528 28500 3534
rect 28448 3470 28500 3476
rect 28540 3528 28592 3534
rect 28540 3470 28592 3476
rect 28460 2961 28488 3470
rect 28552 3194 28580 3470
rect 28540 3188 28592 3194
rect 28540 3130 28592 3136
rect 28446 2952 28502 2961
rect 28446 2887 28502 2896
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 27804 1352 27856 1358
rect 27632 1300 27804 1306
rect 27632 1294 27856 1300
rect 28080 1352 28132 1358
rect 28080 1294 28132 1300
rect 28356 1352 28408 1358
rect 28356 1294 28408 1300
rect 27632 1278 27844 1294
rect 27344 876 27396 882
rect 27344 818 27396 824
rect 26516 808 26568 814
rect 26516 750 26568 756
rect 27816 678 27844 1278
rect 28552 1018 28580 2382
rect 28644 1766 28672 7142
rect 28828 3602 28856 7686
rect 28908 6656 28960 6662
rect 28960 6604 29040 6610
rect 28908 6598 29040 6604
rect 28920 6582 29040 6598
rect 29012 5114 29040 6582
rect 29104 5778 29132 9522
rect 29182 9344 29238 9353
rect 29182 9279 29238 9288
rect 29196 8634 29224 9279
rect 29288 9178 29316 13466
rect 29380 12481 29408 15864
rect 29552 15846 29604 15852
rect 29642 15872 29698 15881
rect 29642 15807 29698 15816
rect 29656 15706 29684 15807
rect 29644 15700 29696 15706
rect 29644 15642 29696 15648
rect 29748 15638 29776 16918
rect 29840 16674 29868 17274
rect 29932 16794 29960 20198
rect 30012 19712 30064 19718
rect 30012 19654 30064 19660
rect 30024 18578 30052 19654
rect 30208 18970 30236 20334
rect 30288 19712 30340 19718
rect 30288 19654 30340 19660
rect 30300 19446 30328 19654
rect 30288 19440 30340 19446
rect 30288 19382 30340 19388
rect 30196 18964 30248 18970
rect 30196 18906 30248 18912
rect 30286 18728 30342 18737
rect 30286 18663 30342 18672
rect 30024 18550 30236 18578
rect 30104 18420 30156 18426
rect 30104 18362 30156 18368
rect 30012 18080 30064 18086
rect 30012 18022 30064 18028
rect 30024 17134 30052 18022
rect 30012 17128 30064 17134
rect 30012 17070 30064 17076
rect 30012 16992 30064 16998
rect 30012 16934 30064 16940
rect 29920 16788 29972 16794
rect 29920 16730 29972 16736
rect 29840 16646 29960 16674
rect 29826 16416 29882 16425
rect 29826 16351 29882 16360
rect 29736 15632 29788 15638
rect 29550 15600 29606 15609
rect 29736 15574 29788 15580
rect 29550 15535 29606 15544
rect 29458 15328 29514 15337
rect 29458 15263 29514 15272
rect 29472 14958 29500 15263
rect 29460 14952 29512 14958
rect 29460 14894 29512 14900
rect 29460 14544 29512 14550
rect 29460 14486 29512 14492
rect 29472 13954 29500 14486
rect 29564 14074 29592 15535
rect 29644 15156 29696 15162
rect 29644 15098 29696 15104
rect 29552 14068 29604 14074
rect 29552 14010 29604 14016
rect 29472 13938 29592 13954
rect 29656 13938 29684 15098
rect 29472 13932 29604 13938
rect 29472 13926 29552 13932
rect 29552 13874 29604 13880
rect 29644 13932 29696 13938
rect 29644 13874 29696 13880
rect 29460 12640 29512 12646
rect 29460 12582 29512 12588
rect 29366 12472 29422 12481
rect 29366 12407 29422 12416
rect 29472 10606 29500 12582
rect 29564 12434 29592 13874
rect 29644 13796 29696 13802
rect 29644 13738 29696 13744
rect 29656 12714 29684 13738
rect 29748 13530 29776 15574
rect 29840 14074 29868 16351
rect 29932 15586 29960 16646
rect 30024 16182 30052 16934
rect 30012 16176 30064 16182
rect 30012 16118 30064 16124
rect 30024 16017 30052 16118
rect 30010 16008 30066 16017
rect 30010 15943 30066 15952
rect 30012 15904 30064 15910
rect 30012 15846 30064 15852
rect 30024 15745 30052 15846
rect 30010 15736 30066 15745
rect 30010 15671 30066 15680
rect 29932 15570 30052 15586
rect 29932 15564 30064 15570
rect 29932 15558 30012 15564
rect 30012 15506 30064 15512
rect 29920 15088 29972 15094
rect 29920 15030 29972 15036
rect 29932 14618 29960 15030
rect 29920 14612 29972 14618
rect 29920 14554 29972 14560
rect 29920 14408 29972 14414
rect 29920 14350 29972 14356
rect 29828 14068 29880 14074
rect 29828 14010 29880 14016
rect 29828 13728 29880 13734
rect 29828 13670 29880 13676
rect 29736 13524 29788 13530
rect 29736 13466 29788 13472
rect 29840 13326 29868 13670
rect 29828 13320 29880 13326
rect 29828 13262 29880 13268
rect 29644 12708 29696 12714
rect 29644 12650 29696 12656
rect 29736 12640 29788 12646
rect 29736 12582 29788 12588
rect 29564 12406 29684 12434
rect 29552 11824 29604 11830
rect 29552 11766 29604 11772
rect 29564 11540 29592 11766
rect 29656 11694 29684 12406
rect 29748 12306 29776 12582
rect 29736 12300 29788 12306
rect 29736 12242 29788 12248
rect 29644 11688 29696 11694
rect 29644 11630 29696 11636
rect 29644 11552 29696 11558
rect 29564 11512 29644 11540
rect 29644 11494 29696 11500
rect 29552 11348 29604 11354
rect 29552 11290 29604 11296
rect 29564 10606 29592 11290
rect 29748 10674 29776 12242
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 29460 10600 29512 10606
rect 29460 10542 29512 10548
rect 29552 10600 29604 10606
rect 29552 10542 29604 10548
rect 29368 10464 29420 10470
rect 29368 10406 29420 10412
rect 29380 9382 29408 10406
rect 29460 9716 29512 9722
rect 29460 9658 29512 9664
rect 29564 9674 29592 10542
rect 29368 9376 29420 9382
rect 29368 9318 29420 9324
rect 29276 9172 29328 9178
rect 29276 9114 29328 9120
rect 29380 8974 29408 9318
rect 29368 8968 29420 8974
rect 29274 8936 29330 8945
rect 29330 8916 29368 8922
rect 29330 8910 29420 8916
rect 29330 8894 29408 8910
rect 29274 8871 29330 8880
rect 29368 8832 29420 8838
rect 29368 8774 29420 8780
rect 29184 8628 29236 8634
rect 29184 8570 29236 8576
rect 29196 8378 29224 8570
rect 29196 8350 29316 8378
rect 29184 8288 29236 8294
rect 29184 8230 29236 8236
rect 29092 5772 29144 5778
rect 29092 5714 29144 5720
rect 29104 5234 29132 5714
rect 29092 5228 29144 5234
rect 29092 5170 29144 5176
rect 29012 5086 29132 5114
rect 29000 5024 29052 5030
rect 29000 4966 29052 4972
rect 28816 3596 28868 3602
rect 28816 3538 28868 3544
rect 28722 3088 28778 3097
rect 28722 3023 28778 3032
rect 28736 1834 28764 3023
rect 28814 1864 28870 1873
rect 28724 1828 28776 1834
rect 28814 1799 28870 1808
rect 28724 1770 28776 1776
rect 28828 1766 28856 1799
rect 28632 1760 28684 1766
rect 28632 1702 28684 1708
rect 28816 1760 28868 1766
rect 28816 1702 28868 1708
rect 28540 1012 28592 1018
rect 28540 954 28592 960
rect 28644 814 28672 1702
rect 29012 1562 29040 4966
rect 29104 4010 29132 5086
rect 29196 4078 29224 8230
rect 29288 7342 29316 8350
rect 29380 8022 29408 8774
rect 29368 8016 29420 8022
rect 29368 7958 29420 7964
rect 29276 7336 29328 7342
rect 29276 7278 29328 7284
rect 29288 5914 29316 7278
rect 29276 5908 29328 5914
rect 29276 5850 29328 5856
rect 29276 5568 29328 5574
rect 29276 5510 29328 5516
rect 29184 4072 29236 4078
rect 29184 4014 29236 4020
rect 29092 4004 29144 4010
rect 29092 3946 29144 3952
rect 29196 3738 29224 4014
rect 29184 3732 29236 3738
rect 29184 3674 29236 3680
rect 29092 3528 29144 3534
rect 29092 3470 29144 3476
rect 29104 1766 29132 3470
rect 29092 1760 29144 1766
rect 29092 1702 29144 1708
rect 29000 1556 29052 1562
rect 29000 1498 29052 1504
rect 29288 882 29316 5510
rect 29380 5370 29408 7958
rect 29472 7342 29500 9658
rect 29564 9646 29684 9674
rect 29552 8968 29604 8974
rect 29552 8910 29604 8916
rect 29564 7954 29592 8910
rect 29552 7948 29604 7954
rect 29552 7890 29604 7896
rect 29460 7336 29512 7342
rect 29460 7278 29512 7284
rect 29472 5914 29500 7278
rect 29550 6896 29606 6905
rect 29550 6831 29606 6840
rect 29564 6730 29592 6831
rect 29552 6724 29604 6730
rect 29552 6666 29604 6672
rect 29656 6610 29684 9646
rect 29840 9489 29868 13262
rect 29932 12986 29960 14350
rect 30024 13297 30052 15506
rect 30010 13288 30066 13297
rect 30010 13223 30066 13232
rect 29920 12980 29972 12986
rect 29920 12922 29972 12928
rect 29918 12064 29974 12073
rect 29918 11999 29974 12008
rect 29932 11257 29960 11999
rect 29918 11248 29974 11257
rect 29918 11183 29974 11192
rect 29826 9480 29882 9489
rect 29826 9415 29882 9424
rect 29840 9110 29868 9415
rect 29828 9104 29880 9110
rect 29828 9046 29880 9052
rect 29932 8922 29960 11183
rect 30012 11076 30064 11082
rect 30012 11018 30064 11024
rect 30024 9042 30052 11018
rect 30116 11014 30144 18362
rect 30208 11218 30236 18550
rect 30300 18426 30328 18663
rect 30288 18420 30340 18426
rect 30288 18362 30340 18368
rect 30300 14958 30328 18362
rect 30380 18352 30432 18358
rect 30380 18294 30432 18300
rect 30392 18057 30420 18294
rect 30378 18048 30434 18057
rect 30378 17983 30434 17992
rect 30378 17640 30434 17649
rect 30378 17575 30380 17584
rect 30432 17575 30434 17584
rect 30380 17546 30432 17552
rect 30378 17096 30434 17105
rect 30378 17031 30434 17040
rect 30392 16794 30420 17031
rect 30380 16788 30432 16794
rect 30380 16730 30432 16736
rect 30380 15972 30432 15978
rect 30380 15914 30432 15920
rect 30392 15162 30420 15914
rect 30380 15156 30432 15162
rect 30380 15098 30432 15104
rect 30378 15056 30434 15065
rect 30378 14991 30434 15000
rect 30288 14952 30340 14958
rect 30288 14894 30340 14900
rect 30288 14816 30340 14822
rect 30288 14758 30340 14764
rect 30300 13802 30328 14758
rect 30392 13870 30420 14991
rect 30380 13864 30432 13870
rect 30380 13806 30432 13812
rect 30288 13796 30340 13802
rect 30288 13738 30340 13744
rect 30378 13696 30434 13705
rect 30378 13631 30434 13640
rect 30288 13184 30340 13190
rect 30288 13126 30340 13132
rect 30300 12850 30328 13126
rect 30392 12986 30420 13631
rect 30380 12980 30432 12986
rect 30380 12922 30432 12928
rect 30288 12844 30340 12850
rect 30288 12786 30340 12792
rect 30380 12776 30432 12782
rect 30380 12718 30432 12724
rect 30392 11694 30420 12718
rect 30380 11688 30432 11694
rect 30380 11630 30432 11636
rect 30288 11552 30340 11558
rect 30288 11494 30340 11500
rect 30196 11212 30248 11218
rect 30196 11154 30248 11160
rect 30104 11008 30156 11014
rect 30104 10950 30156 10956
rect 30300 10554 30328 11494
rect 30392 11354 30420 11630
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 30116 10526 30328 10554
rect 30116 10470 30144 10526
rect 30104 10464 30156 10470
rect 30104 10406 30156 10412
rect 30288 10464 30340 10470
rect 30288 10406 30340 10412
rect 30116 9382 30144 10406
rect 30300 10198 30328 10406
rect 30288 10192 30340 10198
rect 30288 10134 30340 10140
rect 30300 9722 30328 10134
rect 30380 9920 30432 9926
rect 30380 9862 30432 9868
rect 30288 9716 30340 9722
rect 30288 9658 30340 9664
rect 30104 9376 30156 9382
rect 30104 9318 30156 9324
rect 30288 9376 30340 9382
rect 30288 9318 30340 9324
rect 30012 9036 30064 9042
rect 30012 8978 30064 8984
rect 29932 8894 30052 8922
rect 30024 8838 30052 8894
rect 30012 8832 30064 8838
rect 30012 8774 30064 8780
rect 29826 8528 29882 8537
rect 29826 8463 29882 8472
rect 29736 7200 29788 7206
rect 29736 7142 29788 7148
rect 29564 6582 29684 6610
rect 29460 5908 29512 5914
rect 29460 5850 29512 5856
rect 29368 5364 29420 5370
rect 29368 5306 29420 5312
rect 29366 5264 29422 5273
rect 29366 5199 29422 5208
rect 29380 2106 29408 5199
rect 29458 5128 29514 5137
rect 29458 5063 29514 5072
rect 29472 5030 29500 5063
rect 29460 5024 29512 5030
rect 29460 4966 29512 4972
rect 29458 4040 29514 4049
rect 29458 3975 29514 3984
rect 29472 3942 29500 3975
rect 29460 3936 29512 3942
rect 29460 3878 29512 3884
rect 29472 2106 29500 3878
rect 29564 3398 29592 6582
rect 29644 6112 29696 6118
rect 29644 6054 29696 6060
rect 29656 4826 29684 6054
rect 29644 4820 29696 4826
rect 29644 4762 29696 4768
rect 29552 3392 29604 3398
rect 29552 3334 29604 3340
rect 29748 2514 29776 7142
rect 29840 3738 29868 8463
rect 29920 7948 29972 7954
rect 29920 7890 29972 7896
rect 29828 3732 29880 3738
rect 29828 3674 29880 3680
rect 29932 3058 29960 7890
rect 30012 6996 30064 7002
rect 30012 6938 30064 6944
rect 29920 3052 29972 3058
rect 29920 2994 29972 3000
rect 29920 2916 29972 2922
rect 29920 2858 29972 2864
rect 29736 2508 29788 2514
rect 29736 2450 29788 2456
rect 29368 2100 29420 2106
rect 29368 2042 29420 2048
rect 29460 2100 29512 2106
rect 29460 2042 29512 2048
rect 29472 1426 29500 2042
rect 29460 1420 29512 1426
rect 29460 1362 29512 1368
rect 29472 1018 29500 1362
rect 29932 1358 29960 2858
rect 30024 2650 30052 6938
rect 30116 3602 30144 9318
rect 30196 9104 30248 9110
rect 30196 9046 30248 9052
rect 30208 8430 30236 9046
rect 30196 8424 30248 8430
rect 30196 8366 30248 8372
rect 30194 7848 30250 7857
rect 30194 7783 30250 7792
rect 30104 3596 30156 3602
rect 30104 3538 30156 3544
rect 30208 3194 30236 7783
rect 30300 6866 30328 9318
rect 30392 8498 30420 9862
rect 30484 9178 30512 20878
rect 30656 20324 30708 20330
rect 30656 20266 30708 20272
rect 30564 20052 30616 20058
rect 30564 19994 30616 20000
rect 30576 10810 30604 19994
rect 30668 17762 30696 20266
rect 30758 20156 31066 20165
rect 30758 20154 30764 20156
rect 30820 20154 30844 20156
rect 30900 20154 30924 20156
rect 30980 20154 31004 20156
rect 31060 20154 31066 20156
rect 30820 20102 30822 20154
rect 31002 20102 31004 20154
rect 30758 20100 30764 20102
rect 30820 20100 30844 20102
rect 30900 20100 30924 20102
rect 30980 20100 31004 20102
rect 31060 20100 31066 20102
rect 30758 20091 31066 20100
rect 30758 19068 31066 19077
rect 30758 19066 30764 19068
rect 30820 19066 30844 19068
rect 30900 19066 30924 19068
rect 30980 19066 31004 19068
rect 31060 19066 31066 19068
rect 30820 19014 30822 19066
rect 31002 19014 31004 19066
rect 30758 19012 30764 19014
rect 30820 19012 30844 19014
rect 30900 19012 30924 19014
rect 30980 19012 31004 19014
rect 31060 19012 31066 19014
rect 30758 19003 31066 19012
rect 30758 17980 31066 17989
rect 30758 17978 30764 17980
rect 30820 17978 30844 17980
rect 30900 17978 30924 17980
rect 30980 17978 31004 17980
rect 31060 17978 31066 17980
rect 30820 17926 30822 17978
rect 31002 17926 31004 17978
rect 30758 17924 30764 17926
rect 30820 17924 30844 17926
rect 30900 17924 30924 17926
rect 30980 17924 31004 17926
rect 31060 17924 31066 17926
rect 30758 17915 31066 17924
rect 31128 17762 31156 21490
rect 30668 17734 30788 17762
rect 30656 17536 30708 17542
rect 30656 17478 30708 17484
rect 30564 10804 30616 10810
rect 30564 10746 30616 10752
rect 30668 9654 30696 17478
rect 30760 17105 30788 17734
rect 31036 17734 31156 17762
rect 30746 17096 30802 17105
rect 30746 17031 30802 17040
rect 31036 16998 31064 17734
rect 31116 17128 31168 17134
rect 31116 17070 31168 17076
rect 31024 16992 31076 16998
rect 31024 16934 31076 16940
rect 30758 16892 31066 16901
rect 30758 16890 30764 16892
rect 30820 16890 30844 16892
rect 30900 16890 30924 16892
rect 30980 16890 31004 16892
rect 31060 16890 31066 16892
rect 30820 16838 30822 16890
rect 31002 16838 31004 16890
rect 30758 16836 30764 16838
rect 30820 16836 30844 16838
rect 30900 16836 30924 16838
rect 30980 16836 31004 16838
rect 31060 16836 31066 16838
rect 30758 16827 31066 16836
rect 31024 16788 31076 16794
rect 31024 16730 31076 16736
rect 31036 15910 31064 16730
rect 31024 15904 31076 15910
rect 31024 15846 31076 15852
rect 30758 15804 31066 15813
rect 30758 15802 30764 15804
rect 30820 15802 30844 15804
rect 30900 15802 30924 15804
rect 30980 15802 31004 15804
rect 31060 15802 31066 15804
rect 30820 15750 30822 15802
rect 31002 15750 31004 15802
rect 30758 15748 30764 15750
rect 30820 15748 30844 15750
rect 30900 15748 30924 15750
rect 30980 15748 31004 15750
rect 31060 15748 31066 15750
rect 30758 15739 31066 15748
rect 31024 15700 31076 15706
rect 31024 15642 31076 15648
rect 30932 15632 30984 15638
rect 30746 15600 30802 15609
rect 30932 15574 30984 15580
rect 30746 15535 30802 15544
rect 30760 14958 30788 15535
rect 30748 14952 30800 14958
rect 30748 14894 30800 14900
rect 30944 14822 30972 15574
rect 31036 15042 31064 15642
rect 31128 15162 31156 17070
rect 31220 15706 31248 21966
rect 31300 18624 31352 18630
rect 31300 18566 31352 18572
rect 31208 15700 31260 15706
rect 31208 15642 31260 15648
rect 31208 15428 31260 15434
rect 31208 15370 31260 15376
rect 31116 15156 31168 15162
rect 31116 15098 31168 15104
rect 31036 15014 31156 15042
rect 30932 14816 30984 14822
rect 30932 14758 30984 14764
rect 30758 14716 31066 14725
rect 30758 14714 30764 14716
rect 30820 14714 30844 14716
rect 30900 14714 30924 14716
rect 30980 14714 31004 14716
rect 31060 14714 31066 14716
rect 30820 14662 30822 14714
rect 31002 14662 31004 14714
rect 30758 14660 30764 14662
rect 30820 14660 30844 14662
rect 30900 14660 30924 14662
rect 30980 14660 31004 14662
rect 31060 14660 31066 14662
rect 30758 14651 31066 14660
rect 30748 14612 30800 14618
rect 30748 14554 30800 14560
rect 30760 14006 30788 14554
rect 31128 14074 31156 15014
rect 31116 14068 31168 14074
rect 31116 14010 31168 14016
rect 30748 14000 30800 14006
rect 30748 13942 30800 13948
rect 30758 13628 31066 13637
rect 30758 13626 30764 13628
rect 30820 13626 30844 13628
rect 30900 13626 30924 13628
rect 30980 13626 31004 13628
rect 31060 13626 31066 13628
rect 30820 13574 30822 13626
rect 31002 13574 31004 13626
rect 30758 13572 30764 13574
rect 30820 13572 30844 13574
rect 30900 13572 30924 13574
rect 30980 13572 31004 13574
rect 31060 13572 31066 13574
rect 30758 13563 31066 13572
rect 30758 12540 31066 12549
rect 30758 12538 30764 12540
rect 30820 12538 30844 12540
rect 30900 12538 30924 12540
rect 30980 12538 31004 12540
rect 31060 12538 31066 12540
rect 30820 12486 30822 12538
rect 31002 12486 31004 12538
rect 30758 12484 30764 12486
rect 30820 12484 30844 12486
rect 30900 12484 30924 12486
rect 30980 12484 31004 12486
rect 31060 12484 31066 12486
rect 30758 12475 31066 12484
rect 30758 11452 31066 11461
rect 30758 11450 30764 11452
rect 30820 11450 30844 11452
rect 30900 11450 30924 11452
rect 30980 11450 31004 11452
rect 31060 11450 31066 11452
rect 30820 11398 30822 11450
rect 31002 11398 31004 11450
rect 30758 11396 30764 11398
rect 30820 11396 30844 11398
rect 30900 11396 30924 11398
rect 30980 11396 31004 11398
rect 31060 11396 31066 11398
rect 30758 11387 31066 11396
rect 30758 10364 31066 10373
rect 30758 10362 30764 10364
rect 30820 10362 30844 10364
rect 30900 10362 30924 10364
rect 30980 10362 31004 10364
rect 31060 10362 31066 10364
rect 30820 10310 30822 10362
rect 31002 10310 31004 10362
rect 30758 10308 30764 10310
rect 30820 10308 30844 10310
rect 30900 10308 30924 10310
rect 30980 10308 31004 10310
rect 31060 10308 31066 10310
rect 30758 10299 31066 10308
rect 30656 9648 30708 9654
rect 30656 9590 30708 9596
rect 30758 9276 31066 9285
rect 30758 9274 30764 9276
rect 30820 9274 30844 9276
rect 30900 9274 30924 9276
rect 30980 9274 31004 9276
rect 31060 9274 31066 9276
rect 30820 9222 30822 9274
rect 31002 9222 31004 9274
rect 30758 9220 30764 9222
rect 30820 9220 30844 9222
rect 30900 9220 30924 9222
rect 30980 9220 31004 9222
rect 31060 9220 31066 9222
rect 30758 9211 31066 9220
rect 30472 9172 30524 9178
rect 30472 9114 30524 9120
rect 30472 8832 30524 8838
rect 30472 8774 30524 8780
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 30380 7744 30432 7750
rect 30380 7686 30432 7692
rect 30288 6860 30340 6866
rect 30288 6802 30340 6808
rect 30392 4146 30420 7686
rect 30380 4140 30432 4146
rect 30380 4082 30432 4088
rect 30484 4026 30512 8774
rect 31220 8362 31248 15370
rect 31312 11694 31340 18566
rect 31390 18320 31446 18329
rect 31390 18255 31446 18264
rect 31404 13938 31432 18255
rect 31392 13932 31444 13938
rect 31392 13874 31444 13880
rect 31300 11688 31352 11694
rect 31300 11630 31352 11636
rect 31208 8356 31260 8362
rect 31208 8298 31260 8304
rect 30758 8188 31066 8197
rect 30758 8186 30764 8188
rect 30820 8186 30844 8188
rect 30900 8186 30924 8188
rect 30980 8186 31004 8188
rect 31060 8186 31066 8188
rect 30820 8134 30822 8186
rect 31002 8134 31004 8186
rect 30758 8132 30764 8134
rect 30820 8132 30844 8134
rect 30900 8132 30924 8134
rect 30980 8132 31004 8134
rect 31060 8132 31066 8134
rect 30758 8123 31066 8132
rect 30758 7100 31066 7109
rect 30758 7098 30764 7100
rect 30820 7098 30844 7100
rect 30900 7098 30924 7100
rect 30980 7098 31004 7100
rect 31060 7098 31066 7100
rect 30820 7046 30822 7098
rect 31002 7046 31004 7098
rect 30758 7044 30764 7046
rect 30820 7044 30844 7046
rect 30900 7044 30924 7046
rect 30980 7044 31004 7046
rect 31060 7044 31066 7046
rect 30758 7035 31066 7044
rect 30758 6012 31066 6021
rect 30758 6010 30764 6012
rect 30820 6010 30844 6012
rect 30900 6010 30924 6012
rect 30980 6010 31004 6012
rect 31060 6010 31066 6012
rect 30820 5958 30822 6010
rect 31002 5958 31004 6010
rect 30758 5956 30764 5958
rect 30820 5956 30844 5958
rect 30900 5956 30924 5958
rect 30980 5956 31004 5958
rect 31060 5956 31066 5958
rect 30758 5947 31066 5956
rect 30758 4924 31066 4933
rect 30758 4922 30764 4924
rect 30820 4922 30844 4924
rect 30900 4922 30924 4924
rect 30980 4922 31004 4924
rect 31060 4922 31066 4924
rect 30820 4870 30822 4922
rect 31002 4870 31004 4922
rect 30758 4868 30764 4870
rect 30820 4868 30844 4870
rect 30900 4868 30924 4870
rect 30980 4868 31004 4870
rect 31060 4868 31066 4870
rect 30758 4859 31066 4868
rect 30392 3998 30512 4026
rect 30196 3188 30248 3194
rect 30196 3130 30248 3136
rect 30392 2922 30420 3998
rect 30758 3836 31066 3845
rect 30758 3834 30764 3836
rect 30820 3834 30844 3836
rect 30900 3834 30924 3836
rect 30980 3834 31004 3836
rect 31060 3834 31066 3836
rect 30820 3782 30822 3834
rect 31002 3782 31004 3834
rect 30758 3780 30764 3782
rect 30820 3780 30844 3782
rect 30900 3780 30924 3782
rect 30980 3780 31004 3782
rect 31060 3780 31066 3782
rect 30758 3771 31066 3780
rect 30380 2916 30432 2922
rect 30380 2858 30432 2864
rect 30758 2748 31066 2757
rect 30758 2746 30764 2748
rect 30820 2746 30844 2748
rect 30900 2746 30924 2748
rect 30980 2746 31004 2748
rect 31060 2746 31066 2748
rect 30820 2694 30822 2746
rect 31002 2694 31004 2746
rect 30758 2692 30764 2694
rect 30820 2692 30844 2694
rect 30900 2692 30924 2694
rect 30980 2692 31004 2694
rect 31060 2692 31066 2694
rect 30758 2683 31066 2692
rect 30012 2644 30064 2650
rect 30012 2586 30064 2592
rect 30758 1660 31066 1669
rect 30758 1658 30764 1660
rect 30820 1658 30844 1660
rect 30900 1658 30924 1660
rect 30980 1658 31004 1660
rect 31060 1658 31066 1660
rect 30820 1606 30822 1658
rect 31002 1606 31004 1658
rect 30758 1604 30764 1606
rect 30820 1604 30844 1606
rect 30900 1604 30924 1606
rect 30980 1604 31004 1606
rect 31060 1604 31066 1606
rect 30758 1595 31066 1604
rect 29920 1352 29972 1358
rect 29920 1294 29972 1300
rect 29460 1012 29512 1018
rect 29460 954 29512 960
rect 29276 876 29328 882
rect 29276 818 29328 824
rect 28632 808 28684 814
rect 28632 750 28684 756
rect 29182 776 29238 785
rect 29182 711 29238 720
rect 29196 678 29224 711
rect 25688 672 25740 678
rect 25688 614 25740 620
rect 26056 672 26108 678
rect 26056 614 26108 620
rect 26240 672 26292 678
rect 26240 614 26292 620
rect 27804 672 27856 678
rect 27804 614 27856 620
rect 29184 672 29236 678
rect 29184 614 29236 620
rect 25700 406 25728 614
rect 26068 474 26096 614
rect 26056 468 26108 474
rect 26056 410 26108 416
rect 25688 400 25740 406
rect 24950 368 25006 377
rect 25688 342 25740 348
rect 24950 303 25006 312
rect 26252 202 26280 614
rect 30758 572 31066 581
rect 30758 570 30764 572
rect 30820 570 30844 572
rect 30900 570 30924 572
rect 30980 570 31004 572
rect 31060 570 31066 572
rect 30820 518 30822 570
rect 31002 518 31004 570
rect 30758 516 30764 518
rect 30820 516 30844 518
rect 30900 516 30924 518
rect 30980 516 31004 518
rect 31060 516 31066 518
rect 30758 507 31066 516
rect 26240 196 26292 202
rect 26240 138 26292 144
rect 24858 96 24914 105
rect 15566 31 15622 40
rect 16396 60 16448 66
rect 12440 2 12492 8
rect 24858 31 24914 40
rect 16396 2 16448 8
<< via2 >>
rect 846 18264 902 18320
rect 2502 21936 2558 21992
rect 1674 17992 1730 18048
rect 1674 17620 1676 17640
rect 1676 17620 1728 17640
rect 1728 17620 1730 17640
rect 1674 17584 1730 17620
rect 1766 14864 1822 14920
rect 1490 12416 1546 12472
rect 2042 16496 2098 16552
rect 2042 15544 2098 15600
rect 2134 15000 2190 15056
rect 2318 19080 2374 19136
rect 1950 14456 2006 14512
rect 2778 17584 2834 17640
rect 2502 15408 2558 15464
rect 1858 13912 1914 13968
rect 2226 13268 2228 13288
rect 2228 13268 2280 13288
rect 2280 13268 2282 13288
rect 2226 13232 2282 13268
rect 1950 11192 2006 11248
rect 1398 6704 1454 6760
rect 1582 6976 1638 7032
rect 938 3848 994 3904
rect 1582 5752 1638 5808
rect 1306 3984 1362 4040
rect 1674 5616 1730 5672
rect 938 1672 994 1728
rect 2318 9968 2374 10024
rect 2226 7792 2282 7848
rect 2134 6316 2190 6352
rect 2134 6296 2136 6316
rect 2136 6296 2188 6316
rect 2188 6296 2190 6316
rect 2042 5072 2098 5128
rect 2134 4120 2190 4176
rect 1766 1808 1822 1864
rect 2778 16768 2834 16824
rect 3514 20984 3570 21040
rect 4199 21786 4255 21788
rect 4279 21786 4335 21788
rect 4359 21786 4415 21788
rect 4439 21786 4495 21788
rect 4199 21734 4245 21786
rect 4245 21734 4255 21786
rect 4279 21734 4309 21786
rect 4309 21734 4321 21786
rect 4321 21734 4335 21786
rect 4359 21734 4373 21786
rect 4373 21734 4385 21786
rect 4385 21734 4415 21786
rect 4439 21734 4449 21786
rect 4449 21734 4495 21786
rect 4199 21732 4255 21734
rect 4279 21732 4335 21734
rect 4359 21732 4415 21734
rect 4439 21732 4495 21734
rect 4066 21120 4122 21176
rect 4618 20712 4674 20768
rect 4199 20698 4255 20700
rect 4279 20698 4335 20700
rect 4359 20698 4415 20700
rect 4439 20698 4495 20700
rect 4199 20646 4245 20698
rect 4245 20646 4255 20698
rect 4279 20646 4309 20698
rect 4309 20646 4321 20698
rect 4321 20646 4335 20698
rect 4359 20646 4373 20698
rect 4373 20646 4385 20698
rect 4385 20646 4415 20698
rect 4439 20646 4449 20698
rect 4449 20646 4495 20698
rect 4199 20644 4255 20646
rect 4279 20644 4335 20646
rect 4359 20644 4415 20646
rect 4439 20644 4495 20646
rect 4526 20440 4582 20496
rect 3422 19896 3478 19952
rect 3054 16088 3110 16144
rect 3054 15816 3110 15872
rect 2962 10648 3018 10704
rect 3606 19760 3662 19816
rect 3698 17720 3754 17776
rect 4199 19610 4255 19612
rect 4279 19610 4335 19612
rect 4359 19610 4415 19612
rect 4439 19610 4495 19612
rect 4199 19558 4245 19610
rect 4245 19558 4255 19610
rect 4279 19558 4309 19610
rect 4309 19558 4321 19610
rect 4321 19558 4335 19610
rect 4359 19558 4373 19610
rect 4373 19558 4385 19610
rect 4385 19558 4415 19610
rect 4439 19558 4449 19610
rect 4449 19558 4495 19610
rect 4199 19556 4255 19558
rect 4279 19556 4335 19558
rect 4359 19556 4415 19558
rect 4439 19556 4495 19558
rect 4066 18808 4122 18864
rect 4199 18522 4255 18524
rect 4279 18522 4335 18524
rect 4359 18522 4415 18524
rect 4439 18522 4495 18524
rect 4199 18470 4245 18522
rect 4245 18470 4255 18522
rect 4279 18470 4309 18522
rect 4309 18470 4321 18522
rect 4321 18470 4335 18522
rect 4359 18470 4373 18522
rect 4373 18470 4385 18522
rect 4385 18470 4415 18522
rect 4439 18470 4449 18522
rect 4449 18470 4495 18522
rect 4199 18468 4255 18470
rect 4279 18468 4335 18470
rect 4359 18468 4415 18470
rect 4439 18468 4495 18470
rect 3974 18128 4030 18184
rect 4894 20340 4896 20360
rect 4896 20340 4948 20360
rect 4948 20340 4950 20360
rect 4894 20304 4950 20340
rect 5078 20576 5134 20632
rect 3790 17176 3846 17232
rect 4199 17434 4255 17436
rect 4279 17434 4335 17436
rect 4359 17434 4415 17436
rect 4439 17434 4495 17436
rect 4199 17382 4245 17434
rect 4245 17382 4255 17434
rect 4279 17382 4309 17434
rect 4309 17382 4321 17434
rect 4321 17382 4335 17434
rect 4359 17382 4373 17434
rect 4373 17382 4385 17434
rect 4385 17382 4415 17434
rect 4439 17382 4449 17434
rect 4449 17382 4495 17434
rect 4199 17380 4255 17382
rect 4279 17380 4335 17382
rect 4359 17380 4415 17382
rect 4439 17380 4495 17382
rect 4199 16346 4255 16348
rect 4279 16346 4335 16348
rect 4359 16346 4415 16348
rect 4439 16346 4495 16348
rect 4199 16294 4245 16346
rect 4245 16294 4255 16346
rect 4279 16294 4309 16346
rect 4309 16294 4321 16346
rect 4321 16294 4335 16346
rect 4359 16294 4373 16346
rect 4373 16294 4385 16346
rect 4385 16294 4415 16346
rect 4439 16294 4449 16346
rect 4449 16294 4495 16346
rect 4199 16292 4255 16294
rect 4279 16292 4335 16294
rect 4359 16292 4415 16294
rect 4439 16292 4495 16294
rect 4199 15258 4255 15260
rect 4279 15258 4335 15260
rect 4359 15258 4415 15260
rect 4439 15258 4495 15260
rect 4199 15206 4245 15258
rect 4245 15206 4255 15258
rect 4279 15206 4309 15258
rect 4309 15206 4321 15258
rect 4321 15206 4335 15258
rect 4359 15206 4373 15258
rect 4373 15206 4385 15258
rect 4385 15206 4415 15258
rect 4439 15206 4449 15258
rect 4449 15206 4495 15258
rect 4199 15204 4255 15206
rect 4279 15204 4335 15206
rect 4359 15204 4415 15206
rect 4439 15204 4495 15206
rect 3422 12860 3424 12880
rect 3424 12860 3476 12880
rect 3476 12860 3478 12880
rect 3422 12824 3478 12860
rect 3422 12724 3424 12744
rect 3424 12724 3476 12744
rect 3476 12724 3478 12744
rect 3422 12688 3478 12724
rect 3698 13912 3754 13968
rect 3514 11756 3570 11792
rect 3514 11736 3516 11756
rect 3516 11736 3568 11756
rect 3568 11736 3570 11756
rect 4986 18944 5042 19000
rect 6550 21800 6606 21856
rect 5814 21664 5870 21720
rect 5814 20848 5870 20904
rect 6458 20884 6460 20904
rect 6460 20884 6512 20904
rect 6512 20884 6514 20904
rect 6458 20848 6514 20884
rect 6642 20848 6698 20904
rect 5354 18672 5410 18728
rect 5630 19624 5686 19680
rect 5814 19488 5870 19544
rect 5814 19080 5870 19136
rect 5354 17992 5410 18048
rect 4894 16088 4950 16144
rect 4199 14170 4255 14172
rect 4279 14170 4335 14172
rect 4359 14170 4415 14172
rect 4439 14170 4495 14172
rect 4199 14118 4245 14170
rect 4245 14118 4255 14170
rect 4279 14118 4309 14170
rect 4309 14118 4321 14170
rect 4321 14118 4335 14170
rect 4359 14118 4373 14170
rect 4373 14118 4385 14170
rect 4385 14118 4415 14170
rect 4439 14118 4449 14170
rect 4449 14118 4495 14170
rect 4199 14116 4255 14118
rect 4279 14116 4335 14118
rect 4359 14116 4415 14118
rect 4439 14116 4495 14118
rect 4158 13504 4214 13560
rect 4199 13082 4255 13084
rect 4279 13082 4335 13084
rect 4359 13082 4415 13084
rect 4439 13082 4495 13084
rect 4199 13030 4245 13082
rect 4245 13030 4255 13082
rect 4279 13030 4309 13082
rect 4309 13030 4321 13082
rect 4321 13030 4335 13082
rect 4359 13030 4373 13082
rect 4373 13030 4385 13082
rect 4385 13030 4415 13082
rect 4439 13030 4449 13082
rect 4449 13030 4495 13082
rect 4199 13028 4255 13030
rect 4279 13028 4335 13030
rect 4359 13028 4415 13030
rect 4439 13028 4495 13030
rect 5262 14320 5318 14376
rect 4199 11994 4255 11996
rect 4279 11994 4335 11996
rect 4359 11994 4415 11996
rect 4439 11994 4495 11996
rect 4199 11942 4245 11994
rect 4245 11942 4255 11994
rect 4279 11942 4309 11994
rect 4309 11942 4321 11994
rect 4321 11942 4335 11994
rect 4359 11942 4373 11994
rect 4373 11942 4385 11994
rect 4385 11942 4415 11994
rect 4439 11942 4449 11994
rect 4449 11942 4495 11994
rect 4199 11940 4255 11942
rect 4279 11940 4335 11942
rect 4359 11940 4415 11942
rect 4439 11940 4495 11942
rect 5814 17740 5870 17776
rect 5814 17720 5816 17740
rect 5816 17720 5868 17740
rect 5868 17720 5870 17740
rect 5722 17448 5778 17504
rect 5446 16088 5502 16144
rect 5446 15272 5502 15328
rect 5722 15156 5778 15192
rect 5722 15136 5724 15156
rect 5724 15136 5776 15156
rect 5776 15136 5778 15156
rect 5906 14048 5962 14104
rect 5170 12144 5226 12200
rect 4199 10906 4255 10908
rect 4279 10906 4335 10908
rect 4359 10906 4415 10908
rect 4439 10906 4495 10908
rect 4199 10854 4245 10906
rect 4245 10854 4255 10906
rect 4279 10854 4309 10906
rect 4309 10854 4321 10906
rect 4321 10854 4335 10906
rect 4359 10854 4373 10906
rect 4373 10854 4385 10906
rect 4385 10854 4415 10906
rect 4439 10854 4449 10906
rect 4449 10854 4495 10906
rect 4199 10852 4255 10854
rect 4279 10852 4335 10854
rect 4359 10852 4415 10854
rect 4439 10852 4495 10854
rect 4199 9818 4255 9820
rect 4279 9818 4335 9820
rect 4359 9818 4415 9820
rect 4439 9818 4495 9820
rect 4199 9766 4245 9818
rect 4245 9766 4255 9818
rect 4279 9766 4309 9818
rect 4309 9766 4321 9818
rect 4321 9766 4335 9818
rect 4359 9766 4373 9818
rect 4373 9766 4385 9818
rect 4385 9766 4415 9818
rect 4439 9766 4449 9818
rect 4449 9766 4495 9818
rect 4199 9764 4255 9766
rect 4279 9764 4335 9766
rect 4359 9764 4415 9766
rect 4439 9764 4495 9766
rect 5078 10804 5134 10840
rect 5078 10784 5080 10804
rect 5080 10784 5132 10804
rect 5132 10784 5134 10804
rect 5354 10512 5410 10568
rect 3330 8916 3332 8936
rect 3332 8916 3384 8936
rect 3384 8916 3386 8936
rect 3330 8880 3386 8916
rect 4199 8730 4255 8732
rect 4279 8730 4335 8732
rect 4359 8730 4415 8732
rect 4439 8730 4495 8732
rect 4199 8678 4245 8730
rect 4245 8678 4255 8730
rect 4279 8678 4309 8730
rect 4309 8678 4321 8730
rect 4321 8678 4335 8730
rect 4359 8678 4373 8730
rect 4373 8678 4385 8730
rect 4385 8678 4415 8730
rect 4439 8678 4449 8730
rect 4449 8678 4495 8730
rect 4199 8676 4255 8678
rect 4279 8676 4335 8678
rect 4359 8676 4415 8678
rect 4439 8676 4495 8678
rect 2410 8200 2466 8256
rect 2686 8064 2742 8120
rect 2870 7248 2926 7304
rect 2778 6840 2834 6896
rect 2502 5888 2558 5944
rect 2778 5208 2834 5264
rect 3146 6976 3202 7032
rect 2778 3984 2834 4040
rect 2962 4020 2964 4040
rect 2964 4020 3016 4040
rect 3016 4020 3018 4040
rect 2962 3984 3018 4020
rect 2778 3712 2834 3768
rect 3054 3712 3110 3768
rect 3054 2916 3110 2952
rect 3054 2896 3056 2916
rect 3056 2896 3108 2916
rect 3108 2896 3110 2916
rect 3882 6840 3938 6896
rect 3422 4564 3424 4584
rect 3424 4564 3476 4584
rect 3476 4564 3478 4584
rect 3422 4528 3478 4564
rect 3514 2760 3570 2816
rect 3514 2644 3570 2680
rect 3514 2624 3516 2644
rect 3516 2624 3568 2644
rect 3568 2624 3570 2644
rect 4199 7642 4255 7644
rect 4279 7642 4335 7644
rect 4359 7642 4415 7644
rect 4439 7642 4495 7644
rect 4199 7590 4245 7642
rect 4245 7590 4255 7642
rect 4279 7590 4309 7642
rect 4309 7590 4321 7642
rect 4321 7590 4335 7642
rect 4359 7590 4373 7642
rect 4373 7590 4385 7642
rect 4385 7590 4415 7642
rect 4439 7590 4449 7642
rect 4449 7590 4495 7642
rect 4199 7588 4255 7590
rect 4279 7588 4335 7590
rect 4359 7588 4415 7590
rect 4439 7588 4495 7590
rect 4434 7148 4436 7168
rect 4436 7148 4488 7168
rect 4488 7148 4490 7168
rect 4434 7112 4490 7148
rect 4199 6554 4255 6556
rect 4279 6554 4335 6556
rect 4359 6554 4415 6556
rect 4439 6554 4495 6556
rect 4199 6502 4245 6554
rect 4245 6502 4255 6554
rect 4279 6502 4309 6554
rect 4309 6502 4321 6554
rect 4321 6502 4335 6554
rect 4359 6502 4373 6554
rect 4373 6502 4385 6554
rect 4385 6502 4415 6554
rect 4439 6502 4449 6554
rect 4449 6502 4495 6554
rect 4199 6500 4255 6502
rect 4279 6500 4335 6502
rect 4359 6500 4415 6502
rect 4439 6500 4495 6502
rect 3698 3984 3754 4040
rect 4199 5466 4255 5468
rect 4279 5466 4335 5468
rect 4359 5466 4415 5468
rect 4439 5466 4495 5468
rect 4199 5414 4245 5466
rect 4245 5414 4255 5466
rect 4279 5414 4309 5466
rect 4309 5414 4321 5466
rect 4321 5414 4335 5466
rect 4359 5414 4373 5466
rect 4373 5414 4385 5466
rect 4385 5414 4415 5466
rect 4439 5414 4449 5466
rect 4449 5414 4495 5466
rect 4199 5412 4255 5414
rect 4279 5412 4335 5414
rect 4359 5412 4415 5414
rect 4439 5412 4495 5414
rect 4618 6976 4674 7032
rect 4199 4378 4255 4380
rect 4279 4378 4335 4380
rect 4359 4378 4415 4380
rect 4439 4378 4495 4380
rect 4199 4326 4245 4378
rect 4245 4326 4255 4378
rect 4279 4326 4309 4378
rect 4309 4326 4321 4378
rect 4321 4326 4335 4378
rect 4359 4326 4373 4378
rect 4373 4326 4385 4378
rect 4385 4326 4415 4378
rect 4439 4326 4449 4378
rect 4449 4326 4495 4378
rect 4199 4324 4255 4326
rect 4279 4324 4335 4326
rect 4359 4324 4415 4326
rect 4439 4324 4495 4326
rect 4618 3848 4674 3904
rect 3790 2388 3792 2408
rect 3792 2388 3844 2408
rect 3844 2388 3846 2408
rect 3790 2352 3846 2388
rect 4526 3440 4582 3496
rect 4199 3290 4255 3292
rect 4279 3290 4335 3292
rect 4359 3290 4415 3292
rect 4439 3290 4495 3292
rect 4199 3238 4245 3290
rect 4245 3238 4255 3290
rect 4279 3238 4309 3290
rect 4309 3238 4321 3290
rect 4321 3238 4335 3290
rect 4359 3238 4373 3290
rect 4373 3238 4385 3290
rect 4385 3238 4415 3290
rect 4439 3238 4449 3290
rect 4449 3238 4495 3290
rect 4199 3236 4255 3238
rect 4279 3236 4335 3238
rect 4359 3236 4415 3238
rect 4439 3236 4495 3238
rect 4158 3032 4214 3088
rect 3974 2624 4030 2680
rect 4250 2508 4306 2544
rect 4250 2488 4252 2508
rect 4252 2488 4304 2508
rect 4304 2488 4306 2508
rect 4199 2202 4255 2204
rect 4279 2202 4335 2204
rect 4359 2202 4415 2204
rect 4439 2202 4495 2204
rect 4199 2150 4245 2202
rect 4245 2150 4255 2202
rect 4279 2150 4309 2202
rect 4309 2150 4321 2202
rect 4321 2150 4335 2202
rect 4359 2150 4373 2202
rect 4373 2150 4385 2202
rect 4385 2150 4415 2202
rect 4439 2150 4449 2202
rect 4449 2150 4495 2202
rect 4199 2148 4255 2150
rect 4279 2148 4335 2150
rect 4359 2148 4415 2150
rect 4439 2148 4495 2150
rect 4342 1964 4398 2000
rect 4342 1944 4344 1964
rect 4344 1944 4396 1964
rect 4396 1944 4398 1964
rect 3606 1400 3662 1456
rect 4434 1672 4490 1728
rect 4250 1400 4306 1456
rect 4434 1400 4490 1456
rect 4250 1300 4252 1320
rect 4252 1300 4304 1320
rect 4304 1300 4306 1320
rect 4250 1264 4306 1300
rect 4199 1114 4255 1116
rect 4279 1114 4335 1116
rect 4359 1114 4415 1116
rect 4439 1114 4495 1116
rect 4199 1062 4245 1114
rect 4245 1062 4255 1114
rect 4279 1062 4309 1114
rect 4309 1062 4321 1114
rect 4321 1062 4335 1114
rect 4359 1062 4373 1114
rect 4373 1062 4385 1114
rect 4385 1062 4415 1114
rect 4439 1062 4449 1114
rect 4449 1062 4495 1114
rect 4199 1060 4255 1062
rect 4279 1060 4335 1062
rect 4359 1060 4415 1062
rect 4439 1060 4495 1062
rect 4066 856 4122 912
rect 4618 720 4674 776
rect 5170 6704 5226 6760
rect 4986 4392 5042 4448
rect 4986 3848 5042 3904
rect 5078 2760 5134 2816
rect 5722 11464 5778 11520
rect 6090 20304 6146 20360
rect 6182 14728 6238 14784
rect 6458 18400 6514 18456
rect 6090 12960 6146 13016
rect 6458 17992 6514 18048
rect 9126 22208 9182 22264
rect 14370 22228 14426 22264
rect 22282 22244 22284 22264
rect 22284 22244 22336 22264
rect 22336 22244 22338 22264
rect 14370 22208 14372 22228
rect 14372 22208 14424 22228
rect 14424 22208 14426 22228
rect 9034 22072 9090 22128
rect 8666 21664 8722 21720
rect 7010 21392 7066 21448
rect 7102 21120 7158 21176
rect 7194 19760 7250 19816
rect 6918 18944 6974 19000
rect 6734 18400 6790 18456
rect 6826 17312 6882 17368
rect 6826 17040 6882 17096
rect 6550 16652 6606 16688
rect 6550 16632 6552 16652
rect 6552 16632 6604 16652
rect 6604 16632 6606 16652
rect 6826 15272 6882 15328
rect 7102 17076 7104 17096
rect 7104 17076 7156 17096
rect 7156 17076 7158 17096
rect 7102 17040 7158 17076
rect 7010 15952 7066 16008
rect 7102 15816 7158 15872
rect 8390 21256 8446 21312
rect 7994 21242 8050 21244
rect 8074 21242 8130 21244
rect 8154 21242 8210 21244
rect 8234 21242 8290 21244
rect 7994 21190 8040 21242
rect 8040 21190 8050 21242
rect 8074 21190 8104 21242
rect 8104 21190 8116 21242
rect 8116 21190 8130 21242
rect 8154 21190 8168 21242
rect 8168 21190 8180 21242
rect 8180 21190 8210 21242
rect 8234 21190 8244 21242
rect 8244 21190 8290 21242
rect 7994 21188 8050 21190
rect 8074 21188 8130 21190
rect 8154 21188 8210 21190
rect 8234 21188 8290 21190
rect 8482 21120 8538 21176
rect 7378 17720 7434 17776
rect 7010 15272 7066 15328
rect 6642 14048 6698 14104
rect 6642 13504 6698 13560
rect 6550 13368 6606 13424
rect 7378 15136 7434 15192
rect 7194 14728 7250 14784
rect 6366 12688 6422 12744
rect 5814 9016 5870 9072
rect 6366 9560 6422 9616
rect 7654 18944 7710 19000
rect 8482 20712 8538 20768
rect 8850 21256 8906 21312
rect 9494 21800 9550 21856
rect 9218 21256 9274 21312
rect 7994 20154 8050 20156
rect 8074 20154 8130 20156
rect 8154 20154 8210 20156
rect 8234 20154 8290 20156
rect 7994 20102 8040 20154
rect 8040 20102 8050 20154
rect 8074 20102 8104 20154
rect 8104 20102 8116 20154
rect 8116 20102 8130 20154
rect 8154 20102 8168 20154
rect 8168 20102 8180 20154
rect 8180 20102 8210 20154
rect 8234 20102 8244 20154
rect 8244 20102 8290 20154
rect 7994 20100 8050 20102
rect 8074 20100 8130 20102
rect 8154 20100 8210 20102
rect 8234 20100 8290 20102
rect 8206 19760 8262 19816
rect 7994 19066 8050 19068
rect 8074 19066 8130 19068
rect 8154 19066 8210 19068
rect 8234 19066 8290 19068
rect 7994 19014 8040 19066
rect 8040 19014 8050 19066
rect 8074 19014 8104 19066
rect 8104 19014 8116 19066
rect 8116 19014 8130 19066
rect 8154 19014 8168 19066
rect 8168 19014 8180 19066
rect 8180 19014 8210 19066
rect 8234 19014 8244 19066
rect 8244 19014 8290 19066
rect 7994 19012 8050 19014
rect 8074 19012 8130 19014
rect 8154 19012 8210 19014
rect 8234 19012 8290 19014
rect 8666 19352 8722 19408
rect 9402 20304 9458 20360
rect 8942 19352 8998 19408
rect 8942 19216 8998 19272
rect 8666 18808 8722 18864
rect 8850 18808 8906 18864
rect 7654 18400 7710 18456
rect 7746 17992 7802 18048
rect 7562 15136 7618 15192
rect 7562 15000 7618 15056
rect 7654 13640 7710 13696
rect 7994 17978 8050 17980
rect 8074 17978 8130 17980
rect 8154 17978 8210 17980
rect 8234 17978 8290 17980
rect 7994 17926 8040 17978
rect 8040 17926 8050 17978
rect 8074 17926 8104 17978
rect 8104 17926 8116 17978
rect 8116 17926 8130 17978
rect 8154 17926 8168 17978
rect 8168 17926 8180 17978
rect 8180 17926 8210 17978
rect 8234 17926 8244 17978
rect 8244 17926 8290 17978
rect 7994 17924 8050 17926
rect 8074 17924 8130 17926
rect 8154 17924 8210 17926
rect 8234 17924 8290 17926
rect 8206 17720 8262 17776
rect 8574 17856 8630 17912
rect 8758 18400 8814 18456
rect 8942 18536 8998 18592
rect 9586 19624 9642 19680
rect 9678 18944 9734 19000
rect 9310 18808 9366 18864
rect 9402 18400 9458 18456
rect 9402 17856 9458 17912
rect 7994 16890 8050 16892
rect 8074 16890 8130 16892
rect 8154 16890 8210 16892
rect 8234 16890 8290 16892
rect 7994 16838 8040 16890
rect 8040 16838 8050 16890
rect 8074 16838 8104 16890
rect 8104 16838 8116 16890
rect 8116 16838 8130 16890
rect 8154 16838 8168 16890
rect 8168 16838 8180 16890
rect 8180 16838 8210 16890
rect 8234 16838 8244 16890
rect 8244 16838 8290 16890
rect 7994 16836 8050 16838
rect 8074 16836 8130 16838
rect 8154 16836 8210 16838
rect 8234 16836 8290 16838
rect 8666 16904 8722 16960
rect 8574 16768 8630 16824
rect 8482 16632 8538 16688
rect 8298 15952 8354 16008
rect 7994 15802 8050 15804
rect 8074 15802 8130 15804
rect 8154 15802 8210 15804
rect 8234 15802 8290 15804
rect 7994 15750 8040 15802
rect 8040 15750 8050 15802
rect 8074 15750 8104 15802
rect 8104 15750 8116 15802
rect 8116 15750 8130 15802
rect 8154 15750 8168 15802
rect 8168 15750 8180 15802
rect 8180 15750 8210 15802
rect 8234 15750 8244 15802
rect 8244 15750 8290 15802
rect 7994 15748 8050 15750
rect 8074 15748 8130 15750
rect 8154 15748 8210 15750
rect 8234 15748 8290 15750
rect 7930 15000 7986 15056
rect 7994 14714 8050 14716
rect 8074 14714 8130 14716
rect 8154 14714 8210 14716
rect 8234 14714 8290 14716
rect 7994 14662 8040 14714
rect 8040 14662 8050 14714
rect 8074 14662 8104 14714
rect 8104 14662 8116 14714
rect 8116 14662 8130 14714
rect 8154 14662 8168 14714
rect 8168 14662 8180 14714
rect 8180 14662 8210 14714
rect 8234 14662 8244 14714
rect 8244 14662 8290 14714
rect 7994 14660 8050 14662
rect 8074 14660 8130 14662
rect 8154 14660 8210 14662
rect 8234 14660 8290 14662
rect 7994 13626 8050 13628
rect 8074 13626 8130 13628
rect 8154 13626 8210 13628
rect 8234 13626 8290 13628
rect 7994 13574 8040 13626
rect 8040 13574 8050 13626
rect 8074 13574 8104 13626
rect 8104 13574 8116 13626
rect 8116 13574 8130 13626
rect 8154 13574 8168 13626
rect 8168 13574 8180 13626
rect 8180 13574 8210 13626
rect 8234 13574 8244 13626
rect 8244 13574 8290 13626
rect 7994 13572 8050 13574
rect 8074 13572 8130 13574
rect 8154 13572 8210 13574
rect 8234 13572 8290 13574
rect 9034 16360 9090 16416
rect 8666 14728 8722 14784
rect 8390 12960 8446 13016
rect 7994 12538 8050 12540
rect 8074 12538 8130 12540
rect 8154 12538 8210 12540
rect 8234 12538 8290 12540
rect 7994 12486 8040 12538
rect 8040 12486 8050 12538
rect 8074 12486 8104 12538
rect 8104 12486 8116 12538
rect 8116 12486 8130 12538
rect 8154 12486 8168 12538
rect 8168 12486 8180 12538
rect 8180 12486 8210 12538
rect 8234 12486 8244 12538
rect 8244 12486 8290 12538
rect 7994 12484 8050 12486
rect 8074 12484 8130 12486
rect 8154 12484 8210 12486
rect 8234 12484 8290 12486
rect 7838 11464 7894 11520
rect 7994 11450 8050 11452
rect 8074 11450 8130 11452
rect 8154 11450 8210 11452
rect 8234 11450 8290 11452
rect 7994 11398 8040 11450
rect 8040 11398 8050 11450
rect 8074 11398 8104 11450
rect 8104 11398 8116 11450
rect 8116 11398 8130 11450
rect 8154 11398 8168 11450
rect 8168 11398 8180 11450
rect 8180 11398 8210 11450
rect 8234 11398 8244 11450
rect 8244 11398 8290 11450
rect 7994 11396 8050 11398
rect 8074 11396 8130 11398
rect 8154 11396 8210 11398
rect 8234 11396 8290 11398
rect 6090 9152 6146 9208
rect 5630 7112 5686 7168
rect 5814 6840 5870 6896
rect 6366 7792 6422 7848
rect 6366 6840 6422 6896
rect 5630 5480 5686 5536
rect 5814 6024 5870 6080
rect 5906 4664 5962 4720
rect 5630 4020 5632 4040
rect 5632 4020 5684 4040
rect 5684 4020 5686 4040
rect 5630 3984 5686 4020
rect 5630 3576 5686 3632
rect 5446 3304 5502 3360
rect 5538 2644 5594 2680
rect 5538 2624 5540 2644
rect 5540 2624 5592 2644
rect 5592 2624 5594 2644
rect 5078 1672 5134 1728
rect 6090 6432 6146 6488
rect 6182 4392 6238 4448
rect 5170 1128 5226 1184
rect 5446 992 5502 1048
rect 3974 40 4030 96
rect 5814 1672 5870 1728
rect 6090 2216 6146 2272
rect 5906 1556 5962 1592
rect 5906 1536 5908 1556
rect 5908 1536 5960 1556
rect 5960 1536 5962 1556
rect 6274 1808 6330 1864
rect 6734 7404 6790 7440
rect 6734 7384 6736 7404
rect 6736 7384 6788 7404
rect 6788 7384 6790 7404
rect 7194 9036 7250 9072
rect 7194 9016 7196 9036
rect 7196 9016 7248 9036
rect 7248 9016 7250 9036
rect 7286 6432 7342 6488
rect 7470 10104 7526 10160
rect 7470 9152 7526 9208
rect 7994 10362 8050 10364
rect 8074 10362 8130 10364
rect 8154 10362 8210 10364
rect 8234 10362 8290 10364
rect 7994 10310 8040 10362
rect 8040 10310 8050 10362
rect 8074 10310 8104 10362
rect 8104 10310 8116 10362
rect 8116 10310 8130 10362
rect 8154 10310 8168 10362
rect 8168 10310 8180 10362
rect 8180 10310 8210 10362
rect 8234 10310 8244 10362
rect 8244 10310 8290 10362
rect 7994 10308 8050 10310
rect 8074 10308 8130 10310
rect 8154 10308 8210 10310
rect 8234 10308 8290 10310
rect 8666 13912 8722 13968
rect 8850 13776 8906 13832
rect 8482 10920 8538 10976
rect 8390 9560 8446 9616
rect 9494 16632 9550 16688
rect 9126 15272 9182 15328
rect 9126 14320 9182 14376
rect 9678 16088 9734 16144
rect 9586 15272 9642 15328
rect 9862 20032 9918 20088
rect 9402 13812 9404 13832
rect 9404 13812 9456 13832
rect 9456 13812 9458 13832
rect 9402 13776 9458 13812
rect 9586 13404 9588 13424
rect 9588 13404 9640 13424
rect 9640 13404 9642 13424
rect 9586 13368 9642 13404
rect 10966 21936 11022 21992
rect 11426 21936 11482 21992
rect 10506 20712 10562 20768
rect 10506 20440 10562 20496
rect 10414 20032 10470 20088
rect 10506 19896 10562 19952
rect 10230 18808 10286 18864
rect 10138 17584 10194 17640
rect 10046 14728 10102 14784
rect 10138 13368 10194 13424
rect 10138 12960 10194 13016
rect 9678 12280 9734 12336
rect 9678 12008 9734 12064
rect 9954 11328 10010 11384
rect 8666 10376 8722 10432
rect 7994 9274 8050 9276
rect 8074 9274 8130 9276
rect 8154 9274 8210 9276
rect 8234 9274 8290 9276
rect 7994 9222 8040 9274
rect 8040 9222 8050 9274
rect 8074 9222 8104 9274
rect 8104 9222 8116 9274
rect 8116 9222 8130 9274
rect 8154 9222 8168 9274
rect 8168 9222 8180 9274
rect 8180 9222 8210 9274
rect 8234 9222 8244 9274
rect 8244 9222 8290 9274
rect 7994 9220 8050 9222
rect 8074 9220 8130 9222
rect 8154 9220 8210 9222
rect 8234 9220 8290 9222
rect 7470 8472 7526 8528
rect 7010 5888 7066 5944
rect 6734 5480 6790 5536
rect 6918 2760 6974 2816
rect 6642 2624 6698 2680
rect 8482 8916 8484 8936
rect 8484 8916 8536 8936
rect 8536 8916 8538 8936
rect 8482 8880 8538 8916
rect 9862 10920 9918 10976
rect 9586 10784 9642 10840
rect 9218 8472 9274 8528
rect 7654 8084 7710 8120
rect 7654 8064 7656 8084
rect 7656 8064 7708 8084
rect 7708 8064 7710 8084
rect 7994 8186 8050 8188
rect 8074 8186 8130 8188
rect 8154 8186 8210 8188
rect 8234 8186 8290 8188
rect 7994 8134 8040 8186
rect 8040 8134 8050 8186
rect 8074 8134 8104 8186
rect 8104 8134 8116 8186
rect 8116 8134 8130 8186
rect 8154 8134 8168 8186
rect 8168 8134 8180 8186
rect 8180 8134 8210 8186
rect 8234 8134 8244 8186
rect 8244 8134 8290 8186
rect 7994 8132 8050 8134
rect 8074 8132 8130 8134
rect 8154 8132 8210 8134
rect 8234 8132 8290 8134
rect 7838 7112 7894 7168
rect 7746 6296 7802 6352
rect 7654 6060 7656 6080
rect 7656 6060 7708 6080
rect 7708 6060 7710 6080
rect 7654 6024 7710 6060
rect 7994 7098 8050 7100
rect 8074 7098 8130 7100
rect 8154 7098 8210 7100
rect 8234 7098 8290 7100
rect 7994 7046 8040 7098
rect 8040 7046 8050 7098
rect 8074 7046 8104 7098
rect 8104 7046 8116 7098
rect 8116 7046 8130 7098
rect 8154 7046 8168 7098
rect 8168 7046 8180 7098
rect 8180 7046 8210 7098
rect 8234 7046 8244 7098
rect 8244 7046 8290 7098
rect 7994 7044 8050 7046
rect 8074 7044 8130 7046
rect 8154 7044 8210 7046
rect 8234 7044 8290 7046
rect 8390 6160 8446 6216
rect 7994 6010 8050 6012
rect 8074 6010 8130 6012
rect 8154 6010 8210 6012
rect 8234 6010 8290 6012
rect 7994 5958 8040 6010
rect 8040 5958 8050 6010
rect 8074 5958 8104 6010
rect 8104 5958 8116 6010
rect 8116 5958 8130 6010
rect 8154 5958 8168 6010
rect 8168 5958 8180 6010
rect 8180 5958 8210 6010
rect 8234 5958 8244 6010
rect 8244 5958 8290 6010
rect 7994 5956 8050 5958
rect 8074 5956 8130 5958
rect 8154 5956 8210 5958
rect 8234 5956 8290 5958
rect 7994 4922 8050 4924
rect 8074 4922 8130 4924
rect 8154 4922 8210 4924
rect 8234 4922 8290 4924
rect 7994 4870 8040 4922
rect 8040 4870 8050 4922
rect 8074 4870 8104 4922
rect 8104 4870 8116 4922
rect 8116 4870 8130 4922
rect 8154 4870 8168 4922
rect 8168 4870 8180 4922
rect 8180 4870 8210 4922
rect 8234 4870 8244 4922
rect 8244 4870 8290 4922
rect 7994 4868 8050 4870
rect 8074 4868 8130 4870
rect 8154 4868 8210 4870
rect 8234 4868 8290 4870
rect 7378 2216 7434 2272
rect 7994 3834 8050 3836
rect 8074 3834 8130 3836
rect 8154 3834 8210 3836
rect 8234 3834 8290 3836
rect 7994 3782 8040 3834
rect 8040 3782 8050 3834
rect 8074 3782 8104 3834
rect 8104 3782 8116 3834
rect 8116 3782 8130 3834
rect 8154 3782 8168 3834
rect 8168 3782 8180 3834
rect 8180 3782 8210 3834
rect 8234 3782 8244 3834
rect 8244 3782 8290 3834
rect 7994 3780 8050 3782
rect 8074 3780 8130 3782
rect 8154 3780 8210 3782
rect 8234 3780 8290 3782
rect 7994 2746 8050 2748
rect 8074 2746 8130 2748
rect 8154 2746 8210 2748
rect 8234 2746 8290 2748
rect 7994 2694 8040 2746
rect 8040 2694 8050 2746
rect 8074 2694 8104 2746
rect 8104 2694 8116 2746
rect 8116 2694 8130 2746
rect 8154 2694 8168 2746
rect 8168 2694 8180 2746
rect 8180 2694 8210 2746
rect 8234 2694 8244 2746
rect 8244 2694 8290 2746
rect 7994 2692 8050 2694
rect 8074 2692 8130 2694
rect 8154 2692 8210 2694
rect 8234 2692 8290 2694
rect 9862 9560 9918 9616
rect 9678 7792 9734 7848
rect 8942 5208 8998 5264
rect 8850 4528 8906 4584
rect 7994 1658 8050 1660
rect 8074 1658 8130 1660
rect 8154 1658 8210 1660
rect 8234 1658 8290 1660
rect 7994 1606 8040 1658
rect 8040 1606 8050 1658
rect 8074 1606 8104 1658
rect 8104 1606 8116 1658
rect 8116 1606 8130 1658
rect 8154 1606 8168 1658
rect 8168 1606 8180 1658
rect 8180 1606 8210 1658
rect 8234 1606 8244 1658
rect 8244 1606 8290 1658
rect 7994 1604 8050 1606
rect 8074 1604 8130 1606
rect 8154 1604 8210 1606
rect 8234 1604 8290 1606
rect 7746 1536 7802 1592
rect 8298 992 8354 1048
rect 8942 3304 8998 3360
rect 9310 3440 9366 3496
rect 9126 1808 9182 1864
rect 9310 1808 9366 1864
rect 10598 17448 10654 17504
rect 10414 16768 10470 16824
rect 10322 15680 10378 15736
rect 10506 14864 10562 14920
rect 10874 21256 10930 21312
rect 10874 20712 10930 20768
rect 10874 19488 10930 19544
rect 11789 21786 11845 21788
rect 11869 21786 11925 21788
rect 11949 21786 12005 21788
rect 12029 21786 12085 21788
rect 11789 21734 11835 21786
rect 11835 21734 11845 21786
rect 11869 21734 11899 21786
rect 11899 21734 11911 21786
rect 11911 21734 11925 21786
rect 11949 21734 11963 21786
rect 11963 21734 11975 21786
rect 11975 21734 12005 21786
rect 12029 21734 12039 21786
rect 12039 21734 12085 21786
rect 11789 21732 11845 21734
rect 11869 21732 11925 21734
rect 11949 21732 12005 21734
rect 12029 21732 12085 21734
rect 12162 21664 12218 21720
rect 11518 20712 11574 20768
rect 12162 20984 12218 21040
rect 11789 20698 11845 20700
rect 11869 20698 11925 20700
rect 11949 20698 12005 20700
rect 12029 20698 12085 20700
rect 11789 20646 11835 20698
rect 11835 20646 11845 20698
rect 11869 20646 11899 20698
rect 11899 20646 11911 20698
rect 11911 20646 11925 20698
rect 11949 20646 11963 20698
rect 11963 20646 11975 20698
rect 11975 20646 12005 20698
rect 12029 20646 12039 20698
rect 12039 20646 12085 20698
rect 11789 20644 11845 20646
rect 11869 20644 11925 20646
rect 11949 20644 12005 20646
rect 12029 20644 12085 20646
rect 10966 18536 11022 18592
rect 11789 19610 11845 19612
rect 11869 19610 11925 19612
rect 11949 19610 12005 19612
rect 12029 19610 12085 19612
rect 11789 19558 11835 19610
rect 11835 19558 11845 19610
rect 11869 19558 11899 19610
rect 11899 19558 11911 19610
rect 11911 19558 11925 19610
rect 11949 19558 11963 19610
rect 11963 19558 11975 19610
rect 11975 19558 12005 19610
rect 12029 19558 12039 19610
rect 12039 19558 12085 19610
rect 11789 19556 11845 19558
rect 11869 19556 11925 19558
rect 11949 19556 12005 19558
rect 12029 19556 12085 19558
rect 11702 19080 11758 19136
rect 10690 14864 10746 14920
rect 10322 12144 10378 12200
rect 10322 11328 10378 11384
rect 10782 14184 10838 14240
rect 11058 16088 11114 16144
rect 11789 18522 11845 18524
rect 11869 18522 11925 18524
rect 11949 18522 12005 18524
rect 12029 18522 12085 18524
rect 11789 18470 11835 18522
rect 11835 18470 11845 18522
rect 11869 18470 11899 18522
rect 11899 18470 11911 18522
rect 11911 18470 11925 18522
rect 11949 18470 11963 18522
rect 11963 18470 11975 18522
rect 11975 18470 12005 18522
rect 12029 18470 12039 18522
rect 12039 18470 12085 18522
rect 11789 18468 11845 18470
rect 11869 18468 11925 18470
rect 11949 18468 12005 18470
rect 12029 18468 12085 18470
rect 11789 17434 11845 17436
rect 11869 17434 11925 17436
rect 11949 17434 12005 17436
rect 12029 17434 12085 17436
rect 11789 17382 11835 17434
rect 11835 17382 11845 17434
rect 11869 17382 11899 17434
rect 11899 17382 11911 17434
rect 11911 17382 11925 17434
rect 11949 17382 11963 17434
rect 11963 17382 11975 17434
rect 11975 17382 12005 17434
rect 12029 17382 12039 17434
rect 12039 17382 12085 17434
rect 11789 17380 11845 17382
rect 11869 17380 11925 17382
rect 11949 17380 12005 17382
rect 12029 17380 12085 17382
rect 11702 16632 11758 16688
rect 11150 15680 11206 15736
rect 11058 15408 11114 15464
rect 11150 15272 11206 15328
rect 11058 15136 11114 15192
rect 10598 13132 10600 13152
rect 10600 13132 10652 13152
rect 10652 13132 10654 13152
rect 10598 13096 10654 13132
rect 10598 11464 10654 11520
rect 11150 14592 11206 14648
rect 12254 17176 12310 17232
rect 11789 16346 11845 16348
rect 11869 16346 11925 16348
rect 11949 16346 12005 16348
rect 12029 16346 12085 16348
rect 11789 16294 11835 16346
rect 11835 16294 11845 16346
rect 11869 16294 11899 16346
rect 11899 16294 11911 16346
rect 11911 16294 11925 16346
rect 11949 16294 11963 16346
rect 11963 16294 11975 16346
rect 11975 16294 12005 16346
rect 12029 16294 12039 16346
rect 12039 16294 12085 16346
rect 11789 16292 11845 16294
rect 11869 16292 11925 16294
rect 11949 16292 12005 16294
rect 12029 16292 12085 16294
rect 12346 16088 12402 16144
rect 11789 15258 11845 15260
rect 11869 15258 11925 15260
rect 11949 15258 12005 15260
rect 12029 15258 12085 15260
rect 11789 15206 11835 15258
rect 11835 15206 11845 15258
rect 11869 15206 11899 15258
rect 11899 15206 11911 15258
rect 11911 15206 11925 15258
rect 11949 15206 11963 15258
rect 11963 15206 11975 15258
rect 11975 15206 12005 15258
rect 12029 15206 12039 15258
rect 12039 15206 12085 15258
rect 11789 15204 11845 15206
rect 11869 15204 11925 15206
rect 11949 15204 12005 15206
rect 12029 15204 12085 15206
rect 11150 13640 11206 13696
rect 11058 13504 11114 13560
rect 11789 14170 11845 14172
rect 11869 14170 11925 14172
rect 11949 14170 12005 14172
rect 12029 14170 12085 14172
rect 11789 14118 11835 14170
rect 11835 14118 11845 14170
rect 11869 14118 11899 14170
rect 11899 14118 11911 14170
rect 11911 14118 11925 14170
rect 11949 14118 11963 14170
rect 11963 14118 11975 14170
rect 11975 14118 12005 14170
rect 12029 14118 12039 14170
rect 12039 14118 12085 14170
rect 11789 14116 11845 14118
rect 11869 14116 11925 14118
rect 11949 14116 12005 14118
rect 12029 14116 12085 14118
rect 11886 13912 11942 13968
rect 14002 21972 14004 21992
rect 14004 21972 14056 21992
rect 14056 21972 14058 21992
rect 14002 21936 14058 21972
rect 14094 20984 14150 21040
rect 22282 22208 22338 22244
rect 23754 22244 23756 22264
rect 23756 22244 23808 22264
rect 23808 22244 23810 22264
rect 14646 20984 14702 21040
rect 13358 20168 13414 20224
rect 13818 20712 13874 20768
rect 13910 20032 13966 20088
rect 11334 12960 11390 13016
rect 11150 12824 11206 12880
rect 10782 11464 10838 11520
rect 10598 10648 10654 10704
rect 11150 12300 11206 12336
rect 11150 12280 11152 12300
rect 11152 12280 11204 12300
rect 11204 12280 11206 12300
rect 10966 11600 11022 11656
rect 10874 9696 10930 9752
rect 10690 9288 10746 9344
rect 11789 13082 11845 13084
rect 11869 13082 11925 13084
rect 11949 13082 12005 13084
rect 12029 13082 12085 13084
rect 11789 13030 11835 13082
rect 11835 13030 11845 13082
rect 11869 13030 11899 13082
rect 11899 13030 11911 13082
rect 11911 13030 11925 13082
rect 11949 13030 11963 13082
rect 11963 13030 11975 13082
rect 11975 13030 12005 13082
rect 12029 13030 12039 13082
rect 12039 13030 12085 13082
rect 11789 13028 11845 13030
rect 11869 13028 11925 13030
rect 11949 13028 12005 13030
rect 12029 13028 12085 13030
rect 11610 12416 11666 12472
rect 11426 10376 11482 10432
rect 11426 8472 11482 8528
rect 10874 8200 10930 8256
rect 10506 8064 10562 8120
rect 10598 6024 10654 6080
rect 10690 5616 10746 5672
rect 10782 5072 10838 5128
rect 12162 12552 12218 12608
rect 11978 12144 12034 12200
rect 11789 11994 11845 11996
rect 11869 11994 11925 11996
rect 11949 11994 12005 11996
rect 12029 11994 12085 11996
rect 11789 11942 11835 11994
rect 11835 11942 11845 11994
rect 11869 11942 11899 11994
rect 11899 11942 11911 11994
rect 11911 11942 11925 11994
rect 11949 11942 11963 11994
rect 11963 11942 11975 11994
rect 11975 11942 12005 11994
rect 12029 11942 12039 11994
rect 12039 11942 12085 11994
rect 11789 11940 11845 11942
rect 11869 11940 11925 11942
rect 11949 11940 12005 11942
rect 12029 11940 12085 11942
rect 12162 11872 12218 11928
rect 13174 16224 13230 16280
rect 12990 15816 13046 15872
rect 12806 14900 12808 14920
rect 12808 14900 12860 14920
rect 12860 14900 12862 14920
rect 12806 14864 12862 14900
rect 13266 15544 13322 15600
rect 13174 14592 13230 14648
rect 12714 12416 12770 12472
rect 12346 12008 12402 12064
rect 11794 11076 11850 11112
rect 11794 11056 11796 11076
rect 11796 11056 11848 11076
rect 11848 11056 11850 11076
rect 11789 10906 11845 10908
rect 11869 10906 11925 10908
rect 11949 10906 12005 10908
rect 12029 10906 12085 10908
rect 11789 10854 11835 10906
rect 11835 10854 11845 10906
rect 11869 10854 11899 10906
rect 11899 10854 11911 10906
rect 11911 10854 11925 10906
rect 11949 10854 11963 10906
rect 11963 10854 11975 10906
rect 11975 10854 12005 10906
rect 12029 10854 12039 10906
rect 12039 10854 12085 10906
rect 11789 10852 11845 10854
rect 11869 10852 11925 10854
rect 11949 10852 12005 10854
rect 12029 10852 12085 10854
rect 11789 9818 11845 9820
rect 11869 9818 11925 9820
rect 11949 9818 12005 9820
rect 12029 9818 12085 9820
rect 11789 9766 11835 9818
rect 11835 9766 11845 9818
rect 11869 9766 11899 9818
rect 11899 9766 11911 9818
rect 11911 9766 11925 9818
rect 11949 9766 11963 9818
rect 11963 9766 11975 9818
rect 11975 9766 12005 9818
rect 12029 9766 12039 9818
rect 12039 9766 12085 9818
rect 11789 9764 11845 9766
rect 11869 9764 11925 9766
rect 11949 9764 12005 9766
rect 12029 9764 12085 9766
rect 11789 8730 11845 8732
rect 11869 8730 11925 8732
rect 11949 8730 12005 8732
rect 12029 8730 12085 8732
rect 11789 8678 11835 8730
rect 11835 8678 11845 8730
rect 11869 8678 11899 8730
rect 11899 8678 11911 8730
rect 11911 8678 11925 8730
rect 11949 8678 11963 8730
rect 11963 8678 11975 8730
rect 11975 8678 12005 8730
rect 12029 8678 12039 8730
rect 12039 8678 12085 8730
rect 11789 8676 11845 8678
rect 11869 8676 11925 8678
rect 11949 8676 12005 8678
rect 12029 8676 12085 8678
rect 12070 8064 12126 8120
rect 12346 9152 12402 9208
rect 12254 8472 12310 8528
rect 11789 7642 11845 7644
rect 11869 7642 11925 7644
rect 11949 7642 12005 7644
rect 12029 7642 12085 7644
rect 11789 7590 11835 7642
rect 11835 7590 11845 7642
rect 11869 7590 11899 7642
rect 11899 7590 11911 7642
rect 11911 7590 11925 7642
rect 11949 7590 11963 7642
rect 11963 7590 11975 7642
rect 11975 7590 12005 7642
rect 12029 7590 12039 7642
rect 12039 7590 12085 7642
rect 11789 7588 11845 7590
rect 11869 7588 11925 7590
rect 11949 7588 12005 7590
rect 12029 7588 12085 7590
rect 11610 7112 11666 7168
rect 12622 11872 12678 11928
rect 12622 10240 12678 10296
rect 12530 9560 12586 9616
rect 11058 6704 11114 6760
rect 11789 6554 11845 6556
rect 11869 6554 11925 6556
rect 11949 6554 12005 6556
rect 12029 6554 12085 6556
rect 11789 6502 11835 6554
rect 11835 6502 11845 6554
rect 11869 6502 11899 6554
rect 11899 6502 11911 6554
rect 11911 6502 11925 6554
rect 11949 6502 11963 6554
rect 11963 6502 11975 6554
rect 11975 6502 12005 6554
rect 12029 6502 12039 6554
rect 12039 6502 12085 6554
rect 11789 6500 11845 6502
rect 11869 6500 11925 6502
rect 11949 6500 12005 6502
rect 12029 6500 12085 6502
rect 13542 19624 13598 19680
rect 13634 19352 13690 19408
rect 14002 19352 14058 19408
rect 13450 18944 13506 19000
rect 13542 18400 13598 18456
rect 14278 18672 14334 18728
rect 13542 15020 13598 15056
rect 13542 15000 13544 15020
rect 13544 15000 13596 15020
rect 13596 15000 13598 15020
rect 13818 14320 13874 14376
rect 13450 12552 13506 12608
rect 13450 11872 13506 11928
rect 11150 4800 11206 4856
rect 10414 3984 10470 4040
rect 9678 1128 9734 1184
rect 11426 6024 11482 6080
rect 12346 5752 12402 5808
rect 11789 5466 11845 5468
rect 11869 5466 11925 5468
rect 11949 5466 12005 5468
rect 12029 5466 12085 5468
rect 11789 5414 11835 5466
rect 11835 5414 11845 5466
rect 11869 5414 11899 5466
rect 11899 5414 11911 5466
rect 11911 5414 11925 5466
rect 11949 5414 11963 5466
rect 11963 5414 11975 5466
rect 11975 5414 12005 5466
rect 12029 5414 12039 5466
rect 12039 5414 12085 5466
rect 11789 5412 11845 5414
rect 11869 5412 11925 5414
rect 11949 5412 12005 5414
rect 12029 5412 12085 5414
rect 11978 4800 12034 4856
rect 11789 4378 11845 4380
rect 11869 4378 11925 4380
rect 11949 4378 12005 4380
rect 12029 4378 12085 4380
rect 11789 4326 11835 4378
rect 11835 4326 11845 4378
rect 11869 4326 11899 4378
rect 11899 4326 11911 4378
rect 11911 4326 11925 4378
rect 11949 4326 11963 4378
rect 11963 4326 11975 4378
rect 11975 4326 12005 4378
rect 12029 4326 12039 4378
rect 12039 4326 12085 4378
rect 11789 4324 11845 4326
rect 11869 4324 11925 4326
rect 11949 4324 12005 4326
rect 12029 4324 12085 4326
rect 11789 3290 11845 3292
rect 11869 3290 11925 3292
rect 11949 3290 12005 3292
rect 12029 3290 12085 3292
rect 11789 3238 11835 3290
rect 11835 3238 11845 3290
rect 11869 3238 11899 3290
rect 11899 3238 11911 3290
rect 11911 3238 11925 3290
rect 11949 3238 11963 3290
rect 11963 3238 11975 3290
rect 11975 3238 12005 3290
rect 12029 3238 12039 3290
rect 12039 3238 12085 3290
rect 11789 3236 11845 3238
rect 11869 3236 11925 3238
rect 11949 3236 12005 3238
rect 12029 3236 12085 3238
rect 12806 6160 12862 6216
rect 11789 2202 11845 2204
rect 11869 2202 11925 2204
rect 11949 2202 12005 2204
rect 12029 2202 12085 2204
rect 11789 2150 11835 2202
rect 11835 2150 11845 2202
rect 11869 2150 11899 2202
rect 11899 2150 11911 2202
rect 11911 2150 11925 2202
rect 11949 2150 11963 2202
rect 11963 2150 11975 2202
rect 11975 2150 12005 2202
rect 12029 2150 12039 2202
rect 12039 2150 12085 2202
rect 11789 2148 11845 2150
rect 11869 2148 11925 2150
rect 11949 2148 12005 2150
rect 12029 2148 12085 2150
rect 12254 1808 12310 1864
rect 11426 1400 11482 1456
rect 7994 570 8050 572
rect 8074 570 8130 572
rect 8154 570 8210 572
rect 8234 570 8290 572
rect 7994 518 8040 570
rect 8040 518 8050 570
rect 8074 518 8104 570
rect 8104 518 8116 570
rect 8116 518 8130 570
rect 8154 518 8168 570
rect 8168 518 8180 570
rect 8180 518 8210 570
rect 8234 518 8244 570
rect 8244 518 8290 570
rect 7994 516 8050 518
rect 8074 516 8130 518
rect 8154 516 8210 518
rect 8234 516 8290 518
rect 9218 312 9274 368
rect 11789 1114 11845 1116
rect 11869 1114 11925 1116
rect 11949 1114 12005 1116
rect 12029 1114 12085 1116
rect 11789 1062 11835 1114
rect 11835 1062 11845 1114
rect 11869 1062 11899 1114
rect 11899 1062 11911 1114
rect 11911 1062 11925 1114
rect 11949 1062 11963 1114
rect 11963 1062 11975 1114
rect 11975 1062 12005 1114
rect 12029 1062 12039 1114
rect 12039 1062 12085 1114
rect 11789 1060 11845 1062
rect 11869 1060 11925 1062
rect 11949 1060 12005 1062
rect 12029 1060 12085 1062
rect 13726 13796 13782 13832
rect 13726 13776 13728 13796
rect 13728 13776 13780 13796
rect 13780 13776 13782 13796
rect 13726 13232 13782 13288
rect 13726 12008 13782 12064
rect 13174 10376 13230 10432
rect 13174 9288 13230 9344
rect 13082 8336 13138 8392
rect 14094 12144 14150 12200
rect 13726 7948 13782 7984
rect 13726 7928 13728 7948
rect 13728 7928 13780 7948
rect 13780 7928 13782 7948
rect 14554 18808 14610 18864
rect 15382 21256 15438 21312
rect 15198 20460 15254 20496
rect 15198 20440 15200 20460
rect 15200 20440 15252 20460
rect 15252 20440 15254 20460
rect 15106 19352 15162 19408
rect 15014 19216 15070 19272
rect 15106 19116 15108 19136
rect 15108 19116 15160 19136
rect 15160 19116 15162 19136
rect 15106 19080 15162 19116
rect 15106 18944 15162 19000
rect 14554 16632 14610 16688
rect 14462 16224 14518 16280
rect 14462 15156 14518 15192
rect 14462 15136 14464 15156
rect 14464 15136 14516 15156
rect 14516 15136 14518 15156
rect 14554 14864 14610 14920
rect 15382 19896 15438 19952
rect 16118 21256 16174 21312
rect 15584 21242 15640 21244
rect 15664 21242 15720 21244
rect 15744 21242 15800 21244
rect 15824 21242 15880 21244
rect 15584 21190 15630 21242
rect 15630 21190 15640 21242
rect 15664 21190 15694 21242
rect 15694 21190 15706 21242
rect 15706 21190 15720 21242
rect 15744 21190 15758 21242
rect 15758 21190 15770 21242
rect 15770 21190 15800 21242
rect 15824 21190 15834 21242
rect 15834 21190 15880 21242
rect 15584 21188 15640 21190
rect 15664 21188 15720 21190
rect 15744 21188 15800 21190
rect 15824 21188 15880 21190
rect 16762 21664 16818 21720
rect 15750 20440 15806 20496
rect 15584 20154 15640 20156
rect 15664 20154 15720 20156
rect 15744 20154 15800 20156
rect 15824 20154 15880 20156
rect 15584 20102 15630 20154
rect 15630 20102 15640 20154
rect 15664 20102 15694 20154
rect 15694 20102 15706 20154
rect 15706 20102 15720 20154
rect 15744 20102 15758 20154
rect 15758 20102 15770 20154
rect 15770 20102 15800 20154
rect 15824 20102 15834 20154
rect 15834 20102 15880 20154
rect 15584 20100 15640 20102
rect 15664 20100 15720 20102
rect 15744 20100 15800 20102
rect 15824 20100 15880 20102
rect 15750 19488 15806 19544
rect 15584 19066 15640 19068
rect 15664 19066 15720 19068
rect 15744 19066 15800 19068
rect 15824 19066 15880 19068
rect 15584 19014 15630 19066
rect 15630 19014 15640 19066
rect 15664 19014 15694 19066
rect 15694 19014 15706 19066
rect 15706 19014 15720 19066
rect 15744 19014 15758 19066
rect 15758 19014 15770 19066
rect 15770 19014 15800 19066
rect 15824 19014 15834 19066
rect 15834 19014 15880 19066
rect 15584 19012 15640 19014
rect 15664 19012 15720 19014
rect 15744 19012 15800 19014
rect 15824 19012 15880 19014
rect 15584 17978 15640 17980
rect 15664 17978 15720 17980
rect 15744 17978 15800 17980
rect 15824 17978 15880 17980
rect 15584 17926 15630 17978
rect 15630 17926 15640 17978
rect 15664 17926 15694 17978
rect 15694 17926 15706 17978
rect 15706 17926 15720 17978
rect 15744 17926 15758 17978
rect 15758 17926 15770 17978
rect 15770 17926 15800 17978
rect 15824 17926 15834 17978
rect 15834 17926 15880 17978
rect 15584 17924 15640 17926
rect 15664 17924 15720 17926
rect 15744 17924 15800 17926
rect 15824 17924 15880 17926
rect 15474 17584 15530 17640
rect 15198 16904 15254 16960
rect 15106 14456 15162 14512
rect 15584 16890 15640 16892
rect 15664 16890 15720 16892
rect 15744 16890 15800 16892
rect 15824 16890 15880 16892
rect 15584 16838 15630 16890
rect 15630 16838 15640 16890
rect 15664 16838 15694 16890
rect 15694 16838 15706 16890
rect 15706 16838 15720 16890
rect 15744 16838 15758 16890
rect 15758 16838 15770 16890
rect 15770 16838 15800 16890
rect 15824 16838 15834 16890
rect 15834 16838 15880 16890
rect 15584 16836 15640 16838
rect 15664 16836 15720 16838
rect 15744 16836 15800 16838
rect 15824 16836 15880 16838
rect 16210 20168 16266 20224
rect 16210 19624 16266 19680
rect 16118 18128 16174 18184
rect 16486 19080 16542 19136
rect 16394 18264 16450 18320
rect 16210 17040 16266 17096
rect 15106 13912 15162 13968
rect 15584 15802 15640 15804
rect 15664 15802 15720 15804
rect 15744 15802 15800 15804
rect 15824 15802 15880 15804
rect 15584 15750 15630 15802
rect 15630 15750 15640 15802
rect 15664 15750 15694 15802
rect 15694 15750 15706 15802
rect 15706 15750 15720 15802
rect 15744 15750 15758 15802
rect 15758 15750 15770 15802
rect 15770 15750 15800 15802
rect 15824 15750 15834 15802
rect 15834 15750 15880 15802
rect 15584 15748 15640 15750
rect 15664 15748 15720 15750
rect 15744 15748 15800 15750
rect 15824 15748 15880 15750
rect 16118 16496 16174 16552
rect 15584 14714 15640 14716
rect 15664 14714 15720 14716
rect 15744 14714 15800 14716
rect 15824 14714 15880 14716
rect 15584 14662 15630 14714
rect 15630 14662 15640 14714
rect 15664 14662 15694 14714
rect 15694 14662 15706 14714
rect 15706 14662 15720 14714
rect 15744 14662 15758 14714
rect 15758 14662 15770 14714
rect 15770 14662 15800 14714
rect 15824 14662 15834 14714
rect 15834 14662 15880 14714
rect 15584 14660 15640 14662
rect 15664 14660 15720 14662
rect 15744 14660 15800 14662
rect 15824 14660 15880 14662
rect 15584 13626 15640 13628
rect 15664 13626 15720 13628
rect 15744 13626 15800 13628
rect 15824 13626 15880 13628
rect 15584 13574 15630 13626
rect 15630 13574 15640 13626
rect 15664 13574 15694 13626
rect 15694 13574 15706 13626
rect 15706 13574 15720 13626
rect 15744 13574 15758 13626
rect 15758 13574 15770 13626
rect 15770 13574 15800 13626
rect 15824 13574 15834 13626
rect 15834 13574 15880 13626
rect 15584 13572 15640 13574
rect 15664 13572 15720 13574
rect 15744 13572 15800 13574
rect 15824 13572 15880 13574
rect 15584 12538 15640 12540
rect 15664 12538 15720 12540
rect 15744 12538 15800 12540
rect 15824 12538 15880 12540
rect 15584 12486 15630 12538
rect 15630 12486 15640 12538
rect 15664 12486 15694 12538
rect 15694 12486 15706 12538
rect 15706 12486 15720 12538
rect 15744 12486 15758 12538
rect 15758 12486 15770 12538
rect 15770 12486 15800 12538
rect 15824 12486 15834 12538
rect 15834 12486 15880 12538
rect 15584 12484 15640 12486
rect 15664 12484 15720 12486
rect 15744 12484 15800 12486
rect 15824 12484 15880 12486
rect 16118 14320 16174 14376
rect 15106 8336 15162 8392
rect 14370 8200 14426 8256
rect 13726 6840 13782 6896
rect 14186 7656 14242 7712
rect 13910 6860 13966 6896
rect 13910 6840 13912 6860
rect 13912 6840 13964 6860
rect 13964 6840 13966 6860
rect 12806 2352 12862 2408
rect 6642 176 6698 232
rect 14646 6160 14702 6216
rect 14922 7112 14978 7168
rect 15842 12180 15844 12200
rect 15844 12180 15896 12200
rect 15896 12180 15898 12200
rect 15842 12144 15898 12180
rect 15584 11450 15640 11452
rect 15664 11450 15720 11452
rect 15744 11450 15800 11452
rect 15824 11450 15880 11452
rect 15584 11398 15630 11450
rect 15630 11398 15640 11450
rect 15664 11398 15694 11450
rect 15694 11398 15706 11450
rect 15706 11398 15720 11450
rect 15744 11398 15758 11450
rect 15758 11398 15770 11450
rect 15770 11398 15800 11450
rect 15824 11398 15834 11450
rect 15834 11398 15880 11450
rect 15584 11396 15640 11398
rect 15664 11396 15720 11398
rect 15744 11396 15800 11398
rect 15824 11396 15880 11398
rect 15934 10648 15990 10704
rect 15584 10362 15640 10364
rect 15664 10362 15720 10364
rect 15744 10362 15800 10364
rect 15824 10362 15880 10364
rect 15584 10310 15630 10362
rect 15630 10310 15640 10362
rect 15664 10310 15694 10362
rect 15694 10310 15706 10362
rect 15706 10310 15720 10362
rect 15744 10310 15758 10362
rect 15758 10310 15770 10362
rect 15770 10310 15800 10362
rect 15824 10310 15834 10362
rect 15834 10310 15880 10362
rect 15584 10308 15640 10310
rect 15664 10308 15720 10310
rect 15744 10308 15800 10310
rect 15824 10308 15880 10310
rect 15584 9274 15640 9276
rect 15664 9274 15720 9276
rect 15744 9274 15800 9276
rect 15824 9274 15880 9276
rect 15584 9222 15630 9274
rect 15630 9222 15640 9274
rect 15664 9222 15694 9274
rect 15694 9222 15706 9274
rect 15706 9222 15720 9274
rect 15744 9222 15758 9274
rect 15758 9222 15770 9274
rect 15770 9222 15800 9274
rect 15824 9222 15834 9274
rect 15834 9222 15880 9274
rect 15584 9220 15640 9222
rect 15664 9220 15720 9222
rect 15744 9220 15800 9222
rect 15824 9220 15880 9222
rect 15584 8186 15640 8188
rect 15664 8186 15720 8188
rect 15744 8186 15800 8188
rect 15824 8186 15880 8188
rect 15584 8134 15630 8186
rect 15630 8134 15640 8186
rect 15664 8134 15694 8186
rect 15694 8134 15706 8186
rect 15706 8134 15720 8186
rect 15744 8134 15758 8186
rect 15758 8134 15770 8186
rect 15770 8134 15800 8186
rect 15824 8134 15834 8186
rect 15834 8134 15880 8186
rect 15584 8132 15640 8134
rect 15664 8132 15720 8134
rect 15744 8132 15800 8134
rect 15824 8132 15880 8134
rect 15566 7656 15622 7712
rect 15658 7384 15714 7440
rect 15584 7098 15640 7100
rect 15664 7098 15720 7100
rect 15744 7098 15800 7100
rect 15824 7098 15880 7100
rect 15584 7046 15630 7098
rect 15630 7046 15640 7098
rect 15664 7046 15694 7098
rect 15694 7046 15706 7098
rect 15706 7046 15720 7098
rect 15744 7046 15758 7098
rect 15758 7046 15770 7098
rect 15770 7046 15800 7098
rect 15824 7046 15834 7098
rect 15834 7046 15880 7098
rect 15584 7044 15640 7046
rect 15664 7044 15720 7046
rect 15744 7044 15800 7046
rect 15824 7044 15880 7046
rect 16302 16496 16358 16552
rect 16670 18808 16726 18864
rect 16854 18264 16910 18320
rect 17590 20984 17646 21040
rect 18050 20848 18106 20904
rect 17130 18128 17186 18184
rect 16762 17856 16818 17912
rect 17038 16088 17094 16144
rect 16854 15544 16910 15600
rect 16578 14864 16634 14920
rect 17130 15020 17186 15056
rect 17130 15000 17132 15020
rect 17132 15000 17184 15020
rect 17184 15000 17186 15020
rect 16946 13776 17002 13832
rect 15658 6724 15714 6760
rect 15658 6704 15660 6724
rect 15660 6704 15712 6724
rect 15712 6704 15714 6724
rect 15584 6010 15640 6012
rect 15664 6010 15720 6012
rect 15744 6010 15800 6012
rect 15824 6010 15880 6012
rect 15584 5958 15630 6010
rect 15630 5958 15640 6010
rect 15664 5958 15694 6010
rect 15694 5958 15706 6010
rect 15706 5958 15720 6010
rect 15744 5958 15758 6010
rect 15758 5958 15770 6010
rect 15770 5958 15800 6010
rect 15824 5958 15834 6010
rect 15834 5958 15880 6010
rect 15584 5956 15640 5958
rect 15664 5956 15720 5958
rect 15744 5956 15800 5958
rect 15824 5956 15880 5958
rect 14738 3032 14794 3088
rect 14738 1400 14794 1456
rect 15584 4922 15640 4924
rect 15664 4922 15720 4924
rect 15744 4922 15800 4924
rect 15824 4922 15880 4924
rect 15584 4870 15630 4922
rect 15630 4870 15640 4922
rect 15664 4870 15694 4922
rect 15694 4870 15706 4922
rect 15706 4870 15720 4922
rect 15744 4870 15758 4922
rect 15758 4870 15770 4922
rect 15770 4870 15800 4922
rect 15824 4870 15834 4922
rect 15834 4870 15880 4922
rect 15584 4868 15640 4870
rect 15664 4868 15720 4870
rect 15744 4868 15800 4870
rect 15824 4868 15880 4870
rect 16670 12688 16726 12744
rect 16394 10648 16450 10704
rect 16210 7792 16266 7848
rect 16394 6860 16450 6896
rect 16394 6840 16396 6860
rect 16396 6840 16448 6860
rect 16448 6840 16450 6860
rect 15584 3834 15640 3836
rect 15664 3834 15720 3836
rect 15744 3834 15800 3836
rect 15824 3834 15880 3836
rect 15584 3782 15630 3834
rect 15630 3782 15640 3834
rect 15664 3782 15694 3834
rect 15694 3782 15706 3834
rect 15706 3782 15720 3834
rect 15744 3782 15758 3834
rect 15758 3782 15770 3834
rect 15770 3782 15800 3834
rect 15824 3782 15834 3834
rect 15834 3782 15880 3834
rect 15584 3780 15640 3782
rect 15664 3780 15720 3782
rect 15744 3780 15800 3782
rect 15824 3780 15880 3782
rect 15584 2746 15640 2748
rect 15664 2746 15720 2748
rect 15744 2746 15800 2748
rect 15824 2746 15880 2748
rect 15584 2694 15630 2746
rect 15630 2694 15640 2746
rect 15664 2694 15694 2746
rect 15694 2694 15706 2746
rect 15706 2694 15720 2746
rect 15744 2694 15758 2746
rect 15758 2694 15770 2746
rect 15770 2694 15800 2746
rect 15824 2694 15834 2746
rect 15834 2694 15880 2746
rect 15584 2692 15640 2694
rect 15664 2692 15720 2694
rect 15744 2692 15800 2694
rect 15824 2692 15880 2694
rect 15584 1658 15640 1660
rect 15664 1658 15720 1660
rect 15744 1658 15800 1660
rect 15824 1658 15880 1660
rect 15584 1606 15630 1658
rect 15630 1606 15640 1658
rect 15664 1606 15694 1658
rect 15694 1606 15706 1658
rect 15706 1606 15720 1658
rect 15744 1606 15758 1658
rect 15758 1606 15770 1658
rect 15770 1606 15800 1658
rect 15824 1606 15834 1658
rect 15834 1606 15880 1658
rect 15584 1604 15640 1606
rect 15664 1604 15720 1606
rect 15744 1604 15800 1606
rect 15824 1604 15880 1606
rect 17314 19252 17316 19272
rect 17316 19252 17368 19272
rect 17368 19252 17370 19272
rect 17314 19216 17370 19252
rect 17774 19080 17830 19136
rect 17498 18536 17554 18592
rect 17498 17992 17554 18048
rect 17406 16224 17462 16280
rect 17406 16088 17462 16144
rect 16762 9016 16818 9072
rect 16670 7928 16726 7984
rect 17130 9016 17186 9072
rect 17222 7792 17278 7848
rect 17498 11736 17554 11792
rect 17590 9424 17646 9480
rect 17130 6432 17186 6488
rect 17406 6296 17462 6352
rect 17590 7248 17646 7304
rect 18326 21256 18382 21312
rect 18234 20712 18290 20768
rect 18418 20440 18474 20496
rect 18234 19488 18290 19544
rect 21638 22072 21694 22128
rect 19379 21786 19435 21788
rect 19459 21786 19515 21788
rect 19539 21786 19595 21788
rect 19619 21786 19675 21788
rect 19379 21734 19425 21786
rect 19425 21734 19435 21786
rect 19459 21734 19489 21786
rect 19489 21734 19501 21786
rect 19501 21734 19515 21786
rect 19539 21734 19553 21786
rect 19553 21734 19565 21786
rect 19565 21734 19595 21786
rect 19619 21734 19629 21786
rect 19629 21734 19675 21786
rect 19379 21732 19435 21734
rect 19459 21732 19515 21734
rect 19539 21732 19595 21734
rect 19619 21732 19675 21734
rect 18510 17856 18566 17912
rect 19379 20698 19435 20700
rect 19459 20698 19515 20700
rect 19539 20698 19595 20700
rect 19619 20698 19675 20700
rect 19379 20646 19425 20698
rect 19425 20646 19435 20698
rect 19459 20646 19489 20698
rect 19489 20646 19501 20698
rect 19501 20646 19515 20698
rect 19539 20646 19553 20698
rect 19553 20646 19565 20698
rect 19565 20646 19595 20698
rect 19619 20646 19629 20698
rect 19629 20646 19675 20698
rect 19379 20644 19435 20646
rect 19459 20644 19515 20646
rect 19539 20644 19595 20646
rect 19619 20644 19675 20646
rect 18878 19896 18934 19952
rect 19982 20576 20038 20632
rect 19982 20440 20038 20496
rect 19379 19610 19435 19612
rect 19459 19610 19515 19612
rect 19539 19610 19595 19612
rect 19619 19610 19675 19612
rect 19379 19558 19425 19610
rect 19425 19558 19435 19610
rect 19459 19558 19489 19610
rect 19489 19558 19501 19610
rect 19501 19558 19515 19610
rect 19539 19558 19553 19610
rect 19553 19558 19565 19610
rect 19565 19558 19595 19610
rect 19619 19558 19629 19610
rect 19629 19558 19675 19610
rect 19379 19556 19435 19558
rect 19459 19556 19515 19558
rect 19539 19556 19595 19558
rect 19619 19556 19675 19558
rect 19706 19352 19762 19408
rect 19338 19216 19394 19272
rect 19379 18522 19435 18524
rect 19459 18522 19515 18524
rect 19539 18522 19595 18524
rect 19619 18522 19675 18524
rect 19379 18470 19425 18522
rect 19425 18470 19435 18522
rect 19459 18470 19489 18522
rect 19489 18470 19501 18522
rect 19501 18470 19515 18522
rect 19539 18470 19553 18522
rect 19553 18470 19565 18522
rect 19565 18470 19595 18522
rect 19619 18470 19629 18522
rect 19629 18470 19675 18522
rect 19379 18468 19435 18470
rect 19459 18468 19515 18470
rect 19539 18468 19595 18470
rect 19619 18468 19675 18470
rect 19246 18400 19302 18456
rect 20166 20984 20222 21040
rect 20626 20304 20682 20360
rect 21086 19760 21142 19816
rect 20534 19352 20590 19408
rect 19379 17434 19435 17436
rect 19459 17434 19515 17436
rect 19539 17434 19595 17436
rect 19619 17434 19675 17436
rect 19379 17382 19425 17434
rect 19425 17382 19435 17434
rect 19459 17382 19489 17434
rect 19489 17382 19501 17434
rect 19501 17382 19515 17434
rect 19539 17382 19553 17434
rect 19553 17382 19565 17434
rect 19565 17382 19595 17434
rect 19619 17382 19629 17434
rect 19629 17382 19675 17434
rect 19379 17380 19435 17382
rect 19459 17380 19515 17382
rect 19539 17380 19595 17382
rect 19619 17380 19675 17382
rect 19430 16904 19486 16960
rect 18786 16632 18842 16688
rect 18326 14492 18328 14512
rect 18328 14492 18380 14512
rect 18380 14492 18382 14512
rect 18326 14456 18382 14492
rect 17774 7656 17830 7712
rect 16854 3732 16910 3768
rect 16854 3712 16856 3732
rect 16856 3712 16908 3732
rect 16908 3712 16910 3732
rect 16762 3576 16818 3632
rect 15584 570 15640 572
rect 15664 570 15720 572
rect 15744 570 15800 572
rect 15824 570 15880 572
rect 15584 518 15630 570
rect 15630 518 15640 570
rect 15664 518 15694 570
rect 15694 518 15706 570
rect 15706 518 15720 570
rect 15744 518 15758 570
rect 15758 518 15770 570
rect 15770 518 15800 570
rect 15824 518 15834 570
rect 15834 518 15880 570
rect 15584 516 15640 518
rect 15664 516 15720 518
rect 15744 516 15800 518
rect 15824 516 15880 518
rect 15290 40 15346 96
rect 15566 40 15622 96
rect 17866 3576 17922 3632
rect 18142 3848 18198 3904
rect 18050 3032 18106 3088
rect 17866 1400 17922 1456
rect 18786 14456 18842 14512
rect 19379 16346 19435 16348
rect 19459 16346 19515 16348
rect 19539 16346 19595 16348
rect 19619 16346 19675 16348
rect 19379 16294 19425 16346
rect 19425 16294 19435 16346
rect 19459 16294 19489 16346
rect 19489 16294 19501 16346
rect 19501 16294 19515 16346
rect 19539 16294 19553 16346
rect 19553 16294 19565 16346
rect 19565 16294 19595 16346
rect 19619 16294 19629 16346
rect 19629 16294 19675 16346
rect 19379 16292 19435 16294
rect 19459 16292 19515 16294
rect 19539 16292 19595 16294
rect 19619 16292 19675 16294
rect 19379 15258 19435 15260
rect 19459 15258 19515 15260
rect 19539 15258 19595 15260
rect 19619 15258 19675 15260
rect 19379 15206 19425 15258
rect 19425 15206 19435 15258
rect 19459 15206 19489 15258
rect 19489 15206 19501 15258
rect 19501 15206 19515 15258
rect 19539 15206 19553 15258
rect 19553 15206 19565 15258
rect 19565 15206 19595 15258
rect 19619 15206 19629 15258
rect 19629 15206 19675 15258
rect 19379 15204 19435 15206
rect 19459 15204 19515 15206
rect 19539 15204 19595 15206
rect 19619 15204 19675 15206
rect 19379 14170 19435 14172
rect 19459 14170 19515 14172
rect 19539 14170 19595 14172
rect 19619 14170 19675 14172
rect 19379 14118 19425 14170
rect 19425 14118 19435 14170
rect 19459 14118 19489 14170
rect 19489 14118 19501 14170
rect 19501 14118 19515 14170
rect 19539 14118 19553 14170
rect 19553 14118 19565 14170
rect 19565 14118 19595 14170
rect 19619 14118 19629 14170
rect 19629 14118 19675 14170
rect 19379 14116 19435 14118
rect 19459 14116 19515 14118
rect 19539 14116 19595 14118
rect 19619 14116 19675 14118
rect 19338 13776 19394 13832
rect 18970 13368 19026 13424
rect 19706 13776 19762 13832
rect 19379 13082 19435 13084
rect 19459 13082 19515 13084
rect 19539 13082 19595 13084
rect 19619 13082 19675 13084
rect 19379 13030 19425 13082
rect 19425 13030 19435 13082
rect 19459 13030 19489 13082
rect 19489 13030 19501 13082
rect 19501 13030 19515 13082
rect 19539 13030 19553 13082
rect 19553 13030 19565 13082
rect 19565 13030 19595 13082
rect 19619 13030 19629 13082
rect 19629 13030 19675 13082
rect 19379 13028 19435 13030
rect 19459 13028 19515 13030
rect 19539 13028 19595 13030
rect 19619 13028 19675 13030
rect 19982 16768 20038 16824
rect 20350 15408 20406 15464
rect 20074 12724 20076 12744
rect 20076 12724 20128 12744
rect 20128 12724 20130 12744
rect 20074 12688 20130 12724
rect 19379 11994 19435 11996
rect 19459 11994 19515 11996
rect 19539 11994 19595 11996
rect 19619 11994 19675 11996
rect 19379 11942 19425 11994
rect 19425 11942 19435 11994
rect 19459 11942 19489 11994
rect 19489 11942 19501 11994
rect 19501 11942 19515 11994
rect 19539 11942 19553 11994
rect 19553 11942 19565 11994
rect 19565 11942 19595 11994
rect 19619 11942 19629 11994
rect 19629 11942 19675 11994
rect 19379 11940 19435 11942
rect 19459 11940 19515 11942
rect 19539 11940 19595 11942
rect 19619 11940 19675 11942
rect 19379 10906 19435 10908
rect 19459 10906 19515 10908
rect 19539 10906 19595 10908
rect 19619 10906 19675 10908
rect 19379 10854 19425 10906
rect 19425 10854 19435 10906
rect 19459 10854 19489 10906
rect 19489 10854 19501 10906
rect 19501 10854 19515 10906
rect 19539 10854 19553 10906
rect 19553 10854 19565 10906
rect 19565 10854 19595 10906
rect 19619 10854 19629 10906
rect 19629 10854 19675 10906
rect 19379 10852 19435 10854
rect 19459 10852 19515 10854
rect 19539 10852 19595 10854
rect 19619 10852 19675 10854
rect 19379 9818 19435 9820
rect 19459 9818 19515 9820
rect 19539 9818 19595 9820
rect 19619 9818 19675 9820
rect 19379 9766 19425 9818
rect 19425 9766 19435 9818
rect 19459 9766 19489 9818
rect 19489 9766 19501 9818
rect 19501 9766 19515 9818
rect 19539 9766 19553 9818
rect 19553 9766 19565 9818
rect 19565 9766 19595 9818
rect 19619 9766 19629 9818
rect 19629 9766 19675 9818
rect 19379 9764 19435 9766
rect 19459 9764 19515 9766
rect 19539 9764 19595 9766
rect 19619 9764 19675 9766
rect 19379 8730 19435 8732
rect 19459 8730 19515 8732
rect 19539 8730 19595 8732
rect 19619 8730 19675 8732
rect 19379 8678 19425 8730
rect 19425 8678 19435 8730
rect 19459 8678 19489 8730
rect 19489 8678 19501 8730
rect 19501 8678 19515 8730
rect 19539 8678 19553 8730
rect 19553 8678 19565 8730
rect 19565 8678 19595 8730
rect 19619 8678 19629 8730
rect 19629 8678 19675 8730
rect 19379 8676 19435 8678
rect 19459 8676 19515 8678
rect 19539 8676 19595 8678
rect 19619 8676 19675 8678
rect 18878 7656 18934 7712
rect 18602 6840 18658 6896
rect 18970 6432 19026 6488
rect 19379 7642 19435 7644
rect 19459 7642 19515 7644
rect 19539 7642 19595 7644
rect 19619 7642 19675 7644
rect 19379 7590 19425 7642
rect 19425 7590 19435 7642
rect 19459 7590 19489 7642
rect 19489 7590 19501 7642
rect 19501 7590 19515 7642
rect 19539 7590 19553 7642
rect 19553 7590 19565 7642
rect 19565 7590 19595 7642
rect 19619 7590 19629 7642
rect 19629 7590 19675 7642
rect 19379 7588 19435 7590
rect 19459 7588 19515 7590
rect 19539 7588 19595 7590
rect 19619 7588 19675 7590
rect 19246 6704 19302 6760
rect 19379 6554 19435 6556
rect 19459 6554 19515 6556
rect 19539 6554 19595 6556
rect 19619 6554 19675 6556
rect 19379 6502 19425 6554
rect 19425 6502 19435 6554
rect 19459 6502 19489 6554
rect 19489 6502 19501 6554
rect 19501 6502 19515 6554
rect 19539 6502 19553 6554
rect 19553 6502 19565 6554
rect 19565 6502 19595 6554
rect 19619 6502 19629 6554
rect 19629 6502 19675 6554
rect 19379 6500 19435 6502
rect 19459 6500 19515 6502
rect 19539 6500 19595 6502
rect 19619 6500 19675 6502
rect 19379 5466 19435 5468
rect 19459 5466 19515 5468
rect 19539 5466 19595 5468
rect 19619 5466 19675 5468
rect 19379 5414 19425 5466
rect 19425 5414 19435 5466
rect 19459 5414 19489 5466
rect 19489 5414 19501 5466
rect 19501 5414 19515 5466
rect 19539 5414 19553 5466
rect 19553 5414 19565 5466
rect 19565 5414 19595 5466
rect 19619 5414 19629 5466
rect 19629 5414 19675 5466
rect 19379 5412 19435 5414
rect 19459 5412 19515 5414
rect 19539 5412 19595 5414
rect 19619 5412 19675 5414
rect 18878 3712 18934 3768
rect 18970 3440 19026 3496
rect 19246 5072 19302 5128
rect 19379 4378 19435 4380
rect 19459 4378 19515 4380
rect 19539 4378 19595 4380
rect 19619 4378 19675 4380
rect 19379 4326 19425 4378
rect 19425 4326 19435 4378
rect 19459 4326 19489 4378
rect 19489 4326 19501 4378
rect 19501 4326 19515 4378
rect 19539 4326 19553 4378
rect 19553 4326 19565 4378
rect 19565 4326 19595 4378
rect 19619 4326 19629 4378
rect 19629 4326 19675 4378
rect 19379 4324 19435 4326
rect 19459 4324 19515 4326
rect 19539 4324 19595 4326
rect 19619 4324 19675 4326
rect 19379 3290 19435 3292
rect 19459 3290 19515 3292
rect 19539 3290 19595 3292
rect 19619 3290 19675 3292
rect 19379 3238 19425 3290
rect 19425 3238 19435 3290
rect 19459 3238 19489 3290
rect 19489 3238 19501 3290
rect 19501 3238 19515 3290
rect 19539 3238 19553 3290
rect 19553 3238 19565 3290
rect 19565 3238 19595 3290
rect 19619 3238 19629 3290
rect 19629 3238 19675 3290
rect 19379 3236 19435 3238
rect 19459 3236 19515 3238
rect 19539 3236 19595 3238
rect 19619 3236 19675 3238
rect 19338 3052 19394 3088
rect 19338 3032 19340 3052
rect 19340 3032 19392 3052
rect 19392 3032 19394 3052
rect 19379 2202 19435 2204
rect 19459 2202 19515 2204
rect 19539 2202 19595 2204
rect 19619 2202 19675 2204
rect 19379 2150 19425 2202
rect 19425 2150 19435 2202
rect 19459 2150 19489 2202
rect 19489 2150 19501 2202
rect 19501 2150 19515 2202
rect 19539 2150 19553 2202
rect 19553 2150 19565 2202
rect 19565 2150 19595 2202
rect 19619 2150 19629 2202
rect 19629 2150 19675 2202
rect 19379 2148 19435 2150
rect 19459 2148 19515 2150
rect 19539 2148 19595 2150
rect 19619 2148 19675 2150
rect 19338 1536 19394 1592
rect 19379 1114 19435 1116
rect 19459 1114 19515 1116
rect 19539 1114 19595 1116
rect 19619 1114 19675 1116
rect 19379 1062 19425 1114
rect 19425 1062 19435 1114
rect 19459 1062 19489 1114
rect 19489 1062 19501 1114
rect 19501 1062 19515 1114
rect 19539 1062 19553 1114
rect 19553 1062 19565 1114
rect 19565 1062 19595 1114
rect 19619 1062 19629 1114
rect 19629 1062 19675 1114
rect 19379 1060 19435 1062
rect 19459 1060 19515 1062
rect 19539 1060 19595 1062
rect 19619 1060 19675 1062
rect 20258 10124 20314 10160
rect 20258 10104 20260 10124
rect 20260 10104 20312 10124
rect 20312 10104 20314 10124
rect 20718 19624 20774 19680
rect 20718 18264 20774 18320
rect 20718 17720 20774 17776
rect 20626 17176 20682 17232
rect 20902 17992 20958 18048
rect 21086 17720 21142 17776
rect 21178 17448 21234 17504
rect 21178 17196 21234 17232
rect 21178 17176 21180 17196
rect 21180 17176 21232 17196
rect 21232 17176 21234 17196
rect 21086 16652 21142 16688
rect 21086 16632 21088 16652
rect 21088 16632 21140 16652
rect 21140 16632 21142 16652
rect 20718 16496 20774 16552
rect 20534 16088 20590 16144
rect 21914 21800 21970 21856
rect 22098 21664 22154 21720
rect 21822 20848 21878 20904
rect 21822 20576 21878 20632
rect 21914 20304 21970 20360
rect 22282 20304 22338 20360
rect 21822 18400 21878 18456
rect 21638 17312 21694 17368
rect 20902 15136 20958 15192
rect 21546 13776 21602 13832
rect 21638 13096 21694 13152
rect 20626 9968 20682 10024
rect 21638 11600 21694 11656
rect 21086 10648 21142 10704
rect 21086 10104 21142 10160
rect 22558 22072 22614 22128
rect 22558 17856 22614 17912
rect 23294 22072 23350 22128
rect 23174 21242 23230 21244
rect 23254 21242 23310 21244
rect 23334 21242 23390 21244
rect 23414 21242 23470 21244
rect 23174 21190 23220 21242
rect 23220 21190 23230 21242
rect 23254 21190 23284 21242
rect 23284 21190 23296 21242
rect 23296 21190 23310 21242
rect 23334 21190 23348 21242
rect 23348 21190 23360 21242
rect 23360 21190 23390 21242
rect 23414 21190 23424 21242
rect 23424 21190 23470 21242
rect 23174 21188 23230 21190
rect 23254 21188 23310 21190
rect 23334 21188 23390 21190
rect 23414 21188 23470 21190
rect 23174 20154 23230 20156
rect 23254 20154 23310 20156
rect 23334 20154 23390 20156
rect 23414 20154 23470 20156
rect 23174 20102 23220 20154
rect 23220 20102 23230 20154
rect 23254 20102 23284 20154
rect 23284 20102 23296 20154
rect 23296 20102 23310 20154
rect 23334 20102 23348 20154
rect 23348 20102 23360 20154
rect 23360 20102 23390 20154
rect 23414 20102 23424 20154
rect 23424 20102 23470 20154
rect 23174 20100 23230 20102
rect 23254 20100 23310 20102
rect 23334 20100 23390 20102
rect 23414 20100 23470 20102
rect 23386 19896 23442 19952
rect 23570 19760 23626 19816
rect 23754 22208 23810 22244
rect 25042 22092 25098 22128
rect 25042 22072 25044 22092
rect 25044 22072 25096 22092
rect 25096 22072 25098 22092
rect 23754 21800 23810 21856
rect 24674 21664 24730 21720
rect 26330 21936 26386 21992
rect 23938 20848 23994 20904
rect 23846 19896 23902 19952
rect 23846 19624 23902 19680
rect 23174 19066 23230 19068
rect 23254 19066 23310 19068
rect 23334 19066 23390 19068
rect 23414 19066 23470 19068
rect 23174 19014 23220 19066
rect 23220 19014 23230 19066
rect 23254 19014 23284 19066
rect 23284 19014 23296 19066
rect 23296 19014 23310 19066
rect 23334 19014 23348 19066
rect 23348 19014 23360 19066
rect 23360 19014 23390 19066
rect 23414 19014 23424 19066
rect 23424 19014 23470 19066
rect 23174 19012 23230 19014
rect 23254 19012 23310 19014
rect 23334 19012 23390 19014
rect 23414 19012 23470 19014
rect 23386 18808 23442 18864
rect 23662 18400 23718 18456
rect 23386 18128 23442 18184
rect 23570 18148 23626 18184
rect 23570 18128 23572 18148
rect 23572 18128 23624 18148
rect 23624 18128 23626 18148
rect 23174 17978 23230 17980
rect 23254 17978 23310 17980
rect 23334 17978 23390 17980
rect 23414 17978 23470 17980
rect 23174 17926 23220 17978
rect 23220 17926 23230 17978
rect 23254 17926 23284 17978
rect 23284 17926 23296 17978
rect 23296 17926 23310 17978
rect 23334 17926 23348 17978
rect 23348 17926 23360 17978
rect 23360 17926 23390 17978
rect 23414 17926 23424 17978
rect 23424 17926 23470 17978
rect 23174 17924 23230 17926
rect 23254 17924 23310 17926
rect 23334 17924 23390 17926
rect 23414 17924 23470 17926
rect 22742 16768 22798 16824
rect 21914 13912 21970 13968
rect 21914 12688 21970 12744
rect 24858 20576 24914 20632
rect 24214 18844 24216 18864
rect 24216 18844 24268 18864
rect 24268 18844 24270 18864
rect 24214 18808 24270 18844
rect 24490 18400 24546 18456
rect 24398 18300 24400 18320
rect 24400 18300 24452 18320
rect 24452 18300 24454 18320
rect 24398 18264 24454 18300
rect 23018 16904 23074 16960
rect 23174 16890 23230 16892
rect 23254 16890 23310 16892
rect 23334 16890 23390 16892
rect 23414 16890 23470 16892
rect 23174 16838 23220 16890
rect 23220 16838 23230 16890
rect 23254 16838 23284 16890
rect 23284 16838 23296 16890
rect 23296 16838 23310 16890
rect 23334 16838 23348 16890
rect 23348 16838 23360 16890
rect 23360 16838 23390 16890
rect 23414 16838 23424 16890
rect 23424 16838 23470 16890
rect 23174 16836 23230 16838
rect 23254 16836 23310 16838
rect 23334 16836 23390 16838
rect 23414 16836 23470 16838
rect 24030 16496 24086 16552
rect 23174 15802 23230 15804
rect 23254 15802 23310 15804
rect 23334 15802 23390 15804
rect 23414 15802 23470 15804
rect 23174 15750 23220 15802
rect 23220 15750 23230 15802
rect 23254 15750 23284 15802
rect 23284 15750 23296 15802
rect 23296 15750 23310 15802
rect 23334 15750 23348 15802
rect 23348 15750 23360 15802
rect 23360 15750 23390 15802
rect 23414 15750 23424 15802
rect 23424 15750 23470 15802
rect 23174 15748 23230 15750
rect 23254 15748 23310 15750
rect 23334 15748 23390 15750
rect 23414 15748 23470 15750
rect 22650 13912 22706 13968
rect 22926 13912 22982 13968
rect 22374 13368 22430 13424
rect 23174 14714 23230 14716
rect 23254 14714 23310 14716
rect 23334 14714 23390 14716
rect 23414 14714 23470 14716
rect 23174 14662 23220 14714
rect 23220 14662 23230 14714
rect 23254 14662 23284 14714
rect 23284 14662 23296 14714
rect 23296 14662 23310 14714
rect 23334 14662 23348 14714
rect 23348 14662 23360 14714
rect 23360 14662 23390 14714
rect 23414 14662 23424 14714
rect 23424 14662 23470 14714
rect 23174 14660 23230 14662
rect 23254 14660 23310 14662
rect 23334 14660 23390 14662
rect 23414 14660 23470 14662
rect 23846 15156 23902 15192
rect 23846 15136 23848 15156
rect 23848 15136 23900 15156
rect 23900 15136 23902 15156
rect 23846 14456 23902 14512
rect 24766 17856 24822 17912
rect 24582 17040 24638 17096
rect 25134 19252 25136 19272
rect 25136 19252 25188 19272
rect 25188 19252 25190 19272
rect 25134 19216 25190 19252
rect 25318 17720 25374 17776
rect 25226 17312 25282 17368
rect 25318 16124 25320 16144
rect 25320 16124 25372 16144
rect 25372 16124 25374 16144
rect 25318 16088 25374 16124
rect 24766 15816 24822 15872
rect 24490 15680 24546 15736
rect 24398 14592 24454 14648
rect 24398 13932 24454 13968
rect 24398 13912 24400 13932
rect 24400 13912 24452 13932
rect 24452 13912 24454 13932
rect 23570 13640 23626 13696
rect 23174 13626 23230 13628
rect 23254 13626 23310 13628
rect 23334 13626 23390 13628
rect 23414 13626 23470 13628
rect 23174 13574 23220 13626
rect 23220 13574 23230 13626
rect 23254 13574 23284 13626
rect 23284 13574 23296 13626
rect 23296 13574 23310 13626
rect 23334 13574 23348 13626
rect 23348 13574 23360 13626
rect 23360 13574 23390 13626
rect 23414 13574 23424 13626
rect 23424 13574 23470 13626
rect 23174 13572 23230 13574
rect 23254 13572 23310 13574
rect 23334 13572 23390 13574
rect 23414 13572 23470 13574
rect 23938 13524 23994 13560
rect 23938 13504 23940 13524
rect 23940 13504 23992 13524
rect 23992 13504 23994 13524
rect 22926 13096 22982 13152
rect 22834 12824 22890 12880
rect 24398 13368 24454 13424
rect 23754 12724 23756 12744
rect 23756 12724 23808 12744
rect 23808 12724 23810 12744
rect 23754 12688 23810 12724
rect 23174 12538 23230 12540
rect 23254 12538 23310 12540
rect 23334 12538 23390 12540
rect 23414 12538 23470 12540
rect 23174 12486 23220 12538
rect 23220 12486 23230 12538
rect 23254 12486 23284 12538
rect 23284 12486 23296 12538
rect 23296 12486 23310 12538
rect 23334 12486 23348 12538
rect 23348 12486 23360 12538
rect 23360 12486 23390 12538
rect 23414 12486 23424 12538
rect 23424 12486 23470 12538
rect 23174 12484 23230 12486
rect 23254 12484 23310 12486
rect 23334 12484 23390 12486
rect 23414 12484 23470 12486
rect 20626 7248 20682 7304
rect 20166 5208 20222 5264
rect 21178 8608 21234 8664
rect 20994 8336 21050 8392
rect 21270 8336 21326 8392
rect 20626 5788 20628 5808
rect 20628 5788 20680 5808
rect 20680 5788 20682 5808
rect 20626 5752 20682 5788
rect 20626 5636 20682 5672
rect 20626 5616 20628 5636
rect 20628 5616 20680 5636
rect 20680 5616 20682 5636
rect 22006 8492 22062 8528
rect 22006 8472 22008 8492
rect 22008 8472 22060 8492
rect 22060 8472 22062 8492
rect 20994 6160 21050 6216
rect 22190 9968 22246 10024
rect 22466 9832 22522 9888
rect 23174 11450 23230 11452
rect 23254 11450 23310 11452
rect 23334 11450 23390 11452
rect 23414 11450 23470 11452
rect 23174 11398 23220 11450
rect 23220 11398 23230 11450
rect 23254 11398 23284 11450
rect 23284 11398 23296 11450
rect 23296 11398 23310 11450
rect 23334 11398 23348 11450
rect 23348 11398 23360 11450
rect 23360 11398 23390 11450
rect 23414 11398 23424 11450
rect 23424 11398 23470 11450
rect 23174 11396 23230 11398
rect 23254 11396 23310 11398
rect 23334 11396 23390 11398
rect 23414 11396 23470 11398
rect 23478 10512 23534 10568
rect 23174 10362 23230 10364
rect 23254 10362 23310 10364
rect 23334 10362 23390 10364
rect 23414 10362 23470 10364
rect 23174 10310 23220 10362
rect 23220 10310 23230 10362
rect 23254 10310 23284 10362
rect 23284 10310 23296 10362
rect 23296 10310 23310 10362
rect 23334 10310 23348 10362
rect 23348 10310 23360 10362
rect 23360 10310 23390 10362
rect 23414 10310 23424 10362
rect 23424 10310 23470 10362
rect 23174 10308 23230 10310
rect 23254 10308 23310 10310
rect 23334 10308 23390 10310
rect 23414 10308 23470 10310
rect 23478 9460 23480 9480
rect 23480 9460 23532 9480
rect 23532 9460 23534 9480
rect 23478 9424 23534 9460
rect 23570 9288 23626 9344
rect 23174 9274 23230 9276
rect 23254 9274 23310 9276
rect 23334 9274 23390 9276
rect 23414 9274 23470 9276
rect 23174 9222 23220 9274
rect 23220 9222 23230 9274
rect 23254 9222 23284 9274
rect 23284 9222 23296 9274
rect 23296 9222 23310 9274
rect 23334 9222 23348 9274
rect 23348 9222 23360 9274
rect 23360 9222 23390 9274
rect 23414 9222 23424 9274
rect 23424 9222 23470 9274
rect 23174 9220 23230 9222
rect 23254 9220 23310 9222
rect 23334 9220 23390 9222
rect 23414 9220 23470 9222
rect 23754 9560 23810 9616
rect 23018 8608 23074 8664
rect 23174 8186 23230 8188
rect 23254 8186 23310 8188
rect 23334 8186 23390 8188
rect 23414 8186 23470 8188
rect 23174 8134 23220 8186
rect 23220 8134 23230 8186
rect 23254 8134 23284 8186
rect 23284 8134 23296 8186
rect 23296 8134 23310 8186
rect 23334 8134 23348 8186
rect 23348 8134 23360 8186
rect 23360 8134 23390 8186
rect 23414 8134 23424 8186
rect 23424 8134 23470 8186
rect 23174 8132 23230 8134
rect 23254 8132 23310 8134
rect 23334 8132 23390 8134
rect 23414 8132 23470 8134
rect 23174 7098 23230 7100
rect 23254 7098 23310 7100
rect 23334 7098 23390 7100
rect 23414 7098 23470 7100
rect 23174 7046 23220 7098
rect 23220 7046 23230 7098
rect 23254 7046 23284 7098
rect 23284 7046 23296 7098
rect 23296 7046 23310 7098
rect 23334 7046 23348 7098
rect 23348 7046 23360 7098
rect 23360 7046 23390 7098
rect 23414 7046 23424 7098
rect 23424 7046 23470 7098
rect 23174 7044 23230 7046
rect 23254 7044 23310 7046
rect 23334 7044 23390 7046
rect 23414 7044 23470 7046
rect 24214 11600 24270 11656
rect 24030 8880 24086 8936
rect 24122 7404 24178 7440
rect 24122 7384 24124 7404
rect 24124 7384 24176 7404
rect 24176 7384 24178 7404
rect 25962 21684 26018 21720
rect 25962 21664 25964 21684
rect 25964 21664 26016 21684
rect 26016 21664 26018 21684
rect 26146 21120 26202 21176
rect 26238 20848 26294 20904
rect 26969 21786 27025 21788
rect 27049 21786 27105 21788
rect 27129 21786 27185 21788
rect 27209 21786 27265 21788
rect 26969 21734 27015 21786
rect 27015 21734 27025 21786
rect 27049 21734 27079 21786
rect 27079 21734 27091 21786
rect 27091 21734 27105 21786
rect 27129 21734 27143 21786
rect 27143 21734 27155 21786
rect 27155 21734 27185 21786
rect 27209 21734 27219 21786
rect 27219 21734 27265 21786
rect 26969 21732 27025 21734
rect 27049 21732 27105 21734
rect 27129 21732 27185 21734
rect 27209 21732 27265 21734
rect 26698 21528 26754 21584
rect 27802 21392 27858 21448
rect 26238 19488 26294 19544
rect 26054 19352 26110 19408
rect 26238 17992 26294 18048
rect 26054 17720 26110 17776
rect 26054 17448 26110 17504
rect 25870 16088 25926 16144
rect 26969 20698 27025 20700
rect 27049 20698 27105 20700
rect 27129 20698 27185 20700
rect 27209 20698 27265 20700
rect 26969 20646 27015 20698
rect 27015 20646 27025 20698
rect 27049 20646 27079 20698
rect 27079 20646 27091 20698
rect 27091 20646 27105 20698
rect 27129 20646 27143 20698
rect 27143 20646 27155 20698
rect 27155 20646 27185 20698
rect 27209 20646 27219 20698
rect 27219 20646 27265 20698
rect 26969 20644 27025 20646
rect 27049 20644 27105 20646
rect 27129 20644 27185 20646
rect 27209 20644 27265 20646
rect 28170 20440 28226 20496
rect 27618 19916 27674 19952
rect 27618 19896 27620 19916
rect 27620 19896 27672 19916
rect 27672 19896 27674 19916
rect 26969 19610 27025 19612
rect 27049 19610 27105 19612
rect 27129 19610 27185 19612
rect 27209 19610 27265 19612
rect 26969 19558 27015 19610
rect 27015 19558 27025 19610
rect 27049 19558 27079 19610
rect 27079 19558 27091 19610
rect 27091 19558 27105 19610
rect 27129 19558 27143 19610
rect 27143 19558 27155 19610
rect 27155 19558 27185 19610
rect 27209 19558 27219 19610
rect 27219 19558 27265 19610
rect 26969 19556 27025 19558
rect 27049 19556 27105 19558
rect 27129 19556 27185 19558
rect 27209 19556 27265 19558
rect 27250 19372 27306 19408
rect 27250 19352 27252 19372
rect 27252 19352 27304 19372
rect 27304 19352 27306 19372
rect 26606 17856 26662 17912
rect 25686 14456 25742 14512
rect 26330 14900 26332 14920
rect 26332 14900 26384 14920
rect 26384 14900 26386 14920
rect 26330 14864 26386 14900
rect 25962 12144 26018 12200
rect 25410 11736 25466 11792
rect 22558 6704 22614 6760
rect 21822 5616 21878 5672
rect 22006 5616 22062 5672
rect 20350 2372 20406 2408
rect 20350 2352 20352 2372
rect 20352 2352 20404 2372
rect 20404 2352 20406 2372
rect 20994 1672 21050 1728
rect 22742 5752 22798 5808
rect 23174 6010 23230 6012
rect 23254 6010 23310 6012
rect 23334 6010 23390 6012
rect 23414 6010 23470 6012
rect 23174 5958 23220 6010
rect 23220 5958 23230 6010
rect 23254 5958 23284 6010
rect 23284 5958 23296 6010
rect 23296 5958 23310 6010
rect 23334 5958 23348 6010
rect 23348 5958 23360 6010
rect 23360 5958 23390 6010
rect 23414 5958 23424 6010
rect 23424 5958 23470 6010
rect 23174 5956 23230 5958
rect 23254 5956 23310 5958
rect 23334 5956 23390 5958
rect 23414 5956 23470 5958
rect 23174 4922 23230 4924
rect 23254 4922 23310 4924
rect 23334 4922 23390 4924
rect 23414 4922 23470 4924
rect 23174 4870 23220 4922
rect 23220 4870 23230 4922
rect 23254 4870 23284 4922
rect 23284 4870 23296 4922
rect 23296 4870 23310 4922
rect 23334 4870 23348 4922
rect 23348 4870 23360 4922
rect 23360 4870 23390 4922
rect 23414 4870 23424 4922
rect 23424 4870 23470 4922
rect 23174 4868 23230 4870
rect 23254 4868 23310 4870
rect 23334 4868 23390 4870
rect 23414 4868 23470 4870
rect 24122 5888 24178 5944
rect 24674 9560 24730 9616
rect 25962 11736 26018 11792
rect 26146 9424 26202 9480
rect 25410 8336 25466 8392
rect 21638 2388 21640 2408
rect 21640 2388 21692 2408
rect 21692 2388 21694 2408
rect 21638 2352 21694 2388
rect 22926 3848 22982 3904
rect 23174 3834 23230 3836
rect 23254 3834 23310 3836
rect 23334 3834 23390 3836
rect 23414 3834 23470 3836
rect 23174 3782 23220 3834
rect 23220 3782 23230 3834
rect 23254 3782 23284 3834
rect 23284 3782 23296 3834
rect 23296 3782 23310 3834
rect 23334 3782 23348 3834
rect 23348 3782 23360 3834
rect 23360 3782 23390 3834
rect 23414 3782 23424 3834
rect 23424 3782 23470 3834
rect 23174 3780 23230 3782
rect 23254 3780 23310 3782
rect 23334 3780 23390 3782
rect 23414 3780 23470 3782
rect 22926 3032 22982 3088
rect 23174 2746 23230 2748
rect 23254 2746 23310 2748
rect 23334 2746 23390 2748
rect 23414 2746 23470 2748
rect 23174 2694 23220 2746
rect 23220 2694 23230 2746
rect 23254 2694 23284 2746
rect 23284 2694 23296 2746
rect 23296 2694 23310 2746
rect 23334 2694 23348 2746
rect 23348 2694 23360 2746
rect 23360 2694 23390 2746
rect 23414 2694 23424 2746
rect 23424 2694 23470 2746
rect 23174 2692 23230 2694
rect 23254 2692 23310 2694
rect 23334 2692 23390 2694
rect 23414 2692 23470 2694
rect 21638 1672 21694 1728
rect 21362 1128 21418 1184
rect 23386 2216 23442 2272
rect 22834 2080 22890 2136
rect 22834 1536 22890 1592
rect 24030 2644 24086 2680
rect 24030 2624 24032 2644
rect 24032 2624 24084 2644
rect 24084 2624 24086 2644
rect 24858 6160 24914 6216
rect 23174 1658 23230 1660
rect 23254 1658 23310 1660
rect 23334 1658 23390 1660
rect 23414 1658 23470 1660
rect 23174 1606 23220 1658
rect 23220 1606 23230 1658
rect 23254 1606 23284 1658
rect 23284 1606 23296 1658
rect 23296 1606 23310 1658
rect 23334 1606 23348 1658
rect 23348 1606 23360 1658
rect 23360 1606 23390 1658
rect 23414 1606 23424 1658
rect 23424 1606 23470 1658
rect 23174 1604 23230 1606
rect 23254 1604 23310 1606
rect 23334 1604 23390 1606
rect 23414 1604 23470 1606
rect 23754 1672 23810 1728
rect 23754 1420 23810 1456
rect 23754 1400 23756 1420
rect 23756 1400 23808 1420
rect 23808 1400 23810 1420
rect 23478 856 23534 912
rect 23938 1420 23994 1456
rect 23938 1400 23940 1420
rect 23940 1400 23992 1420
rect 23992 1400 23994 1420
rect 23174 570 23230 572
rect 23254 570 23310 572
rect 23334 570 23390 572
rect 23414 570 23470 572
rect 23174 518 23220 570
rect 23220 518 23230 570
rect 23254 518 23284 570
rect 23284 518 23296 570
rect 23296 518 23310 570
rect 23334 518 23348 570
rect 23348 518 23360 570
rect 23360 518 23390 570
rect 23414 518 23424 570
rect 23424 518 23470 570
rect 23174 516 23230 518
rect 23254 516 23310 518
rect 23334 516 23390 518
rect 23414 516 23470 518
rect 24490 2624 24546 2680
rect 26146 9036 26202 9072
rect 26146 9016 26148 9036
rect 26148 9016 26200 9036
rect 26200 9016 26202 9036
rect 26146 7384 26202 7440
rect 26969 18522 27025 18524
rect 27049 18522 27105 18524
rect 27129 18522 27185 18524
rect 27209 18522 27265 18524
rect 26969 18470 27015 18522
rect 27015 18470 27025 18522
rect 27049 18470 27079 18522
rect 27079 18470 27091 18522
rect 27091 18470 27105 18522
rect 27129 18470 27143 18522
rect 27143 18470 27155 18522
rect 27155 18470 27185 18522
rect 27209 18470 27219 18522
rect 27219 18470 27265 18522
rect 26969 18468 27025 18470
rect 27049 18468 27105 18470
rect 27129 18468 27185 18470
rect 27209 18468 27265 18470
rect 26969 17434 27025 17436
rect 27049 17434 27105 17436
rect 27129 17434 27185 17436
rect 27209 17434 27265 17436
rect 26969 17382 27015 17434
rect 27015 17382 27025 17434
rect 27049 17382 27079 17434
rect 27079 17382 27091 17434
rect 27091 17382 27105 17434
rect 27129 17382 27143 17434
rect 27143 17382 27155 17434
rect 27155 17382 27185 17434
rect 27209 17382 27219 17434
rect 27219 17382 27265 17434
rect 26969 17380 27025 17382
rect 27049 17380 27105 17382
rect 27129 17380 27185 17382
rect 27209 17380 27265 17382
rect 26969 16346 27025 16348
rect 27049 16346 27105 16348
rect 27129 16346 27185 16348
rect 27209 16346 27265 16348
rect 26969 16294 27015 16346
rect 27015 16294 27025 16346
rect 27049 16294 27079 16346
rect 27079 16294 27091 16346
rect 27091 16294 27105 16346
rect 27129 16294 27143 16346
rect 27143 16294 27155 16346
rect 27155 16294 27185 16346
rect 27209 16294 27219 16346
rect 27219 16294 27265 16346
rect 26969 16292 27025 16294
rect 27049 16292 27105 16294
rect 27129 16292 27185 16294
rect 27209 16292 27265 16294
rect 26974 16088 27030 16144
rect 26969 15258 27025 15260
rect 27049 15258 27105 15260
rect 27129 15258 27185 15260
rect 27209 15258 27265 15260
rect 26969 15206 27015 15258
rect 27015 15206 27025 15258
rect 27049 15206 27079 15258
rect 27079 15206 27091 15258
rect 27091 15206 27105 15258
rect 27129 15206 27143 15258
rect 27143 15206 27155 15258
rect 27155 15206 27185 15258
rect 27209 15206 27219 15258
rect 27219 15206 27265 15258
rect 26969 15204 27025 15206
rect 27049 15204 27105 15206
rect 27129 15204 27185 15206
rect 27209 15204 27265 15206
rect 27250 14320 27306 14376
rect 26969 14170 27025 14172
rect 27049 14170 27105 14172
rect 27129 14170 27185 14172
rect 27209 14170 27265 14172
rect 26969 14118 27015 14170
rect 27015 14118 27025 14170
rect 27049 14118 27079 14170
rect 27079 14118 27091 14170
rect 27091 14118 27105 14170
rect 27129 14118 27143 14170
rect 27143 14118 27155 14170
rect 27155 14118 27185 14170
rect 27209 14118 27219 14170
rect 27219 14118 27265 14170
rect 26969 14116 27025 14118
rect 27049 14116 27105 14118
rect 27129 14116 27185 14118
rect 27209 14116 27265 14118
rect 27434 16360 27490 16416
rect 27618 18128 27674 18184
rect 27710 16904 27766 16960
rect 27710 15680 27766 15736
rect 27618 15272 27674 15328
rect 26882 13504 26938 13560
rect 26969 13082 27025 13084
rect 27049 13082 27105 13084
rect 27129 13082 27185 13084
rect 27209 13082 27265 13084
rect 26969 13030 27015 13082
rect 27015 13030 27025 13082
rect 27049 13030 27079 13082
rect 27079 13030 27091 13082
rect 27091 13030 27105 13082
rect 27129 13030 27143 13082
rect 27143 13030 27155 13082
rect 27155 13030 27185 13082
rect 27209 13030 27219 13082
rect 27219 13030 27265 13082
rect 26969 13028 27025 13030
rect 27049 13028 27105 13030
rect 27129 13028 27185 13030
rect 27209 13028 27265 13030
rect 27526 12824 27582 12880
rect 27158 12416 27214 12472
rect 26330 11056 26386 11112
rect 26514 8880 26570 8936
rect 18234 176 18290 232
rect 25502 2216 25558 2272
rect 25318 1672 25374 1728
rect 26969 11994 27025 11996
rect 27049 11994 27105 11996
rect 27129 11994 27185 11996
rect 27209 11994 27265 11996
rect 26969 11942 27015 11994
rect 27015 11942 27025 11994
rect 27049 11942 27079 11994
rect 27079 11942 27091 11994
rect 27091 11942 27105 11994
rect 27129 11942 27143 11994
rect 27143 11942 27155 11994
rect 27155 11942 27185 11994
rect 27209 11942 27219 11994
rect 27219 11942 27265 11994
rect 26969 11940 27025 11942
rect 27049 11940 27105 11942
rect 27129 11940 27185 11942
rect 27209 11940 27265 11942
rect 26969 10906 27025 10908
rect 27049 10906 27105 10908
rect 27129 10906 27185 10908
rect 27209 10906 27265 10908
rect 26969 10854 27015 10906
rect 27015 10854 27025 10906
rect 27049 10854 27079 10906
rect 27079 10854 27091 10906
rect 27091 10854 27105 10906
rect 27129 10854 27143 10906
rect 27143 10854 27155 10906
rect 27155 10854 27185 10906
rect 27209 10854 27219 10906
rect 27219 10854 27265 10906
rect 26969 10852 27025 10854
rect 27049 10852 27105 10854
rect 27129 10852 27185 10854
rect 27209 10852 27265 10854
rect 26969 9818 27025 9820
rect 27049 9818 27105 9820
rect 27129 9818 27185 9820
rect 27209 9818 27265 9820
rect 26969 9766 27015 9818
rect 27015 9766 27025 9818
rect 27049 9766 27079 9818
rect 27079 9766 27091 9818
rect 27091 9766 27105 9818
rect 27129 9766 27143 9818
rect 27143 9766 27155 9818
rect 27155 9766 27185 9818
rect 27209 9766 27219 9818
rect 27219 9766 27265 9818
rect 26969 9764 27025 9766
rect 27049 9764 27105 9766
rect 27129 9764 27185 9766
rect 27209 9764 27265 9766
rect 26974 9016 27030 9072
rect 26969 8730 27025 8732
rect 27049 8730 27105 8732
rect 27129 8730 27185 8732
rect 27209 8730 27265 8732
rect 26969 8678 27015 8730
rect 27015 8678 27025 8730
rect 27049 8678 27079 8730
rect 27079 8678 27091 8730
rect 27091 8678 27105 8730
rect 27129 8678 27143 8730
rect 27143 8678 27155 8730
rect 27155 8678 27185 8730
rect 27209 8678 27219 8730
rect 27219 8678 27265 8730
rect 26969 8676 27025 8678
rect 27049 8676 27105 8678
rect 27129 8676 27185 8678
rect 27209 8676 27265 8678
rect 27894 18844 27896 18864
rect 27896 18844 27948 18864
rect 27948 18844 27950 18864
rect 27894 18808 27950 18844
rect 27986 16668 27988 16688
rect 27988 16668 28040 16688
rect 28040 16668 28042 16688
rect 27986 16632 28042 16668
rect 27894 15680 27950 15736
rect 27894 15408 27950 15464
rect 28354 18400 28410 18456
rect 28354 17176 28410 17232
rect 28262 16496 28318 16552
rect 28538 16496 28594 16552
rect 28262 15816 28318 15872
rect 28170 15272 28226 15328
rect 27434 10104 27490 10160
rect 28538 15544 28594 15600
rect 28446 14592 28502 14648
rect 26969 7642 27025 7644
rect 27049 7642 27105 7644
rect 27129 7642 27185 7644
rect 27209 7642 27265 7644
rect 26969 7590 27015 7642
rect 27015 7590 27025 7642
rect 27049 7590 27079 7642
rect 27079 7590 27091 7642
rect 27091 7590 27105 7642
rect 27129 7590 27143 7642
rect 27143 7590 27155 7642
rect 27155 7590 27185 7642
rect 27209 7590 27219 7642
rect 27219 7590 27265 7642
rect 26969 7588 27025 7590
rect 27049 7588 27105 7590
rect 27129 7588 27185 7590
rect 27209 7588 27265 7590
rect 26974 6840 27030 6896
rect 26969 6554 27025 6556
rect 27049 6554 27105 6556
rect 27129 6554 27185 6556
rect 27209 6554 27265 6556
rect 26969 6502 27015 6554
rect 27015 6502 27025 6554
rect 27049 6502 27079 6554
rect 27079 6502 27091 6554
rect 27091 6502 27105 6554
rect 27129 6502 27143 6554
rect 27143 6502 27155 6554
rect 27155 6502 27185 6554
rect 27209 6502 27219 6554
rect 27219 6502 27265 6554
rect 26969 6500 27025 6502
rect 27049 6500 27105 6502
rect 27129 6500 27185 6502
rect 27209 6500 27265 6502
rect 26790 5888 26846 5944
rect 26969 5466 27025 5468
rect 27049 5466 27105 5468
rect 27129 5466 27185 5468
rect 27209 5466 27265 5468
rect 26969 5414 27015 5466
rect 27015 5414 27025 5466
rect 27049 5414 27079 5466
rect 27079 5414 27091 5466
rect 27091 5414 27105 5466
rect 27129 5414 27143 5466
rect 27143 5414 27155 5466
rect 27155 5414 27185 5466
rect 27209 5414 27219 5466
rect 27219 5414 27265 5466
rect 26969 5412 27025 5414
rect 27049 5412 27105 5414
rect 27129 5412 27185 5414
rect 27209 5412 27265 5414
rect 27158 4700 27160 4720
rect 27160 4700 27212 4720
rect 27212 4700 27214 4720
rect 27158 4664 27214 4700
rect 26969 4378 27025 4380
rect 27049 4378 27105 4380
rect 27129 4378 27185 4380
rect 27209 4378 27265 4380
rect 26969 4326 27015 4378
rect 27015 4326 27025 4378
rect 27049 4326 27079 4378
rect 27079 4326 27091 4378
rect 27091 4326 27105 4378
rect 27129 4326 27143 4378
rect 27143 4326 27155 4378
rect 27155 4326 27185 4378
rect 27209 4326 27219 4378
rect 27219 4326 27265 4378
rect 26969 4324 27025 4326
rect 27049 4324 27105 4326
rect 27129 4324 27185 4326
rect 27209 4324 27265 4326
rect 26330 2488 26386 2544
rect 26054 2080 26110 2136
rect 26422 1400 26478 1456
rect 25962 1128 26018 1184
rect 26606 1264 26662 1320
rect 27250 3440 27306 3496
rect 26969 3290 27025 3292
rect 27049 3290 27105 3292
rect 27129 3290 27185 3292
rect 27209 3290 27265 3292
rect 26969 3238 27015 3290
rect 27015 3238 27025 3290
rect 27049 3238 27079 3290
rect 27079 3238 27091 3290
rect 27091 3238 27105 3290
rect 27129 3238 27143 3290
rect 27143 3238 27155 3290
rect 27155 3238 27185 3290
rect 27209 3238 27219 3290
rect 27219 3238 27265 3290
rect 26969 3236 27025 3238
rect 27049 3236 27105 3238
rect 27129 3236 27185 3238
rect 27209 3236 27265 3238
rect 27894 7248 27950 7304
rect 28906 19352 28962 19408
rect 28998 19080 29054 19136
rect 28998 18808 29054 18864
rect 29182 18808 29238 18864
rect 28630 14864 28686 14920
rect 28538 13912 28594 13968
rect 28538 13776 28594 13832
rect 28906 17720 28962 17776
rect 28998 17040 29054 17096
rect 29642 19760 29698 19816
rect 29642 18944 29698 19000
rect 30764 21242 30820 21244
rect 30844 21242 30900 21244
rect 30924 21242 30980 21244
rect 31004 21242 31060 21244
rect 30764 21190 30810 21242
rect 30810 21190 30820 21242
rect 30844 21190 30874 21242
rect 30874 21190 30886 21242
rect 30886 21190 30900 21242
rect 30924 21190 30938 21242
rect 30938 21190 30950 21242
rect 30950 21190 30980 21242
rect 31004 21190 31014 21242
rect 31014 21190 31060 21242
rect 30764 21188 30820 21190
rect 30844 21188 30900 21190
rect 30924 21188 30980 21190
rect 31004 21188 31060 21190
rect 29642 16768 29698 16824
rect 29550 16632 29606 16688
rect 29458 16224 29514 16280
rect 29366 16088 29422 16144
rect 28814 11736 28870 11792
rect 29182 9968 29238 10024
rect 28078 5616 28134 5672
rect 27710 4120 27766 4176
rect 26969 2202 27025 2204
rect 27049 2202 27105 2204
rect 27129 2202 27185 2204
rect 27209 2202 27265 2204
rect 26969 2150 27015 2202
rect 27015 2150 27025 2202
rect 27049 2150 27079 2202
rect 27079 2150 27091 2202
rect 27091 2150 27105 2202
rect 27129 2150 27143 2202
rect 27143 2150 27155 2202
rect 27155 2150 27185 2202
rect 27209 2150 27219 2202
rect 27219 2150 27265 2202
rect 26969 2148 27025 2150
rect 27049 2148 27105 2150
rect 27129 2148 27185 2150
rect 27209 2148 27265 2150
rect 27526 1944 27582 2000
rect 26969 1114 27025 1116
rect 27049 1114 27105 1116
rect 27129 1114 27185 1116
rect 27209 1114 27265 1116
rect 26969 1062 27015 1114
rect 27015 1062 27025 1114
rect 27049 1062 27079 1114
rect 27079 1062 27091 1114
rect 27091 1062 27105 1114
rect 27129 1062 27143 1114
rect 27143 1062 27155 1114
rect 27155 1062 27185 1114
rect 27209 1062 27219 1114
rect 27219 1062 27265 1114
rect 26969 1060 27025 1062
rect 27049 1060 27105 1062
rect 27129 1060 27185 1062
rect 27209 1060 27265 1062
rect 27802 3576 27858 3632
rect 28446 2896 28502 2952
rect 29182 9288 29238 9344
rect 29642 15816 29698 15872
rect 30286 18672 30342 18728
rect 29826 16360 29882 16416
rect 29550 15544 29606 15600
rect 29458 15272 29514 15328
rect 29366 12416 29422 12472
rect 30010 15952 30066 16008
rect 30010 15680 30066 15736
rect 29274 8880 29330 8936
rect 28722 3032 28778 3088
rect 28814 1808 28870 1864
rect 29550 6840 29606 6896
rect 30010 13232 30066 13288
rect 29918 12008 29974 12064
rect 29918 11192 29974 11248
rect 29826 9424 29882 9480
rect 30378 17992 30434 18048
rect 30378 17604 30434 17640
rect 30378 17584 30380 17604
rect 30380 17584 30432 17604
rect 30432 17584 30434 17604
rect 30378 17040 30434 17096
rect 30378 15000 30434 15056
rect 30378 13640 30434 13696
rect 29826 8472 29882 8528
rect 29366 5208 29422 5264
rect 29458 5072 29514 5128
rect 29458 3984 29514 4040
rect 30194 7792 30250 7848
rect 30764 20154 30820 20156
rect 30844 20154 30900 20156
rect 30924 20154 30980 20156
rect 31004 20154 31060 20156
rect 30764 20102 30810 20154
rect 30810 20102 30820 20154
rect 30844 20102 30874 20154
rect 30874 20102 30886 20154
rect 30886 20102 30900 20154
rect 30924 20102 30938 20154
rect 30938 20102 30950 20154
rect 30950 20102 30980 20154
rect 31004 20102 31014 20154
rect 31014 20102 31060 20154
rect 30764 20100 30820 20102
rect 30844 20100 30900 20102
rect 30924 20100 30980 20102
rect 31004 20100 31060 20102
rect 30764 19066 30820 19068
rect 30844 19066 30900 19068
rect 30924 19066 30980 19068
rect 31004 19066 31060 19068
rect 30764 19014 30810 19066
rect 30810 19014 30820 19066
rect 30844 19014 30874 19066
rect 30874 19014 30886 19066
rect 30886 19014 30900 19066
rect 30924 19014 30938 19066
rect 30938 19014 30950 19066
rect 30950 19014 30980 19066
rect 31004 19014 31014 19066
rect 31014 19014 31060 19066
rect 30764 19012 30820 19014
rect 30844 19012 30900 19014
rect 30924 19012 30980 19014
rect 31004 19012 31060 19014
rect 30764 17978 30820 17980
rect 30844 17978 30900 17980
rect 30924 17978 30980 17980
rect 31004 17978 31060 17980
rect 30764 17926 30810 17978
rect 30810 17926 30820 17978
rect 30844 17926 30874 17978
rect 30874 17926 30886 17978
rect 30886 17926 30900 17978
rect 30924 17926 30938 17978
rect 30938 17926 30950 17978
rect 30950 17926 30980 17978
rect 31004 17926 31014 17978
rect 31014 17926 31060 17978
rect 30764 17924 30820 17926
rect 30844 17924 30900 17926
rect 30924 17924 30980 17926
rect 31004 17924 31060 17926
rect 30746 17040 30802 17096
rect 30764 16890 30820 16892
rect 30844 16890 30900 16892
rect 30924 16890 30980 16892
rect 31004 16890 31060 16892
rect 30764 16838 30810 16890
rect 30810 16838 30820 16890
rect 30844 16838 30874 16890
rect 30874 16838 30886 16890
rect 30886 16838 30900 16890
rect 30924 16838 30938 16890
rect 30938 16838 30950 16890
rect 30950 16838 30980 16890
rect 31004 16838 31014 16890
rect 31014 16838 31060 16890
rect 30764 16836 30820 16838
rect 30844 16836 30900 16838
rect 30924 16836 30980 16838
rect 31004 16836 31060 16838
rect 30764 15802 30820 15804
rect 30844 15802 30900 15804
rect 30924 15802 30980 15804
rect 31004 15802 31060 15804
rect 30764 15750 30810 15802
rect 30810 15750 30820 15802
rect 30844 15750 30874 15802
rect 30874 15750 30886 15802
rect 30886 15750 30900 15802
rect 30924 15750 30938 15802
rect 30938 15750 30950 15802
rect 30950 15750 30980 15802
rect 31004 15750 31014 15802
rect 31014 15750 31060 15802
rect 30764 15748 30820 15750
rect 30844 15748 30900 15750
rect 30924 15748 30980 15750
rect 31004 15748 31060 15750
rect 30746 15544 30802 15600
rect 30764 14714 30820 14716
rect 30844 14714 30900 14716
rect 30924 14714 30980 14716
rect 31004 14714 31060 14716
rect 30764 14662 30810 14714
rect 30810 14662 30820 14714
rect 30844 14662 30874 14714
rect 30874 14662 30886 14714
rect 30886 14662 30900 14714
rect 30924 14662 30938 14714
rect 30938 14662 30950 14714
rect 30950 14662 30980 14714
rect 31004 14662 31014 14714
rect 31014 14662 31060 14714
rect 30764 14660 30820 14662
rect 30844 14660 30900 14662
rect 30924 14660 30980 14662
rect 31004 14660 31060 14662
rect 30764 13626 30820 13628
rect 30844 13626 30900 13628
rect 30924 13626 30980 13628
rect 31004 13626 31060 13628
rect 30764 13574 30810 13626
rect 30810 13574 30820 13626
rect 30844 13574 30874 13626
rect 30874 13574 30886 13626
rect 30886 13574 30900 13626
rect 30924 13574 30938 13626
rect 30938 13574 30950 13626
rect 30950 13574 30980 13626
rect 31004 13574 31014 13626
rect 31014 13574 31060 13626
rect 30764 13572 30820 13574
rect 30844 13572 30900 13574
rect 30924 13572 30980 13574
rect 31004 13572 31060 13574
rect 30764 12538 30820 12540
rect 30844 12538 30900 12540
rect 30924 12538 30980 12540
rect 31004 12538 31060 12540
rect 30764 12486 30810 12538
rect 30810 12486 30820 12538
rect 30844 12486 30874 12538
rect 30874 12486 30886 12538
rect 30886 12486 30900 12538
rect 30924 12486 30938 12538
rect 30938 12486 30950 12538
rect 30950 12486 30980 12538
rect 31004 12486 31014 12538
rect 31014 12486 31060 12538
rect 30764 12484 30820 12486
rect 30844 12484 30900 12486
rect 30924 12484 30980 12486
rect 31004 12484 31060 12486
rect 30764 11450 30820 11452
rect 30844 11450 30900 11452
rect 30924 11450 30980 11452
rect 31004 11450 31060 11452
rect 30764 11398 30810 11450
rect 30810 11398 30820 11450
rect 30844 11398 30874 11450
rect 30874 11398 30886 11450
rect 30886 11398 30900 11450
rect 30924 11398 30938 11450
rect 30938 11398 30950 11450
rect 30950 11398 30980 11450
rect 31004 11398 31014 11450
rect 31014 11398 31060 11450
rect 30764 11396 30820 11398
rect 30844 11396 30900 11398
rect 30924 11396 30980 11398
rect 31004 11396 31060 11398
rect 30764 10362 30820 10364
rect 30844 10362 30900 10364
rect 30924 10362 30980 10364
rect 31004 10362 31060 10364
rect 30764 10310 30810 10362
rect 30810 10310 30820 10362
rect 30844 10310 30874 10362
rect 30874 10310 30886 10362
rect 30886 10310 30900 10362
rect 30924 10310 30938 10362
rect 30938 10310 30950 10362
rect 30950 10310 30980 10362
rect 31004 10310 31014 10362
rect 31014 10310 31060 10362
rect 30764 10308 30820 10310
rect 30844 10308 30900 10310
rect 30924 10308 30980 10310
rect 31004 10308 31060 10310
rect 30764 9274 30820 9276
rect 30844 9274 30900 9276
rect 30924 9274 30980 9276
rect 31004 9274 31060 9276
rect 30764 9222 30810 9274
rect 30810 9222 30820 9274
rect 30844 9222 30874 9274
rect 30874 9222 30886 9274
rect 30886 9222 30900 9274
rect 30924 9222 30938 9274
rect 30938 9222 30950 9274
rect 30950 9222 30980 9274
rect 31004 9222 31014 9274
rect 31014 9222 31060 9274
rect 30764 9220 30820 9222
rect 30844 9220 30900 9222
rect 30924 9220 30980 9222
rect 31004 9220 31060 9222
rect 31390 18264 31446 18320
rect 30764 8186 30820 8188
rect 30844 8186 30900 8188
rect 30924 8186 30980 8188
rect 31004 8186 31060 8188
rect 30764 8134 30810 8186
rect 30810 8134 30820 8186
rect 30844 8134 30874 8186
rect 30874 8134 30886 8186
rect 30886 8134 30900 8186
rect 30924 8134 30938 8186
rect 30938 8134 30950 8186
rect 30950 8134 30980 8186
rect 31004 8134 31014 8186
rect 31014 8134 31060 8186
rect 30764 8132 30820 8134
rect 30844 8132 30900 8134
rect 30924 8132 30980 8134
rect 31004 8132 31060 8134
rect 30764 7098 30820 7100
rect 30844 7098 30900 7100
rect 30924 7098 30980 7100
rect 31004 7098 31060 7100
rect 30764 7046 30810 7098
rect 30810 7046 30820 7098
rect 30844 7046 30874 7098
rect 30874 7046 30886 7098
rect 30886 7046 30900 7098
rect 30924 7046 30938 7098
rect 30938 7046 30950 7098
rect 30950 7046 30980 7098
rect 31004 7046 31014 7098
rect 31014 7046 31060 7098
rect 30764 7044 30820 7046
rect 30844 7044 30900 7046
rect 30924 7044 30980 7046
rect 31004 7044 31060 7046
rect 30764 6010 30820 6012
rect 30844 6010 30900 6012
rect 30924 6010 30980 6012
rect 31004 6010 31060 6012
rect 30764 5958 30810 6010
rect 30810 5958 30820 6010
rect 30844 5958 30874 6010
rect 30874 5958 30886 6010
rect 30886 5958 30900 6010
rect 30924 5958 30938 6010
rect 30938 5958 30950 6010
rect 30950 5958 30980 6010
rect 31004 5958 31014 6010
rect 31014 5958 31060 6010
rect 30764 5956 30820 5958
rect 30844 5956 30900 5958
rect 30924 5956 30980 5958
rect 31004 5956 31060 5958
rect 30764 4922 30820 4924
rect 30844 4922 30900 4924
rect 30924 4922 30980 4924
rect 31004 4922 31060 4924
rect 30764 4870 30810 4922
rect 30810 4870 30820 4922
rect 30844 4870 30874 4922
rect 30874 4870 30886 4922
rect 30886 4870 30900 4922
rect 30924 4870 30938 4922
rect 30938 4870 30950 4922
rect 30950 4870 30980 4922
rect 31004 4870 31014 4922
rect 31014 4870 31060 4922
rect 30764 4868 30820 4870
rect 30844 4868 30900 4870
rect 30924 4868 30980 4870
rect 31004 4868 31060 4870
rect 30764 3834 30820 3836
rect 30844 3834 30900 3836
rect 30924 3834 30980 3836
rect 31004 3834 31060 3836
rect 30764 3782 30810 3834
rect 30810 3782 30820 3834
rect 30844 3782 30874 3834
rect 30874 3782 30886 3834
rect 30886 3782 30900 3834
rect 30924 3782 30938 3834
rect 30938 3782 30950 3834
rect 30950 3782 30980 3834
rect 31004 3782 31014 3834
rect 31014 3782 31060 3834
rect 30764 3780 30820 3782
rect 30844 3780 30900 3782
rect 30924 3780 30980 3782
rect 31004 3780 31060 3782
rect 30764 2746 30820 2748
rect 30844 2746 30900 2748
rect 30924 2746 30980 2748
rect 31004 2746 31060 2748
rect 30764 2694 30810 2746
rect 30810 2694 30820 2746
rect 30844 2694 30874 2746
rect 30874 2694 30886 2746
rect 30886 2694 30900 2746
rect 30924 2694 30938 2746
rect 30938 2694 30950 2746
rect 30950 2694 30980 2746
rect 31004 2694 31014 2746
rect 31014 2694 31060 2746
rect 30764 2692 30820 2694
rect 30844 2692 30900 2694
rect 30924 2692 30980 2694
rect 31004 2692 31060 2694
rect 30764 1658 30820 1660
rect 30844 1658 30900 1660
rect 30924 1658 30980 1660
rect 31004 1658 31060 1660
rect 30764 1606 30810 1658
rect 30810 1606 30820 1658
rect 30844 1606 30874 1658
rect 30874 1606 30886 1658
rect 30886 1606 30900 1658
rect 30924 1606 30938 1658
rect 30938 1606 30950 1658
rect 30950 1606 30980 1658
rect 31004 1606 31014 1658
rect 31014 1606 31060 1658
rect 30764 1604 30820 1606
rect 30844 1604 30900 1606
rect 30924 1604 30980 1606
rect 31004 1604 31060 1606
rect 29182 720 29238 776
rect 24950 312 25006 368
rect 30764 570 30820 572
rect 30844 570 30900 572
rect 30924 570 30980 572
rect 31004 570 31060 572
rect 30764 518 30810 570
rect 30810 518 30820 570
rect 30844 518 30874 570
rect 30874 518 30886 570
rect 30886 518 30900 570
rect 30924 518 30938 570
rect 30938 518 30950 570
rect 30950 518 30980 570
rect 31004 518 31014 570
rect 31014 518 31060 570
rect 30764 516 30820 518
rect 30844 516 30900 518
rect 30924 516 30980 518
rect 31004 516 31060 518
rect 24858 40 24914 96
<< metal3 >>
rect 9121 22266 9187 22269
rect 2822 22264 9187 22266
rect 2822 22208 9126 22264
rect 9182 22208 9187 22264
rect 2822 22206 9187 22208
rect 2822 22132 2882 22206
rect 9121 22203 9187 22206
rect 14365 22268 14431 22269
rect 14365 22264 14412 22268
rect 14476 22266 14482 22268
rect 22277 22266 22343 22269
rect 23749 22266 23815 22269
rect 14365 22208 14370 22264
rect 14365 22204 14412 22208
rect 14476 22206 14522 22266
rect 22277 22264 23815 22266
rect 22277 22208 22282 22264
rect 22338 22208 23754 22264
rect 23810 22208 23815 22264
rect 22277 22206 23815 22208
rect 14476 22204 14482 22206
rect 14365 22203 14431 22204
rect 22277 22203 22343 22206
rect 23749 22203 23815 22206
rect 2814 22068 2820 22132
rect 2884 22068 2890 22132
rect 9029 22130 9095 22133
rect 21633 22130 21699 22133
rect 22553 22130 22619 22133
rect 9029 22128 17970 22130
rect 9029 22072 9034 22128
rect 9090 22072 17970 22128
rect 9029 22070 17970 22072
rect 9029 22067 9095 22070
rect 2497 21994 2563 21997
rect 10961 21996 11027 21997
rect 10910 21994 10916 21996
rect 2497 21992 2790 21994
rect 2497 21936 2502 21992
rect 2558 21936 2790 21992
rect 2497 21934 2790 21936
rect 10870 21934 10916 21994
rect 10980 21992 11027 21996
rect 11022 21936 11027 21992
rect 2497 21931 2563 21934
rect 2730 21586 2790 21934
rect 10910 21932 10916 21934
rect 10980 21932 11027 21936
rect 10961 21931 11027 21932
rect 11421 21994 11487 21997
rect 13997 21994 14063 21997
rect 11421 21992 12082 21994
rect 11421 21936 11426 21992
rect 11482 21962 12082 21992
rect 13126 21992 14063 21994
rect 13126 21962 14002 21992
rect 11482 21936 12020 21962
rect 11421 21934 12020 21936
rect 11421 21931 11487 21934
rect 12014 21898 12020 21934
rect 12084 21898 12090 21962
rect 13118 21898 13124 21962
rect 13188 21936 14002 21962
rect 14058 21936 14063 21992
rect 13188 21934 14063 21936
rect 17910 21994 17970 22070
rect 21633 22128 22619 22130
rect 21633 22072 21638 22128
rect 21694 22072 22558 22128
rect 22614 22072 22619 22128
rect 21633 22070 22619 22072
rect 21633 22067 21699 22070
rect 22553 22067 22619 22070
rect 23289 22130 23355 22133
rect 25037 22130 25103 22133
rect 23289 22128 25103 22130
rect 23289 22072 23294 22128
rect 23350 22072 25042 22128
rect 25098 22072 25103 22128
rect 23289 22070 25103 22072
rect 23289 22067 23355 22070
rect 25037 22067 25103 22070
rect 26325 21994 26391 21997
rect 17910 21992 26391 21994
rect 17910 21936 26330 21992
rect 26386 21936 26391 21992
rect 17910 21934 26391 21936
rect 13188 21898 13194 21934
rect 13997 21931 14063 21934
rect 26325 21931 26391 21934
rect 6545 21858 6611 21861
rect 9489 21858 9555 21861
rect 6545 21856 9555 21858
rect 6545 21800 6550 21856
rect 6606 21800 9494 21856
rect 9550 21800 9555 21856
rect 6545 21798 9555 21800
rect 6545 21795 6611 21798
rect 9489 21795 9555 21798
rect 21909 21860 21975 21861
rect 21909 21856 21956 21860
rect 22020 21858 22026 21860
rect 21909 21800 21914 21856
rect 21909 21796 21956 21800
rect 22020 21798 22066 21858
rect 22020 21796 22026 21798
rect 23606 21796 23612 21860
rect 23676 21858 23682 21860
rect 23749 21858 23815 21861
rect 23676 21856 23815 21858
rect 23676 21800 23754 21856
rect 23810 21800 23815 21856
rect 23676 21798 23815 21800
rect 23676 21796 23682 21798
rect 21909 21795 21975 21796
rect 23749 21795 23815 21798
rect 4189 21792 4505 21793
rect 4189 21728 4195 21792
rect 4259 21728 4275 21792
rect 4339 21728 4355 21792
rect 4419 21728 4435 21792
rect 4499 21728 4505 21792
rect 4189 21727 4505 21728
rect 11779 21792 12095 21793
rect 11779 21728 11785 21792
rect 11849 21728 11865 21792
rect 11929 21728 11945 21792
rect 12009 21728 12025 21792
rect 12089 21728 12095 21792
rect 11779 21727 12095 21728
rect 19369 21792 19685 21793
rect 19369 21728 19375 21792
rect 19439 21728 19455 21792
rect 19519 21728 19535 21792
rect 19599 21728 19615 21792
rect 19679 21728 19685 21792
rect 19369 21727 19685 21728
rect 26959 21792 27275 21793
rect 26959 21728 26965 21792
rect 27029 21728 27045 21792
rect 27109 21728 27125 21792
rect 27189 21728 27205 21792
rect 27269 21728 27275 21792
rect 26959 21727 27275 21728
rect 5809 21722 5875 21725
rect 8661 21722 8727 21725
rect 5809 21720 8727 21722
rect 5809 21664 5814 21720
rect 5870 21664 8666 21720
rect 8722 21664 8727 21720
rect 5809 21662 8727 21664
rect 5809 21659 5875 21662
rect 8661 21659 8727 21662
rect 12157 21722 12223 21725
rect 16757 21722 16823 21725
rect 12157 21720 16823 21722
rect 12157 21664 12162 21720
rect 12218 21664 16762 21720
rect 16818 21664 16823 21720
rect 12157 21662 16823 21664
rect 12157 21659 12223 21662
rect 16757 21659 16823 21662
rect 22093 21722 22159 21725
rect 24669 21722 24735 21725
rect 25957 21722 26023 21725
rect 22093 21720 26023 21722
rect 22093 21664 22098 21720
rect 22154 21664 24674 21720
rect 24730 21664 25962 21720
rect 26018 21664 26023 21720
rect 22093 21662 26023 21664
rect 22093 21659 22159 21662
rect 24669 21659 24735 21662
rect 25957 21659 26023 21662
rect 26693 21586 26759 21589
rect 2730 21584 26759 21586
rect 2730 21528 26698 21584
rect 26754 21528 26759 21584
rect 2730 21526 26759 21528
rect 26693 21523 26759 21526
rect 7005 21450 7071 21453
rect 27797 21450 27863 21453
rect 7005 21448 27863 21450
rect 7005 21392 7010 21448
rect 7066 21392 27802 21448
rect 27858 21392 27863 21448
rect 7005 21390 27863 21392
rect 7005 21387 7071 21390
rect 27797 21387 27863 21390
rect 8385 21314 8451 21317
rect 8845 21314 8911 21317
rect 8385 21312 8911 21314
rect 8385 21256 8390 21312
rect 8446 21256 8850 21312
rect 8906 21256 8911 21312
rect 8385 21254 8911 21256
rect 8385 21251 8451 21254
rect 8845 21251 8911 21254
rect 9213 21314 9279 21317
rect 10174 21314 10180 21316
rect 9213 21312 10180 21314
rect 9213 21256 9218 21312
rect 9274 21256 10180 21312
rect 9213 21254 10180 21256
rect 9213 21251 9279 21254
rect 10174 21252 10180 21254
rect 10244 21252 10250 21316
rect 10869 21314 10935 21317
rect 15377 21314 15443 21317
rect 10869 21312 15443 21314
rect 10869 21256 10874 21312
rect 10930 21256 15382 21312
rect 15438 21256 15443 21312
rect 10869 21254 15443 21256
rect 10869 21251 10935 21254
rect 15377 21251 15443 21254
rect 16113 21314 16179 21317
rect 18321 21314 18387 21317
rect 16113 21312 18387 21314
rect 16113 21256 16118 21312
rect 16174 21256 18326 21312
rect 18382 21256 18387 21312
rect 16113 21254 18387 21256
rect 16113 21251 16179 21254
rect 18321 21251 18387 21254
rect 7984 21248 8300 21249
rect 7984 21184 7990 21248
rect 8054 21184 8070 21248
rect 8134 21184 8150 21248
rect 8214 21184 8230 21248
rect 8294 21184 8300 21248
rect 7984 21183 8300 21184
rect 15574 21248 15890 21249
rect 15574 21184 15580 21248
rect 15644 21184 15660 21248
rect 15724 21184 15740 21248
rect 15804 21184 15820 21248
rect 15884 21184 15890 21248
rect 15574 21183 15890 21184
rect 23164 21248 23480 21249
rect 23164 21184 23170 21248
rect 23234 21184 23250 21248
rect 23314 21184 23330 21248
rect 23394 21184 23410 21248
rect 23474 21184 23480 21248
rect 23164 21183 23480 21184
rect 30754 21248 31070 21249
rect 30754 21184 30760 21248
rect 30824 21184 30840 21248
rect 30904 21184 30920 21248
rect 30984 21184 31000 21248
rect 31064 21184 31070 21248
rect 30754 21183 31070 21184
rect 4061 21178 4127 21181
rect 7097 21178 7163 21181
rect 4061 21176 7163 21178
rect 4061 21120 4066 21176
rect 4122 21120 7102 21176
rect 7158 21120 7163 21176
rect 4061 21118 7163 21120
rect 4061 21115 4127 21118
rect 7097 21115 7163 21118
rect 8477 21178 8543 21181
rect 26141 21178 26207 21181
rect 26366 21178 26372 21180
rect 8477 21176 12450 21178
rect 8477 21120 8482 21176
rect 8538 21120 12450 21176
rect 8477 21118 12450 21120
rect 8477 21115 8543 21118
rect 3509 21042 3575 21045
rect 12157 21042 12223 21045
rect 3509 21040 12223 21042
rect 3509 20984 3514 21040
rect 3570 20984 12162 21040
rect 12218 20984 12223 21040
rect 3509 20982 12223 20984
rect 12390 21042 12450 21118
rect 26141 21176 26372 21178
rect 26141 21120 26146 21176
rect 26202 21120 26372 21176
rect 26141 21118 26372 21120
rect 26141 21115 26207 21118
rect 26366 21116 26372 21118
rect 26436 21116 26442 21180
rect 14089 21042 14155 21045
rect 12390 21040 14155 21042
rect 12390 20984 14094 21040
rect 14150 20984 14155 21040
rect 12390 20982 14155 20984
rect 3509 20979 3575 20982
rect 12157 20979 12223 20982
rect 14089 20979 14155 20982
rect 14641 21042 14707 21045
rect 17585 21042 17651 21045
rect 14641 21040 17651 21042
rect 14641 20984 14646 21040
rect 14702 20984 17590 21040
rect 17646 20984 17651 21040
rect 14641 20982 17651 20984
rect 14641 20979 14707 20982
rect 17585 20979 17651 20982
rect 20161 21042 20227 21045
rect 25630 21042 25636 21044
rect 20161 21040 25636 21042
rect 20161 20984 20166 21040
rect 20222 20984 25636 21040
rect 20161 20982 25636 20984
rect 20161 20979 20227 20982
rect 25630 20980 25636 20982
rect 25700 20980 25706 21044
rect 5809 20906 5875 20909
rect 6453 20906 6519 20909
rect 5809 20904 6519 20906
rect 5809 20848 5814 20904
rect 5870 20848 6458 20904
rect 6514 20848 6519 20904
rect 5809 20846 6519 20848
rect 5809 20843 5875 20846
rect 6453 20843 6519 20846
rect 6637 20906 6703 20909
rect 18045 20906 18111 20909
rect 6637 20904 18111 20906
rect 6637 20848 6642 20904
rect 6698 20848 18050 20904
rect 18106 20848 18111 20904
rect 6637 20846 18111 20848
rect 6637 20843 6703 20846
rect 18045 20843 18111 20846
rect 21817 20906 21883 20909
rect 23933 20906 23999 20909
rect 26233 20906 26299 20909
rect 27654 20906 27660 20908
rect 21817 20904 27660 20906
rect 21817 20848 21822 20904
rect 21878 20848 23938 20904
rect 23994 20848 26238 20904
rect 26294 20848 27660 20904
rect 21817 20846 27660 20848
rect 21817 20843 21883 20846
rect 23933 20843 23999 20846
rect 26233 20843 26299 20846
rect 27654 20844 27660 20846
rect 27724 20844 27730 20908
rect 4613 20770 4679 20773
rect 8477 20770 8543 20773
rect 4613 20768 8543 20770
rect 4613 20712 4618 20768
rect 4674 20712 8482 20768
rect 8538 20712 8543 20768
rect 4613 20710 8543 20712
rect 4613 20707 4679 20710
rect 8477 20707 8543 20710
rect 8886 20708 8892 20772
rect 8956 20770 8962 20772
rect 10501 20770 10567 20773
rect 8956 20768 10567 20770
rect 8956 20712 10506 20768
rect 10562 20712 10567 20768
rect 8956 20710 10567 20712
rect 8956 20708 8962 20710
rect 10501 20707 10567 20710
rect 10869 20770 10935 20773
rect 11513 20770 11579 20773
rect 10869 20768 11579 20770
rect 10869 20712 10874 20768
rect 10930 20712 11518 20768
rect 11574 20712 11579 20768
rect 10869 20710 11579 20712
rect 10869 20707 10935 20710
rect 11513 20707 11579 20710
rect 13813 20770 13879 20773
rect 18229 20770 18295 20773
rect 24342 20770 24348 20772
rect 13813 20768 18295 20770
rect 13813 20712 13818 20768
rect 13874 20712 18234 20768
rect 18290 20712 18295 20768
rect 13813 20710 18295 20712
rect 13813 20707 13879 20710
rect 18229 20707 18295 20710
rect 20118 20710 24348 20770
rect 4189 20704 4505 20705
rect 4189 20640 4195 20704
rect 4259 20640 4275 20704
rect 4339 20640 4355 20704
rect 4419 20640 4435 20704
rect 4499 20640 4505 20704
rect 4189 20639 4505 20640
rect 11779 20704 12095 20705
rect 11779 20640 11785 20704
rect 11849 20640 11865 20704
rect 11929 20640 11945 20704
rect 12009 20640 12025 20704
rect 12089 20640 12095 20704
rect 11779 20639 12095 20640
rect 19369 20704 19685 20705
rect 19369 20640 19375 20704
rect 19439 20640 19455 20704
rect 19519 20640 19535 20704
rect 19599 20640 19615 20704
rect 19679 20640 19685 20704
rect 19369 20639 19685 20640
rect 5073 20634 5139 20637
rect 9622 20634 9628 20636
rect 5073 20632 9628 20634
rect 5073 20576 5078 20632
rect 5134 20576 9628 20632
rect 5073 20574 9628 20576
rect 5073 20571 5139 20574
rect 9622 20572 9628 20574
rect 9692 20572 9698 20636
rect 10358 20572 10364 20636
rect 10428 20572 10434 20636
rect 14222 20572 14228 20636
rect 14292 20634 14298 20636
rect 19977 20634 20043 20637
rect 20118 20634 20178 20710
rect 24342 20708 24348 20710
rect 24412 20708 24418 20772
rect 26959 20704 27275 20705
rect 26959 20640 26965 20704
rect 27029 20640 27045 20704
rect 27109 20640 27125 20704
rect 27189 20640 27205 20704
rect 27269 20640 27275 20704
rect 26959 20639 27275 20640
rect 14292 20574 19258 20634
rect 14292 20572 14298 20574
rect 4521 20498 4587 20501
rect 10366 20498 10426 20572
rect 4521 20496 10426 20498
rect 4521 20440 4526 20496
rect 4582 20440 10426 20496
rect 4521 20438 10426 20440
rect 10501 20498 10567 20501
rect 15193 20498 15259 20501
rect 10501 20496 15259 20498
rect 10501 20440 10506 20496
rect 10562 20440 15198 20496
rect 15254 20440 15259 20496
rect 10501 20438 15259 20440
rect 4521 20435 4587 20438
rect 10501 20435 10567 20438
rect 15193 20435 15259 20438
rect 15745 20498 15811 20501
rect 18413 20498 18479 20501
rect 15745 20496 18479 20498
rect 15745 20440 15750 20496
rect 15806 20440 18418 20496
rect 18474 20440 18479 20496
rect 15745 20438 18479 20440
rect 19198 20498 19258 20574
rect 19977 20632 20178 20634
rect 19977 20576 19982 20632
rect 20038 20576 20178 20632
rect 19977 20574 20178 20576
rect 21817 20634 21883 20637
rect 24853 20634 24919 20637
rect 21817 20632 24919 20634
rect 21817 20576 21822 20632
rect 21878 20576 24858 20632
rect 24914 20576 24919 20632
rect 21817 20574 24919 20576
rect 19977 20571 20043 20574
rect 21817 20571 21883 20574
rect 24853 20571 24919 20574
rect 19977 20498 20043 20501
rect 28165 20498 28231 20501
rect 19198 20496 20043 20498
rect 19198 20440 19982 20496
rect 20038 20440 20043 20496
rect 19198 20438 20043 20440
rect 15745 20435 15811 20438
rect 18413 20435 18479 20438
rect 19977 20435 20043 20438
rect 20854 20496 28231 20498
rect 20854 20440 28170 20496
rect 28226 20440 28231 20496
rect 20854 20438 28231 20440
rect 4889 20362 4955 20365
rect 6085 20362 6151 20365
rect 9397 20362 9463 20365
rect 20621 20362 20687 20365
rect 4889 20360 8586 20362
rect 4889 20304 4894 20360
rect 4950 20304 6090 20360
rect 6146 20304 8586 20360
rect 4889 20302 8586 20304
rect 4889 20299 4955 20302
rect 6085 20299 6151 20302
rect 8526 20226 8586 20302
rect 9397 20360 20687 20362
rect 9397 20304 9402 20360
rect 9458 20304 20626 20360
rect 20682 20304 20687 20360
rect 9397 20302 20687 20304
rect 9397 20299 9463 20302
rect 20621 20299 20687 20302
rect 13353 20226 13419 20229
rect 8526 20224 13419 20226
rect 8526 20168 13358 20224
rect 13414 20168 13419 20224
rect 8526 20166 13419 20168
rect 13353 20163 13419 20166
rect 16205 20226 16271 20229
rect 20854 20226 20914 20438
rect 28165 20435 28231 20438
rect 21909 20362 21975 20365
rect 22277 20362 22343 20365
rect 21909 20360 22343 20362
rect 21909 20304 21914 20360
rect 21970 20304 22282 20360
rect 22338 20304 22343 20360
rect 21909 20302 22343 20304
rect 21909 20299 21975 20302
rect 22277 20299 22343 20302
rect 16205 20224 20914 20226
rect 16205 20168 16210 20224
rect 16266 20168 20914 20224
rect 16205 20166 20914 20168
rect 16205 20163 16271 20166
rect 7984 20160 8300 20161
rect 7984 20096 7990 20160
rect 8054 20096 8070 20160
rect 8134 20096 8150 20160
rect 8214 20096 8230 20160
rect 8294 20096 8300 20160
rect 7984 20095 8300 20096
rect 15574 20160 15890 20161
rect 15574 20096 15580 20160
rect 15644 20096 15660 20160
rect 15724 20096 15740 20160
rect 15804 20096 15820 20160
rect 15884 20096 15890 20160
rect 15574 20095 15890 20096
rect 23164 20160 23480 20161
rect 23164 20096 23170 20160
rect 23234 20096 23250 20160
rect 23314 20096 23330 20160
rect 23394 20096 23410 20160
rect 23474 20096 23480 20160
rect 23164 20095 23480 20096
rect 30754 20160 31070 20161
rect 30754 20096 30760 20160
rect 30824 20096 30840 20160
rect 30904 20096 30920 20160
rect 30984 20096 31000 20160
rect 31064 20096 31070 20160
rect 30754 20095 31070 20096
rect 9438 20028 9444 20092
rect 9508 20090 9514 20092
rect 9857 20090 9923 20093
rect 9508 20088 9923 20090
rect 9508 20032 9862 20088
rect 9918 20032 9923 20088
rect 9508 20030 9923 20032
rect 9508 20028 9514 20030
rect 9857 20027 9923 20030
rect 10409 20090 10475 20093
rect 13905 20090 13971 20093
rect 10409 20088 13971 20090
rect 10409 20032 10414 20088
rect 10470 20032 13910 20088
rect 13966 20032 13971 20088
rect 10409 20030 13971 20032
rect 10409 20027 10475 20030
rect 13905 20027 13971 20030
rect 3417 19954 3483 19957
rect 10501 19954 10567 19957
rect 15377 19954 15443 19957
rect 3417 19952 10567 19954
rect 3417 19896 3422 19952
rect 3478 19896 10506 19952
rect 10562 19896 10567 19952
rect 3417 19894 10567 19896
rect 3417 19891 3483 19894
rect 10501 19891 10567 19894
rect 10734 19952 15443 19954
rect 10734 19896 15382 19952
rect 15438 19896 15443 19952
rect 10734 19894 15443 19896
rect 3601 19818 3667 19821
rect 7189 19818 7255 19821
rect 3601 19816 7255 19818
rect 3601 19760 3606 19816
rect 3662 19760 7194 19816
rect 7250 19760 7255 19816
rect 3601 19758 7255 19760
rect 3601 19755 3667 19758
rect 7189 19755 7255 19758
rect 8201 19818 8267 19821
rect 9254 19818 9260 19820
rect 8201 19816 9260 19818
rect 8201 19760 8206 19816
rect 8262 19760 9260 19816
rect 8201 19758 9260 19760
rect 8201 19755 8267 19758
rect 9254 19756 9260 19758
rect 9324 19756 9330 19820
rect 9622 19756 9628 19820
rect 9692 19818 9698 19820
rect 10734 19818 10794 19894
rect 15377 19891 15443 19894
rect 18873 19954 18939 19957
rect 23381 19954 23447 19957
rect 18873 19952 23447 19954
rect 18873 19896 18878 19952
rect 18934 19896 23386 19952
rect 23442 19896 23447 19952
rect 18873 19894 23447 19896
rect 18873 19891 18939 19894
rect 23381 19891 23447 19894
rect 23841 19954 23907 19957
rect 27613 19954 27679 19957
rect 23841 19952 27679 19954
rect 23841 19896 23846 19952
rect 23902 19896 27618 19952
rect 27674 19896 27679 19952
rect 23841 19894 27679 19896
rect 23841 19891 23907 19894
rect 27613 19891 27679 19894
rect 21081 19818 21147 19821
rect 9692 19758 10794 19818
rect 10918 19816 21147 19818
rect 10918 19760 21086 19816
rect 21142 19760 21147 19816
rect 10918 19758 21147 19760
rect 9692 19756 9698 19758
rect 5625 19682 5691 19685
rect 9581 19682 9647 19685
rect 5625 19680 9647 19682
rect 5625 19624 5630 19680
rect 5686 19624 9586 19680
rect 9642 19624 9647 19680
rect 5625 19622 9647 19624
rect 5625 19619 5691 19622
rect 9581 19619 9647 19622
rect 4189 19616 4505 19617
rect 4189 19552 4195 19616
rect 4259 19552 4275 19616
rect 4339 19552 4355 19616
rect 4419 19552 4435 19616
rect 4499 19552 4505 19616
rect 4189 19551 4505 19552
rect 10918 19549 10978 19758
rect 21081 19755 21147 19758
rect 23565 19818 23631 19821
rect 29637 19818 29703 19821
rect 23565 19816 29703 19818
rect 23565 19760 23570 19816
rect 23626 19760 29642 19816
rect 29698 19760 29703 19816
rect 23565 19758 29703 19760
rect 23565 19755 23631 19758
rect 29637 19755 29703 19758
rect 13537 19682 13603 19685
rect 16205 19682 16271 19685
rect 13537 19680 16271 19682
rect 13537 19624 13542 19680
rect 13598 19624 16210 19680
rect 16266 19624 16271 19680
rect 13537 19622 16271 19624
rect 13537 19619 13603 19622
rect 16205 19619 16271 19622
rect 20713 19682 20779 19685
rect 23841 19682 23907 19685
rect 20713 19680 23907 19682
rect 20713 19624 20718 19680
rect 20774 19624 23846 19680
rect 23902 19624 23907 19680
rect 20713 19622 23907 19624
rect 20713 19619 20779 19622
rect 23841 19619 23907 19622
rect 11779 19616 12095 19617
rect 11779 19552 11785 19616
rect 11849 19552 11865 19616
rect 11929 19552 11945 19616
rect 12009 19552 12025 19616
rect 12089 19552 12095 19616
rect 11779 19551 12095 19552
rect 19369 19616 19685 19617
rect 19369 19552 19375 19616
rect 19439 19552 19455 19616
rect 19519 19552 19535 19616
rect 19599 19552 19615 19616
rect 19679 19552 19685 19616
rect 19369 19551 19685 19552
rect 26959 19616 27275 19617
rect 26959 19552 26965 19616
rect 27029 19552 27045 19616
rect 27109 19552 27125 19616
rect 27189 19552 27205 19616
rect 27269 19552 27275 19616
rect 26959 19551 27275 19552
rect 5809 19546 5875 19549
rect 10869 19546 10978 19549
rect 5809 19544 10978 19546
rect 5809 19488 5814 19544
rect 5870 19488 10874 19544
rect 10930 19488 10978 19544
rect 5809 19486 10978 19488
rect 15745 19546 15811 19549
rect 18229 19546 18295 19549
rect 26233 19546 26299 19549
rect 15745 19544 18295 19546
rect 15745 19488 15750 19544
rect 15806 19488 18234 19544
rect 18290 19488 18295 19544
rect 15745 19486 18295 19488
rect 5809 19483 5875 19486
rect 10869 19483 10935 19486
rect 15745 19483 15811 19486
rect 18229 19483 18295 19486
rect 19934 19544 26299 19546
rect 19934 19488 26238 19544
rect 26294 19488 26299 19544
rect 19934 19486 26299 19488
rect 8518 19410 8524 19412
rect 8342 19350 8524 19410
rect 4654 19212 4660 19276
rect 4724 19274 4730 19276
rect 8342 19274 8402 19350
rect 8518 19348 8524 19350
rect 8588 19348 8594 19412
rect 8661 19410 8727 19413
rect 8937 19410 9003 19413
rect 8661 19408 9003 19410
rect 8661 19352 8666 19408
rect 8722 19352 8942 19408
rect 8998 19352 9003 19408
rect 8661 19350 9003 19352
rect 8661 19347 8727 19350
rect 8937 19347 9003 19350
rect 9254 19348 9260 19412
rect 9324 19410 9330 19412
rect 13629 19410 13695 19413
rect 9324 19408 13695 19410
rect 9324 19352 13634 19408
rect 13690 19352 13695 19408
rect 9324 19350 13695 19352
rect 9324 19348 9330 19350
rect 13629 19347 13695 19350
rect 13997 19412 14063 19413
rect 13997 19408 14044 19412
rect 14108 19410 14114 19412
rect 15101 19410 15167 19413
rect 19701 19410 19767 19413
rect 19934 19410 19994 19486
rect 26233 19483 26299 19486
rect 13997 19352 14002 19408
rect 13997 19348 14044 19352
rect 14108 19350 14154 19410
rect 15101 19408 15210 19410
rect 15101 19352 15106 19408
rect 15162 19352 15210 19408
rect 14108 19348 14114 19350
rect 13997 19347 14063 19348
rect 15101 19347 15210 19352
rect 19701 19408 19994 19410
rect 19701 19352 19706 19408
rect 19762 19352 19994 19408
rect 19701 19350 19994 19352
rect 20529 19410 20595 19413
rect 26049 19410 26115 19413
rect 20529 19408 26115 19410
rect 20529 19352 20534 19408
rect 20590 19352 26054 19408
rect 26110 19352 26115 19408
rect 20529 19350 26115 19352
rect 19701 19347 19767 19350
rect 20529 19347 20595 19350
rect 26049 19347 26115 19350
rect 27245 19410 27311 19413
rect 28901 19410 28967 19413
rect 27245 19408 28967 19410
rect 27245 19352 27250 19408
rect 27306 19352 28906 19408
rect 28962 19352 28967 19408
rect 27245 19350 28967 19352
rect 27245 19347 27311 19350
rect 28901 19347 28967 19350
rect 4724 19214 8402 19274
rect 8937 19274 9003 19277
rect 15009 19274 15075 19277
rect 15150 19276 15210 19347
rect 8937 19272 15075 19274
rect 8937 19216 8942 19272
rect 8998 19216 15014 19272
rect 15070 19216 15075 19272
rect 8937 19214 15075 19216
rect 4724 19212 4730 19214
rect 8937 19211 9003 19214
rect 15009 19211 15075 19214
rect 15142 19212 15148 19276
rect 15212 19212 15218 19276
rect 17309 19274 17375 19277
rect 19333 19274 19399 19277
rect 17309 19272 19399 19274
rect 17309 19216 17314 19272
rect 17370 19216 19338 19272
rect 19394 19216 19399 19272
rect 17309 19214 19399 19216
rect 17309 19211 17375 19214
rect 19333 19211 19399 19214
rect 22870 19212 22876 19276
rect 22940 19274 22946 19276
rect 25129 19274 25195 19277
rect 25262 19274 25268 19276
rect 22940 19214 23674 19274
rect 22940 19212 22946 19214
rect 2313 19138 2379 19141
rect 5809 19138 5875 19141
rect 11462 19138 11468 19140
rect 2313 19136 5875 19138
rect 2313 19080 2318 19136
rect 2374 19080 5814 19136
rect 5870 19080 5875 19136
rect 2313 19078 5875 19080
rect 2313 19075 2379 19078
rect 5809 19075 5875 19078
rect 8526 19078 11468 19138
rect 7984 19072 8300 19073
rect 7984 19008 7990 19072
rect 8054 19008 8070 19072
rect 8134 19008 8150 19072
rect 8214 19008 8230 19072
rect 8294 19008 8300 19072
rect 7984 19007 8300 19008
rect 4981 19002 5047 19005
rect 6913 19002 6979 19005
rect 4981 19000 6979 19002
rect 4981 18944 4986 19000
rect 5042 18944 6918 19000
rect 6974 18944 6979 19000
rect 4981 18942 6979 18944
rect 4981 18939 5047 18942
rect 6913 18939 6979 18942
rect 7649 19002 7715 19005
rect 7782 19002 7788 19004
rect 7649 19000 7788 19002
rect 7649 18944 7654 19000
rect 7710 18944 7788 19000
rect 7649 18942 7788 18944
rect 7649 18939 7715 18942
rect 7782 18940 7788 18942
rect 7852 18940 7858 19004
rect 4061 18866 4127 18869
rect 8526 18866 8586 19078
rect 11462 19076 11468 19078
rect 11532 19076 11538 19140
rect 11697 19138 11763 19141
rect 12198 19138 12204 19140
rect 11697 19136 12204 19138
rect 11697 19080 11702 19136
rect 11758 19080 12204 19136
rect 11697 19078 12204 19080
rect 11697 19075 11763 19078
rect 12198 19076 12204 19078
rect 12268 19138 12274 19140
rect 15101 19138 15167 19141
rect 16481 19140 16547 19141
rect 12268 19136 15167 19138
rect 12268 19080 15106 19136
rect 15162 19080 15167 19136
rect 12268 19078 15167 19080
rect 12268 19076 12274 19078
rect 15101 19075 15167 19078
rect 16430 19076 16436 19140
rect 16500 19138 16547 19140
rect 16500 19136 16592 19138
rect 16542 19080 16592 19136
rect 16500 19078 16592 19080
rect 16500 19076 16547 19078
rect 16982 19076 16988 19140
rect 17052 19138 17058 19140
rect 17769 19138 17835 19141
rect 17052 19136 17835 19138
rect 17052 19080 17774 19136
rect 17830 19080 17835 19136
rect 17052 19078 17835 19080
rect 23614 19138 23674 19214
rect 25129 19272 25268 19274
rect 25129 19216 25134 19272
rect 25190 19216 25268 19272
rect 25129 19214 25268 19216
rect 25129 19211 25195 19214
rect 25262 19212 25268 19214
rect 25332 19212 25338 19276
rect 26734 19138 26740 19140
rect 23614 19078 26740 19138
rect 17052 19076 17058 19078
rect 16481 19075 16547 19076
rect 17769 19075 17835 19078
rect 26734 19076 26740 19078
rect 26804 19076 26810 19140
rect 28993 19138 29059 19141
rect 29310 19138 29316 19140
rect 28993 19136 29316 19138
rect 28993 19080 28998 19136
rect 29054 19080 29316 19136
rect 28993 19078 29316 19080
rect 28993 19075 29059 19078
rect 29310 19076 29316 19078
rect 29380 19076 29386 19140
rect 15574 19072 15890 19073
rect 15574 19008 15580 19072
rect 15644 19008 15660 19072
rect 15724 19008 15740 19072
rect 15804 19008 15820 19072
rect 15884 19008 15890 19072
rect 15574 19007 15890 19008
rect 23164 19072 23480 19073
rect 23164 19008 23170 19072
rect 23234 19008 23250 19072
rect 23314 19008 23330 19072
rect 23394 19008 23410 19072
rect 23474 19008 23480 19072
rect 23164 19007 23480 19008
rect 30754 19072 31070 19073
rect 30754 19008 30760 19072
rect 30824 19008 30840 19072
rect 30904 19008 30920 19072
rect 30984 19008 31000 19072
rect 31064 19008 31070 19072
rect 30754 19007 31070 19008
rect 9254 19002 9260 19004
rect 8664 18942 9260 19002
rect 8664 18869 8724 18942
rect 9254 18940 9260 18942
rect 9324 18940 9330 19004
rect 9673 19002 9739 19005
rect 13445 19002 13511 19005
rect 9673 19000 13511 19002
rect 9673 18944 9678 19000
rect 9734 18944 13450 19000
rect 13506 18944 13511 19000
rect 9673 18942 13511 18944
rect 9673 18939 9739 18942
rect 13445 18939 13511 18942
rect 15101 19002 15167 19005
rect 15326 19002 15332 19004
rect 15101 19000 15332 19002
rect 15101 18944 15106 19000
rect 15162 18944 15332 19000
rect 15101 18942 15332 18944
rect 15101 18939 15167 18942
rect 15326 18940 15332 18942
rect 15396 18940 15402 19004
rect 29637 19002 29703 19005
rect 23982 19000 29703 19002
rect 23982 18944 29642 19000
rect 29698 18944 29703 19000
rect 23982 18942 29703 18944
rect 4061 18864 8586 18866
rect 4061 18808 4066 18864
rect 4122 18808 8586 18864
rect 4061 18806 8586 18808
rect 8661 18864 8727 18869
rect 8661 18808 8666 18864
rect 8722 18808 8727 18864
rect 4061 18803 4127 18806
rect 8661 18803 8727 18808
rect 8845 18866 8911 18869
rect 9305 18866 9371 18869
rect 8845 18864 9371 18866
rect 8845 18808 8850 18864
rect 8906 18808 9310 18864
rect 9366 18808 9371 18864
rect 8845 18806 9371 18808
rect 8845 18803 8911 18806
rect 9305 18803 9371 18806
rect 10225 18866 10291 18869
rect 14549 18866 14615 18869
rect 10225 18864 14615 18866
rect 10225 18808 10230 18864
rect 10286 18808 14554 18864
rect 14610 18808 14615 18864
rect 10225 18806 14615 18808
rect 10225 18803 10291 18806
rect 14549 18803 14615 18806
rect 16062 18804 16068 18868
rect 16132 18866 16138 18868
rect 16665 18866 16731 18869
rect 16132 18864 16731 18866
rect 16132 18808 16670 18864
rect 16726 18808 16731 18864
rect 16132 18806 16731 18808
rect 16132 18804 16138 18806
rect 16665 18803 16731 18806
rect 23381 18866 23447 18869
rect 23982 18866 24042 18942
rect 29637 18939 29703 18942
rect 23381 18864 24042 18866
rect 23381 18808 23386 18864
rect 23442 18808 24042 18864
rect 23381 18806 24042 18808
rect 24209 18866 24275 18869
rect 27889 18866 27955 18869
rect 24209 18864 27955 18866
rect 24209 18808 24214 18864
rect 24270 18808 27894 18864
rect 27950 18808 27955 18864
rect 24209 18806 27955 18808
rect 23381 18803 23447 18806
rect 24209 18803 24275 18806
rect 27889 18803 27955 18806
rect 28993 18866 29059 18869
rect 29177 18866 29243 18869
rect 28993 18864 29243 18866
rect 28993 18808 28998 18864
rect 29054 18808 29182 18864
rect 29238 18808 29243 18864
rect 28993 18806 29243 18808
rect 28993 18803 29059 18806
rect 29177 18803 29243 18806
rect 5349 18730 5415 18733
rect 12566 18730 12572 18732
rect 5349 18728 12572 18730
rect 5349 18672 5354 18728
rect 5410 18672 12572 18728
rect 5349 18670 12572 18672
rect 5349 18667 5415 18670
rect 12566 18668 12572 18670
rect 12636 18668 12642 18732
rect 14273 18730 14339 18733
rect 30281 18730 30347 18733
rect 14273 18728 30347 18730
rect 14273 18672 14278 18728
rect 14334 18672 30286 18728
rect 30342 18672 30347 18728
rect 14273 18670 30347 18672
rect 14273 18667 14339 18670
rect 30281 18667 30347 18670
rect 8937 18594 9003 18597
rect 10961 18594 11027 18597
rect 17493 18594 17559 18597
rect 8937 18592 11027 18594
rect 8937 18536 8942 18592
rect 8998 18536 10966 18592
rect 11022 18536 11027 18592
rect 8937 18534 11027 18536
rect 8937 18531 9003 18534
rect 10961 18531 11027 18534
rect 12390 18592 17559 18594
rect 12390 18536 17498 18592
rect 17554 18536 17559 18592
rect 12390 18534 17559 18536
rect 4189 18528 4505 18529
rect 4189 18464 4195 18528
rect 4259 18464 4275 18528
rect 4339 18464 4355 18528
rect 4419 18464 4435 18528
rect 4499 18464 4505 18528
rect 4189 18463 4505 18464
rect 11779 18528 12095 18529
rect 11779 18464 11785 18528
rect 11849 18464 11865 18528
rect 11929 18464 11945 18528
rect 12009 18464 12025 18528
rect 12089 18464 12095 18528
rect 11779 18463 12095 18464
rect 5942 18396 5948 18460
rect 6012 18458 6018 18460
rect 6453 18458 6519 18461
rect 6012 18456 6519 18458
rect 6012 18400 6458 18456
rect 6514 18400 6519 18456
rect 6012 18398 6519 18400
rect 6012 18396 6018 18398
rect 6453 18395 6519 18398
rect 6729 18458 6795 18461
rect 7649 18460 7715 18461
rect 7414 18458 7420 18460
rect 6729 18456 7420 18458
rect 6729 18400 6734 18456
rect 6790 18400 7420 18456
rect 6729 18398 7420 18400
rect 6729 18395 6795 18398
rect 7414 18396 7420 18398
rect 7484 18396 7490 18460
rect 7598 18396 7604 18460
rect 7668 18458 7715 18460
rect 8753 18458 8819 18461
rect 9397 18458 9463 18461
rect 7668 18456 7760 18458
rect 7710 18400 7760 18456
rect 7668 18398 7760 18400
rect 8753 18456 9463 18458
rect 8753 18400 8758 18456
rect 8814 18400 9402 18456
rect 9458 18400 9463 18456
rect 8753 18398 9463 18400
rect 7668 18396 7715 18398
rect 7649 18395 7715 18396
rect 8753 18395 8819 18398
rect 9397 18395 9463 18398
rect 841 18322 907 18325
rect 12390 18322 12450 18534
rect 17493 18531 17559 18534
rect 22502 18532 22508 18596
rect 22572 18594 22578 18596
rect 22572 18534 24778 18594
rect 22572 18532 22578 18534
rect 19369 18528 19685 18529
rect 19369 18464 19375 18528
rect 19439 18464 19455 18528
rect 19519 18464 19535 18528
rect 19599 18464 19615 18528
rect 19679 18464 19685 18528
rect 19369 18463 19685 18464
rect 13537 18458 13603 18461
rect 19241 18458 19307 18461
rect 21817 18458 21883 18461
rect 23657 18458 23723 18461
rect 13537 18456 19307 18458
rect 13537 18400 13542 18456
rect 13598 18400 19246 18456
rect 19302 18400 19307 18456
rect 13537 18398 19307 18400
rect 13537 18395 13603 18398
rect 19241 18395 19307 18398
rect 20486 18456 23723 18458
rect 20486 18400 21822 18456
rect 21878 18400 23662 18456
rect 23718 18400 23723 18456
rect 20486 18398 23723 18400
rect 841 18320 12450 18322
rect 841 18264 846 18320
rect 902 18264 12450 18320
rect 841 18262 12450 18264
rect 841 18259 907 18262
rect 13670 18260 13676 18324
rect 13740 18322 13746 18324
rect 16389 18322 16455 18325
rect 13740 18320 16455 18322
rect 13740 18264 16394 18320
rect 16450 18264 16455 18320
rect 13740 18262 16455 18264
rect 13740 18260 13746 18262
rect 16389 18259 16455 18262
rect 16849 18322 16915 18325
rect 20486 18322 20546 18398
rect 21817 18395 21883 18398
rect 23657 18395 23723 18398
rect 24158 18396 24164 18460
rect 24228 18458 24234 18460
rect 24485 18458 24551 18461
rect 24228 18456 24551 18458
rect 24228 18400 24490 18456
rect 24546 18400 24551 18456
rect 24228 18398 24551 18400
rect 24228 18396 24234 18398
rect 24485 18395 24551 18398
rect 16849 18320 20546 18322
rect 16849 18264 16854 18320
rect 16910 18264 20546 18320
rect 16849 18262 20546 18264
rect 20713 18322 20779 18325
rect 24393 18322 24459 18325
rect 20713 18320 24459 18322
rect 20713 18264 20718 18320
rect 20774 18264 24398 18320
rect 24454 18264 24459 18320
rect 20713 18262 24459 18264
rect 24718 18322 24778 18534
rect 26959 18528 27275 18529
rect 26959 18464 26965 18528
rect 27029 18464 27045 18528
rect 27109 18464 27125 18528
rect 27189 18464 27205 18528
rect 27269 18464 27275 18528
rect 26959 18463 27275 18464
rect 28349 18460 28415 18461
rect 28349 18458 28396 18460
rect 28304 18456 28396 18458
rect 28304 18400 28354 18456
rect 28304 18398 28396 18400
rect 28349 18396 28396 18398
rect 28460 18396 28466 18460
rect 28349 18395 28415 18396
rect 31385 18322 31451 18325
rect 24718 18320 31451 18322
rect 24718 18264 31390 18320
rect 31446 18264 31451 18320
rect 24718 18262 31451 18264
rect 16849 18259 16915 18262
rect 20713 18259 20779 18262
rect 24393 18259 24459 18262
rect 31385 18259 31451 18262
rect 3969 18186 4035 18189
rect 3969 18184 8586 18186
rect 3969 18128 3974 18184
rect 4030 18128 8586 18184
rect 3969 18126 8586 18128
rect 3969 18123 4035 18126
rect 1669 18050 1735 18053
rect 5349 18052 5415 18053
rect 6453 18052 6519 18053
rect 5206 18050 5212 18052
rect 1669 18048 5212 18050
rect 1669 17992 1674 18048
rect 1730 17992 5212 18048
rect 1669 17990 5212 17992
rect 1669 17987 1735 17990
rect 5206 17988 5212 17990
rect 5276 17988 5282 18052
rect 5349 18048 5396 18052
rect 5460 18050 5466 18052
rect 6453 18050 6500 18052
rect 5349 17992 5354 18048
rect 5349 17988 5396 17992
rect 5460 17990 5506 18050
rect 6408 18048 6500 18050
rect 6408 17992 6458 18048
rect 6408 17990 6500 17992
rect 5460 17988 5466 17990
rect 6453 17988 6500 17990
rect 6564 17988 6570 18052
rect 7046 17988 7052 18052
rect 7116 18050 7122 18052
rect 7741 18050 7807 18053
rect 7116 18048 7807 18050
rect 7116 17992 7746 18048
rect 7802 17992 7807 18048
rect 7116 17990 7807 17992
rect 8526 18050 8586 18126
rect 9438 18124 9444 18188
rect 9508 18186 9514 18188
rect 16113 18186 16179 18189
rect 9508 18184 16179 18186
rect 9508 18128 16118 18184
rect 16174 18128 16179 18184
rect 9508 18126 16179 18128
rect 9508 18124 9514 18126
rect 16113 18123 16179 18126
rect 17125 18186 17191 18189
rect 23381 18186 23447 18189
rect 17125 18184 23447 18186
rect 17125 18128 17130 18184
rect 17186 18128 23386 18184
rect 23442 18128 23447 18184
rect 17125 18126 23447 18128
rect 17125 18123 17191 18126
rect 23381 18123 23447 18126
rect 23565 18186 23631 18189
rect 27613 18186 27679 18189
rect 23565 18184 27679 18186
rect 23565 18128 23570 18184
rect 23626 18128 27618 18184
rect 27674 18128 27679 18184
rect 23565 18126 27679 18128
rect 23565 18123 23631 18126
rect 27613 18123 27679 18126
rect 15142 18050 15148 18052
rect 8526 17990 15148 18050
rect 7116 17988 7122 17990
rect 5349 17987 5415 17988
rect 6453 17987 6519 17988
rect 7741 17987 7807 17990
rect 15142 17988 15148 17990
rect 15212 17988 15218 18052
rect 17493 18050 17559 18053
rect 20897 18050 20963 18053
rect 17493 18048 20963 18050
rect 17493 17992 17498 18048
rect 17554 17992 20902 18048
rect 20958 17992 20963 18048
rect 17493 17990 20963 17992
rect 17493 17987 17559 17990
rect 20897 17987 20963 17990
rect 24158 17988 24164 18052
rect 24228 18050 24234 18052
rect 26233 18050 26299 18053
rect 24228 18048 26299 18050
rect 24228 17992 26238 18048
rect 26294 17992 26299 18048
rect 24228 17990 26299 17992
rect 24228 17988 24234 17990
rect 26233 17987 26299 17990
rect 30373 18052 30439 18053
rect 30373 18048 30420 18052
rect 30484 18050 30490 18052
rect 30373 17992 30378 18048
rect 30373 17988 30420 17992
rect 30484 17990 30530 18050
rect 30484 17988 30490 17990
rect 30373 17987 30439 17988
rect 7984 17984 8300 17985
rect 7984 17920 7990 17984
rect 8054 17920 8070 17984
rect 8134 17920 8150 17984
rect 8214 17920 8230 17984
rect 8294 17920 8300 17984
rect 7984 17919 8300 17920
rect 15574 17984 15890 17985
rect 15574 17920 15580 17984
rect 15644 17920 15660 17984
rect 15724 17920 15740 17984
rect 15804 17920 15820 17984
rect 15884 17920 15890 17984
rect 15574 17919 15890 17920
rect 23164 17984 23480 17985
rect 23164 17920 23170 17984
rect 23234 17920 23250 17984
rect 23314 17920 23330 17984
rect 23394 17920 23410 17984
rect 23474 17920 23480 17984
rect 23164 17919 23480 17920
rect 30754 17984 31070 17985
rect 30754 17920 30760 17984
rect 30824 17920 30840 17984
rect 30904 17920 30920 17984
rect 30984 17920 31000 17984
rect 31064 17920 31070 17984
rect 30754 17919 31070 17920
rect 8569 17914 8635 17917
rect 9397 17914 9463 17917
rect 8569 17912 9463 17914
rect 8569 17856 8574 17912
rect 8630 17856 9402 17912
rect 9458 17856 9463 17912
rect 8569 17854 9463 17856
rect 8569 17851 8635 17854
rect 9397 17851 9463 17854
rect 16062 17852 16068 17916
rect 16132 17914 16138 17916
rect 16757 17914 16823 17917
rect 16132 17912 16823 17914
rect 16132 17856 16762 17912
rect 16818 17856 16823 17912
rect 16132 17854 16823 17856
rect 16132 17852 16138 17854
rect 16757 17851 16823 17854
rect 18505 17914 18571 17917
rect 22553 17914 22619 17917
rect 18505 17912 22619 17914
rect 18505 17856 18510 17912
rect 18566 17856 22558 17912
rect 22614 17856 22619 17912
rect 18505 17854 22619 17856
rect 18505 17851 18571 17854
rect 22553 17851 22619 17854
rect 24761 17914 24827 17917
rect 26601 17914 26667 17917
rect 24761 17912 26667 17914
rect 24761 17856 24766 17912
rect 24822 17856 26606 17912
rect 26662 17856 26667 17912
rect 24761 17854 26667 17856
rect 24761 17851 24827 17854
rect 26601 17851 26667 17854
rect 3693 17778 3759 17781
rect 5809 17778 5875 17781
rect 7373 17778 7439 17781
rect 3693 17776 7439 17778
rect 3693 17720 3698 17776
rect 3754 17720 5814 17776
rect 5870 17720 7378 17776
rect 7434 17720 7439 17776
rect 3693 17718 7439 17720
rect 3693 17715 3759 17718
rect 5809 17715 5875 17718
rect 7373 17715 7439 17718
rect 8201 17778 8267 17781
rect 20713 17778 20779 17781
rect 8201 17776 20779 17778
rect 8201 17720 8206 17776
rect 8262 17720 20718 17776
rect 20774 17720 20779 17776
rect 8201 17718 20779 17720
rect 8201 17715 8267 17718
rect 20713 17715 20779 17718
rect 21081 17778 21147 17781
rect 25313 17778 25379 17781
rect 21081 17776 25379 17778
rect 21081 17720 21086 17776
rect 21142 17720 25318 17776
rect 25374 17720 25379 17776
rect 21081 17718 25379 17720
rect 21081 17715 21147 17718
rect 25313 17715 25379 17718
rect 26049 17778 26115 17781
rect 28901 17778 28967 17781
rect 26049 17776 28967 17778
rect 26049 17720 26054 17776
rect 26110 17720 28906 17776
rect 28962 17720 28967 17776
rect 26049 17718 28967 17720
rect 26049 17715 26115 17718
rect 28901 17715 28967 17718
rect 1669 17642 1735 17645
rect 2773 17642 2839 17645
rect 10133 17642 10199 17645
rect 15469 17642 15535 17645
rect 29494 17642 29500 17644
rect 1669 17640 10199 17642
rect 1669 17584 1674 17640
rect 1730 17584 2778 17640
rect 2834 17584 10138 17640
rect 10194 17584 10199 17640
rect 1669 17582 10199 17584
rect 1669 17579 1735 17582
rect 2773 17579 2839 17582
rect 10133 17579 10199 17582
rect 10734 17582 12450 17642
rect 5717 17506 5783 17509
rect 10593 17506 10659 17509
rect 5717 17504 10659 17506
rect 5717 17448 5722 17504
rect 5778 17448 10598 17504
rect 10654 17448 10659 17504
rect 5717 17446 10659 17448
rect 5717 17443 5783 17446
rect 10593 17443 10659 17446
rect 4189 17440 4505 17441
rect 4189 17376 4195 17440
rect 4259 17376 4275 17440
rect 4339 17376 4355 17440
rect 4419 17376 4435 17440
rect 4499 17376 4505 17440
rect 4189 17375 4505 17376
rect 6821 17370 6887 17373
rect 10734 17370 10794 17582
rect 11779 17440 12095 17441
rect 11779 17376 11785 17440
rect 11849 17376 11865 17440
rect 11929 17376 11945 17440
rect 12009 17376 12025 17440
rect 12089 17376 12095 17440
rect 11779 17375 12095 17376
rect 6821 17368 10794 17370
rect 6821 17312 6826 17368
rect 6882 17312 10794 17368
rect 6821 17310 10794 17312
rect 6821 17307 6887 17310
rect 3785 17234 3851 17237
rect 12249 17234 12315 17237
rect 3785 17232 12315 17234
rect 3785 17176 3790 17232
rect 3846 17176 12254 17232
rect 12310 17176 12315 17232
rect 3785 17174 12315 17176
rect 12390 17234 12450 17582
rect 15469 17640 29500 17642
rect 15469 17584 15474 17640
rect 15530 17584 29500 17640
rect 15469 17582 29500 17584
rect 15469 17579 15535 17582
rect 29494 17580 29500 17582
rect 29564 17642 29570 17644
rect 30373 17642 30439 17645
rect 29564 17640 30439 17642
rect 29564 17584 30378 17640
rect 30434 17584 30439 17640
rect 29564 17582 30439 17584
rect 29564 17580 29570 17582
rect 30373 17579 30439 17582
rect 21173 17506 21239 17509
rect 26049 17506 26115 17509
rect 21173 17504 26115 17506
rect 21173 17448 21178 17504
rect 21234 17448 26054 17504
rect 26110 17448 26115 17504
rect 21173 17446 26115 17448
rect 21173 17443 21239 17446
rect 26049 17443 26115 17446
rect 19369 17440 19685 17441
rect 19369 17376 19375 17440
rect 19439 17376 19455 17440
rect 19519 17376 19535 17440
rect 19599 17376 19615 17440
rect 19679 17376 19685 17440
rect 19369 17375 19685 17376
rect 26959 17440 27275 17441
rect 26959 17376 26965 17440
rect 27029 17376 27045 17440
rect 27109 17376 27125 17440
rect 27189 17376 27205 17440
rect 27269 17376 27275 17440
rect 26959 17375 27275 17376
rect 21633 17370 21699 17373
rect 25221 17370 25287 17373
rect 21633 17368 25287 17370
rect 21633 17312 21638 17368
rect 21694 17312 25226 17368
rect 25282 17312 25287 17368
rect 21633 17310 25287 17312
rect 21633 17307 21699 17310
rect 25221 17307 25287 17310
rect 20621 17234 20687 17237
rect 12390 17232 20687 17234
rect 12390 17176 20626 17232
rect 20682 17176 20687 17232
rect 12390 17174 20687 17176
rect 3785 17171 3851 17174
rect 12249 17171 12315 17174
rect 20621 17171 20687 17174
rect 21173 17234 21239 17237
rect 28349 17234 28415 17237
rect 21173 17232 28415 17234
rect 21173 17176 21178 17232
rect 21234 17176 28354 17232
rect 28410 17176 28415 17232
rect 21173 17174 28415 17176
rect 21173 17171 21239 17174
rect 28349 17171 28415 17174
rect 6821 17096 6887 17101
rect 6821 17040 6826 17096
rect 6882 17040 6887 17096
rect 6821 17035 6887 17040
rect 7097 17098 7163 17101
rect 16205 17098 16271 17101
rect 24577 17098 24643 17101
rect 7097 17096 12450 17098
rect 7097 17040 7102 17096
rect 7158 17040 12450 17096
rect 7097 17038 12450 17040
rect 7097 17035 7163 17038
rect 2773 16826 2839 16829
rect 6824 16826 6884 17035
rect 8661 16964 8727 16965
rect 8661 16962 8708 16964
rect 8616 16960 8708 16962
rect 8616 16904 8666 16960
rect 8616 16902 8708 16904
rect 8661 16900 8708 16902
rect 8772 16900 8778 16964
rect 12390 16962 12450 17038
rect 16205 17096 24643 17098
rect 16205 17040 16210 17096
rect 16266 17040 24582 17096
rect 24638 17040 24643 17096
rect 16205 17038 24643 17040
rect 16205 17035 16271 17038
rect 24577 17035 24643 17038
rect 28993 17098 29059 17101
rect 30373 17098 30439 17101
rect 30741 17098 30807 17101
rect 28993 17096 30439 17098
rect 28993 17040 28998 17096
rect 29054 17040 30378 17096
rect 30434 17040 30439 17096
rect 28993 17038 30439 17040
rect 28993 17035 29059 17038
rect 30373 17035 30439 17038
rect 30606 17096 30807 17098
rect 30606 17040 30746 17096
rect 30802 17040 30807 17096
rect 30606 17038 30807 17040
rect 15193 16962 15259 16965
rect 12390 16960 15259 16962
rect 12390 16904 15198 16960
rect 15254 16904 15259 16960
rect 12390 16902 15259 16904
rect 8661 16899 8727 16900
rect 15193 16899 15259 16902
rect 19425 16962 19491 16965
rect 23013 16962 23079 16965
rect 19425 16960 23079 16962
rect 19425 16904 19430 16960
rect 19486 16904 23018 16960
rect 23074 16904 23079 16960
rect 19425 16902 23079 16904
rect 19425 16899 19491 16902
rect 23013 16899 23079 16902
rect 27470 16900 27476 16964
rect 27540 16962 27546 16964
rect 27705 16962 27771 16965
rect 27540 16960 27771 16962
rect 27540 16904 27710 16960
rect 27766 16904 27771 16960
rect 27540 16902 27771 16904
rect 27540 16900 27546 16902
rect 27705 16899 27771 16902
rect 7984 16896 8300 16897
rect 7984 16832 7990 16896
rect 8054 16832 8070 16896
rect 8134 16832 8150 16896
rect 8214 16832 8230 16896
rect 8294 16832 8300 16896
rect 7984 16831 8300 16832
rect 15574 16896 15890 16897
rect 15574 16832 15580 16896
rect 15644 16832 15660 16896
rect 15724 16832 15740 16896
rect 15804 16832 15820 16896
rect 15884 16832 15890 16896
rect 15574 16831 15890 16832
rect 23164 16896 23480 16897
rect 23164 16832 23170 16896
rect 23234 16832 23250 16896
rect 23314 16832 23330 16896
rect 23394 16832 23410 16896
rect 23474 16832 23480 16896
rect 23164 16831 23480 16832
rect 2773 16824 6884 16826
rect 2773 16768 2778 16824
rect 2834 16768 6884 16824
rect 2773 16766 6884 16768
rect 8569 16826 8635 16829
rect 10409 16826 10475 16829
rect 8569 16824 10475 16826
rect 8569 16768 8574 16824
rect 8630 16768 10414 16824
rect 10470 16768 10475 16824
rect 8569 16766 10475 16768
rect 2773 16763 2839 16766
rect 8569 16763 8635 16766
rect 10409 16763 10475 16766
rect 19977 16826 20043 16829
rect 22737 16826 22803 16829
rect 19977 16824 22803 16826
rect 19977 16768 19982 16824
rect 20038 16768 22742 16824
rect 22798 16768 22803 16824
rect 19977 16766 22803 16768
rect 19977 16763 20043 16766
rect 22737 16763 22803 16766
rect 26182 16764 26188 16828
rect 26252 16826 26258 16828
rect 29637 16826 29703 16829
rect 26252 16824 29703 16826
rect 26252 16768 29642 16824
rect 29698 16768 29703 16824
rect 26252 16766 29703 16768
rect 26252 16764 26258 16766
rect 29637 16763 29703 16766
rect 6545 16690 6611 16693
rect 8477 16690 8543 16693
rect 9489 16690 9555 16693
rect 6545 16688 8218 16690
rect 6545 16632 6550 16688
rect 6606 16632 8218 16688
rect 6545 16630 8218 16632
rect 6545 16627 6611 16630
rect 2037 16554 2103 16557
rect 8158 16554 8218 16630
rect 8477 16688 9555 16690
rect 8477 16632 8482 16688
rect 8538 16632 9494 16688
rect 9550 16632 9555 16688
rect 8477 16630 9555 16632
rect 8477 16627 8543 16630
rect 9489 16627 9555 16630
rect 10726 16628 10732 16692
rect 10796 16690 10802 16692
rect 11697 16690 11763 16693
rect 10796 16688 11763 16690
rect 10796 16632 11702 16688
rect 11758 16632 11763 16688
rect 10796 16630 11763 16632
rect 10796 16628 10802 16630
rect 11697 16627 11763 16630
rect 14549 16690 14615 16693
rect 18781 16690 18847 16693
rect 14549 16688 18847 16690
rect 14549 16632 14554 16688
rect 14610 16632 18786 16688
rect 18842 16632 18847 16688
rect 14549 16630 18847 16632
rect 14549 16627 14615 16630
rect 18781 16627 18847 16630
rect 21081 16690 21147 16693
rect 27981 16690 28047 16693
rect 21081 16688 28047 16690
rect 21081 16632 21086 16688
rect 21142 16632 27986 16688
rect 28042 16632 28047 16688
rect 21081 16630 28047 16632
rect 21081 16627 21147 16630
rect 27981 16627 28047 16630
rect 29545 16690 29611 16693
rect 29678 16690 29684 16692
rect 29545 16688 29684 16690
rect 29545 16632 29550 16688
rect 29606 16632 29684 16688
rect 29545 16630 29684 16632
rect 29545 16627 29611 16630
rect 29678 16628 29684 16630
rect 29748 16628 29754 16692
rect 16113 16554 16179 16557
rect 2037 16552 8034 16554
rect 2037 16496 2042 16552
rect 2098 16496 8034 16552
rect 2037 16494 8034 16496
rect 8158 16552 16179 16554
rect 8158 16496 16118 16552
rect 16174 16496 16179 16552
rect 8158 16494 16179 16496
rect 2037 16491 2103 16494
rect 7974 16418 8034 16494
rect 16113 16491 16179 16494
rect 16297 16554 16363 16557
rect 20713 16554 20779 16557
rect 16297 16552 20779 16554
rect 16297 16496 16302 16552
rect 16358 16496 20718 16552
rect 20774 16496 20779 16552
rect 16297 16494 20779 16496
rect 16297 16491 16363 16494
rect 20713 16491 20779 16494
rect 24025 16554 24091 16557
rect 28257 16554 28323 16557
rect 24025 16552 28323 16554
rect 24025 16496 24030 16552
rect 24086 16496 28262 16552
rect 28318 16496 28323 16552
rect 24025 16494 28323 16496
rect 24025 16491 24091 16494
rect 28257 16491 28323 16494
rect 28533 16554 28599 16557
rect 30606 16554 30666 17038
rect 30741 17035 30807 17038
rect 30754 16896 31070 16897
rect 30754 16832 30760 16896
rect 30824 16832 30840 16896
rect 30904 16832 30920 16896
rect 30984 16832 31000 16896
rect 31064 16832 31070 16896
rect 30754 16831 31070 16832
rect 28533 16552 30666 16554
rect 28533 16496 28538 16552
rect 28594 16496 30666 16552
rect 28533 16494 30666 16496
rect 28533 16491 28599 16494
rect 8518 16418 8524 16420
rect 7974 16358 8524 16418
rect 8518 16356 8524 16358
rect 8588 16356 8594 16420
rect 9029 16418 9095 16421
rect 9438 16418 9444 16420
rect 9029 16416 9444 16418
rect 9029 16360 9034 16416
rect 9090 16360 9444 16416
rect 9029 16358 9444 16360
rect 9029 16355 9095 16358
rect 9438 16356 9444 16358
rect 9508 16356 9514 16420
rect 27429 16418 27495 16421
rect 29821 16418 29887 16421
rect 27429 16416 29887 16418
rect 27429 16360 27434 16416
rect 27490 16360 29826 16416
rect 29882 16360 29887 16416
rect 27429 16358 29887 16360
rect 27429 16355 27495 16358
rect 29821 16355 29887 16358
rect 4189 16352 4505 16353
rect 4189 16288 4195 16352
rect 4259 16288 4275 16352
rect 4339 16288 4355 16352
rect 4419 16288 4435 16352
rect 4499 16288 4505 16352
rect 4189 16287 4505 16288
rect 11779 16352 12095 16353
rect 11779 16288 11785 16352
rect 11849 16288 11865 16352
rect 11929 16288 11945 16352
rect 12009 16288 12025 16352
rect 12089 16288 12095 16352
rect 11779 16287 12095 16288
rect 19369 16352 19685 16353
rect 19369 16288 19375 16352
rect 19439 16288 19455 16352
rect 19519 16288 19535 16352
rect 19599 16288 19615 16352
rect 19679 16288 19685 16352
rect 19369 16287 19685 16288
rect 26959 16352 27275 16353
rect 26959 16288 26965 16352
rect 27029 16288 27045 16352
rect 27109 16288 27125 16352
rect 27189 16288 27205 16352
rect 27269 16288 27275 16352
rect 26959 16287 27275 16288
rect 13169 16282 13235 16285
rect 14457 16282 14523 16285
rect 17401 16282 17467 16285
rect 24158 16282 24164 16284
rect 4616 16222 9874 16282
rect 3049 16146 3115 16149
rect 4616 16146 4676 16222
rect 3049 16144 4676 16146
rect 3049 16088 3054 16144
rect 3110 16088 4676 16144
rect 3049 16086 4676 16088
rect 4889 16146 4955 16149
rect 5441 16146 5507 16149
rect 9673 16146 9739 16149
rect 4889 16144 5274 16146
rect 4889 16088 4894 16144
rect 4950 16088 5274 16144
rect 4889 16086 5274 16088
rect 3049 16083 3115 16086
rect 4889 16083 4955 16086
rect 5214 16010 5274 16086
rect 5441 16144 9739 16146
rect 5441 16088 5446 16144
rect 5502 16088 9678 16144
rect 9734 16088 9739 16144
rect 5441 16086 9739 16088
rect 5441 16083 5507 16086
rect 9673 16083 9739 16086
rect 7005 16010 7071 16013
rect 5214 16008 7071 16010
rect 5214 15952 7010 16008
rect 7066 15952 7071 16008
rect 5214 15950 7071 15952
rect 7005 15947 7071 15950
rect 8293 16010 8359 16013
rect 9814 16010 9874 16222
rect 13169 16280 17467 16282
rect 13169 16224 13174 16280
rect 13230 16224 14462 16280
rect 14518 16224 17406 16280
rect 17462 16224 17467 16280
rect 13169 16222 17467 16224
rect 13169 16219 13235 16222
rect 14457 16219 14523 16222
rect 17401 16219 17467 16222
rect 19750 16222 24164 16282
rect 11053 16146 11119 16149
rect 12341 16146 12407 16149
rect 11053 16144 12407 16146
rect 11053 16088 11058 16144
rect 11114 16088 12346 16144
rect 12402 16088 12407 16144
rect 11053 16086 12407 16088
rect 11053 16083 11119 16086
rect 12341 16083 12407 16086
rect 17033 16146 17099 16149
rect 17401 16146 17467 16149
rect 19750 16146 19810 16222
rect 24158 16220 24164 16222
rect 24228 16220 24234 16284
rect 29453 16282 29519 16285
rect 29318 16280 29519 16282
rect 29318 16224 29458 16280
rect 29514 16224 29519 16280
rect 29318 16222 29519 16224
rect 29318 16149 29378 16222
rect 29453 16219 29519 16222
rect 17033 16144 19810 16146
rect 17033 16088 17038 16144
rect 17094 16088 17406 16144
rect 17462 16088 19810 16144
rect 17033 16086 19810 16088
rect 20529 16146 20595 16149
rect 25313 16146 25379 16149
rect 20529 16144 25379 16146
rect 20529 16088 20534 16144
rect 20590 16088 25318 16144
rect 25374 16088 25379 16144
rect 20529 16086 25379 16088
rect 17033 16083 17099 16086
rect 17401 16083 17467 16086
rect 20529 16083 20595 16086
rect 25313 16083 25379 16086
rect 25865 16146 25931 16149
rect 26969 16146 27035 16149
rect 25865 16144 27035 16146
rect 25865 16088 25870 16144
rect 25926 16088 26974 16144
rect 27030 16088 27035 16144
rect 25865 16086 27035 16088
rect 29318 16144 29427 16149
rect 29318 16088 29366 16144
rect 29422 16088 29427 16144
rect 29318 16086 29427 16088
rect 25865 16083 25931 16086
rect 26969 16083 27035 16086
rect 29361 16083 29427 16086
rect 30005 16010 30071 16013
rect 8293 16008 9506 16010
rect 8293 15952 8298 16008
rect 8354 15952 9506 16008
rect 8293 15950 9506 15952
rect 9814 16008 30071 16010
rect 9814 15952 30010 16008
rect 30066 15952 30071 16008
rect 9814 15950 30071 15952
rect 8293 15947 8359 15950
rect 3049 15874 3115 15877
rect 7097 15874 7163 15877
rect 3049 15872 7163 15874
rect 3049 15816 3054 15872
rect 3110 15816 7102 15872
rect 7158 15816 7163 15872
rect 3049 15814 7163 15816
rect 9446 15874 9506 15950
rect 30005 15947 30071 15950
rect 12985 15874 13051 15877
rect 9446 15872 13051 15874
rect 9446 15816 12990 15872
rect 13046 15816 13051 15872
rect 9446 15814 13051 15816
rect 3049 15811 3115 15814
rect 7097 15811 7163 15814
rect 12985 15811 13051 15814
rect 24761 15874 24827 15877
rect 28257 15874 28323 15877
rect 24761 15872 28323 15874
rect 24761 15816 24766 15872
rect 24822 15816 28262 15872
rect 28318 15816 28323 15872
rect 24761 15814 28323 15816
rect 24761 15811 24827 15814
rect 28257 15811 28323 15814
rect 29310 15812 29316 15876
rect 29380 15874 29386 15876
rect 29637 15874 29703 15877
rect 29380 15872 29703 15874
rect 29380 15816 29642 15872
rect 29698 15816 29703 15872
rect 29380 15814 29703 15816
rect 29380 15812 29386 15814
rect 29637 15811 29703 15814
rect 7984 15808 8300 15809
rect 7984 15744 7990 15808
rect 8054 15744 8070 15808
rect 8134 15744 8150 15808
rect 8214 15744 8230 15808
rect 8294 15744 8300 15808
rect 7984 15743 8300 15744
rect 15574 15808 15890 15809
rect 15574 15744 15580 15808
rect 15644 15744 15660 15808
rect 15724 15744 15740 15808
rect 15804 15744 15820 15808
rect 15884 15744 15890 15808
rect 15574 15743 15890 15744
rect 23164 15808 23480 15809
rect 23164 15744 23170 15808
rect 23234 15744 23250 15808
rect 23314 15744 23330 15808
rect 23394 15744 23410 15808
rect 23474 15744 23480 15808
rect 23164 15743 23480 15744
rect 30754 15808 31070 15809
rect 30754 15744 30760 15808
rect 30824 15744 30840 15808
rect 30904 15744 30920 15808
rect 30984 15744 31000 15808
rect 31064 15744 31070 15808
rect 30754 15743 31070 15744
rect 10317 15738 10383 15741
rect 11145 15738 11211 15741
rect 24485 15738 24551 15741
rect 27705 15738 27771 15741
rect 10317 15736 13508 15738
rect 10317 15680 10322 15736
rect 10378 15680 11150 15736
rect 11206 15680 13508 15736
rect 10317 15678 13508 15680
rect 10317 15675 10383 15678
rect 11145 15675 11211 15678
rect 2037 15602 2103 15605
rect 13261 15602 13327 15605
rect 2037 15600 13327 15602
rect 2037 15544 2042 15600
rect 2098 15544 13266 15600
rect 13322 15544 13327 15600
rect 2037 15542 13327 15544
rect 2037 15539 2103 15542
rect 13261 15539 13327 15542
rect 2497 15466 2563 15469
rect 9438 15466 9444 15468
rect 2497 15464 9444 15466
rect 2497 15408 2502 15464
rect 2558 15408 9444 15464
rect 2497 15406 9444 15408
rect 2497 15403 2563 15406
rect 9438 15404 9444 15406
rect 9508 15404 9514 15468
rect 9622 15404 9628 15468
rect 9692 15466 9698 15468
rect 11053 15466 11119 15469
rect 9692 15464 11119 15466
rect 9692 15408 11058 15464
rect 11114 15408 11119 15464
rect 9692 15406 11119 15408
rect 13448 15466 13508 15678
rect 24485 15736 27771 15738
rect 24485 15680 24490 15736
rect 24546 15680 27710 15736
rect 27766 15680 27771 15736
rect 24485 15678 27771 15680
rect 24485 15675 24551 15678
rect 27705 15675 27771 15678
rect 27889 15738 27955 15741
rect 30005 15738 30071 15741
rect 27889 15736 30071 15738
rect 27889 15680 27894 15736
rect 27950 15680 30010 15736
rect 30066 15680 30071 15736
rect 27889 15678 30071 15680
rect 27889 15675 27955 15678
rect 30005 15675 30071 15678
rect 16849 15602 16915 15605
rect 28533 15602 28599 15605
rect 16849 15600 28599 15602
rect 16849 15544 16854 15600
rect 16910 15544 28538 15600
rect 28594 15544 28599 15600
rect 16849 15542 28599 15544
rect 16849 15539 16915 15542
rect 20345 15466 20411 15469
rect 27889 15466 27955 15469
rect 13448 15464 27955 15466
rect 13448 15408 20350 15464
rect 20406 15408 27894 15464
rect 27950 15408 27955 15464
rect 13448 15406 27955 15408
rect 9692 15404 9698 15406
rect 11053 15403 11119 15406
rect 20345 15403 20411 15406
rect 27889 15403 27955 15406
rect 5441 15330 5507 15333
rect 6821 15330 6887 15333
rect 5441 15328 6887 15330
rect 5441 15272 5446 15328
rect 5502 15272 6826 15328
rect 6882 15272 6887 15328
rect 5441 15270 6887 15272
rect 5441 15267 5507 15270
rect 6821 15267 6887 15270
rect 7005 15330 7071 15333
rect 9121 15330 9187 15333
rect 7005 15328 9187 15330
rect 7005 15272 7010 15328
rect 7066 15272 9126 15328
rect 9182 15272 9187 15328
rect 7005 15270 9187 15272
rect 7005 15267 7071 15270
rect 9121 15267 9187 15270
rect 9581 15330 9647 15333
rect 11145 15330 11211 15333
rect 9581 15328 11211 15330
rect 9581 15272 9586 15328
rect 9642 15272 11150 15328
rect 11206 15272 11211 15328
rect 9581 15270 11211 15272
rect 9581 15267 9647 15270
rect 11145 15267 11211 15270
rect 27613 15328 27679 15333
rect 27613 15272 27618 15328
rect 27674 15272 27679 15328
rect 27613 15267 27679 15272
rect 28030 15330 28090 15542
rect 28533 15539 28599 15542
rect 29545 15602 29611 15605
rect 29678 15602 29684 15604
rect 29545 15600 29684 15602
rect 29545 15544 29550 15600
rect 29606 15544 29684 15600
rect 29545 15542 29684 15544
rect 29545 15539 29611 15542
rect 29678 15540 29684 15542
rect 29748 15540 29754 15604
rect 30414 15540 30420 15604
rect 30484 15602 30490 15604
rect 30741 15602 30807 15605
rect 30484 15600 30807 15602
rect 30484 15544 30746 15600
rect 30802 15544 30807 15600
rect 30484 15542 30807 15544
rect 30484 15540 30490 15542
rect 30741 15539 30807 15542
rect 29126 15466 29132 15468
rect 28950 15406 29132 15466
rect 28165 15330 28231 15333
rect 28030 15328 28231 15330
rect 28030 15272 28170 15328
rect 28226 15272 28231 15328
rect 28030 15270 28231 15272
rect 28165 15267 28231 15270
rect 4189 15264 4505 15265
rect 4189 15200 4195 15264
rect 4259 15200 4275 15264
rect 4339 15200 4355 15264
rect 4419 15200 4435 15264
rect 4499 15200 4505 15264
rect 4189 15199 4505 15200
rect 11779 15264 12095 15265
rect 11779 15200 11785 15264
rect 11849 15200 11865 15264
rect 11929 15200 11945 15264
rect 12009 15200 12025 15264
rect 12089 15200 12095 15264
rect 11779 15199 12095 15200
rect 19369 15264 19685 15265
rect 19369 15200 19375 15264
rect 19439 15200 19455 15264
rect 19519 15200 19535 15264
rect 19599 15200 19615 15264
rect 19679 15200 19685 15264
rect 19369 15199 19685 15200
rect 26959 15264 27275 15265
rect 26959 15200 26965 15264
rect 27029 15200 27045 15264
rect 27109 15200 27125 15264
rect 27189 15200 27205 15264
rect 27269 15200 27275 15264
rect 26959 15199 27275 15200
rect 5717 15194 5783 15197
rect 7373 15194 7439 15197
rect 5717 15192 7439 15194
rect 5717 15136 5722 15192
rect 5778 15136 7378 15192
rect 7434 15136 7439 15192
rect 5717 15134 7439 15136
rect 5717 15131 5783 15134
rect 7373 15131 7439 15134
rect 7557 15194 7623 15197
rect 11053 15194 11119 15197
rect 7557 15192 11119 15194
rect 7557 15136 7562 15192
rect 7618 15136 11058 15192
rect 11114 15136 11119 15192
rect 7557 15134 11119 15136
rect 7557 15131 7623 15134
rect 11053 15131 11119 15134
rect 14457 15194 14523 15197
rect 15142 15194 15148 15196
rect 14457 15192 15148 15194
rect 14457 15136 14462 15192
rect 14518 15136 15148 15192
rect 14457 15134 15148 15136
rect 14457 15131 14523 15134
rect 15142 15132 15148 15134
rect 15212 15132 15218 15196
rect 20897 15194 20963 15197
rect 23841 15194 23907 15197
rect 20897 15192 23907 15194
rect 20897 15136 20902 15192
rect 20958 15136 23846 15192
rect 23902 15136 23907 15192
rect 20897 15134 23907 15136
rect 27616 15194 27676 15267
rect 28950 15194 29010 15406
rect 29126 15404 29132 15406
rect 29196 15404 29202 15468
rect 29453 15332 29519 15333
rect 29453 15330 29500 15332
rect 29408 15328 29500 15330
rect 29408 15272 29458 15328
rect 29408 15270 29500 15272
rect 29453 15268 29500 15270
rect 29564 15268 29570 15332
rect 29453 15267 29519 15268
rect 27616 15134 29010 15194
rect 20897 15131 20963 15134
rect 23841 15131 23907 15134
rect 2129 15058 2195 15061
rect 7557 15058 7623 15061
rect 2129 15056 7623 15058
rect 2129 15000 2134 15056
rect 2190 15000 7562 15056
rect 7618 15000 7623 15056
rect 2129 14998 7623 15000
rect 2129 14995 2195 14998
rect 7557 14995 7623 14998
rect 7925 15058 7991 15061
rect 13537 15058 13603 15061
rect 7925 15056 13603 15058
rect 7925 15000 7930 15056
rect 7986 15000 13542 15056
rect 13598 15000 13603 15056
rect 7925 14998 13603 15000
rect 7925 14995 7991 14998
rect 13537 14995 13603 14998
rect 17125 15058 17191 15061
rect 26182 15058 26188 15060
rect 17125 15056 26188 15058
rect 17125 15000 17130 15056
rect 17186 15000 26188 15056
rect 17125 14998 26188 15000
rect 17125 14995 17191 14998
rect 26182 14996 26188 14998
rect 26252 14996 26258 15060
rect 26734 14996 26740 15060
rect 26804 15058 26810 15060
rect 30373 15058 30439 15061
rect 26804 15056 30439 15058
rect 26804 15000 30378 15056
rect 30434 15000 30439 15056
rect 26804 14998 30439 15000
rect 26804 14996 26810 14998
rect 30373 14995 30439 14998
rect 1761 14922 1827 14925
rect 10501 14922 10567 14925
rect 1761 14920 10567 14922
rect 1761 14864 1766 14920
rect 1822 14864 10506 14920
rect 10562 14864 10567 14920
rect 1761 14862 10567 14864
rect 1761 14859 1827 14862
rect 10501 14859 10567 14862
rect 10685 14922 10751 14925
rect 12801 14922 12867 14925
rect 10685 14920 12867 14922
rect 10685 14864 10690 14920
rect 10746 14864 12806 14920
rect 12862 14864 12867 14920
rect 10685 14862 12867 14864
rect 10685 14859 10751 14862
rect 12801 14859 12867 14862
rect 14549 14922 14615 14925
rect 16573 14922 16639 14925
rect 26325 14922 26391 14925
rect 14549 14920 26391 14922
rect 14549 14864 14554 14920
rect 14610 14864 16578 14920
rect 16634 14864 26330 14920
rect 26386 14864 26391 14920
rect 14549 14862 26391 14864
rect 14549 14859 14615 14862
rect 16573 14859 16639 14862
rect 26325 14859 26391 14862
rect 27654 14860 27660 14924
rect 27724 14922 27730 14924
rect 28625 14922 28691 14925
rect 27724 14920 28691 14922
rect 27724 14864 28630 14920
rect 28686 14864 28691 14920
rect 27724 14862 28691 14864
rect 27724 14860 27730 14862
rect 28625 14859 28691 14862
rect 6177 14786 6243 14789
rect 7189 14786 7255 14789
rect 6177 14784 7255 14786
rect 6177 14728 6182 14784
rect 6238 14728 7194 14784
rect 7250 14728 7255 14784
rect 6177 14726 7255 14728
rect 6177 14723 6243 14726
rect 7189 14723 7255 14726
rect 7414 14724 7420 14788
rect 7484 14724 7490 14788
rect 8661 14786 8727 14789
rect 10041 14786 10107 14789
rect 8661 14784 10107 14786
rect 8661 14728 8666 14784
rect 8722 14728 10046 14784
rect 10102 14728 10107 14784
rect 8661 14726 10107 14728
rect 1945 14514 2011 14517
rect 7422 14514 7482 14724
rect 8661 14723 8727 14726
rect 10041 14723 10107 14726
rect 7984 14720 8300 14721
rect 7984 14656 7990 14720
rect 8054 14656 8070 14720
rect 8134 14656 8150 14720
rect 8214 14656 8230 14720
rect 8294 14656 8300 14720
rect 7984 14655 8300 14656
rect 15574 14720 15890 14721
rect 15574 14656 15580 14720
rect 15644 14656 15660 14720
rect 15724 14656 15740 14720
rect 15804 14656 15820 14720
rect 15884 14656 15890 14720
rect 15574 14655 15890 14656
rect 23164 14720 23480 14721
rect 23164 14656 23170 14720
rect 23234 14656 23250 14720
rect 23314 14656 23330 14720
rect 23394 14656 23410 14720
rect 23474 14656 23480 14720
rect 23164 14655 23480 14656
rect 30754 14720 31070 14721
rect 30754 14656 30760 14720
rect 30824 14656 30840 14720
rect 30904 14656 30920 14720
rect 30984 14656 31000 14720
rect 31064 14656 31070 14720
rect 30754 14655 31070 14656
rect 11145 14650 11211 14653
rect 13169 14650 13235 14653
rect 11145 14648 13235 14650
rect 11145 14592 11150 14648
rect 11206 14592 13174 14648
rect 13230 14592 13235 14648
rect 11145 14590 13235 14592
rect 11145 14587 11211 14590
rect 13169 14587 13235 14590
rect 24393 14650 24459 14653
rect 28441 14650 28507 14653
rect 24393 14648 28507 14650
rect 24393 14592 24398 14648
rect 24454 14592 28446 14648
rect 28502 14592 28507 14648
rect 24393 14590 28507 14592
rect 24393 14587 24459 14590
rect 28441 14587 28507 14590
rect 15101 14514 15167 14517
rect 18321 14514 18387 14517
rect 1945 14512 2790 14514
rect 1945 14456 1950 14512
rect 2006 14456 2790 14512
rect 1945 14454 2790 14456
rect 7422 14454 9506 14514
rect 1945 14451 2011 14454
rect 2730 14378 2790 14454
rect 5257 14378 5323 14381
rect 9121 14378 9187 14381
rect 2730 14318 4906 14378
rect 4846 14242 4906 14318
rect 5257 14376 9187 14378
rect 5257 14320 5262 14376
rect 5318 14320 9126 14376
rect 9182 14320 9187 14376
rect 5257 14318 9187 14320
rect 9446 14378 9506 14454
rect 15101 14512 18387 14514
rect 15101 14456 15106 14512
rect 15162 14456 18326 14512
rect 18382 14456 18387 14512
rect 15101 14454 18387 14456
rect 15101 14451 15167 14454
rect 18321 14451 18387 14454
rect 18781 14514 18847 14517
rect 23841 14514 23907 14517
rect 25681 14514 25747 14517
rect 18781 14512 25747 14514
rect 18781 14456 18786 14512
rect 18842 14456 23846 14512
rect 23902 14456 25686 14512
rect 25742 14456 25747 14512
rect 18781 14454 25747 14456
rect 18781 14451 18847 14454
rect 23841 14451 23907 14454
rect 25681 14451 25747 14454
rect 13813 14378 13879 14381
rect 9446 14376 13879 14378
rect 9446 14320 13818 14376
rect 13874 14320 13879 14376
rect 9446 14318 13879 14320
rect 5257 14315 5323 14318
rect 9121 14315 9187 14318
rect 13813 14315 13879 14318
rect 16113 14378 16179 14381
rect 27245 14378 27311 14381
rect 27470 14378 27476 14380
rect 16113 14376 27476 14378
rect 16113 14320 16118 14376
rect 16174 14320 27250 14376
rect 27306 14320 27476 14376
rect 16113 14318 27476 14320
rect 16113 14315 16179 14318
rect 27245 14315 27311 14318
rect 27470 14316 27476 14318
rect 27540 14316 27546 14380
rect 10777 14242 10843 14245
rect 4846 14240 10843 14242
rect 4846 14184 10782 14240
rect 10838 14184 10843 14240
rect 4846 14182 10843 14184
rect 10777 14179 10843 14182
rect 4189 14176 4505 14177
rect 4189 14112 4195 14176
rect 4259 14112 4275 14176
rect 4339 14112 4355 14176
rect 4419 14112 4435 14176
rect 4499 14112 4505 14176
rect 4189 14111 4505 14112
rect 11779 14176 12095 14177
rect 11779 14112 11785 14176
rect 11849 14112 11865 14176
rect 11929 14112 11945 14176
rect 12009 14112 12025 14176
rect 12089 14112 12095 14176
rect 11779 14111 12095 14112
rect 19369 14176 19685 14177
rect 19369 14112 19375 14176
rect 19439 14112 19455 14176
rect 19519 14112 19535 14176
rect 19599 14112 19615 14176
rect 19679 14112 19685 14176
rect 19369 14111 19685 14112
rect 26959 14176 27275 14177
rect 26959 14112 26965 14176
rect 27029 14112 27045 14176
rect 27109 14112 27125 14176
rect 27189 14112 27205 14176
rect 27269 14112 27275 14176
rect 26959 14111 27275 14112
rect 5901 14106 5967 14109
rect 6637 14106 6703 14109
rect 5901 14104 6010 14106
rect 5901 14048 5906 14104
rect 5962 14048 6010 14104
rect 5901 14043 6010 14048
rect 6637 14104 11714 14106
rect 6637 14048 6642 14104
rect 6698 14048 11714 14104
rect 6637 14046 11714 14048
rect 6637 14043 6703 14046
rect 1853 13970 1919 13973
rect 3693 13970 3759 13973
rect 5950 13970 6010 14043
rect 8661 13970 8727 13973
rect 1853 13968 2790 13970
rect 1853 13912 1858 13968
rect 1914 13912 2790 13968
rect 1853 13910 2790 13912
rect 1853 13907 1919 13910
rect 2730 13834 2790 13910
rect 3693 13968 8727 13970
rect 3693 13912 3698 13968
rect 3754 13912 8666 13968
rect 8722 13912 8727 13968
rect 3693 13910 8727 13912
rect 3693 13907 3759 13910
rect 8661 13907 8727 13910
rect 8845 13834 8911 13837
rect 9397 13834 9463 13837
rect 2730 13774 8586 13834
rect 4838 13636 4844 13700
rect 4908 13698 4914 13700
rect 7649 13698 7715 13701
rect 4908 13696 7715 13698
rect 4908 13640 7654 13696
rect 7710 13640 7715 13696
rect 4908 13638 7715 13640
rect 8526 13698 8586 13774
rect 8845 13832 9463 13834
rect 8845 13776 8850 13832
rect 8906 13776 9402 13832
rect 9458 13776 9463 13832
rect 8845 13774 9463 13776
rect 11654 13834 11714 14046
rect 11881 13970 11947 13973
rect 15101 13970 15167 13973
rect 11881 13968 15167 13970
rect 11881 13912 11886 13968
rect 11942 13912 15106 13968
rect 15162 13912 15167 13968
rect 11881 13910 15167 13912
rect 11881 13907 11947 13910
rect 15101 13907 15167 13910
rect 21909 13970 21975 13973
rect 22645 13970 22711 13973
rect 21909 13968 22711 13970
rect 21909 13912 21914 13968
rect 21970 13912 22650 13968
rect 22706 13912 22711 13968
rect 21909 13910 22711 13912
rect 21909 13907 21975 13910
rect 22645 13907 22711 13910
rect 22921 13970 22987 13973
rect 24393 13970 24459 13973
rect 22921 13968 24459 13970
rect 22921 13912 22926 13968
rect 22982 13912 24398 13968
rect 24454 13912 24459 13968
rect 22921 13910 24459 13912
rect 22921 13907 22987 13910
rect 24393 13907 24459 13910
rect 28533 13972 28599 13973
rect 28533 13968 28580 13972
rect 28644 13970 28650 13972
rect 28533 13912 28538 13968
rect 28533 13908 28580 13912
rect 28644 13910 28690 13970
rect 28644 13908 28650 13910
rect 28533 13907 28599 13908
rect 13721 13834 13787 13837
rect 11654 13832 13787 13834
rect 11654 13776 13726 13832
rect 13782 13776 13787 13832
rect 11654 13774 13787 13776
rect 8845 13771 8911 13774
rect 9397 13771 9463 13774
rect 13721 13771 13787 13774
rect 16941 13834 17007 13837
rect 19333 13834 19399 13837
rect 16941 13832 19399 13834
rect 16941 13776 16946 13832
rect 17002 13776 19338 13832
rect 19394 13776 19399 13832
rect 16941 13774 19399 13776
rect 16941 13771 17007 13774
rect 19333 13771 19399 13774
rect 19701 13834 19767 13837
rect 20662 13834 20668 13836
rect 19701 13832 20668 13834
rect 19701 13776 19706 13832
rect 19762 13776 20668 13832
rect 19701 13774 20668 13776
rect 19701 13771 19767 13774
rect 20662 13772 20668 13774
rect 20732 13772 20738 13836
rect 21541 13834 21607 13837
rect 28390 13834 28396 13836
rect 21541 13832 28396 13834
rect 21541 13776 21546 13832
rect 21602 13776 28396 13832
rect 21541 13774 28396 13776
rect 21541 13771 21607 13774
rect 28390 13772 28396 13774
rect 28460 13834 28466 13836
rect 28533 13834 28599 13837
rect 28460 13832 28599 13834
rect 28460 13776 28538 13832
rect 28594 13776 28599 13832
rect 28460 13774 28599 13776
rect 28460 13772 28466 13774
rect 28533 13771 28599 13774
rect 11145 13698 11211 13701
rect 8526 13696 11211 13698
rect 8526 13640 11150 13696
rect 11206 13640 11211 13696
rect 8526 13638 11211 13640
rect 4908 13636 4914 13638
rect 7649 13635 7715 13638
rect 11145 13635 11211 13638
rect 23565 13698 23631 13701
rect 30373 13698 30439 13701
rect 23565 13696 30439 13698
rect 23565 13640 23570 13696
rect 23626 13640 30378 13696
rect 30434 13640 30439 13696
rect 23565 13638 30439 13640
rect 23565 13635 23631 13638
rect 30373 13635 30439 13638
rect 7984 13632 8300 13633
rect 7984 13568 7990 13632
rect 8054 13568 8070 13632
rect 8134 13568 8150 13632
rect 8214 13568 8230 13632
rect 8294 13568 8300 13632
rect 7984 13567 8300 13568
rect 15574 13632 15890 13633
rect 15574 13568 15580 13632
rect 15644 13568 15660 13632
rect 15724 13568 15740 13632
rect 15804 13568 15820 13632
rect 15884 13568 15890 13632
rect 15574 13567 15890 13568
rect 23164 13632 23480 13633
rect 23164 13568 23170 13632
rect 23234 13568 23250 13632
rect 23314 13568 23330 13632
rect 23394 13568 23410 13632
rect 23474 13568 23480 13632
rect 23164 13567 23480 13568
rect 30754 13632 31070 13633
rect 30754 13568 30760 13632
rect 30824 13568 30840 13632
rect 30904 13568 30920 13632
rect 30984 13568 31000 13632
rect 31064 13568 31070 13632
rect 30754 13567 31070 13568
rect 4153 13562 4219 13565
rect 6637 13562 6703 13565
rect 4153 13560 6703 13562
rect 4153 13504 4158 13560
rect 4214 13504 6642 13560
rect 6698 13504 6703 13560
rect 4153 13502 6703 13504
rect 4153 13499 4219 13502
rect 6637 13499 6703 13502
rect 8518 13500 8524 13564
rect 8588 13562 8594 13564
rect 11053 13562 11119 13565
rect 8588 13560 11119 13562
rect 8588 13504 11058 13560
rect 11114 13504 11119 13560
rect 8588 13502 11119 13504
rect 8588 13500 8594 13502
rect 11053 13499 11119 13502
rect 23933 13562 23999 13565
rect 26877 13562 26943 13565
rect 23933 13560 26943 13562
rect 23933 13504 23938 13560
rect 23994 13504 26882 13560
rect 26938 13504 26943 13560
rect 23933 13502 26943 13504
rect 23933 13499 23999 13502
rect 26877 13499 26943 13502
rect 6545 13426 6611 13429
rect 9581 13426 9647 13429
rect 6545 13424 9647 13426
rect 6545 13368 6550 13424
rect 6606 13368 9586 13424
rect 9642 13368 9647 13424
rect 6545 13366 9647 13368
rect 6545 13363 6611 13366
rect 9581 13363 9647 13366
rect 10133 13426 10199 13429
rect 18965 13426 19031 13429
rect 10133 13424 19031 13426
rect 10133 13368 10138 13424
rect 10194 13368 18970 13424
rect 19026 13368 19031 13424
rect 10133 13366 19031 13368
rect 10133 13363 10199 13366
rect 18965 13363 19031 13366
rect 22369 13426 22435 13429
rect 24393 13426 24459 13429
rect 22369 13424 24459 13426
rect 22369 13368 22374 13424
rect 22430 13368 24398 13424
rect 24454 13368 24459 13424
rect 22369 13366 24459 13368
rect 22369 13363 22435 13366
rect 24393 13363 24459 13366
rect 2221 13290 2287 13293
rect 13721 13290 13787 13293
rect 30005 13290 30071 13293
rect 2221 13288 30071 13290
rect 2221 13232 2226 13288
rect 2282 13232 13726 13288
rect 13782 13232 30010 13288
rect 30066 13232 30071 13288
rect 2221 13230 30071 13232
rect 2221 13227 2287 13230
rect 13721 13227 13787 13230
rect 30005 13227 30071 13230
rect 5206 13092 5212 13156
rect 5276 13154 5282 13156
rect 10593 13154 10659 13157
rect 5276 13152 10659 13154
rect 5276 13096 10598 13152
rect 10654 13096 10659 13152
rect 5276 13094 10659 13096
rect 5276 13092 5282 13094
rect 10593 13091 10659 13094
rect 21633 13154 21699 13157
rect 22921 13154 22987 13157
rect 21633 13152 22987 13154
rect 21633 13096 21638 13152
rect 21694 13096 22926 13152
rect 22982 13096 22987 13152
rect 21633 13094 22987 13096
rect 21633 13091 21699 13094
rect 22921 13091 22987 13094
rect 4189 13088 4505 13089
rect 4189 13024 4195 13088
rect 4259 13024 4275 13088
rect 4339 13024 4355 13088
rect 4419 13024 4435 13088
rect 4499 13024 4505 13088
rect 4189 13023 4505 13024
rect 11779 13088 12095 13089
rect 11779 13024 11785 13088
rect 11849 13024 11865 13088
rect 11929 13024 11945 13088
rect 12009 13024 12025 13088
rect 12089 13024 12095 13088
rect 11779 13023 12095 13024
rect 19369 13088 19685 13089
rect 19369 13024 19375 13088
rect 19439 13024 19455 13088
rect 19519 13024 19535 13088
rect 19599 13024 19615 13088
rect 19679 13024 19685 13088
rect 19369 13023 19685 13024
rect 26959 13088 27275 13089
rect 26959 13024 26965 13088
rect 27029 13024 27045 13088
rect 27109 13024 27125 13088
rect 27189 13024 27205 13088
rect 27269 13024 27275 13088
rect 26959 13023 27275 13024
rect 6085 13018 6151 13021
rect 8385 13018 8451 13021
rect 9070 13018 9076 13020
rect 6085 13016 8451 13018
rect 6085 12960 6090 13016
rect 6146 12960 8390 13016
rect 8446 12960 8451 13016
rect 6085 12958 8451 12960
rect 6085 12955 6151 12958
rect 8385 12955 8451 12958
rect 8526 12958 9076 13018
rect 3417 12882 3483 12885
rect 8526 12882 8586 12958
rect 9070 12956 9076 12958
rect 9140 12956 9146 13020
rect 9438 12956 9444 13020
rect 9508 13018 9514 13020
rect 10133 13018 10199 13021
rect 11329 13018 11395 13021
rect 9508 13016 10199 13018
rect 9508 12960 10138 13016
rect 10194 12960 10199 13016
rect 9508 12958 10199 12960
rect 9508 12956 9514 12958
rect 10133 12955 10199 12958
rect 10964 13016 11395 13018
rect 10964 12960 11334 13016
rect 11390 12960 11395 13016
rect 10964 12958 11395 12960
rect 3417 12880 8586 12882
rect 3417 12824 3422 12880
rect 3478 12824 8586 12880
rect 3417 12822 8586 12824
rect 3417 12819 3483 12822
rect 8702 12820 8708 12884
rect 8772 12882 8778 12884
rect 10964 12882 11024 12958
rect 11329 12955 11395 12958
rect 8772 12822 11024 12882
rect 11145 12882 11211 12885
rect 19742 12882 19748 12884
rect 11145 12880 19748 12882
rect 11145 12824 11150 12880
rect 11206 12824 19748 12880
rect 11145 12822 19748 12824
rect 8772 12820 8778 12822
rect 11145 12819 11211 12822
rect 19742 12820 19748 12822
rect 19812 12820 19818 12884
rect 22829 12882 22895 12885
rect 27521 12882 27587 12885
rect 22829 12880 27587 12882
rect 22829 12824 22834 12880
rect 22890 12824 27526 12880
rect 27582 12824 27587 12880
rect 22829 12822 27587 12824
rect 22829 12819 22895 12822
rect 27521 12819 27587 12822
rect 3417 12746 3483 12749
rect 6361 12746 6427 12749
rect 16665 12746 16731 12749
rect 3417 12744 4170 12746
rect 3417 12688 3422 12744
rect 3478 12688 4170 12744
rect 3417 12686 4170 12688
rect 3417 12683 3483 12686
rect 1485 12474 1551 12477
rect 2998 12474 3004 12476
rect 1485 12472 3004 12474
rect 1485 12416 1490 12472
rect 1546 12416 3004 12472
rect 1485 12414 3004 12416
rect 1485 12411 1551 12414
rect 2998 12412 3004 12414
rect 3068 12412 3074 12476
rect 4110 12338 4170 12686
rect 6361 12744 16731 12746
rect 6361 12688 6366 12744
rect 6422 12688 16670 12744
rect 16726 12688 16731 12744
rect 6361 12686 16731 12688
rect 6361 12683 6427 12686
rect 16665 12683 16731 12686
rect 20069 12746 20135 12749
rect 21909 12746 21975 12749
rect 23749 12746 23815 12749
rect 20069 12744 23815 12746
rect 20069 12688 20074 12744
rect 20130 12688 21914 12744
rect 21970 12688 23754 12744
rect 23810 12688 23815 12744
rect 20069 12686 23815 12688
rect 20069 12683 20135 12686
rect 21909 12683 21975 12686
rect 23749 12683 23815 12686
rect 12157 12612 12223 12613
rect 13445 12612 13511 12613
rect 12157 12610 12204 12612
rect 12112 12608 12204 12610
rect 12112 12552 12162 12608
rect 12112 12550 12204 12552
rect 12157 12548 12204 12550
rect 12268 12548 12274 12612
rect 13445 12610 13492 12612
rect 12942 12608 13492 12610
rect 13556 12610 13562 12612
rect 12942 12552 13450 12608
rect 12942 12550 13492 12552
rect 12157 12547 12223 12548
rect 7984 12544 8300 12545
rect 7984 12480 7990 12544
rect 8054 12480 8070 12544
rect 8134 12480 8150 12544
rect 8214 12480 8230 12544
rect 8294 12480 8300 12544
rect 7984 12479 8300 12480
rect 11605 12474 11671 12477
rect 12709 12474 12775 12477
rect 11605 12472 12775 12474
rect 11605 12416 11610 12472
rect 11666 12416 12714 12472
rect 12770 12416 12775 12472
rect 11605 12414 12775 12416
rect 11605 12411 11671 12414
rect 12709 12411 12775 12414
rect 5390 12338 5396 12340
rect 4110 12278 5396 12338
rect 5390 12276 5396 12278
rect 5460 12276 5466 12340
rect 9673 12338 9739 12341
rect 9806 12338 9812 12340
rect 9673 12336 9812 12338
rect 9673 12280 9678 12336
rect 9734 12280 9812 12336
rect 9673 12278 9812 12280
rect 9673 12275 9739 12278
rect 9806 12276 9812 12278
rect 9876 12276 9882 12340
rect 11145 12338 11211 12341
rect 12942 12338 13002 12550
rect 13445 12548 13492 12550
rect 13556 12550 13638 12610
rect 13556 12548 13562 12550
rect 13445 12547 13511 12548
rect 15574 12544 15890 12545
rect 15574 12480 15580 12544
rect 15644 12480 15660 12544
rect 15724 12480 15740 12544
rect 15804 12480 15820 12544
rect 15884 12480 15890 12544
rect 15574 12479 15890 12480
rect 23164 12544 23480 12545
rect 23164 12480 23170 12544
rect 23234 12480 23250 12544
rect 23314 12480 23330 12544
rect 23394 12480 23410 12544
rect 23474 12480 23480 12544
rect 23164 12479 23480 12480
rect 30754 12544 31070 12545
rect 30754 12480 30760 12544
rect 30824 12480 30840 12544
rect 30904 12480 30920 12544
rect 30984 12480 31000 12544
rect 31064 12480 31070 12544
rect 30754 12479 31070 12480
rect 27153 12474 27219 12477
rect 29361 12474 29427 12477
rect 27153 12472 29427 12474
rect 27153 12416 27158 12472
rect 27214 12416 29366 12472
rect 29422 12416 29427 12472
rect 27153 12414 29427 12416
rect 27153 12411 27219 12414
rect 29361 12411 29427 12414
rect 11145 12336 13002 12338
rect 11145 12280 11150 12336
rect 11206 12280 13002 12336
rect 11145 12278 13002 12280
rect 11145 12275 11211 12278
rect 5165 12202 5231 12205
rect 10317 12202 10383 12205
rect 5165 12200 10383 12202
rect 5165 12144 5170 12200
rect 5226 12144 10322 12200
rect 10378 12144 10383 12200
rect 5165 12142 10383 12144
rect 5165 12139 5231 12142
rect 10317 12139 10383 12142
rect 10726 12140 10732 12204
rect 10796 12140 10802 12204
rect 11973 12202 12039 12205
rect 14089 12202 14155 12205
rect 11973 12200 14155 12202
rect 11973 12144 11978 12200
rect 12034 12144 14094 12200
rect 14150 12144 14155 12200
rect 11973 12142 14155 12144
rect 9673 12066 9739 12069
rect 10734 12066 10794 12140
rect 11973 12139 12039 12142
rect 14089 12139 14155 12142
rect 15837 12202 15903 12205
rect 25957 12202 26023 12205
rect 15837 12200 26023 12202
rect 15837 12144 15842 12200
rect 15898 12144 25962 12200
rect 26018 12144 26023 12200
rect 15837 12142 26023 12144
rect 15837 12139 15903 12142
rect 25957 12139 26023 12142
rect 9673 12064 10794 12066
rect 9673 12008 9678 12064
rect 9734 12008 10794 12064
rect 9673 12006 10794 12008
rect 12341 12066 12407 12069
rect 13721 12066 13787 12069
rect 12341 12064 13787 12066
rect 12341 12008 12346 12064
rect 12402 12008 13726 12064
rect 13782 12008 13787 12064
rect 12341 12006 13787 12008
rect 9673 12003 9739 12006
rect 12341 12003 12407 12006
rect 13721 12003 13787 12006
rect 29126 12004 29132 12068
rect 29196 12066 29202 12068
rect 29913 12066 29979 12069
rect 29196 12064 29979 12066
rect 29196 12008 29918 12064
rect 29974 12008 29979 12064
rect 29196 12006 29979 12008
rect 29196 12004 29202 12006
rect 29913 12003 29979 12006
rect 4189 12000 4505 12001
rect 4189 11936 4195 12000
rect 4259 11936 4275 12000
rect 4339 11936 4355 12000
rect 4419 11936 4435 12000
rect 4499 11936 4505 12000
rect 4189 11935 4505 11936
rect 11779 12000 12095 12001
rect 11779 11936 11785 12000
rect 11849 11936 11865 12000
rect 11929 11936 11945 12000
rect 12009 11936 12025 12000
rect 12089 11936 12095 12000
rect 11779 11935 12095 11936
rect 19369 12000 19685 12001
rect 19369 11936 19375 12000
rect 19439 11936 19455 12000
rect 19519 11936 19535 12000
rect 19599 11936 19615 12000
rect 19679 11936 19685 12000
rect 19369 11935 19685 11936
rect 26959 12000 27275 12001
rect 26959 11936 26965 12000
rect 27029 11936 27045 12000
rect 27109 11936 27125 12000
rect 27189 11936 27205 12000
rect 27269 11936 27275 12000
rect 26959 11935 27275 11936
rect 12157 11930 12223 11933
rect 12617 11930 12683 11933
rect 13445 11930 13511 11933
rect 12157 11928 13511 11930
rect 12157 11872 12162 11928
rect 12218 11872 12622 11928
rect 12678 11872 13450 11928
rect 13506 11872 13511 11928
rect 12157 11870 13511 11872
rect 12157 11867 12223 11870
rect 12617 11867 12683 11870
rect 13445 11867 13511 11870
rect 3509 11794 3575 11797
rect 14038 11794 14044 11796
rect 3509 11792 14044 11794
rect 3509 11736 3514 11792
rect 3570 11736 14044 11792
rect 3509 11734 14044 11736
rect 3509 11731 3575 11734
rect 14038 11732 14044 11734
rect 14108 11732 14114 11796
rect 17493 11794 17559 11797
rect 25405 11794 25471 11797
rect 17493 11792 25471 11794
rect 17493 11736 17498 11792
rect 17554 11736 25410 11792
rect 25466 11736 25471 11792
rect 17493 11734 25471 11736
rect 17493 11731 17559 11734
rect 25405 11731 25471 11734
rect 25957 11794 26023 11797
rect 28809 11794 28875 11797
rect 25957 11792 28875 11794
rect 25957 11736 25962 11792
rect 26018 11736 28814 11792
rect 28870 11736 28875 11792
rect 25957 11734 28875 11736
rect 25957 11731 26023 11734
rect 28809 11731 28875 11734
rect 5390 11596 5396 11660
rect 5460 11658 5466 11660
rect 5460 11598 10058 11658
rect 5460 11596 5466 11598
rect 5717 11522 5783 11525
rect 7833 11522 7899 11525
rect 5717 11520 7899 11522
rect 5717 11464 5722 11520
rect 5778 11464 7838 11520
rect 7894 11464 7899 11520
rect 5717 11462 7899 11464
rect 9998 11522 10058 11598
rect 10174 11596 10180 11660
rect 10244 11658 10250 11660
rect 10961 11658 11027 11661
rect 16062 11658 16068 11660
rect 10244 11656 11027 11658
rect 10244 11600 10966 11656
rect 11022 11600 11027 11656
rect 10244 11598 11027 11600
rect 10244 11596 10250 11598
rect 10961 11595 11027 11598
rect 11102 11598 16068 11658
rect 10593 11522 10659 11525
rect 9998 11520 10659 11522
rect 9998 11464 10598 11520
rect 10654 11464 10659 11520
rect 9998 11462 10659 11464
rect 5717 11459 5783 11462
rect 7833 11459 7899 11462
rect 10593 11459 10659 11462
rect 10777 11522 10843 11525
rect 11102 11522 11162 11598
rect 16062 11596 16068 11598
rect 16132 11596 16138 11660
rect 21633 11658 21699 11661
rect 24209 11658 24275 11661
rect 21633 11656 24275 11658
rect 21633 11600 21638 11656
rect 21694 11600 24214 11656
rect 24270 11600 24275 11656
rect 21633 11598 24275 11600
rect 21633 11595 21699 11598
rect 24209 11595 24275 11598
rect 10777 11520 11162 11522
rect 10777 11464 10782 11520
rect 10838 11464 11162 11520
rect 10777 11462 11162 11464
rect 10777 11459 10843 11462
rect 7984 11456 8300 11457
rect 7984 11392 7990 11456
rect 8054 11392 8070 11456
rect 8134 11392 8150 11456
rect 8214 11392 8230 11456
rect 8294 11392 8300 11456
rect 7984 11391 8300 11392
rect 15574 11456 15890 11457
rect 15574 11392 15580 11456
rect 15644 11392 15660 11456
rect 15724 11392 15740 11456
rect 15804 11392 15820 11456
rect 15884 11392 15890 11456
rect 15574 11391 15890 11392
rect 23164 11456 23480 11457
rect 23164 11392 23170 11456
rect 23234 11392 23250 11456
rect 23314 11392 23330 11456
rect 23394 11392 23410 11456
rect 23474 11392 23480 11456
rect 23164 11391 23480 11392
rect 30754 11456 31070 11457
rect 30754 11392 30760 11456
rect 30824 11392 30840 11456
rect 30904 11392 30920 11456
rect 30984 11392 31000 11456
rect 31064 11392 31070 11456
rect 30754 11391 31070 11392
rect 9949 11386 10015 11389
rect 10317 11386 10383 11389
rect 9949 11384 10383 11386
rect 9949 11328 9954 11384
rect 10010 11328 10322 11384
rect 10378 11328 10383 11384
rect 9949 11326 10383 11328
rect 9949 11323 10015 11326
rect 10317 11323 10383 11326
rect 1945 11250 2011 11253
rect 29913 11250 29979 11253
rect 1945 11248 29979 11250
rect 1945 11192 1950 11248
rect 2006 11192 29918 11248
rect 29974 11192 29979 11248
rect 1945 11190 29979 11192
rect 1945 11187 2011 11190
rect 29913 11187 29979 11190
rect 11789 11114 11855 11117
rect 8342 11112 11855 11114
rect 8342 11056 11794 11112
rect 11850 11056 11855 11112
rect 8342 11054 11855 11056
rect 6678 10916 6684 10980
rect 6748 10978 6754 10980
rect 8342 10978 8402 11054
rect 11789 11051 11855 11054
rect 20662 11052 20668 11116
rect 20732 11114 20738 11116
rect 26325 11114 26391 11117
rect 20732 11112 26391 11114
rect 20732 11056 26330 11112
rect 26386 11056 26391 11112
rect 20732 11054 26391 11056
rect 20732 11052 20738 11054
rect 26325 11051 26391 11054
rect 6748 10918 8402 10978
rect 8477 10978 8543 10981
rect 9857 10980 9923 10981
rect 9622 10978 9628 10980
rect 8477 10976 9628 10978
rect 8477 10920 8482 10976
rect 8538 10920 9628 10976
rect 8477 10918 9628 10920
rect 6748 10916 6754 10918
rect 8477 10915 8543 10918
rect 9622 10916 9628 10918
rect 9692 10916 9698 10980
rect 9806 10916 9812 10980
rect 9876 10978 9923 10980
rect 9876 10976 9968 10978
rect 9918 10920 9968 10976
rect 9876 10918 9968 10920
rect 9876 10916 9923 10918
rect 9857 10915 9923 10916
rect 4189 10912 4505 10913
rect 4189 10848 4195 10912
rect 4259 10848 4275 10912
rect 4339 10848 4355 10912
rect 4419 10848 4435 10912
rect 4499 10848 4505 10912
rect 4189 10847 4505 10848
rect 11779 10912 12095 10913
rect 11779 10848 11785 10912
rect 11849 10848 11865 10912
rect 11929 10848 11945 10912
rect 12009 10848 12025 10912
rect 12089 10848 12095 10912
rect 11779 10847 12095 10848
rect 19369 10912 19685 10913
rect 19369 10848 19375 10912
rect 19439 10848 19455 10912
rect 19519 10848 19535 10912
rect 19599 10848 19615 10912
rect 19679 10848 19685 10912
rect 19369 10847 19685 10848
rect 26959 10912 27275 10913
rect 26959 10848 26965 10912
rect 27029 10848 27045 10912
rect 27109 10848 27125 10912
rect 27189 10848 27205 10912
rect 27269 10848 27275 10912
rect 26959 10847 27275 10848
rect 5073 10842 5139 10845
rect 9581 10842 9647 10845
rect 5073 10840 9647 10842
rect 5073 10784 5078 10840
rect 5134 10784 9586 10840
rect 9642 10784 9647 10840
rect 5073 10782 9647 10784
rect 5073 10779 5139 10782
rect 9581 10779 9647 10782
rect 2957 10706 3023 10709
rect 8886 10706 8892 10708
rect 2957 10704 8892 10706
rect 2957 10648 2962 10704
rect 3018 10648 8892 10704
rect 2957 10646 8892 10648
rect 2957 10643 3023 10646
rect 8886 10644 8892 10646
rect 8956 10644 8962 10708
rect 10593 10706 10659 10709
rect 15929 10706 15995 10709
rect 10593 10704 15995 10706
rect 10593 10648 10598 10704
rect 10654 10648 15934 10704
rect 15990 10648 15995 10704
rect 10593 10646 15995 10648
rect 10593 10643 10659 10646
rect 15929 10643 15995 10646
rect 16389 10706 16455 10709
rect 21081 10706 21147 10709
rect 16389 10704 21147 10706
rect 16389 10648 16394 10704
rect 16450 10648 21086 10704
rect 21142 10648 21147 10704
rect 16389 10646 21147 10648
rect 16389 10643 16455 10646
rect 21081 10643 21147 10646
rect 5349 10570 5415 10573
rect 23473 10570 23539 10573
rect 5349 10568 23539 10570
rect 5349 10512 5354 10568
rect 5410 10512 23478 10568
rect 23534 10512 23539 10568
rect 5349 10510 23539 10512
rect 5349 10507 5415 10510
rect 23473 10507 23539 10510
rect 8661 10434 8727 10437
rect 11421 10434 11487 10437
rect 13169 10434 13235 10437
rect 8661 10432 13235 10434
rect 8661 10376 8666 10432
rect 8722 10376 11426 10432
rect 11482 10376 13174 10432
rect 13230 10376 13235 10432
rect 8661 10374 13235 10376
rect 8661 10371 8727 10374
rect 11421 10371 11487 10374
rect 13169 10371 13235 10374
rect 7984 10368 8300 10369
rect 7984 10304 7990 10368
rect 8054 10304 8070 10368
rect 8134 10304 8150 10368
rect 8214 10304 8230 10368
rect 8294 10304 8300 10368
rect 7984 10303 8300 10304
rect 15574 10368 15890 10369
rect 15574 10304 15580 10368
rect 15644 10304 15660 10368
rect 15724 10304 15740 10368
rect 15804 10304 15820 10368
rect 15884 10304 15890 10368
rect 15574 10303 15890 10304
rect 23164 10368 23480 10369
rect 23164 10304 23170 10368
rect 23234 10304 23250 10368
rect 23314 10304 23330 10368
rect 23394 10304 23410 10368
rect 23474 10304 23480 10368
rect 23164 10303 23480 10304
rect 30754 10368 31070 10369
rect 30754 10304 30760 10368
rect 30824 10304 30840 10368
rect 30904 10304 30920 10368
rect 30984 10304 31000 10368
rect 31064 10304 31070 10368
rect 30754 10303 31070 10304
rect 12617 10298 12683 10301
rect 12390 10296 12683 10298
rect 12390 10240 12622 10296
rect 12678 10240 12683 10296
rect 12390 10238 12683 10240
rect 7465 10162 7531 10165
rect 12390 10162 12450 10238
rect 12617 10235 12683 10238
rect 7465 10160 12450 10162
rect 7465 10104 7470 10160
rect 7526 10104 12450 10160
rect 7465 10102 12450 10104
rect 7465 10099 7531 10102
rect 19742 10100 19748 10164
rect 19812 10162 19818 10164
rect 20253 10162 20319 10165
rect 19812 10160 20319 10162
rect 19812 10104 20258 10160
rect 20314 10104 20319 10160
rect 19812 10102 20319 10104
rect 19812 10100 19818 10102
rect 20253 10099 20319 10102
rect 21081 10162 21147 10165
rect 27429 10162 27495 10165
rect 21081 10160 27495 10162
rect 21081 10104 21086 10160
rect 21142 10104 27434 10160
rect 27490 10104 27495 10160
rect 21081 10102 27495 10104
rect 21081 10099 21147 10102
rect 27429 10099 27495 10102
rect 2313 10026 2379 10029
rect 9254 10026 9260 10028
rect 2313 10024 9260 10026
rect 2313 9968 2318 10024
rect 2374 9968 9260 10024
rect 2313 9966 9260 9968
rect 2313 9963 2379 9966
rect 9254 9964 9260 9966
rect 9324 9964 9330 10028
rect 20621 10026 20687 10029
rect 22185 10026 22251 10029
rect 29177 10026 29243 10029
rect 20621 10024 22110 10026
rect 20621 9968 20626 10024
rect 20682 9968 22110 10024
rect 20621 9966 22110 9968
rect 20621 9963 20687 9966
rect 22050 9890 22110 9966
rect 22185 10024 29243 10026
rect 22185 9968 22190 10024
rect 22246 9968 29182 10024
rect 29238 9968 29243 10024
rect 22185 9966 29243 9968
rect 22185 9963 22251 9966
rect 29177 9963 29243 9966
rect 22461 9890 22527 9893
rect 22050 9888 22527 9890
rect 22050 9832 22466 9888
rect 22522 9832 22527 9888
rect 22050 9830 22527 9832
rect 22461 9827 22527 9830
rect 4189 9824 4505 9825
rect 4189 9760 4195 9824
rect 4259 9760 4275 9824
rect 4339 9760 4355 9824
rect 4419 9760 4435 9824
rect 4499 9760 4505 9824
rect 4189 9759 4505 9760
rect 11779 9824 12095 9825
rect 11779 9760 11785 9824
rect 11849 9760 11865 9824
rect 11929 9760 11945 9824
rect 12009 9760 12025 9824
rect 12089 9760 12095 9824
rect 11779 9759 12095 9760
rect 19369 9824 19685 9825
rect 19369 9760 19375 9824
rect 19439 9760 19455 9824
rect 19519 9760 19535 9824
rect 19599 9760 19615 9824
rect 19679 9760 19685 9824
rect 19369 9759 19685 9760
rect 26959 9824 27275 9825
rect 26959 9760 26965 9824
rect 27029 9760 27045 9824
rect 27109 9760 27125 9824
rect 27189 9760 27205 9824
rect 27269 9760 27275 9824
rect 26959 9759 27275 9760
rect 5574 9692 5580 9756
rect 5644 9754 5650 9756
rect 10869 9754 10935 9757
rect 5644 9752 10935 9754
rect 5644 9696 10874 9752
rect 10930 9696 10935 9752
rect 5644 9694 10935 9696
rect 5644 9692 5650 9694
rect 10869 9691 10935 9694
rect 6361 9618 6427 9621
rect 8385 9618 8451 9621
rect 6361 9616 8451 9618
rect 6361 9560 6366 9616
rect 6422 9560 8390 9616
rect 8446 9560 8451 9616
rect 6361 9558 8451 9560
rect 6361 9555 6427 9558
rect 8385 9555 8451 9558
rect 9857 9618 9923 9621
rect 12525 9618 12591 9621
rect 9857 9616 12591 9618
rect 9857 9560 9862 9616
rect 9918 9560 12530 9616
rect 12586 9560 12591 9616
rect 9857 9558 12591 9560
rect 9857 9555 9923 9558
rect 12525 9555 12591 9558
rect 23749 9618 23815 9621
rect 24669 9618 24735 9621
rect 23749 9616 24735 9618
rect 23749 9560 23754 9616
rect 23810 9560 24674 9616
rect 24730 9560 24735 9616
rect 23749 9558 24735 9560
rect 23749 9555 23815 9558
rect 24669 9555 24735 9558
rect 6862 9420 6868 9484
rect 6932 9482 6938 9484
rect 17585 9482 17651 9485
rect 6932 9480 17651 9482
rect 6932 9424 17590 9480
rect 17646 9424 17651 9480
rect 6932 9422 17651 9424
rect 6932 9420 6938 9422
rect 17585 9419 17651 9422
rect 23473 9482 23539 9485
rect 26141 9482 26207 9485
rect 29821 9482 29887 9485
rect 23473 9480 29887 9482
rect 23473 9424 23478 9480
rect 23534 9424 26146 9480
rect 26202 9424 29826 9480
rect 29882 9424 29887 9480
rect 23473 9422 29887 9424
rect 23473 9419 23539 9422
rect 26141 9419 26207 9422
rect 29821 9419 29887 9422
rect 10685 9346 10751 9349
rect 13169 9346 13235 9349
rect 10685 9344 13235 9346
rect 10685 9288 10690 9344
rect 10746 9288 13174 9344
rect 13230 9288 13235 9344
rect 10685 9286 13235 9288
rect 10685 9283 10751 9286
rect 13169 9283 13235 9286
rect 23565 9346 23631 9349
rect 29177 9346 29243 9349
rect 23565 9344 29243 9346
rect 23565 9288 23570 9344
rect 23626 9288 29182 9344
rect 29238 9288 29243 9344
rect 23565 9286 29243 9288
rect 23565 9283 23631 9286
rect 29177 9283 29243 9286
rect 7984 9280 8300 9281
rect 7984 9216 7990 9280
rect 8054 9216 8070 9280
rect 8134 9216 8150 9280
rect 8214 9216 8230 9280
rect 8294 9216 8300 9280
rect 7984 9215 8300 9216
rect 15574 9280 15890 9281
rect 15574 9216 15580 9280
rect 15644 9216 15660 9280
rect 15724 9216 15740 9280
rect 15804 9216 15820 9280
rect 15884 9216 15890 9280
rect 15574 9215 15890 9216
rect 23164 9280 23480 9281
rect 23164 9216 23170 9280
rect 23234 9216 23250 9280
rect 23314 9216 23330 9280
rect 23394 9216 23410 9280
rect 23474 9216 23480 9280
rect 23164 9215 23480 9216
rect 30754 9280 31070 9281
rect 30754 9216 30760 9280
rect 30824 9216 30840 9280
rect 30904 9216 30920 9280
rect 30984 9216 31000 9280
rect 31064 9216 31070 9280
rect 30754 9215 31070 9216
rect 6085 9210 6151 9213
rect 7465 9210 7531 9213
rect 12341 9210 12407 9213
rect 6085 9208 7531 9210
rect 6085 9152 6090 9208
rect 6146 9152 7470 9208
rect 7526 9152 7531 9208
rect 6085 9150 7531 9152
rect 6085 9147 6151 9150
rect 7465 9147 7531 9150
rect 9630 9208 12407 9210
rect 9630 9152 12346 9208
rect 12402 9152 12407 9208
rect 9630 9150 12407 9152
rect 5809 9074 5875 9077
rect 7189 9074 7255 9077
rect 9630 9074 9690 9150
rect 12341 9147 12407 9150
rect 5809 9072 9690 9074
rect 5809 9016 5814 9072
rect 5870 9016 7194 9072
rect 7250 9016 9690 9072
rect 5809 9014 9690 9016
rect 16757 9074 16823 9077
rect 17125 9074 17191 9077
rect 16757 9072 17191 9074
rect 16757 9016 16762 9072
rect 16818 9016 17130 9072
rect 17186 9016 17191 9072
rect 16757 9014 17191 9016
rect 5809 9011 5875 9014
rect 7189 9011 7255 9014
rect 16757 9011 16823 9014
rect 17125 9011 17191 9014
rect 26141 9074 26207 9077
rect 26969 9074 27035 9077
rect 26141 9072 27035 9074
rect 26141 9016 26146 9072
rect 26202 9016 26974 9072
rect 27030 9016 27035 9072
rect 26141 9014 27035 9016
rect 26141 9011 26207 9014
rect 26969 9011 27035 9014
rect 3325 8938 3391 8941
rect 8477 8938 8543 8941
rect 3325 8936 8543 8938
rect 3325 8880 3330 8936
rect 3386 8880 8482 8936
rect 8538 8880 8543 8936
rect 3325 8878 8543 8880
rect 3325 8875 3391 8878
rect 8477 8875 8543 8878
rect 14038 8876 14044 8940
rect 14108 8938 14114 8940
rect 24025 8938 24091 8941
rect 14108 8936 24091 8938
rect 14108 8880 24030 8936
rect 24086 8880 24091 8936
rect 14108 8878 24091 8880
rect 14108 8876 14114 8878
rect 24025 8875 24091 8878
rect 26509 8938 26575 8941
rect 29269 8938 29335 8941
rect 26509 8936 29335 8938
rect 26509 8880 26514 8936
rect 26570 8880 29274 8936
rect 29330 8880 29335 8936
rect 26509 8878 29335 8880
rect 26509 8875 26575 8878
rect 29269 8875 29335 8878
rect 4189 8736 4505 8737
rect 4189 8672 4195 8736
rect 4259 8672 4275 8736
rect 4339 8672 4355 8736
rect 4419 8672 4435 8736
rect 4499 8672 4505 8736
rect 4189 8671 4505 8672
rect 11779 8736 12095 8737
rect 11779 8672 11785 8736
rect 11849 8672 11865 8736
rect 11929 8672 11945 8736
rect 12009 8672 12025 8736
rect 12089 8672 12095 8736
rect 11779 8671 12095 8672
rect 19369 8736 19685 8737
rect 19369 8672 19375 8736
rect 19439 8672 19455 8736
rect 19519 8672 19535 8736
rect 19599 8672 19615 8736
rect 19679 8672 19685 8736
rect 19369 8671 19685 8672
rect 26959 8736 27275 8737
rect 26959 8672 26965 8736
rect 27029 8672 27045 8736
rect 27109 8672 27125 8736
rect 27189 8672 27205 8736
rect 27269 8672 27275 8736
rect 26959 8671 27275 8672
rect 21173 8666 21239 8669
rect 23013 8666 23079 8669
rect 21173 8664 23079 8666
rect 21173 8608 21178 8664
rect 21234 8608 23018 8664
rect 23074 8608 23079 8664
rect 21173 8606 23079 8608
rect 21173 8603 21239 8606
rect 23013 8603 23079 8606
rect 7465 8530 7531 8533
rect 9213 8530 9279 8533
rect 11421 8530 11487 8533
rect 12249 8530 12315 8533
rect 7465 8528 12315 8530
rect 7465 8472 7470 8528
rect 7526 8472 9218 8528
rect 9274 8472 11426 8528
rect 11482 8472 12254 8528
rect 12310 8472 12315 8528
rect 7465 8470 12315 8472
rect 7465 8467 7531 8470
rect 9213 8467 9279 8470
rect 11421 8467 11487 8470
rect 12249 8467 12315 8470
rect 22001 8530 22067 8533
rect 29821 8530 29887 8533
rect 22001 8528 29887 8530
rect 22001 8472 22006 8528
rect 22062 8472 29826 8528
rect 29882 8472 29887 8528
rect 22001 8470 29887 8472
rect 22001 8467 22067 8470
rect 29821 8467 29887 8470
rect 13077 8394 13143 8397
rect 4110 8392 13143 8394
rect 4110 8336 13082 8392
rect 13138 8336 13143 8392
rect 4110 8334 13143 8336
rect 2405 8258 2471 8261
rect 4110 8258 4170 8334
rect 13077 8331 13143 8334
rect 15101 8394 15167 8397
rect 20989 8394 21055 8397
rect 15101 8392 21055 8394
rect 15101 8336 15106 8392
rect 15162 8336 20994 8392
rect 21050 8336 21055 8392
rect 15101 8334 21055 8336
rect 15101 8331 15167 8334
rect 20989 8331 21055 8334
rect 21265 8394 21331 8397
rect 25405 8394 25471 8397
rect 21265 8392 25471 8394
rect 21265 8336 21270 8392
rect 21326 8336 25410 8392
rect 25466 8336 25471 8392
rect 21265 8334 25471 8336
rect 21265 8331 21331 8334
rect 25405 8331 25471 8334
rect 2405 8256 4170 8258
rect 2405 8200 2410 8256
rect 2466 8200 4170 8256
rect 2405 8198 4170 8200
rect 10869 8258 10935 8261
rect 14365 8258 14431 8261
rect 10869 8256 14431 8258
rect 10869 8200 10874 8256
rect 10930 8200 14370 8256
rect 14426 8200 14431 8256
rect 10869 8198 14431 8200
rect 2405 8195 2471 8198
rect 10869 8195 10935 8198
rect 14365 8195 14431 8198
rect 7984 8192 8300 8193
rect 7984 8128 7990 8192
rect 8054 8128 8070 8192
rect 8134 8128 8150 8192
rect 8214 8128 8230 8192
rect 8294 8128 8300 8192
rect 7984 8127 8300 8128
rect 15574 8192 15890 8193
rect 15574 8128 15580 8192
rect 15644 8128 15660 8192
rect 15724 8128 15740 8192
rect 15804 8128 15820 8192
rect 15884 8128 15890 8192
rect 15574 8127 15890 8128
rect 23164 8192 23480 8193
rect 23164 8128 23170 8192
rect 23234 8128 23250 8192
rect 23314 8128 23330 8192
rect 23394 8128 23410 8192
rect 23474 8128 23480 8192
rect 23164 8127 23480 8128
rect 30754 8192 31070 8193
rect 30754 8128 30760 8192
rect 30824 8128 30840 8192
rect 30904 8128 30920 8192
rect 30984 8128 31000 8192
rect 31064 8128 31070 8192
rect 30754 8127 31070 8128
rect 2681 8122 2747 8125
rect 7649 8122 7715 8125
rect 2681 8120 7715 8122
rect 2681 8064 2686 8120
rect 2742 8064 7654 8120
rect 7710 8064 7715 8120
rect 2681 8062 7715 8064
rect 2681 8059 2747 8062
rect 7649 8059 7715 8062
rect 10501 8122 10567 8125
rect 12065 8122 12131 8125
rect 10501 8120 12131 8122
rect 10501 8064 10506 8120
rect 10562 8064 12070 8120
rect 12126 8064 12131 8120
rect 10501 8062 12131 8064
rect 10501 8059 10567 8062
rect 12065 8059 12131 8062
rect 13721 7986 13787 7989
rect 16665 7986 16731 7989
rect 13721 7984 16731 7986
rect 13721 7928 13726 7984
rect 13782 7928 16670 7984
rect 16726 7928 16731 7984
rect 13721 7926 16731 7928
rect 13721 7923 13787 7926
rect 16665 7923 16731 7926
rect 2221 7850 2287 7853
rect 6361 7850 6427 7853
rect 2221 7848 6427 7850
rect 2221 7792 2226 7848
rect 2282 7792 6366 7848
rect 6422 7792 6427 7848
rect 2221 7790 6427 7792
rect 2221 7787 2287 7790
rect 6361 7787 6427 7790
rect 9673 7850 9739 7853
rect 16205 7850 16271 7853
rect 9673 7848 16271 7850
rect 9673 7792 9678 7848
rect 9734 7792 16210 7848
rect 16266 7792 16271 7848
rect 9673 7790 16271 7792
rect 9673 7787 9739 7790
rect 16205 7787 16271 7790
rect 17217 7850 17283 7853
rect 30189 7850 30255 7853
rect 17217 7848 30255 7850
rect 17217 7792 17222 7848
rect 17278 7792 30194 7848
rect 30250 7792 30255 7848
rect 17217 7790 30255 7792
rect 17217 7787 17283 7790
rect 30189 7787 30255 7790
rect 14181 7714 14247 7717
rect 15561 7714 15627 7717
rect 14181 7712 15627 7714
rect 14181 7656 14186 7712
rect 14242 7656 15566 7712
rect 15622 7656 15627 7712
rect 14181 7654 15627 7656
rect 14181 7651 14247 7654
rect 15561 7651 15627 7654
rect 17769 7714 17835 7717
rect 18873 7714 18939 7717
rect 17769 7712 18939 7714
rect 17769 7656 17774 7712
rect 17830 7656 18878 7712
rect 18934 7656 18939 7712
rect 17769 7654 18939 7656
rect 17769 7651 17835 7654
rect 18873 7651 18939 7654
rect 4189 7648 4505 7649
rect 4189 7584 4195 7648
rect 4259 7584 4275 7648
rect 4339 7584 4355 7648
rect 4419 7584 4435 7648
rect 4499 7584 4505 7648
rect 4189 7583 4505 7584
rect 11779 7648 12095 7649
rect 11779 7584 11785 7648
rect 11849 7584 11865 7648
rect 11929 7584 11945 7648
rect 12009 7584 12025 7648
rect 12089 7584 12095 7648
rect 11779 7583 12095 7584
rect 19369 7648 19685 7649
rect 19369 7584 19375 7648
rect 19439 7584 19455 7648
rect 19519 7584 19535 7648
rect 19599 7584 19615 7648
rect 19679 7584 19685 7648
rect 19369 7583 19685 7584
rect 26959 7648 27275 7649
rect 26959 7584 26965 7648
rect 27029 7584 27045 7648
rect 27109 7584 27125 7648
rect 27189 7584 27205 7648
rect 27269 7584 27275 7648
rect 26959 7583 27275 7584
rect 6729 7442 6795 7445
rect 15653 7442 15719 7445
rect 6729 7440 15719 7442
rect 6729 7384 6734 7440
rect 6790 7384 15658 7440
rect 15714 7384 15719 7440
rect 6729 7382 15719 7384
rect 6729 7379 6795 7382
rect 15653 7379 15719 7382
rect 24117 7442 24183 7445
rect 26141 7442 26207 7445
rect 24117 7440 26207 7442
rect 24117 7384 24122 7440
rect 24178 7384 26146 7440
rect 26202 7384 26207 7440
rect 24117 7382 26207 7384
rect 24117 7379 24183 7382
rect 26141 7379 26207 7382
rect 2865 7306 2931 7309
rect 17585 7306 17651 7309
rect 2865 7304 17651 7306
rect 2865 7248 2870 7304
rect 2926 7248 17590 7304
rect 17646 7248 17651 7304
rect 2865 7246 17651 7248
rect 2865 7243 2931 7246
rect 17585 7243 17651 7246
rect 20621 7306 20687 7309
rect 27889 7306 27955 7309
rect 20621 7304 27955 7306
rect 20621 7248 20626 7304
rect 20682 7248 27894 7304
rect 27950 7248 27955 7304
rect 20621 7246 27955 7248
rect 20621 7243 20687 7246
rect 27889 7243 27955 7246
rect 4429 7170 4495 7173
rect 5625 7170 5691 7173
rect 7833 7170 7899 7173
rect 4429 7168 7899 7170
rect 4429 7112 4434 7168
rect 4490 7112 5630 7168
rect 5686 7112 7838 7168
rect 7894 7112 7899 7168
rect 4429 7110 7899 7112
rect 4429 7107 4495 7110
rect 5625 7107 5691 7110
rect 7833 7107 7899 7110
rect 11605 7170 11671 7173
rect 14917 7170 14983 7173
rect 11605 7168 14983 7170
rect 11605 7112 11610 7168
rect 11666 7112 14922 7168
rect 14978 7112 14983 7168
rect 11605 7110 14983 7112
rect 11605 7107 11671 7110
rect 14917 7107 14983 7110
rect 7984 7104 8300 7105
rect 7984 7040 7990 7104
rect 8054 7040 8070 7104
rect 8134 7040 8150 7104
rect 8214 7040 8230 7104
rect 8294 7040 8300 7104
rect 7984 7039 8300 7040
rect 15574 7104 15890 7105
rect 15574 7040 15580 7104
rect 15644 7040 15660 7104
rect 15724 7040 15740 7104
rect 15804 7040 15820 7104
rect 15884 7040 15890 7104
rect 15574 7039 15890 7040
rect 23164 7104 23480 7105
rect 23164 7040 23170 7104
rect 23234 7040 23250 7104
rect 23314 7040 23330 7104
rect 23394 7040 23410 7104
rect 23474 7040 23480 7104
rect 23164 7039 23480 7040
rect 30754 7104 31070 7105
rect 30754 7040 30760 7104
rect 30824 7040 30840 7104
rect 30904 7040 30920 7104
rect 30984 7040 31000 7104
rect 31064 7040 31070 7104
rect 30754 7039 31070 7040
rect 1577 7034 1643 7037
rect 3141 7034 3207 7037
rect 4613 7034 4679 7037
rect 1577 7032 4679 7034
rect 1577 6976 1582 7032
rect 1638 6976 3146 7032
rect 3202 6976 4618 7032
rect 4674 6976 4679 7032
rect 1577 6974 4679 6976
rect 1577 6971 1643 6974
rect 3141 6971 3207 6974
rect 4613 6971 4679 6974
rect 2773 6900 2839 6901
rect 2773 6896 2820 6900
rect 2884 6898 2890 6900
rect 3877 6898 3943 6901
rect 5809 6898 5875 6901
rect 2773 6840 2778 6896
rect 2773 6836 2820 6840
rect 2884 6838 2930 6898
rect 3877 6896 5875 6898
rect 3877 6840 3882 6896
rect 3938 6840 5814 6896
rect 5870 6840 5875 6896
rect 3877 6838 5875 6840
rect 2884 6836 2890 6838
rect 2773 6835 2839 6836
rect 3877 6835 3943 6838
rect 5809 6835 5875 6838
rect 6361 6898 6427 6901
rect 13721 6898 13787 6901
rect 6361 6896 13787 6898
rect 6361 6840 6366 6896
rect 6422 6840 13726 6896
rect 13782 6840 13787 6896
rect 6361 6838 13787 6840
rect 6361 6835 6427 6838
rect 13721 6835 13787 6838
rect 13905 6898 13971 6901
rect 16389 6898 16455 6901
rect 13905 6896 16455 6898
rect 13905 6840 13910 6896
rect 13966 6840 16394 6896
rect 16450 6840 16455 6896
rect 13905 6838 16455 6840
rect 13905 6835 13971 6838
rect 16389 6835 16455 6838
rect 18597 6898 18663 6901
rect 26969 6898 27035 6901
rect 18597 6896 27035 6898
rect 18597 6840 18602 6896
rect 18658 6840 26974 6896
rect 27030 6840 27035 6896
rect 18597 6838 27035 6840
rect 18597 6835 18663 6838
rect 26969 6835 27035 6838
rect 28574 6836 28580 6900
rect 28644 6898 28650 6900
rect 29545 6898 29611 6901
rect 28644 6896 29611 6898
rect 28644 6840 29550 6896
rect 29606 6840 29611 6896
rect 28644 6838 29611 6840
rect 28644 6836 28650 6838
rect 29545 6835 29611 6838
rect 1393 6762 1459 6765
rect 5165 6762 5231 6765
rect 1393 6760 5231 6762
rect 1393 6704 1398 6760
rect 1454 6704 5170 6760
rect 5226 6704 5231 6760
rect 1393 6702 5231 6704
rect 1393 6699 1459 6702
rect 5165 6699 5231 6702
rect 11053 6762 11119 6765
rect 15653 6762 15719 6765
rect 11053 6760 15719 6762
rect 11053 6704 11058 6760
rect 11114 6704 15658 6760
rect 15714 6704 15719 6760
rect 11053 6702 15719 6704
rect 11053 6699 11119 6702
rect 15653 6699 15719 6702
rect 19241 6762 19307 6765
rect 22553 6762 22619 6765
rect 19241 6760 22619 6762
rect 19241 6704 19246 6760
rect 19302 6704 22558 6760
rect 22614 6704 22619 6760
rect 19241 6702 22619 6704
rect 19241 6699 19307 6702
rect 22553 6699 22619 6702
rect 4189 6560 4505 6561
rect 4189 6496 4195 6560
rect 4259 6496 4275 6560
rect 4339 6496 4355 6560
rect 4419 6496 4435 6560
rect 4499 6496 4505 6560
rect 4189 6495 4505 6496
rect 11779 6560 12095 6561
rect 11779 6496 11785 6560
rect 11849 6496 11865 6560
rect 11929 6496 11945 6560
rect 12009 6496 12025 6560
rect 12089 6496 12095 6560
rect 11779 6495 12095 6496
rect 19369 6560 19685 6561
rect 19369 6496 19375 6560
rect 19439 6496 19455 6560
rect 19519 6496 19535 6560
rect 19599 6496 19615 6560
rect 19679 6496 19685 6560
rect 19369 6495 19685 6496
rect 26959 6560 27275 6561
rect 26959 6496 26965 6560
rect 27029 6496 27045 6560
rect 27109 6496 27125 6560
rect 27189 6496 27205 6560
rect 27269 6496 27275 6560
rect 26959 6495 27275 6496
rect 6085 6490 6151 6493
rect 6862 6490 6868 6492
rect 6085 6488 6868 6490
rect 6085 6432 6090 6488
rect 6146 6432 6868 6488
rect 6085 6430 6868 6432
rect 6085 6427 6151 6430
rect 6862 6428 6868 6430
rect 6932 6428 6938 6492
rect 7281 6490 7347 6493
rect 17125 6490 17191 6493
rect 18965 6490 19031 6493
rect 7281 6488 8034 6490
rect 7281 6432 7286 6488
rect 7342 6432 8034 6488
rect 7281 6430 8034 6432
rect 7281 6427 7347 6430
rect 2129 6354 2195 6357
rect 7741 6354 7807 6357
rect 2129 6352 7807 6354
rect 2129 6296 2134 6352
rect 2190 6296 7746 6352
rect 7802 6296 7807 6352
rect 2129 6294 7807 6296
rect 7974 6354 8034 6430
rect 17125 6488 19031 6490
rect 17125 6432 17130 6488
rect 17186 6432 18970 6488
rect 19026 6432 19031 6488
rect 17125 6430 19031 6432
rect 17125 6427 17191 6430
rect 18965 6427 19031 6430
rect 17401 6354 17467 6357
rect 7974 6352 17467 6354
rect 7974 6296 17406 6352
rect 17462 6296 17467 6352
rect 7974 6294 17467 6296
rect 2129 6291 2195 6294
rect 7741 6291 7807 6294
rect 17401 6291 17467 6294
rect 8385 6218 8451 6221
rect 12801 6218 12867 6221
rect 14641 6218 14707 6221
rect 8385 6216 14707 6218
rect 8385 6160 8390 6216
rect 8446 6160 12806 6216
rect 12862 6160 14646 6216
rect 14702 6160 14707 6216
rect 8385 6158 14707 6160
rect 8385 6155 8451 6158
rect 12801 6155 12867 6158
rect 14641 6155 14707 6158
rect 20989 6218 21055 6221
rect 24853 6218 24919 6221
rect 20989 6216 24919 6218
rect 20989 6160 20994 6216
rect 21050 6160 24858 6216
rect 24914 6160 24919 6216
rect 20989 6158 24919 6160
rect 20989 6155 21055 6158
rect 24853 6155 24919 6158
rect 5809 6082 5875 6085
rect 7649 6082 7715 6085
rect 5809 6080 7715 6082
rect 5809 6024 5814 6080
rect 5870 6024 7654 6080
rect 7710 6024 7715 6080
rect 5809 6022 7715 6024
rect 5809 6019 5875 6022
rect 7649 6019 7715 6022
rect 10593 6082 10659 6085
rect 11421 6082 11487 6085
rect 10593 6080 11487 6082
rect 10593 6024 10598 6080
rect 10654 6024 11426 6080
rect 11482 6024 11487 6080
rect 10593 6022 11487 6024
rect 10593 6019 10659 6022
rect 11421 6019 11487 6022
rect 7984 6016 8300 6017
rect 7984 5952 7990 6016
rect 8054 5952 8070 6016
rect 8134 5952 8150 6016
rect 8214 5952 8230 6016
rect 8294 5952 8300 6016
rect 7984 5951 8300 5952
rect 15574 6016 15890 6017
rect 15574 5952 15580 6016
rect 15644 5952 15660 6016
rect 15724 5952 15740 6016
rect 15804 5952 15820 6016
rect 15884 5952 15890 6016
rect 15574 5951 15890 5952
rect 23164 6016 23480 6017
rect 23164 5952 23170 6016
rect 23234 5952 23250 6016
rect 23314 5952 23330 6016
rect 23394 5952 23410 6016
rect 23474 5952 23480 6016
rect 23164 5951 23480 5952
rect 30754 6016 31070 6017
rect 30754 5952 30760 6016
rect 30824 5952 30840 6016
rect 30904 5952 30920 6016
rect 30984 5952 31000 6016
rect 31064 5952 31070 6016
rect 30754 5951 31070 5952
rect 2497 5946 2563 5949
rect 7005 5946 7071 5949
rect 2497 5944 7071 5946
rect 2497 5888 2502 5944
rect 2558 5888 7010 5944
rect 7066 5888 7071 5944
rect 2497 5886 7071 5888
rect 2497 5883 2563 5886
rect 7005 5883 7071 5886
rect 24117 5946 24183 5949
rect 26785 5946 26851 5949
rect 24117 5944 26851 5946
rect 24117 5888 24122 5944
rect 24178 5888 26790 5944
rect 26846 5888 26851 5944
rect 24117 5886 26851 5888
rect 24117 5883 24183 5886
rect 26785 5883 26851 5886
rect 1577 5810 1643 5813
rect 12341 5810 12407 5813
rect 1577 5808 12407 5810
rect 1577 5752 1582 5808
rect 1638 5752 12346 5808
rect 12402 5752 12407 5808
rect 1577 5750 12407 5752
rect 1577 5747 1643 5750
rect 12341 5747 12407 5750
rect 20621 5810 20687 5813
rect 22737 5810 22803 5813
rect 20621 5808 22803 5810
rect 20621 5752 20626 5808
rect 20682 5752 22742 5808
rect 22798 5752 22803 5808
rect 20621 5750 22803 5752
rect 20621 5747 20687 5750
rect 22737 5747 22803 5750
rect 1669 5674 1735 5677
rect 10685 5674 10751 5677
rect 1669 5672 10751 5674
rect 1669 5616 1674 5672
rect 1730 5616 10690 5672
rect 10746 5616 10751 5672
rect 1669 5614 10751 5616
rect 1669 5611 1735 5614
rect 10685 5611 10751 5614
rect 20621 5674 20687 5677
rect 21817 5674 21883 5677
rect 20621 5672 21883 5674
rect 20621 5616 20626 5672
rect 20682 5616 21822 5672
rect 21878 5616 21883 5672
rect 20621 5614 21883 5616
rect 20621 5611 20687 5614
rect 21817 5611 21883 5614
rect 22001 5674 22067 5677
rect 28073 5674 28139 5677
rect 22001 5672 28139 5674
rect 22001 5616 22006 5672
rect 22062 5616 28078 5672
rect 28134 5616 28139 5672
rect 22001 5614 28139 5616
rect 22001 5611 22067 5614
rect 28073 5611 28139 5614
rect 5625 5538 5691 5541
rect 6729 5538 6795 5541
rect 5625 5536 6795 5538
rect 5625 5480 5630 5536
rect 5686 5480 6734 5536
rect 6790 5480 6795 5536
rect 5625 5478 6795 5480
rect 5625 5475 5691 5478
rect 6729 5475 6795 5478
rect 4189 5472 4505 5473
rect 4189 5408 4195 5472
rect 4259 5408 4275 5472
rect 4339 5408 4355 5472
rect 4419 5408 4435 5472
rect 4499 5408 4505 5472
rect 4189 5407 4505 5408
rect 11779 5472 12095 5473
rect 11779 5408 11785 5472
rect 11849 5408 11865 5472
rect 11929 5408 11945 5472
rect 12009 5408 12025 5472
rect 12089 5408 12095 5472
rect 11779 5407 12095 5408
rect 19369 5472 19685 5473
rect 19369 5408 19375 5472
rect 19439 5408 19455 5472
rect 19519 5408 19535 5472
rect 19599 5408 19615 5472
rect 19679 5408 19685 5472
rect 19369 5407 19685 5408
rect 26959 5472 27275 5473
rect 26959 5408 26965 5472
rect 27029 5408 27045 5472
rect 27109 5408 27125 5472
rect 27189 5408 27205 5472
rect 27269 5408 27275 5472
rect 26959 5407 27275 5408
rect 2773 5266 2839 5269
rect 8937 5266 9003 5269
rect 2773 5264 9003 5266
rect 2773 5208 2778 5264
rect 2834 5208 8942 5264
rect 8998 5208 9003 5264
rect 2773 5206 9003 5208
rect 2773 5203 2839 5206
rect 8937 5203 9003 5206
rect 20161 5266 20227 5269
rect 29361 5266 29427 5269
rect 20161 5264 29427 5266
rect 20161 5208 20166 5264
rect 20222 5208 29366 5264
rect 29422 5208 29427 5264
rect 20161 5206 29427 5208
rect 20161 5203 20227 5206
rect 29361 5203 29427 5206
rect 2037 5130 2103 5133
rect 10777 5130 10843 5133
rect 2037 5128 10843 5130
rect 2037 5072 2042 5128
rect 2098 5072 10782 5128
rect 10838 5072 10843 5128
rect 2037 5070 10843 5072
rect 2037 5067 2103 5070
rect 10777 5067 10843 5070
rect 19241 5130 19307 5133
rect 29453 5130 29519 5133
rect 19241 5128 29519 5130
rect 19241 5072 19246 5128
rect 19302 5072 29458 5128
rect 29514 5072 29519 5128
rect 19241 5070 29519 5072
rect 19241 5067 19307 5070
rect 29453 5067 29519 5070
rect 7984 4928 8300 4929
rect 7984 4864 7990 4928
rect 8054 4864 8070 4928
rect 8134 4864 8150 4928
rect 8214 4864 8230 4928
rect 8294 4864 8300 4928
rect 7984 4863 8300 4864
rect 15574 4928 15890 4929
rect 15574 4864 15580 4928
rect 15644 4864 15660 4928
rect 15724 4864 15740 4928
rect 15804 4864 15820 4928
rect 15884 4864 15890 4928
rect 15574 4863 15890 4864
rect 23164 4928 23480 4929
rect 23164 4864 23170 4928
rect 23234 4864 23250 4928
rect 23314 4864 23330 4928
rect 23394 4864 23410 4928
rect 23474 4864 23480 4928
rect 23164 4863 23480 4864
rect 30754 4928 31070 4929
rect 30754 4864 30760 4928
rect 30824 4864 30840 4928
rect 30904 4864 30920 4928
rect 30984 4864 31000 4928
rect 31064 4864 31070 4928
rect 30754 4863 31070 4864
rect 11145 4858 11211 4861
rect 11973 4858 12039 4861
rect 11145 4856 12039 4858
rect 11145 4800 11150 4856
rect 11206 4800 11978 4856
rect 12034 4800 12039 4856
rect 11145 4798 12039 4800
rect 11145 4795 11211 4798
rect 11973 4795 12039 4798
rect 5901 4722 5967 4725
rect 27153 4722 27219 4725
rect 5901 4720 27219 4722
rect 5901 4664 5906 4720
rect 5962 4664 27158 4720
rect 27214 4664 27219 4720
rect 5901 4662 27219 4664
rect 5901 4659 5967 4662
rect 27153 4659 27219 4662
rect 3417 4586 3483 4589
rect 8845 4586 8911 4589
rect 3417 4584 8911 4586
rect 3417 4528 3422 4584
rect 3478 4528 8850 4584
rect 8906 4528 8911 4584
rect 3417 4526 8911 4528
rect 3417 4523 3483 4526
rect 8845 4523 8911 4526
rect 4981 4450 5047 4453
rect 6177 4450 6243 4453
rect 4981 4448 6243 4450
rect 4981 4392 4986 4448
rect 5042 4392 6182 4448
rect 6238 4392 6243 4448
rect 4981 4390 6243 4392
rect 4981 4387 5047 4390
rect 6177 4387 6243 4390
rect 4189 4384 4505 4385
rect 4189 4320 4195 4384
rect 4259 4320 4275 4384
rect 4339 4320 4355 4384
rect 4419 4320 4435 4384
rect 4499 4320 4505 4384
rect 4189 4319 4505 4320
rect 11779 4384 12095 4385
rect 11779 4320 11785 4384
rect 11849 4320 11865 4384
rect 11929 4320 11945 4384
rect 12009 4320 12025 4384
rect 12089 4320 12095 4384
rect 11779 4319 12095 4320
rect 19369 4384 19685 4385
rect 19369 4320 19375 4384
rect 19439 4320 19455 4384
rect 19519 4320 19535 4384
rect 19599 4320 19615 4384
rect 19679 4320 19685 4384
rect 19369 4319 19685 4320
rect 26959 4384 27275 4385
rect 26959 4320 26965 4384
rect 27029 4320 27045 4384
rect 27109 4320 27125 4384
rect 27189 4320 27205 4384
rect 27269 4320 27275 4384
rect 26959 4319 27275 4320
rect 2129 4178 2195 4181
rect 27705 4178 27771 4181
rect 2129 4176 27771 4178
rect 2129 4120 2134 4176
rect 2190 4120 27710 4176
rect 27766 4120 27771 4176
rect 2129 4118 27771 4120
rect 2129 4115 2195 4118
rect 27705 4115 27771 4118
rect 1301 4042 1367 4045
rect 2773 4042 2839 4045
rect 2957 4044 3023 4045
rect 2957 4042 3004 4044
rect 1301 4040 2839 4042
rect 1301 3984 1306 4040
rect 1362 3984 2778 4040
rect 2834 3984 2839 4040
rect 1301 3982 2839 3984
rect 2912 4040 3004 4042
rect 2912 3984 2962 4040
rect 2912 3982 3004 3984
rect 1301 3979 1367 3982
rect 2773 3979 2839 3982
rect 2957 3980 3004 3982
rect 3068 3980 3074 4044
rect 3693 4042 3759 4045
rect 5625 4042 5691 4045
rect 10409 4042 10475 4045
rect 29453 4042 29519 4045
rect 3693 4040 5691 4042
rect 3693 3984 3698 4040
rect 3754 3984 5630 4040
rect 5686 3984 5691 4040
rect 3693 3982 5691 3984
rect 2957 3979 3023 3980
rect 3693 3979 3759 3982
rect 5625 3979 5691 3982
rect 5766 4040 29519 4042
rect 5766 3984 10414 4040
rect 10470 3984 29458 4040
rect 29514 3984 29519 4040
rect 5766 3982 29519 3984
rect 933 3906 999 3909
rect 4613 3906 4679 3909
rect 4981 3906 5047 3909
rect 5766 3906 5826 3982
rect 10409 3979 10475 3982
rect 29453 3979 29519 3982
rect 933 3904 4679 3906
rect 933 3848 938 3904
rect 994 3848 4618 3904
rect 4674 3848 4679 3904
rect 933 3846 4679 3848
rect 933 3843 999 3846
rect 4613 3843 4679 3846
rect 4846 3904 5826 3906
rect 4846 3848 4986 3904
rect 5042 3848 5826 3904
rect 4846 3846 5826 3848
rect 18137 3906 18203 3909
rect 22921 3906 22987 3909
rect 18137 3904 22987 3906
rect 18137 3848 18142 3904
rect 18198 3848 22926 3904
rect 22982 3848 22987 3904
rect 18137 3846 22987 3848
rect 2773 3770 2839 3773
rect 3049 3770 3115 3773
rect 4846 3770 4906 3846
rect 4981 3843 5047 3846
rect 18137 3843 18203 3846
rect 22921 3843 22987 3846
rect 7984 3840 8300 3841
rect 7984 3776 7990 3840
rect 8054 3776 8070 3840
rect 8134 3776 8150 3840
rect 8214 3776 8230 3840
rect 8294 3776 8300 3840
rect 7984 3775 8300 3776
rect 15574 3840 15890 3841
rect 15574 3776 15580 3840
rect 15644 3776 15660 3840
rect 15724 3776 15740 3840
rect 15804 3776 15820 3840
rect 15884 3776 15890 3840
rect 15574 3775 15890 3776
rect 23164 3840 23480 3841
rect 23164 3776 23170 3840
rect 23234 3776 23250 3840
rect 23314 3776 23330 3840
rect 23394 3776 23410 3840
rect 23474 3776 23480 3840
rect 23164 3775 23480 3776
rect 30754 3840 31070 3841
rect 30754 3776 30760 3840
rect 30824 3776 30840 3840
rect 30904 3776 30920 3840
rect 30984 3776 31000 3840
rect 31064 3776 31070 3840
rect 30754 3775 31070 3776
rect 2773 3768 4906 3770
rect 2773 3712 2778 3768
rect 2834 3712 3054 3768
rect 3110 3712 4906 3768
rect 2773 3710 4906 3712
rect 16849 3770 16915 3773
rect 18873 3770 18939 3773
rect 16849 3768 18939 3770
rect 16849 3712 16854 3768
rect 16910 3712 18878 3768
rect 18934 3712 18939 3768
rect 16849 3710 18939 3712
rect 2773 3707 2839 3710
rect 3049 3707 3115 3710
rect 16849 3707 16915 3710
rect 18873 3707 18939 3710
rect 5625 3634 5691 3637
rect 16757 3634 16823 3637
rect 5625 3632 16823 3634
rect 5625 3576 5630 3632
rect 5686 3576 16762 3632
rect 16818 3576 16823 3632
rect 5625 3574 16823 3576
rect 5625 3571 5691 3574
rect 16757 3571 16823 3574
rect 17861 3634 17927 3637
rect 27797 3634 27863 3637
rect 17861 3632 27863 3634
rect 17861 3576 17866 3632
rect 17922 3576 27802 3632
rect 27858 3576 27863 3632
rect 17861 3574 27863 3576
rect 17861 3571 17927 3574
rect 27797 3571 27863 3574
rect 4521 3498 4587 3501
rect 9305 3498 9371 3501
rect 4521 3496 9371 3498
rect 4521 3440 4526 3496
rect 4582 3440 9310 3496
rect 9366 3440 9371 3496
rect 4521 3438 9371 3440
rect 4521 3435 4587 3438
rect 9305 3435 9371 3438
rect 18965 3498 19031 3501
rect 27245 3498 27311 3501
rect 18965 3496 27311 3498
rect 18965 3440 18970 3496
rect 19026 3440 27250 3496
rect 27306 3440 27311 3496
rect 18965 3438 27311 3440
rect 18965 3435 19031 3438
rect 27245 3435 27311 3438
rect 5441 3362 5507 3365
rect 8937 3362 9003 3365
rect 5441 3360 9003 3362
rect 5441 3304 5446 3360
rect 5502 3304 8942 3360
rect 8998 3304 9003 3360
rect 5441 3302 9003 3304
rect 5441 3299 5507 3302
rect 8937 3299 9003 3302
rect 4189 3296 4505 3297
rect 4189 3232 4195 3296
rect 4259 3232 4275 3296
rect 4339 3232 4355 3296
rect 4419 3232 4435 3296
rect 4499 3232 4505 3296
rect 4189 3231 4505 3232
rect 11779 3296 12095 3297
rect 11779 3232 11785 3296
rect 11849 3232 11865 3296
rect 11929 3232 11945 3296
rect 12009 3232 12025 3296
rect 12089 3232 12095 3296
rect 11779 3231 12095 3232
rect 19369 3296 19685 3297
rect 19369 3232 19375 3296
rect 19439 3232 19455 3296
rect 19519 3232 19535 3296
rect 19599 3232 19615 3296
rect 19679 3232 19685 3296
rect 19369 3231 19685 3232
rect 26959 3296 27275 3297
rect 26959 3232 26965 3296
rect 27029 3232 27045 3296
rect 27109 3232 27125 3296
rect 27189 3232 27205 3296
rect 27269 3232 27275 3296
rect 26959 3231 27275 3232
rect 4153 3090 4219 3093
rect 14733 3090 14799 3093
rect 4153 3088 14799 3090
rect 4153 3032 4158 3088
rect 4214 3032 14738 3088
rect 14794 3032 14799 3088
rect 4153 3030 14799 3032
rect 4153 3027 4219 3030
rect 14733 3027 14799 3030
rect 18045 3090 18111 3093
rect 19333 3090 19399 3093
rect 18045 3088 19399 3090
rect 18045 3032 18050 3088
rect 18106 3032 19338 3088
rect 19394 3032 19399 3088
rect 18045 3030 19399 3032
rect 18045 3027 18111 3030
rect 19333 3027 19399 3030
rect 22921 3090 22987 3093
rect 28717 3090 28783 3093
rect 22921 3088 28783 3090
rect 22921 3032 22926 3088
rect 22982 3032 28722 3088
rect 28778 3032 28783 3088
rect 22921 3030 28783 3032
rect 22921 3027 22987 3030
rect 28717 3027 28783 3030
rect 3049 2954 3115 2957
rect 28441 2954 28507 2957
rect 3049 2952 28507 2954
rect 3049 2896 3054 2952
rect 3110 2896 28446 2952
rect 28502 2896 28507 2952
rect 3049 2894 28507 2896
rect 3049 2891 3115 2894
rect 28441 2891 28507 2894
rect 3509 2818 3575 2821
rect 5073 2818 5139 2821
rect 6913 2818 6979 2821
rect 3509 2816 6979 2818
rect 3509 2760 3514 2816
rect 3570 2760 5078 2816
rect 5134 2760 6918 2816
rect 6974 2760 6979 2816
rect 3509 2758 6979 2760
rect 3509 2755 3575 2758
rect 5073 2755 5139 2758
rect 6913 2755 6979 2758
rect 7984 2752 8300 2753
rect 7984 2688 7990 2752
rect 8054 2688 8070 2752
rect 8134 2688 8150 2752
rect 8214 2688 8230 2752
rect 8294 2688 8300 2752
rect 7984 2687 8300 2688
rect 15574 2752 15890 2753
rect 15574 2688 15580 2752
rect 15644 2688 15660 2752
rect 15724 2688 15740 2752
rect 15804 2688 15820 2752
rect 15884 2688 15890 2752
rect 15574 2687 15890 2688
rect 23164 2752 23480 2753
rect 23164 2688 23170 2752
rect 23234 2688 23250 2752
rect 23314 2688 23330 2752
rect 23394 2688 23410 2752
rect 23474 2688 23480 2752
rect 23164 2687 23480 2688
rect 30754 2752 31070 2753
rect 30754 2688 30760 2752
rect 30824 2688 30840 2752
rect 30904 2688 30920 2752
rect 30984 2688 31000 2752
rect 31064 2688 31070 2752
rect 30754 2687 31070 2688
rect 3509 2682 3575 2685
rect 3969 2682 4035 2685
rect 5533 2684 5599 2685
rect 6637 2684 6703 2685
rect 5533 2682 5580 2684
rect 3509 2680 4035 2682
rect 3509 2624 3514 2680
rect 3570 2624 3974 2680
rect 4030 2624 4035 2680
rect 3509 2622 4035 2624
rect 5488 2680 5580 2682
rect 5488 2624 5538 2680
rect 5488 2622 5580 2624
rect 3509 2619 3575 2622
rect 3969 2619 4035 2622
rect 5533 2620 5580 2622
rect 5644 2620 5650 2684
rect 6637 2680 6684 2684
rect 6748 2682 6754 2684
rect 24025 2682 24091 2685
rect 24485 2682 24551 2685
rect 6637 2624 6642 2680
rect 6637 2620 6684 2624
rect 6748 2622 6794 2682
rect 24025 2680 24551 2682
rect 24025 2624 24030 2680
rect 24086 2624 24490 2680
rect 24546 2624 24551 2680
rect 24025 2622 24551 2624
rect 6748 2620 6754 2622
rect 5533 2619 5599 2620
rect 6637 2619 6703 2620
rect 24025 2619 24091 2622
rect 24485 2619 24551 2622
rect 4245 2546 4311 2549
rect 26325 2546 26391 2549
rect 4245 2544 26391 2546
rect 4245 2488 4250 2544
rect 4306 2488 26330 2544
rect 26386 2488 26391 2544
rect 4245 2486 26391 2488
rect 4245 2483 4311 2486
rect 26325 2483 26391 2486
rect 3785 2410 3851 2413
rect 12801 2410 12867 2413
rect 3785 2408 12867 2410
rect 3785 2352 3790 2408
rect 3846 2352 12806 2408
rect 12862 2352 12867 2408
rect 3785 2350 12867 2352
rect 3785 2347 3851 2350
rect 12801 2347 12867 2350
rect 20345 2410 20411 2413
rect 21633 2410 21699 2413
rect 20345 2408 21699 2410
rect 20345 2352 20350 2408
rect 20406 2352 21638 2408
rect 21694 2352 21699 2408
rect 20345 2350 21699 2352
rect 20345 2347 20411 2350
rect 21633 2347 21699 2350
rect 6085 2274 6151 2277
rect 7373 2274 7439 2277
rect 6085 2272 7439 2274
rect 6085 2216 6090 2272
rect 6146 2216 7378 2272
rect 7434 2216 7439 2272
rect 6085 2214 7439 2216
rect 6085 2211 6151 2214
rect 7373 2211 7439 2214
rect 23381 2274 23447 2277
rect 25497 2274 25563 2277
rect 23381 2272 25563 2274
rect 23381 2216 23386 2272
rect 23442 2216 25502 2272
rect 25558 2216 25563 2272
rect 23381 2214 25563 2216
rect 23381 2211 23447 2214
rect 25497 2211 25563 2214
rect 4189 2208 4505 2209
rect 4189 2144 4195 2208
rect 4259 2144 4275 2208
rect 4339 2144 4355 2208
rect 4419 2144 4435 2208
rect 4499 2144 4505 2208
rect 4189 2143 4505 2144
rect 11779 2208 12095 2209
rect 11779 2144 11785 2208
rect 11849 2144 11865 2208
rect 11929 2144 11945 2208
rect 12009 2144 12025 2208
rect 12089 2144 12095 2208
rect 11779 2143 12095 2144
rect 19369 2208 19685 2209
rect 19369 2144 19375 2208
rect 19439 2144 19455 2208
rect 19519 2144 19535 2208
rect 19599 2144 19615 2208
rect 19679 2144 19685 2208
rect 19369 2143 19685 2144
rect 26959 2208 27275 2209
rect 26959 2144 26965 2208
rect 27029 2144 27045 2208
rect 27109 2144 27125 2208
rect 27189 2144 27205 2208
rect 27269 2144 27275 2208
rect 26959 2143 27275 2144
rect 22829 2138 22895 2141
rect 26049 2138 26115 2141
rect 22829 2136 26115 2138
rect 22829 2080 22834 2136
rect 22890 2080 26054 2136
rect 26110 2080 26115 2136
rect 22829 2078 26115 2080
rect 22829 2075 22895 2078
rect 26049 2075 26115 2078
rect 4337 2002 4403 2005
rect 27521 2002 27587 2005
rect 4337 2000 27587 2002
rect 4337 1944 4342 2000
rect 4398 1944 27526 2000
rect 27582 1944 27587 2000
rect 4337 1942 27587 1944
rect 4337 1939 4403 1942
rect 27521 1939 27587 1942
rect 1761 1866 1827 1869
rect 6269 1866 6335 1869
rect 9121 1866 9187 1869
rect 1761 1864 6335 1866
rect 1761 1808 1766 1864
rect 1822 1808 6274 1864
rect 6330 1808 6335 1864
rect 1761 1806 6335 1808
rect 1761 1803 1827 1806
rect 6269 1803 6335 1806
rect 7790 1864 9187 1866
rect 7790 1808 9126 1864
rect 9182 1808 9187 1864
rect 7790 1806 9187 1808
rect 933 1730 999 1733
rect 4429 1730 4495 1733
rect 933 1728 4495 1730
rect 933 1672 938 1728
rect 994 1672 4434 1728
rect 4490 1672 4495 1728
rect 933 1670 4495 1672
rect 933 1667 999 1670
rect 4429 1667 4495 1670
rect 5073 1730 5139 1733
rect 5390 1730 5396 1732
rect 5073 1728 5396 1730
rect 5073 1672 5078 1728
rect 5134 1672 5396 1728
rect 5073 1670 5396 1672
rect 5073 1667 5139 1670
rect 5390 1668 5396 1670
rect 5460 1668 5466 1732
rect 5809 1730 5875 1733
rect 7790 1730 7850 1806
rect 9121 1803 9187 1806
rect 9305 1866 9371 1869
rect 12249 1866 12315 1869
rect 28809 1866 28875 1869
rect 9305 1864 28875 1866
rect 9305 1808 9310 1864
rect 9366 1808 12254 1864
rect 12310 1808 28814 1864
rect 28870 1808 28875 1864
rect 9305 1806 28875 1808
rect 9305 1803 9371 1806
rect 12249 1803 12315 1806
rect 28809 1803 28875 1806
rect 5809 1728 7850 1730
rect 5809 1672 5814 1728
rect 5870 1672 7850 1728
rect 5809 1670 7850 1672
rect 20989 1730 21055 1733
rect 21633 1730 21699 1733
rect 20989 1728 21699 1730
rect 20989 1672 20994 1728
rect 21050 1672 21638 1728
rect 21694 1672 21699 1728
rect 20989 1670 21699 1672
rect 5809 1667 5875 1670
rect 20989 1667 21055 1670
rect 21633 1667 21699 1670
rect 23749 1730 23815 1733
rect 25313 1730 25379 1733
rect 23749 1728 25379 1730
rect 23749 1672 23754 1728
rect 23810 1672 25318 1728
rect 25374 1672 25379 1728
rect 23749 1670 25379 1672
rect 23749 1667 23815 1670
rect 25313 1667 25379 1670
rect 7984 1664 8300 1665
rect 7984 1600 7990 1664
rect 8054 1600 8070 1664
rect 8134 1600 8150 1664
rect 8214 1600 8230 1664
rect 8294 1600 8300 1664
rect 7984 1599 8300 1600
rect 15574 1664 15890 1665
rect 15574 1600 15580 1664
rect 15644 1600 15660 1664
rect 15724 1600 15740 1664
rect 15804 1600 15820 1664
rect 15884 1600 15890 1664
rect 15574 1599 15890 1600
rect 23164 1664 23480 1665
rect 23164 1600 23170 1664
rect 23234 1600 23250 1664
rect 23314 1600 23330 1664
rect 23394 1600 23410 1664
rect 23474 1600 23480 1664
rect 23164 1599 23480 1600
rect 30754 1664 31070 1665
rect 30754 1600 30760 1664
rect 30824 1600 30840 1664
rect 30904 1600 30920 1664
rect 30984 1600 31000 1664
rect 31064 1600 31070 1664
rect 30754 1599 31070 1600
rect 5901 1594 5967 1597
rect 7741 1594 7807 1597
rect 19333 1594 19399 1597
rect 22829 1594 22895 1597
rect 5901 1592 7807 1594
rect 5901 1536 5906 1592
rect 5962 1536 7746 1592
rect 7802 1536 7807 1592
rect 5901 1534 7807 1536
rect 5901 1531 5967 1534
rect 7741 1531 7807 1534
rect 17726 1592 22895 1594
rect 17726 1536 19338 1592
rect 19394 1536 22834 1592
rect 22890 1536 22895 1592
rect 17726 1534 22895 1536
rect 3601 1458 3667 1461
rect 4245 1458 4311 1461
rect 3601 1456 4311 1458
rect 3601 1400 3606 1456
rect 3662 1400 4250 1456
rect 4306 1400 4311 1456
rect 3601 1398 4311 1400
rect 3601 1395 3667 1398
rect 4245 1395 4311 1398
rect 4429 1458 4495 1461
rect 11421 1458 11487 1461
rect 4429 1456 11487 1458
rect 4429 1400 4434 1456
rect 4490 1400 11426 1456
rect 11482 1400 11487 1456
rect 4429 1398 11487 1400
rect 4429 1395 4495 1398
rect 11421 1395 11487 1398
rect 14733 1458 14799 1461
rect 17726 1458 17786 1534
rect 19333 1531 19399 1534
rect 22829 1531 22895 1534
rect 14733 1456 17786 1458
rect 14733 1400 14738 1456
rect 14794 1400 17786 1456
rect 14733 1398 17786 1400
rect 17861 1458 17927 1461
rect 23749 1458 23815 1461
rect 17861 1456 23815 1458
rect 17861 1400 17866 1456
rect 17922 1400 23754 1456
rect 23810 1400 23815 1456
rect 17861 1398 23815 1400
rect 14733 1395 14799 1398
rect 17861 1395 17927 1398
rect 23749 1395 23815 1398
rect 23933 1458 23999 1461
rect 26417 1458 26483 1461
rect 23933 1456 26483 1458
rect 23933 1400 23938 1456
rect 23994 1400 26422 1456
rect 26478 1400 26483 1456
rect 23933 1398 26483 1400
rect 23933 1395 23999 1398
rect 26417 1395 26483 1398
rect 4245 1322 4311 1325
rect 26601 1322 26667 1325
rect 4245 1320 26667 1322
rect 4245 1264 4250 1320
rect 4306 1264 26606 1320
rect 26662 1264 26667 1320
rect 4245 1262 26667 1264
rect 4245 1259 4311 1262
rect 26601 1259 26667 1262
rect 5165 1186 5231 1189
rect 9673 1186 9739 1189
rect 5165 1184 9739 1186
rect 5165 1128 5170 1184
rect 5226 1128 9678 1184
rect 9734 1128 9739 1184
rect 5165 1126 9739 1128
rect 5165 1123 5231 1126
rect 9673 1123 9739 1126
rect 21357 1186 21423 1189
rect 25957 1186 26023 1189
rect 21357 1184 26023 1186
rect 21357 1128 21362 1184
rect 21418 1128 25962 1184
rect 26018 1128 26023 1184
rect 21357 1126 26023 1128
rect 21357 1123 21423 1126
rect 25957 1123 26023 1126
rect 4189 1120 4505 1121
rect 4189 1056 4195 1120
rect 4259 1056 4275 1120
rect 4339 1056 4355 1120
rect 4419 1056 4435 1120
rect 4499 1056 4505 1120
rect 4189 1055 4505 1056
rect 11779 1120 12095 1121
rect 11779 1056 11785 1120
rect 11849 1056 11865 1120
rect 11929 1056 11945 1120
rect 12009 1056 12025 1120
rect 12089 1056 12095 1120
rect 11779 1055 12095 1056
rect 19369 1120 19685 1121
rect 19369 1056 19375 1120
rect 19439 1056 19455 1120
rect 19519 1056 19535 1120
rect 19599 1056 19615 1120
rect 19679 1056 19685 1120
rect 19369 1055 19685 1056
rect 26959 1120 27275 1121
rect 26959 1056 26965 1120
rect 27029 1056 27045 1120
rect 27109 1056 27125 1120
rect 27189 1056 27205 1120
rect 27269 1056 27275 1120
rect 26959 1055 27275 1056
rect 5441 1050 5507 1053
rect 8293 1050 8359 1053
rect 5441 1048 8359 1050
rect 5441 992 5446 1048
rect 5502 992 8298 1048
rect 8354 992 8359 1048
rect 5441 990 8359 992
rect 5441 987 5507 990
rect 8293 987 8359 990
rect 4061 914 4127 917
rect 23473 914 23539 917
rect 4061 912 23539 914
rect 4061 856 4066 912
rect 4122 856 23478 912
rect 23534 856 23539 912
rect 4061 854 23539 856
rect 4061 851 4127 854
rect 23473 851 23539 854
rect 4613 778 4679 781
rect 29177 778 29243 781
rect 4613 776 29243 778
rect 4613 720 4618 776
rect 4674 720 29182 776
rect 29238 720 29243 776
rect 4613 718 29243 720
rect 4613 715 4679 718
rect 29177 715 29243 718
rect 7984 576 8300 577
rect 7984 512 7990 576
rect 8054 512 8070 576
rect 8134 512 8150 576
rect 8214 512 8230 576
rect 8294 512 8300 576
rect 7984 511 8300 512
rect 15574 576 15890 577
rect 15574 512 15580 576
rect 15644 512 15660 576
rect 15724 512 15740 576
rect 15804 512 15820 576
rect 15884 512 15890 576
rect 15574 511 15890 512
rect 23164 576 23480 577
rect 23164 512 23170 576
rect 23234 512 23250 576
rect 23314 512 23330 576
rect 23394 512 23410 576
rect 23474 512 23480 576
rect 23164 511 23480 512
rect 30754 576 31070 577
rect 30754 512 30760 576
rect 30824 512 30840 576
rect 30904 512 30920 576
rect 30984 512 31000 576
rect 31064 512 31070 576
rect 30754 511 31070 512
rect 9213 370 9279 373
rect 24945 370 25011 373
rect 9213 368 25011 370
rect 9213 312 9218 368
rect 9274 312 24950 368
rect 25006 312 25011 368
rect 9213 310 25011 312
rect 9213 307 9279 310
rect 24945 307 25011 310
rect 6637 234 6703 237
rect 18229 234 18295 237
rect 6637 232 18295 234
rect 6637 176 6642 232
rect 6698 176 18234 232
rect 18290 176 18295 232
rect 6637 174 18295 176
rect 6637 171 6703 174
rect 18229 171 18295 174
rect 3969 98 4035 101
rect 15285 98 15351 101
rect 3969 96 15351 98
rect 3969 40 3974 96
rect 4030 40 15290 96
rect 15346 40 15351 96
rect 3969 38 15351 40
rect 3969 35 4035 38
rect 15285 35 15351 38
rect 15561 98 15627 101
rect 24853 98 24919 101
rect 15561 96 24919 98
rect 15561 40 15566 96
rect 15622 40 24858 96
rect 24914 40 24919 96
rect 15561 38 24919 40
rect 15561 35 15627 38
rect 24853 35 24919 38
<< via3 >>
rect 14412 22264 14476 22268
rect 14412 22208 14426 22264
rect 14426 22208 14476 22264
rect 14412 22204 14476 22208
rect 2820 22068 2884 22132
rect 10916 21992 10980 21996
rect 10916 21936 10966 21992
rect 10966 21936 10980 21992
rect 10916 21932 10980 21936
rect 12020 21898 12084 21962
rect 13124 21898 13188 21962
rect 21956 21856 22020 21860
rect 21956 21800 21970 21856
rect 21970 21800 22020 21856
rect 21956 21796 22020 21800
rect 23612 21796 23676 21860
rect 4195 21788 4259 21792
rect 4195 21732 4199 21788
rect 4199 21732 4255 21788
rect 4255 21732 4259 21788
rect 4195 21728 4259 21732
rect 4275 21788 4339 21792
rect 4275 21732 4279 21788
rect 4279 21732 4335 21788
rect 4335 21732 4339 21788
rect 4275 21728 4339 21732
rect 4355 21788 4419 21792
rect 4355 21732 4359 21788
rect 4359 21732 4415 21788
rect 4415 21732 4419 21788
rect 4355 21728 4419 21732
rect 4435 21788 4499 21792
rect 4435 21732 4439 21788
rect 4439 21732 4495 21788
rect 4495 21732 4499 21788
rect 4435 21728 4499 21732
rect 11785 21788 11849 21792
rect 11785 21732 11789 21788
rect 11789 21732 11845 21788
rect 11845 21732 11849 21788
rect 11785 21728 11849 21732
rect 11865 21788 11929 21792
rect 11865 21732 11869 21788
rect 11869 21732 11925 21788
rect 11925 21732 11929 21788
rect 11865 21728 11929 21732
rect 11945 21788 12009 21792
rect 11945 21732 11949 21788
rect 11949 21732 12005 21788
rect 12005 21732 12009 21788
rect 11945 21728 12009 21732
rect 12025 21788 12089 21792
rect 12025 21732 12029 21788
rect 12029 21732 12085 21788
rect 12085 21732 12089 21788
rect 12025 21728 12089 21732
rect 19375 21788 19439 21792
rect 19375 21732 19379 21788
rect 19379 21732 19435 21788
rect 19435 21732 19439 21788
rect 19375 21728 19439 21732
rect 19455 21788 19519 21792
rect 19455 21732 19459 21788
rect 19459 21732 19515 21788
rect 19515 21732 19519 21788
rect 19455 21728 19519 21732
rect 19535 21788 19599 21792
rect 19535 21732 19539 21788
rect 19539 21732 19595 21788
rect 19595 21732 19599 21788
rect 19535 21728 19599 21732
rect 19615 21788 19679 21792
rect 19615 21732 19619 21788
rect 19619 21732 19675 21788
rect 19675 21732 19679 21788
rect 19615 21728 19679 21732
rect 26965 21788 27029 21792
rect 26965 21732 26969 21788
rect 26969 21732 27025 21788
rect 27025 21732 27029 21788
rect 26965 21728 27029 21732
rect 27045 21788 27109 21792
rect 27045 21732 27049 21788
rect 27049 21732 27105 21788
rect 27105 21732 27109 21788
rect 27045 21728 27109 21732
rect 27125 21788 27189 21792
rect 27125 21732 27129 21788
rect 27129 21732 27185 21788
rect 27185 21732 27189 21788
rect 27125 21728 27189 21732
rect 27205 21788 27269 21792
rect 27205 21732 27209 21788
rect 27209 21732 27265 21788
rect 27265 21732 27269 21788
rect 27205 21728 27269 21732
rect 10180 21252 10244 21316
rect 7990 21244 8054 21248
rect 7990 21188 7994 21244
rect 7994 21188 8050 21244
rect 8050 21188 8054 21244
rect 7990 21184 8054 21188
rect 8070 21244 8134 21248
rect 8070 21188 8074 21244
rect 8074 21188 8130 21244
rect 8130 21188 8134 21244
rect 8070 21184 8134 21188
rect 8150 21244 8214 21248
rect 8150 21188 8154 21244
rect 8154 21188 8210 21244
rect 8210 21188 8214 21244
rect 8150 21184 8214 21188
rect 8230 21244 8294 21248
rect 8230 21188 8234 21244
rect 8234 21188 8290 21244
rect 8290 21188 8294 21244
rect 8230 21184 8294 21188
rect 15580 21244 15644 21248
rect 15580 21188 15584 21244
rect 15584 21188 15640 21244
rect 15640 21188 15644 21244
rect 15580 21184 15644 21188
rect 15660 21244 15724 21248
rect 15660 21188 15664 21244
rect 15664 21188 15720 21244
rect 15720 21188 15724 21244
rect 15660 21184 15724 21188
rect 15740 21244 15804 21248
rect 15740 21188 15744 21244
rect 15744 21188 15800 21244
rect 15800 21188 15804 21244
rect 15740 21184 15804 21188
rect 15820 21244 15884 21248
rect 15820 21188 15824 21244
rect 15824 21188 15880 21244
rect 15880 21188 15884 21244
rect 15820 21184 15884 21188
rect 23170 21244 23234 21248
rect 23170 21188 23174 21244
rect 23174 21188 23230 21244
rect 23230 21188 23234 21244
rect 23170 21184 23234 21188
rect 23250 21244 23314 21248
rect 23250 21188 23254 21244
rect 23254 21188 23310 21244
rect 23310 21188 23314 21244
rect 23250 21184 23314 21188
rect 23330 21244 23394 21248
rect 23330 21188 23334 21244
rect 23334 21188 23390 21244
rect 23390 21188 23394 21244
rect 23330 21184 23394 21188
rect 23410 21244 23474 21248
rect 23410 21188 23414 21244
rect 23414 21188 23470 21244
rect 23470 21188 23474 21244
rect 23410 21184 23474 21188
rect 30760 21244 30824 21248
rect 30760 21188 30764 21244
rect 30764 21188 30820 21244
rect 30820 21188 30824 21244
rect 30760 21184 30824 21188
rect 30840 21244 30904 21248
rect 30840 21188 30844 21244
rect 30844 21188 30900 21244
rect 30900 21188 30904 21244
rect 30840 21184 30904 21188
rect 30920 21244 30984 21248
rect 30920 21188 30924 21244
rect 30924 21188 30980 21244
rect 30980 21188 30984 21244
rect 30920 21184 30984 21188
rect 31000 21244 31064 21248
rect 31000 21188 31004 21244
rect 31004 21188 31060 21244
rect 31060 21188 31064 21244
rect 31000 21184 31064 21188
rect 26372 21116 26436 21180
rect 25636 20980 25700 21044
rect 27660 20844 27724 20908
rect 8892 20708 8956 20772
rect 4195 20700 4259 20704
rect 4195 20644 4199 20700
rect 4199 20644 4255 20700
rect 4255 20644 4259 20700
rect 4195 20640 4259 20644
rect 4275 20700 4339 20704
rect 4275 20644 4279 20700
rect 4279 20644 4335 20700
rect 4335 20644 4339 20700
rect 4275 20640 4339 20644
rect 4355 20700 4419 20704
rect 4355 20644 4359 20700
rect 4359 20644 4415 20700
rect 4415 20644 4419 20700
rect 4355 20640 4419 20644
rect 4435 20700 4499 20704
rect 4435 20644 4439 20700
rect 4439 20644 4495 20700
rect 4495 20644 4499 20700
rect 4435 20640 4499 20644
rect 11785 20700 11849 20704
rect 11785 20644 11789 20700
rect 11789 20644 11845 20700
rect 11845 20644 11849 20700
rect 11785 20640 11849 20644
rect 11865 20700 11929 20704
rect 11865 20644 11869 20700
rect 11869 20644 11925 20700
rect 11925 20644 11929 20700
rect 11865 20640 11929 20644
rect 11945 20700 12009 20704
rect 11945 20644 11949 20700
rect 11949 20644 12005 20700
rect 12005 20644 12009 20700
rect 11945 20640 12009 20644
rect 12025 20700 12089 20704
rect 12025 20644 12029 20700
rect 12029 20644 12085 20700
rect 12085 20644 12089 20700
rect 12025 20640 12089 20644
rect 19375 20700 19439 20704
rect 19375 20644 19379 20700
rect 19379 20644 19435 20700
rect 19435 20644 19439 20700
rect 19375 20640 19439 20644
rect 19455 20700 19519 20704
rect 19455 20644 19459 20700
rect 19459 20644 19515 20700
rect 19515 20644 19519 20700
rect 19455 20640 19519 20644
rect 19535 20700 19599 20704
rect 19535 20644 19539 20700
rect 19539 20644 19595 20700
rect 19595 20644 19599 20700
rect 19535 20640 19599 20644
rect 19615 20700 19679 20704
rect 19615 20644 19619 20700
rect 19619 20644 19675 20700
rect 19675 20644 19679 20700
rect 19615 20640 19679 20644
rect 9628 20572 9692 20636
rect 10364 20572 10428 20636
rect 14228 20572 14292 20636
rect 24348 20708 24412 20772
rect 26965 20700 27029 20704
rect 26965 20644 26969 20700
rect 26969 20644 27025 20700
rect 27025 20644 27029 20700
rect 26965 20640 27029 20644
rect 27045 20700 27109 20704
rect 27045 20644 27049 20700
rect 27049 20644 27105 20700
rect 27105 20644 27109 20700
rect 27045 20640 27109 20644
rect 27125 20700 27189 20704
rect 27125 20644 27129 20700
rect 27129 20644 27185 20700
rect 27185 20644 27189 20700
rect 27125 20640 27189 20644
rect 27205 20700 27269 20704
rect 27205 20644 27209 20700
rect 27209 20644 27265 20700
rect 27265 20644 27269 20700
rect 27205 20640 27269 20644
rect 7990 20156 8054 20160
rect 7990 20100 7994 20156
rect 7994 20100 8050 20156
rect 8050 20100 8054 20156
rect 7990 20096 8054 20100
rect 8070 20156 8134 20160
rect 8070 20100 8074 20156
rect 8074 20100 8130 20156
rect 8130 20100 8134 20156
rect 8070 20096 8134 20100
rect 8150 20156 8214 20160
rect 8150 20100 8154 20156
rect 8154 20100 8210 20156
rect 8210 20100 8214 20156
rect 8150 20096 8214 20100
rect 8230 20156 8294 20160
rect 8230 20100 8234 20156
rect 8234 20100 8290 20156
rect 8290 20100 8294 20156
rect 8230 20096 8294 20100
rect 15580 20156 15644 20160
rect 15580 20100 15584 20156
rect 15584 20100 15640 20156
rect 15640 20100 15644 20156
rect 15580 20096 15644 20100
rect 15660 20156 15724 20160
rect 15660 20100 15664 20156
rect 15664 20100 15720 20156
rect 15720 20100 15724 20156
rect 15660 20096 15724 20100
rect 15740 20156 15804 20160
rect 15740 20100 15744 20156
rect 15744 20100 15800 20156
rect 15800 20100 15804 20156
rect 15740 20096 15804 20100
rect 15820 20156 15884 20160
rect 15820 20100 15824 20156
rect 15824 20100 15880 20156
rect 15880 20100 15884 20156
rect 15820 20096 15884 20100
rect 23170 20156 23234 20160
rect 23170 20100 23174 20156
rect 23174 20100 23230 20156
rect 23230 20100 23234 20156
rect 23170 20096 23234 20100
rect 23250 20156 23314 20160
rect 23250 20100 23254 20156
rect 23254 20100 23310 20156
rect 23310 20100 23314 20156
rect 23250 20096 23314 20100
rect 23330 20156 23394 20160
rect 23330 20100 23334 20156
rect 23334 20100 23390 20156
rect 23390 20100 23394 20156
rect 23330 20096 23394 20100
rect 23410 20156 23474 20160
rect 23410 20100 23414 20156
rect 23414 20100 23470 20156
rect 23470 20100 23474 20156
rect 23410 20096 23474 20100
rect 30760 20156 30824 20160
rect 30760 20100 30764 20156
rect 30764 20100 30820 20156
rect 30820 20100 30824 20156
rect 30760 20096 30824 20100
rect 30840 20156 30904 20160
rect 30840 20100 30844 20156
rect 30844 20100 30900 20156
rect 30900 20100 30904 20156
rect 30840 20096 30904 20100
rect 30920 20156 30984 20160
rect 30920 20100 30924 20156
rect 30924 20100 30980 20156
rect 30980 20100 30984 20156
rect 30920 20096 30984 20100
rect 31000 20156 31064 20160
rect 31000 20100 31004 20156
rect 31004 20100 31060 20156
rect 31060 20100 31064 20156
rect 31000 20096 31064 20100
rect 9444 20028 9508 20092
rect 9260 19756 9324 19820
rect 9628 19756 9692 19820
rect 4195 19612 4259 19616
rect 4195 19556 4199 19612
rect 4199 19556 4255 19612
rect 4255 19556 4259 19612
rect 4195 19552 4259 19556
rect 4275 19612 4339 19616
rect 4275 19556 4279 19612
rect 4279 19556 4335 19612
rect 4335 19556 4339 19612
rect 4275 19552 4339 19556
rect 4355 19612 4419 19616
rect 4355 19556 4359 19612
rect 4359 19556 4415 19612
rect 4415 19556 4419 19612
rect 4355 19552 4419 19556
rect 4435 19612 4499 19616
rect 4435 19556 4439 19612
rect 4439 19556 4495 19612
rect 4495 19556 4499 19612
rect 4435 19552 4499 19556
rect 11785 19612 11849 19616
rect 11785 19556 11789 19612
rect 11789 19556 11845 19612
rect 11845 19556 11849 19612
rect 11785 19552 11849 19556
rect 11865 19612 11929 19616
rect 11865 19556 11869 19612
rect 11869 19556 11925 19612
rect 11925 19556 11929 19612
rect 11865 19552 11929 19556
rect 11945 19612 12009 19616
rect 11945 19556 11949 19612
rect 11949 19556 12005 19612
rect 12005 19556 12009 19612
rect 11945 19552 12009 19556
rect 12025 19612 12089 19616
rect 12025 19556 12029 19612
rect 12029 19556 12085 19612
rect 12085 19556 12089 19612
rect 12025 19552 12089 19556
rect 19375 19612 19439 19616
rect 19375 19556 19379 19612
rect 19379 19556 19435 19612
rect 19435 19556 19439 19612
rect 19375 19552 19439 19556
rect 19455 19612 19519 19616
rect 19455 19556 19459 19612
rect 19459 19556 19515 19612
rect 19515 19556 19519 19612
rect 19455 19552 19519 19556
rect 19535 19612 19599 19616
rect 19535 19556 19539 19612
rect 19539 19556 19595 19612
rect 19595 19556 19599 19612
rect 19535 19552 19599 19556
rect 19615 19612 19679 19616
rect 19615 19556 19619 19612
rect 19619 19556 19675 19612
rect 19675 19556 19679 19612
rect 19615 19552 19679 19556
rect 26965 19612 27029 19616
rect 26965 19556 26969 19612
rect 26969 19556 27025 19612
rect 27025 19556 27029 19612
rect 26965 19552 27029 19556
rect 27045 19612 27109 19616
rect 27045 19556 27049 19612
rect 27049 19556 27105 19612
rect 27105 19556 27109 19612
rect 27045 19552 27109 19556
rect 27125 19612 27189 19616
rect 27125 19556 27129 19612
rect 27129 19556 27185 19612
rect 27185 19556 27189 19612
rect 27125 19552 27189 19556
rect 27205 19612 27269 19616
rect 27205 19556 27209 19612
rect 27209 19556 27265 19612
rect 27265 19556 27269 19612
rect 27205 19552 27269 19556
rect 4660 19212 4724 19276
rect 8524 19348 8588 19412
rect 9260 19348 9324 19412
rect 14044 19408 14108 19412
rect 14044 19352 14058 19408
rect 14058 19352 14108 19408
rect 14044 19348 14108 19352
rect 15148 19212 15212 19276
rect 22876 19212 22940 19276
rect 7990 19068 8054 19072
rect 7990 19012 7994 19068
rect 7994 19012 8050 19068
rect 8050 19012 8054 19068
rect 7990 19008 8054 19012
rect 8070 19068 8134 19072
rect 8070 19012 8074 19068
rect 8074 19012 8130 19068
rect 8130 19012 8134 19068
rect 8070 19008 8134 19012
rect 8150 19068 8214 19072
rect 8150 19012 8154 19068
rect 8154 19012 8210 19068
rect 8210 19012 8214 19068
rect 8150 19008 8214 19012
rect 8230 19068 8294 19072
rect 8230 19012 8234 19068
rect 8234 19012 8290 19068
rect 8290 19012 8294 19068
rect 8230 19008 8294 19012
rect 7788 18940 7852 19004
rect 11468 19076 11532 19140
rect 12204 19076 12268 19140
rect 16436 19136 16500 19140
rect 16436 19080 16486 19136
rect 16486 19080 16500 19136
rect 16436 19076 16500 19080
rect 16988 19076 17052 19140
rect 25268 19212 25332 19276
rect 26740 19076 26804 19140
rect 29316 19076 29380 19140
rect 15580 19068 15644 19072
rect 15580 19012 15584 19068
rect 15584 19012 15640 19068
rect 15640 19012 15644 19068
rect 15580 19008 15644 19012
rect 15660 19068 15724 19072
rect 15660 19012 15664 19068
rect 15664 19012 15720 19068
rect 15720 19012 15724 19068
rect 15660 19008 15724 19012
rect 15740 19068 15804 19072
rect 15740 19012 15744 19068
rect 15744 19012 15800 19068
rect 15800 19012 15804 19068
rect 15740 19008 15804 19012
rect 15820 19068 15884 19072
rect 15820 19012 15824 19068
rect 15824 19012 15880 19068
rect 15880 19012 15884 19068
rect 15820 19008 15884 19012
rect 23170 19068 23234 19072
rect 23170 19012 23174 19068
rect 23174 19012 23230 19068
rect 23230 19012 23234 19068
rect 23170 19008 23234 19012
rect 23250 19068 23314 19072
rect 23250 19012 23254 19068
rect 23254 19012 23310 19068
rect 23310 19012 23314 19068
rect 23250 19008 23314 19012
rect 23330 19068 23394 19072
rect 23330 19012 23334 19068
rect 23334 19012 23390 19068
rect 23390 19012 23394 19068
rect 23330 19008 23394 19012
rect 23410 19068 23474 19072
rect 23410 19012 23414 19068
rect 23414 19012 23470 19068
rect 23470 19012 23474 19068
rect 23410 19008 23474 19012
rect 30760 19068 30824 19072
rect 30760 19012 30764 19068
rect 30764 19012 30820 19068
rect 30820 19012 30824 19068
rect 30760 19008 30824 19012
rect 30840 19068 30904 19072
rect 30840 19012 30844 19068
rect 30844 19012 30900 19068
rect 30900 19012 30904 19068
rect 30840 19008 30904 19012
rect 30920 19068 30984 19072
rect 30920 19012 30924 19068
rect 30924 19012 30980 19068
rect 30980 19012 30984 19068
rect 30920 19008 30984 19012
rect 31000 19068 31064 19072
rect 31000 19012 31004 19068
rect 31004 19012 31060 19068
rect 31060 19012 31064 19068
rect 31000 19008 31064 19012
rect 9260 18940 9324 19004
rect 15332 18940 15396 19004
rect 16068 18804 16132 18868
rect 12572 18668 12636 18732
rect 4195 18524 4259 18528
rect 4195 18468 4199 18524
rect 4199 18468 4255 18524
rect 4255 18468 4259 18524
rect 4195 18464 4259 18468
rect 4275 18524 4339 18528
rect 4275 18468 4279 18524
rect 4279 18468 4335 18524
rect 4335 18468 4339 18524
rect 4275 18464 4339 18468
rect 4355 18524 4419 18528
rect 4355 18468 4359 18524
rect 4359 18468 4415 18524
rect 4415 18468 4419 18524
rect 4355 18464 4419 18468
rect 4435 18524 4499 18528
rect 4435 18468 4439 18524
rect 4439 18468 4495 18524
rect 4495 18468 4499 18524
rect 4435 18464 4499 18468
rect 11785 18524 11849 18528
rect 11785 18468 11789 18524
rect 11789 18468 11845 18524
rect 11845 18468 11849 18524
rect 11785 18464 11849 18468
rect 11865 18524 11929 18528
rect 11865 18468 11869 18524
rect 11869 18468 11925 18524
rect 11925 18468 11929 18524
rect 11865 18464 11929 18468
rect 11945 18524 12009 18528
rect 11945 18468 11949 18524
rect 11949 18468 12005 18524
rect 12005 18468 12009 18524
rect 11945 18464 12009 18468
rect 12025 18524 12089 18528
rect 12025 18468 12029 18524
rect 12029 18468 12085 18524
rect 12085 18468 12089 18524
rect 12025 18464 12089 18468
rect 5948 18396 6012 18460
rect 7420 18396 7484 18460
rect 7604 18456 7668 18460
rect 7604 18400 7654 18456
rect 7654 18400 7668 18456
rect 7604 18396 7668 18400
rect 22508 18532 22572 18596
rect 19375 18524 19439 18528
rect 19375 18468 19379 18524
rect 19379 18468 19435 18524
rect 19435 18468 19439 18524
rect 19375 18464 19439 18468
rect 19455 18524 19519 18528
rect 19455 18468 19459 18524
rect 19459 18468 19515 18524
rect 19515 18468 19519 18524
rect 19455 18464 19519 18468
rect 19535 18524 19599 18528
rect 19535 18468 19539 18524
rect 19539 18468 19595 18524
rect 19595 18468 19599 18524
rect 19535 18464 19599 18468
rect 19615 18524 19679 18528
rect 19615 18468 19619 18524
rect 19619 18468 19675 18524
rect 19675 18468 19679 18524
rect 19615 18464 19679 18468
rect 13676 18260 13740 18324
rect 24164 18396 24228 18460
rect 26965 18524 27029 18528
rect 26965 18468 26969 18524
rect 26969 18468 27025 18524
rect 27025 18468 27029 18524
rect 26965 18464 27029 18468
rect 27045 18524 27109 18528
rect 27045 18468 27049 18524
rect 27049 18468 27105 18524
rect 27105 18468 27109 18524
rect 27045 18464 27109 18468
rect 27125 18524 27189 18528
rect 27125 18468 27129 18524
rect 27129 18468 27185 18524
rect 27185 18468 27189 18524
rect 27125 18464 27189 18468
rect 27205 18524 27269 18528
rect 27205 18468 27209 18524
rect 27209 18468 27265 18524
rect 27265 18468 27269 18524
rect 27205 18464 27269 18468
rect 28396 18456 28460 18460
rect 28396 18400 28410 18456
rect 28410 18400 28460 18456
rect 28396 18396 28460 18400
rect 5212 17988 5276 18052
rect 5396 18048 5460 18052
rect 5396 17992 5410 18048
rect 5410 17992 5460 18048
rect 5396 17988 5460 17992
rect 6500 18048 6564 18052
rect 6500 17992 6514 18048
rect 6514 17992 6564 18048
rect 6500 17988 6564 17992
rect 7052 17988 7116 18052
rect 9444 18124 9508 18188
rect 15148 17988 15212 18052
rect 24164 17988 24228 18052
rect 30420 18048 30484 18052
rect 30420 17992 30434 18048
rect 30434 17992 30484 18048
rect 30420 17988 30484 17992
rect 7990 17980 8054 17984
rect 7990 17924 7994 17980
rect 7994 17924 8050 17980
rect 8050 17924 8054 17980
rect 7990 17920 8054 17924
rect 8070 17980 8134 17984
rect 8070 17924 8074 17980
rect 8074 17924 8130 17980
rect 8130 17924 8134 17980
rect 8070 17920 8134 17924
rect 8150 17980 8214 17984
rect 8150 17924 8154 17980
rect 8154 17924 8210 17980
rect 8210 17924 8214 17980
rect 8150 17920 8214 17924
rect 8230 17980 8294 17984
rect 8230 17924 8234 17980
rect 8234 17924 8290 17980
rect 8290 17924 8294 17980
rect 8230 17920 8294 17924
rect 15580 17980 15644 17984
rect 15580 17924 15584 17980
rect 15584 17924 15640 17980
rect 15640 17924 15644 17980
rect 15580 17920 15644 17924
rect 15660 17980 15724 17984
rect 15660 17924 15664 17980
rect 15664 17924 15720 17980
rect 15720 17924 15724 17980
rect 15660 17920 15724 17924
rect 15740 17980 15804 17984
rect 15740 17924 15744 17980
rect 15744 17924 15800 17980
rect 15800 17924 15804 17980
rect 15740 17920 15804 17924
rect 15820 17980 15884 17984
rect 15820 17924 15824 17980
rect 15824 17924 15880 17980
rect 15880 17924 15884 17980
rect 15820 17920 15884 17924
rect 23170 17980 23234 17984
rect 23170 17924 23174 17980
rect 23174 17924 23230 17980
rect 23230 17924 23234 17980
rect 23170 17920 23234 17924
rect 23250 17980 23314 17984
rect 23250 17924 23254 17980
rect 23254 17924 23310 17980
rect 23310 17924 23314 17980
rect 23250 17920 23314 17924
rect 23330 17980 23394 17984
rect 23330 17924 23334 17980
rect 23334 17924 23390 17980
rect 23390 17924 23394 17980
rect 23330 17920 23394 17924
rect 23410 17980 23474 17984
rect 23410 17924 23414 17980
rect 23414 17924 23470 17980
rect 23470 17924 23474 17980
rect 23410 17920 23474 17924
rect 30760 17980 30824 17984
rect 30760 17924 30764 17980
rect 30764 17924 30820 17980
rect 30820 17924 30824 17980
rect 30760 17920 30824 17924
rect 30840 17980 30904 17984
rect 30840 17924 30844 17980
rect 30844 17924 30900 17980
rect 30900 17924 30904 17980
rect 30840 17920 30904 17924
rect 30920 17980 30984 17984
rect 30920 17924 30924 17980
rect 30924 17924 30980 17980
rect 30980 17924 30984 17980
rect 30920 17920 30984 17924
rect 31000 17980 31064 17984
rect 31000 17924 31004 17980
rect 31004 17924 31060 17980
rect 31060 17924 31064 17980
rect 31000 17920 31064 17924
rect 16068 17852 16132 17916
rect 4195 17436 4259 17440
rect 4195 17380 4199 17436
rect 4199 17380 4255 17436
rect 4255 17380 4259 17436
rect 4195 17376 4259 17380
rect 4275 17436 4339 17440
rect 4275 17380 4279 17436
rect 4279 17380 4335 17436
rect 4335 17380 4339 17436
rect 4275 17376 4339 17380
rect 4355 17436 4419 17440
rect 4355 17380 4359 17436
rect 4359 17380 4415 17436
rect 4415 17380 4419 17436
rect 4355 17376 4419 17380
rect 4435 17436 4499 17440
rect 4435 17380 4439 17436
rect 4439 17380 4495 17436
rect 4495 17380 4499 17436
rect 4435 17376 4499 17380
rect 11785 17436 11849 17440
rect 11785 17380 11789 17436
rect 11789 17380 11845 17436
rect 11845 17380 11849 17436
rect 11785 17376 11849 17380
rect 11865 17436 11929 17440
rect 11865 17380 11869 17436
rect 11869 17380 11925 17436
rect 11925 17380 11929 17436
rect 11865 17376 11929 17380
rect 11945 17436 12009 17440
rect 11945 17380 11949 17436
rect 11949 17380 12005 17436
rect 12005 17380 12009 17436
rect 11945 17376 12009 17380
rect 12025 17436 12089 17440
rect 12025 17380 12029 17436
rect 12029 17380 12085 17436
rect 12085 17380 12089 17436
rect 12025 17376 12089 17380
rect 29500 17580 29564 17644
rect 19375 17436 19439 17440
rect 19375 17380 19379 17436
rect 19379 17380 19435 17436
rect 19435 17380 19439 17436
rect 19375 17376 19439 17380
rect 19455 17436 19519 17440
rect 19455 17380 19459 17436
rect 19459 17380 19515 17436
rect 19515 17380 19519 17436
rect 19455 17376 19519 17380
rect 19535 17436 19599 17440
rect 19535 17380 19539 17436
rect 19539 17380 19595 17436
rect 19595 17380 19599 17436
rect 19535 17376 19599 17380
rect 19615 17436 19679 17440
rect 19615 17380 19619 17436
rect 19619 17380 19675 17436
rect 19675 17380 19679 17436
rect 19615 17376 19679 17380
rect 26965 17436 27029 17440
rect 26965 17380 26969 17436
rect 26969 17380 27025 17436
rect 27025 17380 27029 17436
rect 26965 17376 27029 17380
rect 27045 17436 27109 17440
rect 27045 17380 27049 17436
rect 27049 17380 27105 17436
rect 27105 17380 27109 17436
rect 27045 17376 27109 17380
rect 27125 17436 27189 17440
rect 27125 17380 27129 17436
rect 27129 17380 27185 17436
rect 27185 17380 27189 17436
rect 27125 17376 27189 17380
rect 27205 17436 27269 17440
rect 27205 17380 27209 17436
rect 27209 17380 27265 17436
rect 27265 17380 27269 17436
rect 27205 17376 27269 17380
rect 8708 16960 8772 16964
rect 8708 16904 8722 16960
rect 8722 16904 8772 16960
rect 8708 16900 8772 16904
rect 27476 16900 27540 16964
rect 7990 16892 8054 16896
rect 7990 16836 7994 16892
rect 7994 16836 8050 16892
rect 8050 16836 8054 16892
rect 7990 16832 8054 16836
rect 8070 16892 8134 16896
rect 8070 16836 8074 16892
rect 8074 16836 8130 16892
rect 8130 16836 8134 16892
rect 8070 16832 8134 16836
rect 8150 16892 8214 16896
rect 8150 16836 8154 16892
rect 8154 16836 8210 16892
rect 8210 16836 8214 16892
rect 8150 16832 8214 16836
rect 8230 16892 8294 16896
rect 8230 16836 8234 16892
rect 8234 16836 8290 16892
rect 8290 16836 8294 16892
rect 8230 16832 8294 16836
rect 15580 16892 15644 16896
rect 15580 16836 15584 16892
rect 15584 16836 15640 16892
rect 15640 16836 15644 16892
rect 15580 16832 15644 16836
rect 15660 16892 15724 16896
rect 15660 16836 15664 16892
rect 15664 16836 15720 16892
rect 15720 16836 15724 16892
rect 15660 16832 15724 16836
rect 15740 16892 15804 16896
rect 15740 16836 15744 16892
rect 15744 16836 15800 16892
rect 15800 16836 15804 16892
rect 15740 16832 15804 16836
rect 15820 16892 15884 16896
rect 15820 16836 15824 16892
rect 15824 16836 15880 16892
rect 15880 16836 15884 16892
rect 15820 16832 15884 16836
rect 23170 16892 23234 16896
rect 23170 16836 23174 16892
rect 23174 16836 23230 16892
rect 23230 16836 23234 16892
rect 23170 16832 23234 16836
rect 23250 16892 23314 16896
rect 23250 16836 23254 16892
rect 23254 16836 23310 16892
rect 23310 16836 23314 16892
rect 23250 16832 23314 16836
rect 23330 16892 23394 16896
rect 23330 16836 23334 16892
rect 23334 16836 23390 16892
rect 23390 16836 23394 16892
rect 23330 16832 23394 16836
rect 23410 16892 23474 16896
rect 23410 16836 23414 16892
rect 23414 16836 23470 16892
rect 23470 16836 23474 16892
rect 23410 16832 23474 16836
rect 26188 16764 26252 16828
rect 10732 16628 10796 16692
rect 29684 16628 29748 16692
rect 30760 16892 30824 16896
rect 30760 16836 30764 16892
rect 30764 16836 30820 16892
rect 30820 16836 30824 16892
rect 30760 16832 30824 16836
rect 30840 16892 30904 16896
rect 30840 16836 30844 16892
rect 30844 16836 30900 16892
rect 30900 16836 30904 16892
rect 30840 16832 30904 16836
rect 30920 16892 30984 16896
rect 30920 16836 30924 16892
rect 30924 16836 30980 16892
rect 30980 16836 30984 16892
rect 30920 16832 30984 16836
rect 31000 16892 31064 16896
rect 31000 16836 31004 16892
rect 31004 16836 31060 16892
rect 31060 16836 31064 16892
rect 31000 16832 31064 16836
rect 8524 16356 8588 16420
rect 9444 16356 9508 16420
rect 4195 16348 4259 16352
rect 4195 16292 4199 16348
rect 4199 16292 4255 16348
rect 4255 16292 4259 16348
rect 4195 16288 4259 16292
rect 4275 16348 4339 16352
rect 4275 16292 4279 16348
rect 4279 16292 4335 16348
rect 4335 16292 4339 16348
rect 4275 16288 4339 16292
rect 4355 16348 4419 16352
rect 4355 16292 4359 16348
rect 4359 16292 4415 16348
rect 4415 16292 4419 16348
rect 4355 16288 4419 16292
rect 4435 16348 4499 16352
rect 4435 16292 4439 16348
rect 4439 16292 4495 16348
rect 4495 16292 4499 16348
rect 4435 16288 4499 16292
rect 11785 16348 11849 16352
rect 11785 16292 11789 16348
rect 11789 16292 11845 16348
rect 11845 16292 11849 16348
rect 11785 16288 11849 16292
rect 11865 16348 11929 16352
rect 11865 16292 11869 16348
rect 11869 16292 11925 16348
rect 11925 16292 11929 16348
rect 11865 16288 11929 16292
rect 11945 16348 12009 16352
rect 11945 16292 11949 16348
rect 11949 16292 12005 16348
rect 12005 16292 12009 16348
rect 11945 16288 12009 16292
rect 12025 16348 12089 16352
rect 12025 16292 12029 16348
rect 12029 16292 12085 16348
rect 12085 16292 12089 16348
rect 12025 16288 12089 16292
rect 19375 16348 19439 16352
rect 19375 16292 19379 16348
rect 19379 16292 19435 16348
rect 19435 16292 19439 16348
rect 19375 16288 19439 16292
rect 19455 16348 19519 16352
rect 19455 16292 19459 16348
rect 19459 16292 19515 16348
rect 19515 16292 19519 16348
rect 19455 16288 19519 16292
rect 19535 16348 19599 16352
rect 19535 16292 19539 16348
rect 19539 16292 19595 16348
rect 19595 16292 19599 16348
rect 19535 16288 19599 16292
rect 19615 16348 19679 16352
rect 19615 16292 19619 16348
rect 19619 16292 19675 16348
rect 19675 16292 19679 16348
rect 19615 16288 19679 16292
rect 26965 16348 27029 16352
rect 26965 16292 26969 16348
rect 26969 16292 27025 16348
rect 27025 16292 27029 16348
rect 26965 16288 27029 16292
rect 27045 16348 27109 16352
rect 27045 16292 27049 16348
rect 27049 16292 27105 16348
rect 27105 16292 27109 16348
rect 27045 16288 27109 16292
rect 27125 16348 27189 16352
rect 27125 16292 27129 16348
rect 27129 16292 27185 16348
rect 27185 16292 27189 16348
rect 27125 16288 27189 16292
rect 27205 16348 27269 16352
rect 27205 16292 27209 16348
rect 27209 16292 27265 16348
rect 27265 16292 27269 16348
rect 27205 16288 27269 16292
rect 24164 16220 24228 16284
rect 29316 15812 29380 15876
rect 7990 15804 8054 15808
rect 7990 15748 7994 15804
rect 7994 15748 8050 15804
rect 8050 15748 8054 15804
rect 7990 15744 8054 15748
rect 8070 15804 8134 15808
rect 8070 15748 8074 15804
rect 8074 15748 8130 15804
rect 8130 15748 8134 15804
rect 8070 15744 8134 15748
rect 8150 15804 8214 15808
rect 8150 15748 8154 15804
rect 8154 15748 8210 15804
rect 8210 15748 8214 15804
rect 8150 15744 8214 15748
rect 8230 15804 8294 15808
rect 8230 15748 8234 15804
rect 8234 15748 8290 15804
rect 8290 15748 8294 15804
rect 8230 15744 8294 15748
rect 15580 15804 15644 15808
rect 15580 15748 15584 15804
rect 15584 15748 15640 15804
rect 15640 15748 15644 15804
rect 15580 15744 15644 15748
rect 15660 15804 15724 15808
rect 15660 15748 15664 15804
rect 15664 15748 15720 15804
rect 15720 15748 15724 15804
rect 15660 15744 15724 15748
rect 15740 15804 15804 15808
rect 15740 15748 15744 15804
rect 15744 15748 15800 15804
rect 15800 15748 15804 15804
rect 15740 15744 15804 15748
rect 15820 15804 15884 15808
rect 15820 15748 15824 15804
rect 15824 15748 15880 15804
rect 15880 15748 15884 15804
rect 15820 15744 15884 15748
rect 23170 15804 23234 15808
rect 23170 15748 23174 15804
rect 23174 15748 23230 15804
rect 23230 15748 23234 15804
rect 23170 15744 23234 15748
rect 23250 15804 23314 15808
rect 23250 15748 23254 15804
rect 23254 15748 23310 15804
rect 23310 15748 23314 15804
rect 23250 15744 23314 15748
rect 23330 15804 23394 15808
rect 23330 15748 23334 15804
rect 23334 15748 23390 15804
rect 23390 15748 23394 15804
rect 23330 15744 23394 15748
rect 23410 15804 23474 15808
rect 23410 15748 23414 15804
rect 23414 15748 23470 15804
rect 23470 15748 23474 15804
rect 23410 15744 23474 15748
rect 30760 15804 30824 15808
rect 30760 15748 30764 15804
rect 30764 15748 30820 15804
rect 30820 15748 30824 15804
rect 30760 15744 30824 15748
rect 30840 15804 30904 15808
rect 30840 15748 30844 15804
rect 30844 15748 30900 15804
rect 30900 15748 30904 15804
rect 30840 15744 30904 15748
rect 30920 15804 30984 15808
rect 30920 15748 30924 15804
rect 30924 15748 30980 15804
rect 30980 15748 30984 15804
rect 30920 15744 30984 15748
rect 31000 15804 31064 15808
rect 31000 15748 31004 15804
rect 31004 15748 31060 15804
rect 31060 15748 31064 15804
rect 31000 15744 31064 15748
rect 9444 15404 9508 15468
rect 9628 15404 9692 15468
rect 29684 15540 29748 15604
rect 30420 15540 30484 15604
rect 4195 15260 4259 15264
rect 4195 15204 4199 15260
rect 4199 15204 4255 15260
rect 4255 15204 4259 15260
rect 4195 15200 4259 15204
rect 4275 15260 4339 15264
rect 4275 15204 4279 15260
rect 4279 15204 4335 15260
rect 4335 15204 4339 15260
rect 4275 15200 4339 15204
rect 4355 15260 4419 15264
rect 4355 15204 4359 15260
rect 4359 15204 4415 15260
rect 4415 15204 4419 15260
rect 4355 15200 4419 15204
rect 4435 15260 4499 15264
rect 4435 15204 4439 15260
rect 4439 15204 4495 15260
rect 4495 15204 4499 15260
rect 4435 15200 4499 15204
rect 11785 15260 11849 15264
rect 11785 15204 11789 15260
rect 11789 15204 11845 15260
rect 11845 15204 11849 15260
rect 11785 15200 11849 15204
rect 11865 15260 11929 15264
rect 11865 15204 11869 15260
rect 11869 15204 11925 15260
rect 11925 15204 11929 15260
rect 11865 15200 11929 15204
rect 11945 15260 12009 15264
rect 11945 15204 11949 15260
rect 11949 15204 12005 15260
rect 12005 15204 12009 15260
rect 11945 15200 12009 15204
rect 12025 15260 12089 15264
rect 12025 15204 12029 15260
rect 12029 15204 12085 15260
rect 12085 15204 12089 15260
rect 12025 15200 12089 15204
rect 19375 15260 19439 15264
rect 19375 15204 19379 15260
rect 19379 15204 19435 15260
rect 19435 15204 19439 15260
rect 19375 15200 19439 15204
rect 19455 15260 19519 15264
rect 19455 15204 19459 15260
rect 19459 15204 19515 15260
rect 19515 15204 19519 15260
rect 19455 15200 19519 15204
rect 19535 15260 19599 15264
rect 19535 15204 19539 15260
rect 19539 15204 19595 15260
rect 19595 15204 19599 15260
rect 19535 15200 19599 15204
rect 19615 15260 19679 15264
rect 19615 15204 19619 15260
rect 19619 15204 19675 15260
rect 19675 15204 19679 15260
rect 19615 15200 19679 15204
rect 26965 15260 27029 15264
rect 26965 15204 26969 15260
rect 26969 15204 27025 15260
rect 27025 15204 27029 15260
rect 26965 15200 27029 15204
rect 27045 15260 27109 15264
rect 27045 15204 27049 15260
rect 27049 15204 27105 15260
rect 27105 15204 27109 15260
rect 27045 15200 27109 15204
rect 27125 15260 27189 15264
rect 27125 15204 27129 15260
rect 27129 15204 27185 15260
rect 27185 15204 27189 15260
rect 27125 15200 27189 15204
rect 27205 15260 27269 15264
rect 27205 15204 27209 15260
rect 27209 15204 27265 15260
rect 27265 15204 27269 15260
rect 27205 15200 27269 15204
rect 15148 15132 15212 15196
rect 29132 15404 29196 15468
rect 29500 15328 29564 15332
rect 29500 15272 29514 15328
rect 29514 15272 29564 15328
rect 29500 15268 29564 15272
rect 26188 14996 26252 15060
rect 26740 14996 26804 15060
rect 27660 14860 27724 14924
rect 7420 14724 7484 14788
rect 7990 14716 8054 14720
rect 7990 14660 7994 14716
rect 7994 14660 8050 14716
rect 8050 14660 8054 14716
rect 7990 14656 8054 14660
rect 8070 14716 8134 14720
rect 8070 14660 8074 14716
rect 8074 14660 8130 14716
rect 8130 14660 8134 14716
rect 8070 14656 8134 14660
rect 8150 14716 8214 14720
rect 8150 14660 8154 14716
rect 8154 14660 8210 14716
rect 8210 14660 8214 14716
rect 8150 14656 8214 14660
rect 8230 14716 8294 14720
rect 8230 14660 8234 14716
rect 8234 14660 8290 14716
rect 8290 14660 8294 14716
rect 8230 14656 8294 14660
rect 15580 14716 15644 14720
rect 15580 14660 15584 14716
rect 15584 14660 15640 14716
rect 15640 14660 15644 14716
rect 15580 14656 15644 14660
rect 15660 14716 15724 14720
rect 15660 14660 15664 14716
rect 15664 14660 15720 14716
rect 15720 14660 15724 14716
rect 15660 14656 15724 14660
rect 15740 14716 15804 14720
rect 15740 14660 15744 14716
rect 15744 14660 15800 14716
rect 15800 14660 15804 14716
rect 15740 14656 15804 14660
rect 15820 14716 15884 14720
rect 15820 14660 15824 14716
rect 15824 14660 15880 14716
rect 15880 14660 15884 14716
rect 15820 14656 15884 14660
rect 23170 14716 23234 14720
rect 23170 14660 23174 14716
rect 23174 14660 23230 14716
rect 23230 14660 23234 14716
rect 23170 14656 23234 14660
rect 23250 14716 23314 14720
rect 23250 14660 23254 14716
rect 23254 14660 23310 14716
rect 23310 14660 23314 14716
rect 23250 14656 23314 14660
rect 23330 14716 23394 14720
rect 23330 14660 23334 14716
rect 23334 14660 23390 14716
rect 23390 14660 23394 14716
rect 23330 14656 23394 14660
rect 23410 14716 23474 14720
rect 23410 14660 23414 14716
rect 23414 14660 23470 14716
rect 23470 14660 23474 14716
rect 23410 14656 23474 14660
rect 30760 14716 30824 14720
rect 30760 14660 30764 14716
rect 30764 14660 30820 14716
rect 30820 14660 30824 14716
rect 30760 14656 30824 14660
rect 30840 14716 30904 14720
rect 30840 14660 30844 14716
rect 30844 14660 30900 14716
rect 30900 14660 30904 14716
rect 30840 14656 30904 14660
rect 30920 14716 30984 14720
rect 30920 14660 30924 14716
rect 30924 14660 30980 14716
rect 30980 14660 30984 14716
rect 30920 14656 30984 14660
rect 31000 14716 31064 14720
rect 31000 14660 31004 14716
rect 31004 14660 31060 14716
rect 31060 14660 31064 14716
rect 31000 14656 31064 14660
rect 27476 14316 27540 14380
rect 4195 14172 4259 14176
rect 4195 14116 4199 14172
rect 4199 14116 4255 14172
rect 4255 14116 4259 14172
rect 4195 14112 4259 14116
rect 4275 14172 4339 14176
rect 4275 14116 4279 14172
rect 4279 14116 4335 14172
rect 4335 14116 4339 14172
rect 4275 14112 4339 14116
rect 4355 14172 4419 14176
rect 4355 14116 4359 14172
rect 4359 14116 4415 14172
rect 4415 14116 4419 14172
rect 4355 14112 4419 14116
rect 4435 14172 4499 14176
rect 4435 14116 4439 14172
rect 4439 14116 4495 14172
rect 4495 14116 4499 14172
rect 4435 14112 4499 14116
rect 11785 14172 11849 14176
rect 11785 14116 11789 14172
rect 11789 14116 11845 14172
rect 11845 14116 11849 14172
rect 11785 14112 11849 14116
rect 11865 14172 11929 14176
rect 11865 14116 11869 14172
rect 11869 14116 11925 14172
rect 11925 14116 11929 14172
rect 11865 14112 11929 14116
rect 11945 14172 12009 14176
rect 11945 14116 11949 14172
rect 11949 14116 12005 14172
rect 12005 14116 12009 14172
rect 11945 14112 12009 14116
rect 12025 14172 12089 14176
rect 12025 14116 12029 14172
rect 12029 14116 12085 14172
rect 12085 14116 12089 14172
rect 12025 14112 12089 14116
rect 19375 14172 19439 14176
rect 19375 14116 19379 14172
rect 19379 14116 19435 14172
rect 19435 14116 19439 14172
rect 19375 14112 19439 14116
rect 19455 14172 19519 14176
rect 19455 14116 19459 14172
rect 19459 14116 19515 14172
rect 19515 14116 19519 14172
rect 19455 14112 19519 14116
rect 19535 14172 19599 14176
rect 19535 14116 19539 14172
rect 19539 14116 19595 14172
rect 19595 14116 19599 14172
rect 19535 14112 19599 14116
rect 19615 14172 19679 14176
rect 19615 14116 19619 14172
rect 19619 14116 19675 14172
rect 19675 14116 19679 14172
rect 19615 14112 19679 14116
rect 26965 14172 27029 14176
rect 26965 14116 26969 14172
rect 26969 14116 27025 14172
rect 27025 14116 27029 14172
rect 26965 14112 27029 14116
rect 27045 14172 27109 14176
rect 27045 14116 27049 14172
rect 27049 14116 27105 14172
rect 27105 14116 27109 14172
rect 27045 14112 27109 14116
rect 27125 14172 27189 14176
rect 27125 14116 27129 14172
rect 27129 14116 27185 14172
rect 27185 14116 27189 14172
rect 27125 14112 27189 14116
rect 27205 14172 27269 14176
rect 27205 14116 27209 14172
rect 27209 14116 27265 14172
rect 27265 14116 27269 14172
rect 27205 14112 27269 14116
rect 4844 13636 4908 13700
rect 28580 13968 28644 13972
rect 28580 13912 28594 13968
rect 28594 13912 28644 13968
rect 28580 13908 28644 13912
rect 20668 13772 20732 13836
rect 28396 13772 28460 13836
rect 7990 13628 8054 13632
rect 7990 13572 7994 13628
rect 7994 13572 8050 13628
rect 8050 13572 8054 13628
rect 7990 13568 8054 13572
rect 8070 13628 8134 13632
rect 8070 13572 8074 13628
rect 8074 13572 8130 13628
rect 8130 13572 8134 13628
rect 8070 13568 8134 13572
rect 8150 13628 8214 13632
rect 8150 13572 8154 13628
rect 8154 13572 8210 13628
rect 8210 13572 8214 13628
rect 8150 13568 8214 13572
rect 8230 13628 8294 13632
rect 8230 13572 8234 13628
rect 8234 13572 8290 13628
rect 8290 13572 8294 13628
rect 8230 13568 8294 13572
rect 15580 13628 15644 13632
rect 15580 13572 15584 13628
rect 15584 13572 15640 13628
rect 15640 13572 15644 13628
rect 15580 13568 15644 13572
rect 15660 13628 15724 13632
rect 15660 13572 15664 13628
rect 15664 13572 15720 13628
rect 15720 13572 15724 13628
rect 15660 13568 15724 13572
rect 15740 13628 15804 13632
rect 15740 13572 15744 13628
rect 15744 13572 15800 13628
rect 15800 13572 15804 13628
rect 15740 13568 15804 13572
rect 15820 13628 15884 13632
rect 15820 13572 15824 13628
rect 15824 13572 15880 13628
rect 15880 13572 15884 13628
rect 15820 13568 15884 13572
rect 23170 13628 23234 13632
rect 23170 13572 23174 13628
rect 23174 13572 23230 13628
rect 23230 13572 23234 13628
rect 23170 13568 23234 13572
rect 23250 13628 23314 13632
rect 23250 13572 23254 13628
rect 23254 13572 23310 13628
rect 23310 13572 23314 13628
rect 23250 13568 23314 13572
rect 23330 13628 23394 13632
rect 23330 13572 23334 13628
rect 23334 13572 23390 13628
rect 23390 13572 23394 13628
rect 23330 13568 23394 13572
rect 23410 13628 23474 13632
rect 23410 13572 23414 13628
rect 23414 13572 23470 13628
rect 23470 13572 23474 13628
rect 23410 13568 23474 13572
rect 30760 13628 30824 13632
rect 30760 13572 30764 13628
rect 30764 13572 30820 13628
rect 30820 13572 30824 13628
rect 30760 13568 30824 13572
rect 30840 13628 30904 13632
rect 30840 13572 30844 13628
rect 30844 13572 30900 13628
rect 30900 13572 30904 13628
rect 30840 13568 30904 13572
rect 30920 13628 30984 13632
rect 30920 13572 30924 13628
rect 30924 13572 30980 13628
rect 30980 13572 30984 13628
rect 30920 13568 30984 13572
rect 31000 13628 31064 13632
rect 31000 13572 31004 13628
rect 31004 13572 31060 13628
rect 31060 13572 31064 13628
rect 31000 13568 31064 13572
rect 8524 13500 8588 13564
rect 5212 13092 5276 13156
rect 4195 13084 4259 13088
rect 4195 13028 4199 13084
rect 4199 13028 4255 13084
rect 4255 13028 4259 13084
rect 4195 13024 4259 13028
rect 4275 13084 4339 13088
rect 4275 13028 4279 13084
rect 4279 13028 4335 13084
rect 4335 13028 4339 13084
rect 4275 13024 4339 13028
rect 4355 13084 4419 13088
rect 4355 13028 4359 13084
rect 4359 13028 4415 13084
rect 4415 13028 4419 13084
rect 4355 13024 4419 13028
rect 4435 13084 4499 13088
rect 4435 13028 4439 13084
rect 4439 13028 4495 13084
rect 4495 13028 4499 13084
rect 4435 13024 4499 13028
rect 11785 13084 11849 13088
rect 11785 13028 11789 13084
rect 11789 13028 11845 13084
rect 11845 13028 11849 13084
rect 11785 13024 11849 13028
rect 11865 13084 11929 13088
rect 11865 13028 11869 13084
rect 11869 13028 11925 13084
rect 11925 13028 11929 13084
rect 11865 13024 11929 13028
rect 11945 13084 12009 13088
rect 11945 13028 11949 13084
rect 11949 13028 12005 13084
rect 12005 13028 12009 13084
rect 11945 13024 12009 13028
rect 12025 13084 12089 13088
rect 12025 13028 12029 13084
rect 12029 13028 12085 13084
rect 12085 13028 12089 13084
rect 12025 13024 12089 13028
rect 19375 13084 19439 13088
rect 19375 13028 19379 13084
rect 19379 13028 19435 13084
rect 19435 13028 19439 13084
rect 19375 13024 19439 13028
rect 19455 13084 19519 13088
rect 19455 13028 19459 13084
rect 19459 13028 19515 13084
rect 19515 13028 19519 13084
rect 19455 13024 19519 13028
rect 19535 13084 19599 13088
rect 19535 13028 19539 13084
rect 19539 13028 19595 13084
rect 19595 13028 19599 13084
rect 19535 13024 19599 13028
rect 19615 13084 19679 13088
rect 19615 13028 19619 13084
rect 19619 13028 19675 13084
rect 19675 13028 19679 13084
rect 19615 13024 19679 13028
rect 26965 13084 27029 13088
rect 26965 13028 26969 13084
rect 26969 13028 27025 13084
rect 27025 13028 27029 13084
rect 26965 13024 27029 13028
rect 27045 13084 27109 13088
rect 27045 13028 27049 13084
rect 27049 13028 27105 13084
rect 27105 13028 27109 13084
rect 27045 13024 27109 13028
rect 27125 13084 27189 13088
rect 27125 13028 27129 13084
rect 27129 13028 27185 13084
rect 27185 13028 27189 13084
rect 27125 13024 27189 13028
rect 27205 13084 27269 13088
rect 27205 13028 27209 13084
rect 27209 13028 27265 13084
rect 27265 13028 27269 13084
rect 27205 13024 27269 13028
rect 9076 12956 9140 13020
rect 9444 12956 9508 13020
rect 8708 12820 8772 12884
rect 19748 12820 19812 12884
rect 3004 12412 3068 12476
rect 12204 12608 12268 12612
rect 12204 12552 12218 12608
rect 12218 12552 12268 12608
rect 12204 12548 12268 12552
rect 13492 12608 13556 12612
rect 13492 12552 13506 12608
rect 13506 12552 13556 12608
rect 7990 12540 8054 12544
rect 7990 12484 7994 12540
rect 7994 12484 8050 12540
rect 8050 12484 8054 12540
rect 7990 12480 8054 12484
rect 8070 12540 8134 12544
rect 8070 12484 8074 12540
rect 8074 12484 8130 12540
rect 8130 12484 8134 12540
rect 8070 12480 8134 12484
rect 8150 12540 8214 12544
rect 8150 12484 8154 12540
rect 8154 12484 8210 12540
rect 8210 12484 8214 12540
rect 8150 12480 8214 12484
rect 8230 12540 8294 12544
rect 8230 12484 8234 12540
rect 8234 12484 8290 12540
rect 8290 12484 8294 12540
rect 8230 12480 8294 12484
rect 5396 12276 5460 12340
rect 9812 12276 9876 12340
rect 13492 12548 13556 12552
rect 15580 12540 15644 12544
rect 15580 12484 15584 12540
rect 15584 12484 15640 12540
rect 15640 12484 15644 12540
rect 15580 12480 15644 12484
rect 15660 12540 15724 12544
rect 15660 12484 15664 12540
rect 15664 12484 15720 12540
rect 15720 12484 15724 12540
rect 15660 12480 15724 12484
rect 15740 12540 15804 12544
rect 15740 12484 15744 12540
rect 15744 12484 15800 12540
rect 15800 12484 15804 12540
rect 15740 12480 15804 12484
rect 15820 12540 15884 12544
rect 15820 12484 15824 12540
rect 15824 12484 15880 12540
rect 15880 12484 15884 12540
rect 15820 12480 15884 12484
rect 23170 12540 23234 12544
rect 23170 12484 23174 12540
rect 23174 12484 23230 12540
rect 23230 12484 23234 12540
rect 23170 12480 23234 12484
rect 23250 12540 23314 12544
rect 23250 12484 23254 12540
rect 23254 12484 23310 12540
rect 23310 12484 23314 12540
rect 23250 12480 23314 12484
rect 23330 12540 23394 12544
rect 23330 12484 23334 12540
rect 23334 12484 23390 12540
rect 23390 12484 23394 12540
rect 23330 12480 23394 12484
rect 23410 12540 23474 12544
rect 23410 12484 23414 12540
rect 23414 12484 23470 12540
rect 23470 12484 23474 12540
rect 23410 12480 23474 12484
rect 30760 12540 30824 12544
rect 30760 12484 30764 12540
rect 30764 12484 30820 12540
rect 30820 12484 30824 12540
rect 30760 12480 30824 12484
rect 30840 12540 30904 12544
rect 30840 12484 30844 12540
rect 30844 12484 30900 12540
rect 30900 12484 30904 12540
rect 30840 12480 30904 12484
rect 30920 12540 30984 12544
rect 30920 12484 30924 12540
rect 30924 12484 30980 12540
rect 30980 12484 30984 12540
rect 30920 12480 30984 12484
rect 31000 12540 31064 12544
rect 31000 12484 31004 12540
rect 31004 12484 31060 12540
rect 31060 12484 31064 12540
rect 31000 12480 31064 12484
rect 10732 12140 10796 12204
rect 29132 12004 29196 12068
rect 4195 11996 4259 12000
rect 4195 11940 4199 11996
rect 4199 11940 4255 11996
rect 4255 11940 4259 11996
rect 4195 11936 4259 11940
rect 4275 11996 4339 12000
rect 4275 11940 4279 11996
rect 4279 11940 4335 11996
rect 4335 11940 4339 11996
rect 4275 11936 4339 11940
rect 4355 11996 4419 12000
rect 4355 11940 4359 11996
rect 4359 11940 4415 11996
rect 4415 11940 4419 11996
rect 4355 11936 4419 11940
rect 4435 11996 4499 12000
rect 4435 11940 4439 11996
rect 4439 11940 4495 11996
rect 4495 11940 4499 11996
rect 4435 11936 4499 11940
rect 11785 11996 11849 12000
rect 11785 11940 11789 11996
rect 11789 11940 11845 11996
rect 11845 11940 11849 11996
rect 11785 11936 11849 11940
rect 11865 11996 11929 12000
rect 11865 11940 11869 11996
rect 11869 11940 11925 11996
rect 11925 11940 11929 11996
rect 11865 11936 11929 11940
rect 11945 11996 12009 12000
rect 11945 11940 11949 11996
rect 11949 11940 12005 11996
rect 12005 11940 12009 11996
rect 11945 11936 12009 11940
rect 12025 11996 12089 12000
rect 12025 11940 12029 11996
rect 12029 11940 12085 11996
rect 12085 11940 12089 11996
rect 12025 11936 12089 11940
rect 19375 11996 19439 12000
rect 19375 11940 19379 11996
rect 19379 11940 19435 11996
rect 19435 11940 19439 11996
rect 19375 11936 19439 11940
rect 19455 11996 19519 12000
rect 19455 11940 19459 11996
rect 19459 11940 19515 11996
rect 19515 11940 19519 11996
rect 19455 11936 19519 11940
rect 19535 11996 19599 12000
rect 19535 11940 19539 11996
rect 19539 11940 19595 11996
rect 19595 11940 19599 11996
rect 19535 11936 19599 11940
rect 19615 11996 19679 12000
rect 19615 11940 19619 11996
rect 19619 11940 19675 11996
rect 19675 11940 19679 11996
rect 19615 11936 19679 11940
rect 26965 11996 27029 12000
rect 26965 11940 26969 11996
rect 26969 11940 27025 11996
rect 27025 11940 27029 11996
rect 26965 11936 27029 11940
rect 27045 11996 27109 12000
rect 27045 11940 27049 11996
rect 27049 11940 27105 11996
rect 27105 11940 27109 11996
rect 27045 11936 27109 11940
rect 27125 11996 27189 12000
rect 27125 11940 27129 11996
rect 27129 11940 27185 11996
rect 27185 11940 27189 11996
rect 27125 11936 27189 11940
rect 27205 11996 27269 12000
rect 27205 11940 27209 11996
rect 27209 11940 27265 11996
rect 27265 11940 27269 11996
rect 27205 11936 27269 11940
rect 14044 11732 14108 11796
rect 5396 11596 5460 11660
rect 10180 11596 10244 11660
rect 16068 11596 16132 11660
rect 7990 11452 8054 11456
rect 7990 11396 7994 11452
rect 7994 11396 8050 11452
rect 8050 11396 8054 11452
rect 7990 11392 8054 11396
rect 8070 11452 8134 11456
rect 8070 11396 8074 11452
rect 8074 11396 8130 11452
rect 8130 11396 8134 11452
rect 8070 11392 8134 11396
rect 8150 11452 8214 11456
rect 8150 11396 8154 11452
rect 8154 11396 8210 11452
rect 8210 11396 8214 11452
rect 8150 11392 8214 11396
rect 8230 11452 8294 11456
rect 8230 11396 8234 11452
rect 8234 11396 8290 11452
rect 8290 11396 8294 11452
rect 8230 11392 8294 11396
rect 15580 11452 15644 11456
rect 15580 11396 15584 11452
rect 15584 11396 15640 11452
rect 15640 11396 15644 11452
rect 15580 11392 15644 11396
rect 15660 11452 15724 11456
rect 15660 11396 15664 11452
rect 15664 11396 15720 11452
rect 15720 11396 15724 11452
rect 15660 11392 15724 11396
rect 15740 11452 15804 11456
rect 15740 11396 15744 11452
rect 15744 11396 15800 11452
rect 15800 11396 15804 11452
rect 15740 11392 15804 11396
rect 15820 11452 15884 11456
rect 15820 11396 15824 11452
rect 15824 11396 15880 11452
rect 15880 11396 15884 11452
rect 15820 11392 15884 11396
rect 23170 11452 23234 11456
rect 23170 11396 23174 11452
rect 23174 11396 23230 11452
rect 23230 11396 23234 11452
rect 23170 11392 23234 11396
rect 23250 11452 23314 11456
rect 23250 11396 23254 11452
rect 23254 11396 23310 11452
rect 23310 11396 23314 11452
rect 23250 11392 23314 11396
rect 23330 11452 23394 11456
rect 23330 11396 23334 11452
rect 23334 11396 23390 11452
rect 23390 11396 23394 11452
rect 23330 11392 23394 11396
rect 23410 11452 23474 11456
rect 23410 11396 23414 11452
rect 23414 11396 23470 11452
rect 23470 11396 23474 11452
rect 23410 11392 23474 11396
rect 30760 11452 30824 11456
rect 30760 11396 30764 11452
rect 30764 11396 30820 11452
rect 30820 11396 30824 11452
rect 30760 11392 30824 11396
rect 30840 11452 30904 11456
rect 30840 11396 30844 11452
rect 30844 11396 30900 11452
rect 30900 11396 30904 11452
rect 30840 11392 30904 11396
rect 30920 11452 30984 11456
rect 30920 11396 30924 11452
rect 30924 11396 30980 11452
rect 30980 11396 30984 11452
rect 30920 11392 30984 11396
rect 31000 11452 31064 11456
rect 31000 11396 31004 11452
rect 31004 11396 31060 11452
rect 31060 11396 31064 11452
rect 31000 11392 31064 11396
rect 6684 10916 6748 10980
rect 20668 11052 20732 11116
rect 9628 10916 9692 10980
rect 9812 10976 9876 10980
rect 9812 10920 9862 10976
rect 9862 10920 9876 10976
rect 9812 10916 9876 10920
rect 4195 10908 4259 10912
rect 4195 10852 4199 10908
rect 4199 10852 4255 10908
rect 4255 10852 4259 10908
rect 4195 10848 4259 10852
rect 4275 10908 4339 10912
rect 4275 10852 4279 10908
rect 4279 10852 4335 10908
rect 4335 10852 4339 10908
rect 4275 10848 4339 10852
rect 4355 10908 4419 10912
rect 4355 10852 4359 10908
rect 4359 10852 4415 10908
rect 4415 10852 4419 10908
rect 4355 10848 4419 10852
rect 4435 10908 4499 10912
rect 4435 10852 4439 10908
rect 4439 10852 4495 10908
rect 4495 10852 4499 10908
rect 4435 10848 4499 10852
rect 11785 10908 11849 10912
rect 11785 10852 11789 10908
rect 11789 10852 11845 10908
rect 11845 10852 11849 10908
rect 11785 10848 11849 10852
rect 11865 10908 11929 10912
rect 11865 10852 11869 10908
rect 11869 10852 11925 10908
rect 11925 10852 11929 10908
rect 11865 10848 11929 10852
rect 11945 10908 12009 10912
rect 11945 10852 11949 10908
rect 11949 10852 12005 10908
rect 12005 10852 12009 10908
rect 11945 10848 12009 10852
rect 12025 10908 12089 10912
rect 12025 10852 12029 10908
rect 12029 10852 12085 10908
rect 12085 10852 12089 10908
rect 12025 10848 12089 10852
rect 19375 10908 19439 10912
rect 19375 10852 19379 10908
rect 19379 10852 19435 10908
rect 19435 10852 19439 10908
rect 19375 10848 19439 10852
rect 19455 10908 19519 10912
rect 19455 10852 19459 10908
rect 19459 10852 19515 10908
rect 19515 10852 19519 10908
rect 19455 10848 19519 10852
rect 19535 10908 19599 10912
rect 19535 10852 19539 10908
rect 19539 10852 19595 10908
rect 19595 10852 19599 10908
rect 19535 10848 19599 10852
rect 19615 10908 19679 10912
rect 19615 10852 19619 10908
rect 19619 10852 19675 10908
rect 19675 10852 19679 10908
rect 19615 10848 19679 10852
rect 26965 10908 27029 10912
rect 26965 10852 26969 10908
rect 26969 10852 27025 10908
rect 27025 10852 27029 10908
rect 26965 10848 27029 10852
rect 27045 10908 27109 10912
rect 27045 10852 27049 10908
rect 27049 10852 27105 10908
rect 27105 10852 27109 10908
rect 27045 10848 27109 10852
rect 27125 10908 27189 10912
rect 27125 10852 27129 10908
rect 27129 10852 27185 10908
rect 27185 10852 27189 10908
rect 27125 10848 27189 10852
rect 27205 10908 27269 10912
rect 27205 10852 27209 10908
rect 27209 10852 27265 10908
rect 27265 10852 27269 10908
rect 27205 10848 27269 10852
rect 8892 10644 8956 10708
rect 7990 10364 8054 10368
rect 7990 10308 7994 10364
rect 7994 10308 8050 10364
rect 8050 10308 8054 10364
rect 7990 10304 8054 10308
rect 8070 10364 8134 10368
rect 8070 10308 8074 10364
rect 8074 10308 8130 10364
rect 8130 10308 8134 10364
rect 8070 10304 8134 10308
rect 8150 10364 8214 10368
rect 8150 10308 8154 10364
rect 8154 10308 8210 10364
rect 8210 10308 8214 10364
rect 8150 10304 8214 10308
rect 8230 10364 8294 10368
rect 8230 10308 8234 10364
rect 8234 10308 8290 10364
rect 8290 10308 8294 10364
rect 8230 10304 8294 10308
rect 15580 10364 15644 10368
rect 15580 10308 15584 10364
rect 15584 10308 15640 10364
rect 15640 10308 15644 10364
rect 15580 10304 15644 10308
rect 15660 10364 15724 10368
rect 15660 10308 15664 10364
rect 15664 10308 15720 10364
rect 15720 10308 15724 10364
rect 15660 10304 15724 10308
rect 15740 10364 15804 10368
rect 15740 10308 15744 10364
rect 15744 10308 15800 10364
rect 15800 10308 15804 10364
rect 15740 10304 15804 10308
rect 15820 10364 15884 10368
rect 15820 10308 15824 10364
rect 15824 10308 15880 10364
rect 15880 10308 15884 10364
rect 15820 10304 15884 10308
rect 23170 10364 23234 10368
rect 23170 10308 23174 10364
rect 23174 10308 23230 10364
rect 23230 10308 23234 10364
rect 23170 10304 23234 10308
rect 23250 10364 23314 10368
rect 23250 10308 23254 10364
rect 23254 10308 23310 10364
rect 23310 10308 23314 10364
rect 23250 10304 23314 10308
rect 23330 10364 23394 10368
rect 23330 10308 23334 10364
rect 23334 10308 23390 10364
rect 23390 10308 23394 10364
rect 23330 10304 23394 10308
rect 23410 10364 23474 10368
rect 23410 10308 23414 10364
rect 23414 10308 23470 10364
rect 23470 10308 23474 10364
rect 23410 10304 23474 10308
rect 30760 10364 30824 10368
rect 30760 10308 30764 10364
rect 30764 10308 30820 10364
rect 30820 10308 30824 10364
rect 30760 10304 30824 10308
rect 30840 10364 30904 10368
rect 30840 10308 30844 10364
rect 30844 10308 30900 10364
rect 30900 10308 30904 10364
rect 30840 10304 30904 10308
rect 30920 10364 30984 10368
rect 30920 10308 30924 10364
rect 30924 10308 30980 10364
rect 30980 10308 30984 10364
rect 30920 10304 30984 10308
rect 31000 10364 31064 10368
rect 31000 10308 31004 10364
rect 31004 10308 31060 10364
rect 31060 10308 31064 10364
rect 31000 10304 31064 10308
rect 19748 10100 19812 10164
rect 9260 9964 9324 10028
rect 4195 9820 4259 9824
rect 4195 9764 4199 9820
rect 4199 9764 4255 9820
rect 4255 9764 4259 9820
rect 4195 9760 4259 9764
rect 4275 9820 4339 9824
rect 4275 9764 4279 9820
rect 4279 9764 4335 9820
rect 4335 9764 4339 9820
rect 4275 9760 4339 9764
rect 4355 9820 4419 9824
rect 4355 9764 4359 9820
rect 4359 9764 4415 9820
rect 4415 9764 4419 9820
rect 4355 9760 4419 9764
rect 4435 9820 4499 9824
rect 4435 9764 4439 9820
rect 4439 9764 4495 9820
rect 4495 9764 4499 9820
rect 4435 9760 4499 9764
rect 11785 9820 11849 9824
rect 11785 9764 11789 9820
rect 11789 9764 11845 9820
rect 11845 9764 11849 9820
rect 11785 9760 11849 9764
rect 11865 9820 11929 9824
rect 11865 9764 11869 9820
rect 11869 9764 11925 9820
rect 11925 9764 11929 9820
rect 11865 9760 11929 9764
rect 11945 9820 12009 9824
rect 11945 9764 11949 9820
rect 11949 9764 12005 9820
rect 12005 9764 12009 9820
rect 11945 9760 12009 9764
rect 12025 9820 12089 9824
rect 12025 9764 12029 9820
rect 12029 9764 12085 9820
rect 12085 9764 12089 9820
rect 12025 9760 12089 9764
rect 19375 9820 19439 9824
rect 19375 9764 19379 9820
rect 19379 9764 19435 9820
rect 19435 9764 19439 9820
rect 19375 9760 19439 9764
rect 19455 9820 19519 9824
rect 19455 9764 19459 9820
rect 19459 9764 19515 9820
rect 19515 9764 19519 9820
rect 19455 9760 19519 9764
rect 19535 9820 19599 9824
rect 19535 9764 19539 9820
rect 19539 9764 19595 9820
rect 19595 9764 19599 9820
rect 19535 9760 19599 9764
rect 19615 9820 19679 9824
rect 19615 9764 19619 9820
rect 19619 9764 19675 9820
rect 19675 9764 19679 9820
rect 19615 9760 19679 9764
rect 26965 9820 27029 9824
rect 26965 9764 26969 9820
rect 26969 9764 27025 9820
rect 27025 9764 27029 9820
rect 26965 9760 27029 9764
rect 27045 9820 27109 9824
rect 27045 9764 27049 9820
rect 27049 9764 27105 9820
rect 27105 9764 27109 9820
rect 27045 9760 27109 9764
rect 27125 9820 27189 9824
rect 27125 9764 27129 9820
rect 27129 9764 27185 9820
rect 27185 9764 27189 9820
rect 27125 9760 27189 9764
rect 27205 9820 27269 9824
rect 27205 9764 27209 9820
rect 27209 9764 27265 9820
rect 27265 9764 27269 9820
rect 27205 9760 27269 9764
rect 5580 9692 5644 9756
rect 6868 9420 6932 9484
rect 7990 9276 8054 9280
rect 7990 9220 7994 9276
rect 7994 9220 8050 9276
rect 8050 9220 8054 9276
rect 7990 9216 8054 9220
rect 8070 9276 8134 9280
rect 8070 9220 8074 9276
rect 8074 9220 8130 9276
rect 8130 9220 8134 9276
rect 8070 9216 8134 9220
rect 8150 9276 8214 9280
rect 8150 9220 8154 9276
rect 8154 9220 8210 9276
rect 8210 9220 8214 9276
rect 8150 9216 8214 9220
rect 8230 9276 8294 9280
rect 8230 9220 8234 9276
rect 8234 9220 8290 9276
rect 8290 9220 8294 9276
rect 8230 9216 8294 9220
rect 15580 9276 15644 9280
rect 15580 9220 15584 9276
rect 15584 9220 15640 9276
rect 15640 9220 15644 9276
rect 15580 9216 15644 9220
rect 15660 9276 15724 9280
rect 15660 9220 15664 9276
rect 15664 9220 15720 9276
rect 15720 9220 15724 9276
rect 15660 9216 15724 9220
rect 15740 9276 15804 9280
rect 15740 9220 15744 9276
rect 15744 9220 15800 9276
rect 15800 9220 15804 9276
rect 15740 9216 15804 9220
rect 15820 9276 15884 9280
rect 15820 9220 15824 9276
rect 15824 9220 15880 9276
rect 15880 9220 15884 9276
rect 15820 9216 15884 9220
rect 23170 9276 23234 9280
rect 23170 9220 23174 9276
rect 23174 9220 23230 9276
rect 23230 9220 23234 9276
rect 23170 9216 23234 9220
rect 23250 9276 23314 9280
rect 23250 9220 23254 9276
rect 23254 9220 23310 9276
rect 23310 9220 23314 9276
rect 23250 9216 23314 9220
rect 23330 9276 23394 9280
rect 23330 9220 23334 9276
rect 23334 9220 23390 9276
rect 23390 9220 23394 9276
rect 23330 9216 23394 9220
rect 23410 9276 23474 9280
rect 23410 9220 23414 9276
rect 23414 9220 23470 9276
rect 23470 9220 23474 9276
rect 23410 9216 23474 9220
rect 30760 9276 30824 9280
rect 30760 9220 30764 9276
rect 30764 9220 30820 9276
rect 30820 9220 30824 9276
rect 30760 9216 30824 9220
rect 30840 9276 30904 9280
rect 30840 9220 30844 9276
rect 30844 9220 30900 9276
rect 30900 9220 30904 9276
rect 30840 9216 30904 9220
rect 30920 9276 30984 9280
rect 30920 9220 30924 9276
rect 30924 9220 30980 9276
rect 30980 9220 30984 9276
rect 30920 9216 30984 9220
rect 31000 9276 31064 9280
rect 31000 9220 31004 9276
rect 31004 9220 31060 9276
rect 31060 9220 31064 9276
rect 31000 9216 31064 9220
rect 14044 8876 14108 8940
rect 4195 8732 4259 8736
rect 4195 8676 4199 8732
rect 4199 8676 4255 8732
rect 4255 8676 4259 8732
rect 4195 8672 4259 8676
rect 4275 8732 4339 8736
rect 4275 8676 4279 8732
rect 4279 8676 4335 8732
rect 4335 8676 4339 8732
rect 4275 8672 4339 8676
rect 4355 8732 4419 8736
rect 4355 8676 4359 8732
rect 4359 8676 4415 8732
rect 4415 8676 4419 8732
rect 4355 8672 4419 8676
rect 4435 8732 4499 8736
rect 4435 8676 4439 8732
rect 4439 8676 4495 8732
rect 4495 8676 4499 8732
rect 4435 8672 4499 8676
rect 11785 8732 11849 8736
rect 11785 8676 11789 8732
rect 11789 8676 11845 8732
rect 11845 8676 11849 8732
rect 11785 8672 11849 8676
rect 11865 8732 11929 8736
rect 11865 8676 11869 8732
rect 11869 8676 11925 8732
rect 11925 8676 11929 8732
rect 11865 8672 11929 8676
rect 11945 8732 12009 8736
rect 11945 8676 11949 8732
rect 11949 8676 12005 8732
rect 12005 8676 12009 8732
rect 11945 8672 12009 8676
rect 12025 8732 12089 8736
rect 12025 8676 12029 8732
rect 12029 8676 12085 8732
rect 12085 8676 12089 8732
rect 12025 8672 12089 8676
rect 19375 8732 19439 8736
rect 19375 8676 19379 8732
rect 19379 8676 19435 8732
rect 19435 8676 19439 8732
rect 19375 8672 19439 8676
rect 19455 8732 19519 8736
rect 19455 8676 19459 8732
rect 19459 8676 19515 8732
rect 19515 8676 19519 8732
rect 19455 8672 19519 8676
rect 19535 8732 19599 8736
rect 19535 8676 19539 8732
rect 19539 8676 19595 8732
rect 19595 8676 19599 8732
rect 19535 8672 19599 8676
rect 19615 8732 19679 8736
rect 19615 8676 19619 8732
rect 19619 8676 19675 8732
rect 19675 8676 19679 8732
rect 19615 8672 19679 8676
rect 26965 8732 27029 8736
rect 26965 8676 26969 8732
rect 26969 8676 27025 8732
rect 27025 8676 27029 8732
rect 26965 8672 27029 8676
rect 27045 8732 27109 8736
rect 27045 8676 27049 8732
rect 27049 8676 27105 8732
rect 27105 8676 27109 8732
rect 27045 8672 27109 8676
rect 27125 8732 27189 8736
rect 27125 8676 27129 8732
rect 27129 8676 27185 8732
rect 27185 8676 27189 8732
rect 27125 8672 27189 8676
rect 27205 8732 27269 8736
rect 27205 8676 27209 8732
rect 27209 8676 27265 8732
rect 27265 8676 27269 8732
rect 27205 8672 27269 8676
rect 7990 8188 8054 8192
rect 7990 8132 7994 8188
rect 7994 8132 8050 8188
rect 8050 8132 8054 8188
rect 7990 8128 8054 8132
rect 8070 8188 8134 8192
rect 8070 8132 8074 8188
rect 8074 8132 8130 8188
rect 8130 8132 8134 8188
rect 8070 8128 8134 8132
rect 8150 8188 8214 8192
rect 8150 8132 8154 8188
rect 8154 8132 8210 8188
rect 8210 8132 8214 8188
rect 8150 8128 8214 8132
rect 8230 8188 8294 8192
rect 8230 8132 8234 8188
rect 8234 8132 8290 8188
rect 8290 8132 8294 8188
rect 8230 8128 8294 8132
rect 15580 8188 15644 8192
rect 15580 8132 15584 8188
rect 15584 8132 15640 8188
rect 15640 8132 15644 8188
rect 15580 8128 15644 8132
rect 15660 8188 15724 8192
rect 15660 8132 15664 8188
rect 15664 8132 15720 8188
rect 15720 8132 15724 8188
rect 15660 8128 15724 8132
rect 15740 8188 15804 8192
rect 15740 8132 15744 8188
rect 15744 8132 15800 8188
rect 15800 8132 15804 8188
rect 15740 8128 15804 8132
rect 15820 8188 15884 8192
rect 15820 8132 15824 8188
rect 15824 8132 15880 8188
rect 15880 8132 15884 8188
rect 15820 8128 15884 8132
rect 23170 8188 23234 8192
rect 23170 8132 23174 8188
rect 23174 8132 23230 8188
rect 23230 8132 23234 8188
rect 23170 8128 23234 8132
rect 23250 8188 23314 8192
rect 23250 8132 23254 8188
rect 23254 8132 23310 8188
rect 23310 8132 23314 8188
rect 23250 8128 23314 8132
rect 23330 8188 23394 8192
rect 23330 8132 23334 8188
rect 23334 8132 23390 8188
rect 23390 8132 23394 8188
rect 23330 8128 23394 8132
rect 23410 8188 23474 8192
rect 23410 8132 23414 8188
rect 23414 8132 23470 8188
rect 23470 8132 23474 8188
rect 23410 8128 23474 8132
rect 30760 8188 30824 8192
rect 30760 8132 30764 8188
rect 30764 8132 30820 8188
rect 30820 8132 30824 8188
rect 30760 8128 30824 8132
rect 30840 8188 30904 8192
rect 30840 8132 30844 8188
rect 30844 8132 30900 8188
rect 30900 8132 30904 8188
rect 30840 8128 30904 8132
rect 30920 8188 30984 8192
rect 30920 8132 30924 8188
rect 30924 8132 30980 8188
rect 30980 8132 30984 8188
rect 30920 8128 30984 8132
rect 31000 8188 31064 8192
rect 31000 8132 31004 8188
rect 31004 8132 31060 8188
rect 31060 8132 31064 8188
rect 31000 8128 31064 8132
rect 4195 7644 4259 7648
rect 4195 7588 4199 7644
rect 4199 7588 4255 7644
rect 4255 7588 4259 7644
rect 4195 7584 4259 7588
rect 4275 7644 4339 7648
rect 4275 7588 4279 7644
rect 4279 7588 4335 7644
rect 4335 7588 4339 7644
rect 4275 7584 4339 7588
rect 4355 7644 4419 7648
rect 4355 7588 4359 7644
rect 4359 7588 4415 7644
rect 4415 7588 4419 7644
rect 4355 7584 4419 7588
rect 4435 7644 4499 7648
rect 4435 7588 4439 7644
rect 4439 7588 4495 7644
rect 4495 7588 4499 7644
rect 4435 7584 4499 7588
rect 11785 7644 11849 7648
rect 11785 7588 11789 7644
rect 11789 7588 11845 7644
rect 11845 7588 11849 7644
rect 11785 7584 11849 7588
rect 11865 7644 11929 7648
rect 11865 7588 11869 7644
rect 11869 7588 11925 7644
rect 11925 7588 11929 7644
rect 11865 7584 11929 7588
rect 11945 7644 12009 7648
rect 11945 7588 11949 7644
rect 11949 7588 12005 7644
rect 12005 7588 12009 7644
rect 11945 7584 12009 7588
rect 12025 7644 12089 7648
rect 12025 7588 12029 7644
rect 12029 7588 12085 7644
rect 12085 7588 12089 7644
rect 12025 7584 12089 7588
rect 19375 7644 19439 7648
rect 19375 7588 19379 7644
rect 19379 7588 19435 7644
rect 19435 7588 19439 7644
rect 19375 7584 19439 7588
rect 19455 7644 19519 7648
rect 19455 7588 19459 7644
rect 19459 7588 19515 7644
rect 19515 7588 19519 7644
rect 19455 7584 19519 7588
rect 19535 7644 19599 7648
rect 19535 7588 19539 7644
rect 19539 7588 19595 7644
rect 19595 7588 19599 7644
rect 19535 7584 19599 7588
rect 19615 7644 19679 7648
rect 19615 7588 19619 7644
rect 19619 7588 19675 7644
rect 19675 7588 19679 7644
rect 19615 7584 19679 7588
rect 26965 7644 27029 7648
rect 26965 7588 26969 7644
rect 26969 7588 27025 7644
rect 27025 7588 27029 7644
rect 26965 7584 27029 7588
rect 27045 7644 27109 7648
rect 27045 7588 27049 7644
rect 27049 7588 27105 7644
rect 27105 7588 27109 7644
rect 27045 7584 27109 7588
rect 27125 7644 27189 7648
rect 27125 7588 27129 7644
rect 27129 7588 27185 7644
rect 27185 7588 27189 7644
rect 27125 7584 27189 7588
rect 27205 7644 27269 7648
rect 27205 7588 27209 7644
rect 27209 7588 27265 7644
rect 27265 7588 27269 7644
rect 27205 7584 27269 7588
rect 7990 7100 8054 7104
rect 7990 7044 7994 7100
rect 7994 7044 8050 7100
rect 8050 7044 8054 7100
rect 7990 7040 8054 7044
rect 8070 7100 8134 7104
rect 8070 7044 8074 7100
rect 8074 7044 8130 7100
rect 8130 7044 8134 7100
rect 8070 7040 8134 7044
rect 8150 7100 8214 7104
rect 8150 7044 8154 7100
rect 8154 7044 8210 7100
rect 8210 7044 8214 7100
rect 8150 7040 8214 7044
rect 8230 7100 8294 7104
rect 8230 7044 8234 7100
rect 8234 7044 8290 7100
rect 8290 7044 8294 7100
rect 8230 7040 8294 7044
rect 15580 7100 15644 7104
rect 15580 7044 15584 7100
rect 15584 7044 15640 7100
rect 15640 7044 15644 7100
rect 15580 7040 15644 7044
rect 15660 7100 15724 7104
rect 15660 7044 15664 7100
rect 15664 7044 15720 7100
rect 15720 7044 15724 7100
rect 15660 7040 15724 7044
rect 15740 7100 15804 7104
rect 15740 7044 15744 7100
rect 15744 7044 15800 7100
rect 15800 7044 15804 7100
rect 15740 7040 15804 7044
rect 15820 7100 15884 7104
rect 15820 7044 15824 7100
rect 15824 7044 15880 7100
rect 15880 7044 15884 7100
rect 15820 7040 15884 7044
rect 23170 7100 23234 7104
rect 23170 7044 23174 7100
rect 23174 7044 23230 7100
rect 23230 7044 23234 7100
rect 23170 7040 23234 7044
rect 23250 7100 23314 7104
rect 23250 7044 23254 7100
rect 23254 7044 23310 7100
rect 23310 7044 23314 7100
rect 23250 7040 23314 7044
rect 23330 7100 23394 7104
rect 23330 7044 23334 7100
rect 23334 7044 23390 7100
rect 23390 7044 23394 7100
rect 23330 7040 23394 7044
rect 23410 7100 23474 7104
rect 23410 7044 23414 7100
rect 23414 7044 23470 7100
rect 23470 7044 23474 7100
rect 23410 7040 23474 7044
rect 30760 7100 30824 7104
rect 30760 7044 30764 7100
rect 30764 7044 30820 7100
rect 30820 7044 30824 7100
rect 30760 7040 30824 7044
rect 30840 7100 30904 7104
rect 30840 7044 30844 7100
rect 30844 7044 30900 7100
rect 30900 7044 30904 7100
rect 30840 7040 30904 7044
rect 30920 7100 30984 7104
rect 30920 7044 30924 7100
rect 30924 7044 30980 7100
rect 30980 7044 30984 7100
rect 30920 7040 30984 7044
rect 31000 7100 31064 7104
rect 31000 7044 31004 7100
rect 31004 7044 31060 7100
rect 31060 7044 31064 7100
rect 31000 7040 31064 7044
rect 2820 6896 2884 6900
rect 2820 6840 2834 6896
rect 2834 6840 2884 6896
rect 2820 6836 2884 6840
rect 28580 6836 28644 6900
rect 4195 6556 4259 6560
rect 4195 6500 4199 6556
rect 4199 6500 4255 6556
rect 4255 6500 4259 6556
rect 4195 6496 4259 6500
rect 4275 6556 4339 6560
rect 4275 6500 4279 6556
rect 4279 6500 4335 6556
rect 4335 6500 4339 6556
rect 4275 6496 4339 6500
rect 4355 6556 4419 6560
rect 4355 6500 4359 6556
rect 4359 6500 4415 6556
rect 4415 6500 4419 6556
rect 4355 6496 4419 6500
rect 4435 6556 4499 6560
rect 4435 6500 4439 6556
rect 4439 6500 4495 6556
rect 4495 6500 4499 6556
rect 4435 6496 4499 6500
rect 11785 6556 11849 6560
rect 11785 6500 11789 6556
rect 11789 6500 11845 6556
rect 11845 6500 11849 6556
rect 11785 6496 11849 6500
rect 11865 6556 11929 6560
rect 11865 6500 11869 6556
rect 11869 6500 11925 6556
rect 11925 6500 11929 6556
rect 11865 6496 11929 6500
rect 11945 6556 12009 6560
rect 11945 6500 11949 6556
rect 11949 6500 12005 6556
rect 12005 6500 12009 6556
rect 11945 6496 12009 6500
rect 12025 6556 12089 6560
rect 12025 6500 12029 6556
rect 12029 6500 12085 6556
rect 12085 6500 12089 6556
rect 12025 6496 12089 6500
rect 19375 6556 19439 6560
rect 19375 6500 19379 6556
rect 19379 6500 19435 6556
rect 19435 6500 19439 6556
rect 19375 6496 19439 6500
rect 19455 6556 19519 6560
rect 19455 6500 19459 6556
rect 19459 6500 19515 6556
rect 19515 6500 19519 6556
rect 19455 6496 19519 6500
rect 19535 6556 19599 6560
rect 19535 6500 19539 6556
rect 19539 6500 19595 6556
rect 19595 6500 19599 6556
rect 19535 6496 19599 6500
rect 19615 6556 19679 6560
rect 19615 6500 19619 6556
rect 19619 6500 19675 6556
rect 19675 6500 19679 6556
rect 19615 6496 19679 6500
rect 26965 6556 27029 6560
rect 26965 6500 26969 6556
rect 26969 6500 27025 6556
rect 27025 6500 27029 6556
rect 26965 6496 27029 6500
rect 27045 6556 27109 6560
rect 27045 6500 27049 6556
rect 27049 6500 27105 6556
rect 27105 6500 27109 6556
rect 27045 6496 27109 6500
rect 27125 6556 27189 6560
rect 27125 6500 27129 6556
rect 27129 6500 27185 6556
rect 27185 6500 27189 6556
rect 27125 6496 27189 6500
rect 27205 6556 27269 6560
rect 27205 6500 27209 6556
rect 27209 6500 27265 6556
rect 27265 6500 27269 6556
rect 27205 6496 27269 6500
rect 6868 6428 6932 6492
rect 7990 6012 8054 6016
rect 7990 5956 7994 6012
rect 7994 5956 8050 6012
rect 8050 5956 8054 6012
rect 7990 5952 8054 5956
rect 8070 6012 8134 6016
rect 8070 5956 8074 6012
rect 8074 5956 8130 6012
rect 8130 5956 8134 6012
rect 8070 5952 8134 5956
rect 8150 6012 8214 6016
rect 8150 5956 8154 6012
rect 8154 5956 8210 6012
rect 8210 5956 8214 6012
rect 8150 5952 8214 5956
rect 8230 6012 8294 6016
rect 8230 5956 8234 6012
rect 8234 5956 8290 6012
rect 8290 5956 8294 6012
rect 8230 5952 8294 5956
rect 15580 6012 15644 6016
rect 15580 5956 15584 6012
rect 15584 5956 15640 6012
rect 15640 5956 15644 6012
rect 15580 5952 15644 5956
rect 15660 6012 15724 6016
rect 15660 5956 15664 6012
rect 15664 5956 15720 6012
rect 15720 5956 15724 6012
rect 15660 5952 15724 5956
rect 15740 6012 15804 6016
rect 15740 5956 15744 6012
rect 15744 5956 15800 6012
rect 15800 5956 15804 6012
rect 15740 5952 15804 5956
rect 15820 6012 15884 6016
rect 15820 5956 15824 6012
rect 15824 5956 15880 6012
rect 15880 5956 15884 6012
rect 15820 5952 15884 5956
rect 23170 6012 23234 6016
rect 23170 5956 23174 6012
rect 23174 5956 23230 6012
rect 23230 5956 23234 6012
rect 23170 5952 23234 5956
rect 23250 6012 23314 6016
rect 23250 5956 23254 6012
rect 23254 5956 23310 6012
rect 23310 5956 23314 6012
rect 23250 5952 23314 5956
rect 23330 6012 23394 6016
rect 23330 5956 23334 6012
rect 23334 5956 23390 6012
rect 23390 5956 23394 6012
rect 23330 5952 23394 5956
rect 23410 6012 23474 6016
rect 23410 5956 23414 6012
rect 23414 5956 23470 6012
rect 23470 5956 23474 6012
rect 23410 5952 23474 5956
rect 30760 6012 30824 6016
rect 30760 5956 30764 6012
rect 30764 5956 30820 6012
rect 30820 5956 30824 6012
rect 30760 5952 30824 5956
rect 30840 6012 30904 6016
rect 30840 5956 30844 6012
rect 30844 5956 30900 6012
rect 30900 5956 30904 6012
rect 30840 5952 30904 5956
rect 30920 6012 30984 6016
rect 30920 5956 30924 6012
rect 30924 5956 30980 6012
rect 30980 5956 30984 6012
rect 30920 5952 30984 5956
rect 31000 6012 31064 6016
rect 31000 5956 31004 6012
rect 31004 5956 31060 6012
rect 31060 5956 31064 6012
rect 31000 5952 31064 5956
rect 4195 5468 4259 5472
rect 4195 5412 4199 5468
rect 4199 5412 4255 5468
rect 4255 5412 4259 5468
rect 4195 5408 4259 5412
rect 4275 5468 4339 5472
rect 4275 5412 4279 5468
rect 4279 5412 4335 5468
rect 4335 5412 4339 5468
rect 4275 5408 4339 5412
rect 4355 5468 4419 5472
rect 4355 5412 4359 5468
rect 4359 5412 4415 5468
rect 4415 5412 4419 5468
rect 4355 5408 4419 5412
rect 4435 5468 4499 5472
rect 4435 5412 4439 5468
rect 4439 5412 4495 5468
rect 4495 5412 4499 5468
rect 4435 5408 4499 5412
rect 11785 5468 11849 5472
rect 11785 5412 11789 5468
rect 11789 5412 11845 5468
rect 11845 5412 11849 5468
rect 11785 5408 11849 5412
rect 11865 5468 11929 5472
rect 11865 5412 11869 5468
rect 11869 5412 11925 5468
rect 11925 5412 11929 5468
rect 11865 5408 11929 5412
rect 11945 5468 12009 5472
rect 11945 5412 11949 5468
rect 11949 5412 12005 5468
rect 12005 5412 12009 5468
rect 11945 5408 12009 5412
rect 12025 5468 12089 5472
rect 12025 5412 12029 5468
rect 12029 5412 12085 5468
rect 12085 5412 12089 5468
rect 12025 5408 12089 5412
rect 19375 5468 19439 5472
rect 19375 5412 19379 5468
rect 19379 5412 19435 5468
rect 19435 5412 19439 5468
rect 19375 5408 19439 5412
rect 19455 5468 19519 5472
rect 19455 5412 19459 5468
rect 19459 5412 19515 5468
rect 19515 5412 19519 5468
rect 19455 5408 19519 5412
rect 19535 5468 19599 5472
rect 19535 5412 19539 5468
rect 19539 5412 19595 5468
rect 19595 5412 19599 5468
rect 19535 5408 19599 5412
rect 19615 5468 19679 5472
rect 19615 5412 19619 5468
rect 19619 5412 19675 5468
rect 19675 5412 19679 5468
rect 19615 5408 19679 5412
rect 26965 5468 27029 5472
rect 26965 5412 26969 5468
rect 26969 5412 27025 5468
rect 27025 5412 27029 5468
rect 26965 5408 27029 5412
rect 27045 5468 27109 5472
rect 27045 5412 27049 5468
rect 27049 5412 27105 5468
rect 27105 5412 27109 5468
rect 27045 5408 27109 5412
rect 27125 5468 27189 5472
rect 27125 5412 27129 5468
rect 27129 5412 27185 5468
rect 27185 5412 27189 5468
rect 27125 5408 27189 5412
rect 27205 5468 27269 5472
rect 27205 5412 27209 5468
rect 27209 5412 27265 5468
rect 27265 5412 27269 5468
rect 27205 5408 27269 5412
rect 7990 4924 8054 4928
rect 7990 4868 7994 4924
rect 7994 4868 8050 4924
rect 8050 4868 8054 4924
rect 7990 4864 8054 4868
rect 8070 4924 8134 4928
rect 8070 4868 8074 4924
rect 8074 4868 8130 4924
rect 8130 4868 8134 4924
rect 8070 4864 8134 4868
rect 8150 4924 8214 4928
rect 8150 4868 8154 4924
rect 8154 4868 8210 4924
rect 8210 4868 8214 4924
rect 8150 4864 8214 4868
rect 8230 4924 8294 4928
rect 8230 4868 8234 4924
rect 8234 4868 8290 4924
rect 8290 4868 8294 4924
rect 8230 4864 8294 4868
rect 15580 4924 15644 4928
rect 15580 4868 15584 4924
rect 15584 4868 15640 4924
rect 15640 4868 15644 4924
rect 15580 4864 15644 4868
rect 15660 4924 15724 4928
rect 15660 4868 15664 4924
rect 15664 4868 15720 4924
rect 15720 4868 15724 4924
rect 15660 4864 15724 4868
rect 15740 4924 15804 4928
rect 15740 4868 15744 4924
rect 15744 4868 15800 4924
rect 15800 4868 15804 4924
rect 15740 4864 15804 4868
rect 15820 4924 15884 4928
rect 15820 4868 15824 4924
rect 15824 4868 15880 4924
rect 15880 4868 15884 4924
rect 15820 4864 15884 4868
rect 23170 4924 23234 4928
rect 23170 4868 23174 4924
rect 23174 4868 23230 4924
rect 23230 4868 23234 4924
rect 23170 4864 23234 4868
rect 23250 4924 23314 4928
rect 23250 4868 23254 4924
rect 23254 4868 23310 4924
rect 23310 4868 23314 4924
rect 23250 4864 23314 4868
rect 23330 4924 23394 4928
rect 23330 4868 23334 4924
rect 23334 4868 23390 4924
rect 23390 4868 23394 4924
rect 23330 4864 23394 4868
rect 23410 4924 23474 4928
rect 23410 4868 23414 4924
rect 23414 4868 23470 4924
rect 23470 4868 23474 4924
rect 23410 4864 23474 4868
rect 30760 4924 30824 4928
rect 30760 4868 30764 4924
rect 30764 4868 30820 4924
rect 30820 4868 30824 4924
rect 30760 4864 30824 4868
rect 30840 4924 30904 4928
rect 30840 4868 30844 4924
rect 30844 4868 30900 4924
rect 30900 4868 30904 4924
rect 30840 4864 30904 4868
rect 30920 4924 30984 4928
rect 30920 4868 30924 4924
rect 30924 4868 30980 4924
rect 30980 4868 30984 4924
rect 30920 4864 30984 4868
rect 31000 4924 31064 4928
rect 31000 4868 31004 4924
rect 31004 4868 31060 4924
rect 31060 4868 31064 4924
rect 31000 4864 31064 4868
rect 4195 4380 4259 4384
rect 4195 4324 4199 4380
rect 4199 4324 4255 4380
rect 4255 4324 4259 4380
rect 4195 4320 4259 4324
rect 4275 4380 4339 4384
rect 4275 4324 4279 4380
rect 4279 4324 4335 4380
rect 4335 4324 4339 4380
rect 4275 4320 4339 4324
rect 4355 4380 4419 4384
rect 4355 4324 4359 4380
rect 4359 4324 4415 4380
rect 4415 4324 4419 4380
rect 4355 4320 4419 4324
rect 4435 4380 4499 4384
rect 4435 4324 4439 4380
rect 4439 4324 4495 4380
rect 4495 4324 4499 4380
rect 4435 4320 4499 4324
rect 11785 4380 11849 4384
rect 11785 4324 11789 4380
rect 11789 4324 11845 4380
rect 11845 4324 11849 4380
rect 11785 4320 11849 4324
rect 11865 4380 11929 4384
rect 11865 4324 11869 4380
rect 11869 4324 11925 4380
rect 11925 4324 11929 4380
rect 11865 4320 11929 4324
rect 11945 4380 12009 4384
rect 11945 4324 11949 4380
rect 11949 4324 12005 4380
rect 12005 4324 12009 4380
rect 11945 4320 12009 4324
rect 12025 4380 12089 4384
rect 12025 4324 12029 4380
rect 12029 4324 12085 4380
rect 12085 4324 12089 4380
rect 12025 4320 12089 4324
rect 19375 4380 19439 4384
rect 19375 4324 19379 4380
rect 19379 4324 19435 4380
rect 19435 4324 19439 4380
rect 19375 4320 19439 4324
rect 19455 4380 19519 4384
rect 19455 4324 19459 4380
rect 19459 4324 19515 4380
rect 19515 4324 19519 4380
rect 19455 4320 19519 4324
rect 19535 4380 19599 4384
rect 19535 4324 19539 4380
rect 19539 4324 19595 4380
rect 19595 4324 19599 4380
rect 19535 4320 19599 4324
rect 19615 4380 19679 4384
rect 19615 4324 19619 4380
rect 19619 4324 19675 4380
rect 19675 4324 19679 4380
rect 19615 4320 19679 4324
rect 26965 4380 27029 4384
rect 26965 4324 26969 4380
rect 26969 4324 27025 4380
rect 27025 4324 27029 4380
rect 26965 4320 27029 4324
rect 27045 4380 27109 4384
rect 27045 4324 27049 4380
rect 27049 4324 27105 4380
rect 27105 4324 27109 4380
rect 27045 4320 27109 4324
rect 27125 4380 27189 4384
rect 27125 4324 27129 4380
rect 27129 4324 27185 4380
rect 27185 4324 27189 4380
rect 27125 4320 27189 4324
rect 27205 4380 27269 4384
rect 27205 4324 27209 4380
rect 27209 4324 27265 4380
rect 27265 4324 27269 4380
rect 27205 4320 27269 4324
rect 3004 4040 3068 4044
rect 3004 3984 3018 4040
rect 3018 3984 3068 4040
rect 3004 3980 3068 3984
rect 7990 3836 8054 3840
rect 7990 3780 7994 3836
rect 7994 3780 8050 3836
rect 8050 3780 8054 3836
rect 7990 3776 8054 3780
rect 8070 3836 8134 3840
rect 8070 3780 8074 3836
rect 8074 3780 8130 3836
rect 8130 3780 8134 3836
rect 8070 3776 8134 3780
rect 8150 3836 8214 3840
rect 8150 3780 8154 3836
rect 8154 3780 8210 3836
rect 8210 3780 8214 3836
rect 8150 3776 8214 3780
rect 8230 3836 8294 3840
rect 8230 3780 8234 3836
rect 8234 3780 8290 3836
rect 8290 3780 8294 3836
rect 8230 3776 8294 3780
rect 15580 3836 15644 3840
rect 15580 3780 15584 3836
rect 15584 3780 15640 3836
rect 15640 3780 15644 3836
rect 15580 3776 15644 3780
rect 15660 3836 15724 3840
rect 15660 3780 15664 3836
rect 15664 3780 15720 3836
rect 15720 3780 15724 3836
rect 15660 3776 15724 3780
rect 15740 3836 15804 3840
rect 15740 3780 15744 3836
rect 15744 3780 15800 3836
rect 15800 3780 15804 3836
rect 15740 3776 15804 3780
rect 15820 3836 15884 3840
rect 15820 3780 15824 3836
rect 15824 3780 15880 3836
rect 15880 3780 15884 3836
rect 15820 3776 15884 3780
rect 23170 3836 23234 3840
rect 23170 3780 23174 3836
rect 23174 3780 23230 3836
rect 23230 3780 23234 3836
rect 23170 3776 23234 3780
rect 23250 3836 23314 3840
rect 23250 3780 23254 3836
rect 23254 3780 23310 3836
rect 23310 3780 23314 3836
rect 23250 3776 23314 3780
rect 23330 3836 23394 3840
rect 23330 3780 23334 3836
rect 23334 3780 23390 3836
rect 23390 3780 23394 3836
rect 23330 3776 23394 3780
rect 23410 3836 23474 3840
rect 23410 3780 23414 3836
rect 23414 3780 23470 3836
rect 23470 3780 23474 3836
rect 23410 3776 23474 3780
rect 30760 3836 30824 3840
rect 30760 3780 30764 3836
rect 30764 3780 30820 3836
rect 30820 3780 30824 3836
rect 30760 3776 30824 3780
rect 30840 3836 30904 3840
rect 30840 3780 30844 3836
rect 30844 3780 30900 3836
rect 30900 3780 30904 3836
rect 30840 3776 30904 3780
rect 30920 3836 30984 3840
rect 30920 3780 30924 3836
rect 30924 3780 30980 3836
rect 30980 3780 30984 3836
rect 30920 3776 30984 3780
rect 31000 3836 31064 3840
rect 31000 3780 31004 3836
rect 31004 3780 31060 3836
rect 31060 3780 31064 3836
rect 31000 3776 31064 3780
rect 4195 3292 4259 3296
rect 4195 3236 4199 3292
rect 4199 3236 4255 3292
rect 4255 3236 4259 3292
rect 4195 3232 4259 3236
rect 4275 3292 4339 3296
rect 4275 3236 4279 3292
rect 4279 3236 4335 3292
rect 4335 3236 4339 3292
rect 4275 3232 4339 3236
rect 4355 3292 4419 3296
rect 4355 3236 4359 3292
rect 4359 3236 4415 3292
rect 4415 3236 4419 3292
rect 4355 3232 4419 3236
rect 4435 3292 4499 3296
rect 4435 3236 4439 3292
rect 4439 3236 4495 3292
rect 4495 3236 4499 3292
rect 4435 3232 4499 3236
rect 11785 3292 11849 3296
rect 11785 3236 11789 3292
rect 11789 3236 11845 3292
rect 11845 3236 11849 3292
rect 11785 3232 11849 3236
rect 11865 3292 11929 3296
rect 11865 3236 11869 3292
rect 11869 3236 11925 3292
rect 11925 3236 11929 3292
rect 11865 3232 11929 3236
rect 11945 3292 12009 3296
rect 11945 3236 11949 3292
rect 11949 3236 12005 3292
rect 12005 3236 12009 3292
rect 11945 3232 12009 3236
rect 12025 3292 12089 3296
rect 12025 3236 12029 3292
rect 12029 3236 12085 3292
rect 12085 3236 12089 3292
rect 12025 3232 12089 3236
rect 19375 3292 19439 3296
rect 19375 3236 19379 3292
rect 19379 3236 19435 3292
rect 19435 3236 19439 3292
rect 19375 3232 19439 3236
rect 19455 3292 19519 3296
rect 19455 3236 19459 3292
rect 19459 3236 19515 3292
rect 19515 3236 19519 3292
rect 19455 3232 19519 3236
rect 19535 3292 19599 3296
rect 19535 3236 19539 3292
rect 19539 3236 19595 3292
rect 19595 3236 19599 3292
rect 19535 3232 19599 3236
rect 19615 3292 19679 3296
rect 19615 3236 19619 3292
rect 19619 3236 19675 3292
rect 19675 3236 19679 3292
rect 19615 3232 19679 3236
rect 26965 3292 27029 3296
rect 26965 3236 26969 3292
rect 26969 3236 27025 3292
rect 27025 3236 27029 3292
rect 26965 3232 27029 3236
rect 27045 3292 27109 3296
rect 27045 3236 27049 3292
rect 27049 3236 27105 3292
rect 27105 3236 27109 3292
rect 27045 3232 27109 3236
rect 27125 3292 27189 3296
rect 27125 3236 27129 3292
rect 27129 3236 27185 3292
rect 27185 3236 27189 3292
rect 27125 3232 27189 3236
rect 27205 3292 27269 3296
rect 27205 3236 27209 3292
rect 27209 3236 27265 3292
rect 27265 3236 27269 3292
rect 27205 3232 27269 3236
rect 7990 2748 8054 2752
rect 7990 2692 7994 2748
rect 7994 2692 8050 2748
rect 8050 2692 8054 2748
rect 7990 2688 8054 2692
rect 8070 2748 8134 2752
rect 8070 2692 8074 2748
rect 8074 2692 8130 2748
rect 8130 2692 8134 2748
rect 8070 2688 8134 2692
rect 8150 2748 8214 2752
rect 8150 2692 8154 2748
rect 8154 2692 8210 2748
rect 8210 2692 8214 2748
rect 8150 2688 8214 2692
rect 8230 2748 8294 2752
rect 8230 2692 8234 2748
rect 8234 2692 8290 2748
rect 8290 2692 8294 2748
rect 8230 2688 8294 2692
rect 15580 2748 15644 2752
rect 15580 2692 15584 2748
rect 15584 2692 15640 2748
rect 15640 2692 15644 2748
rect 15580 2688 15644 2692
rect 15660 2748 15724 2752
rect 15660 2692 15664 2748
rect 15664 2692 15720 2748
rect 15720 2692 15724 2748
rect 15660 2688 15724 2692
rect 15740 2748 15804 2752
rect 15740 2692 15744 2748
rect 15744 2692 15800 2748
rect 15800 2692 15804 2748
rect 15740 2688 15804 2692
rect 15820 2748 15884 2752
rect 15820 2692 15824 2748
rect 15824 2692 15880 2748
rect 15880 2692 15884 2748
rect 15820 2688 15884 2692
rect 23170 2748 23234 2752
rect 23170 2692 23174 2748
rect 23174 2692 23230 2748
rect 23230 2692 23234 2748
rect 23170 2688 23234 2692
rect 23250 2748 23314 2752
rect 23250 2692 23254 2748
rect 23254 2692 23310 2748
rect 23310 2692 23314 2748
rect 23250 2688 23314 2692
rect 23330 2748 23394 2752
rect 23330 2692 23334 2748
rect 23334 2692 23390 2748
rect 23390 2692 23394 2748
rect 23330 2688 23394 2692
rect 23410 2748 23474 2752
rect 23410 2692 23414 2748
rect 23414 2692 23470 2748
rect 23470 2692 23474 2748
rect 23410 2688 23474 2692
rect 30760 2748 30824 2752
rect 30760 2692 30764 2748
rect 30764 2692 30820 2748
rect 30820 2692 30824 2748
rect 30760 2688 30824 2692
rect 30840 2748 30904 2752
rect 30840 2692 30844 2748
rect 30844 2692 30900 2748
rect 30900 2692 30904 2748
rect 30840 2688 30904 2692
rect 30920 2748 30984 2752
rect 30920 2692 30924 2748
rect 30924 2692 30980 2748
rect 30980 2692 30984 2748
rect 30920 2688 30984 2692
rect 31000 2748 31064 2752
rect 31000 2692 31004 2748
rect 31004 2692 31060 2748
rect 31060 2692 31064 2748
rect 31000 2688 31064 2692
rect 5580 2680 5644 2684
rect 5580 2624 5594 2680
rect 5594 2624 5644 2680
rect 5580 2620 5644 2624
rect 6684 2680 6748 2684
rect 6684 2624 6698 2680
rect 6698 2624 6748 2680
rect 6684 2620 6748 2624
rect 4195 2204 4259 2208
rect 4195 2148 4199 2204
rect 4199 2148 4255 2204
rect 4255 2148 4259 2204
rect 4195 2144 4259 2148
rect 4275 2204 4339 2208
rect 4275 2148 4279 2204
rect 4279 2148 4335 2204
rect 4335 2148 4339 2204
rect 4275 2144 4339 2148
rect 4355 2204 4419 2208
rect 4355 2148 4359 2204
rect 4359 2148 4415 2204
rect 4415 2148 4419 2204
rect 4355 2144 4419 2148
rect 4435 2204 4499 2208
rect 4435 2148 4439 2204
rect 4439 2148 4495 2204
rect 4495 2148 4499 2204
rect 4435 2144 4499 2148
rect 11785 2204 11849 2208
rect 11785 2148 11789 2204
rect 11789 2148 11845 2204
rect 11845 2148 11849 2204
rect 11785 2144 11849 2148
rect 11865 2204 11929 2208
rect 11865 2148 11869 2204
rect 11869 2148 11925 2204
rect 11925 2148 11929 2204
rect 11865 2144 11929 2148
rect 11945 2204 12009 2208
rect 11945 2148 11949 2204
rect 11949 2148 12005 2204
rect 12005 2148 12009 2204
rect 11945 2144 12009 2148
rect 12025 2204 12089 2208
rect 12025 2148 12029 2204
rect 12029 2148 12085 2204
rect 12085 2148 12089 2204
rect 12025 2144 12089 2148
rect 19375 2204 19439 2208
rect 19375 2148 19379 2204
rect 19379 2148 19435 2204
rect 19435 2148 19439 2204
rect 19375 2144 19439 2148
rect 19455 2204 19519 2208
rect 19455 2148 19459 2204
rect 19459 2148 19515 2204
rect 19515 2148 19519 2204
rect 19455 2144 19519 2148
rect 19535 2204 19599 2208
rect 19535 2148 19539 2204
rect 19539 2148 19595 2204
rect 19595 2148 19599 2204
rect 19535 2144 19599 2148
rect 19615 2204 19679 2208
rect 19615 2148 19619 2204
rect 19619 2148 19675 2204
rect 19675 2148 19679 2204
rect 19615 2144 19679 2148
rect 26965 2204 27029 2208
rect 26965 2148 26969 2204
rect 26969 2148 27025 2204
rect 27025 2148 27029 2204
rect 26965 2144 27029 2148
rect 27045 2204 27109 2208
rect 27045 2148 27049 2204
rect 27049 2148 27105 2204
rect 27105 2148 27109 2204
rect 27045 2144 27109 2148
rect 27125 2204 27189 2208
rect 27125 2148 27129 2204
rect 27129 2148 27185 2204
rect 27185 2148 27189 2204
rect 27125 2144 27189 2148
rect 27205 2204 27269 2208
rect 27205 2148 27209 2204
rect 27209 2148 27265 2204
rect 27265 2148 27269 2204
rect 27205 2144 27269 2148
rect 5396 1668 5460 1732
rect 7990 1660 8054 1664
rect 7990 1604 7994 1660
rect 7994 1604 8050 1660
rect 8050 1604 8054 1660
rect 7990 1600 8054 1604
rect 8070 1660 8134 1664
rect 8070 1604 8074 1660
rect 8074 1604 8130 1660
rect 8130 1604 8134 1660
rect 8070 1600 8134 1604
rect 8150 1660 8214 1664
rect 8150 1604 8154 1660
rect 8154 1604 8210 1660
rect 8210 1604 8214 1660
rect 8150 1600 8214 1604
rect 8230 1660 8294 1664
rect 8230 1604 8234 1660
rect 8234 1604 8290 1660
rect 8290 1604 8294 1660
rect 8230 1600 8294 1604
rect 15580 1660 15644 1664
rect 15580 1604 15584 1660
rect 15584 1604 15640 1660
rect 15640 1604 15644 1660
rect 15580 1600 15644 1604
rect 15660 1660 15724 1664
rect 15660 1604 15664 1660
rect 15664 1604 15720 1660
rect 15720 1604 15724 1660
rect 15660 1600 15724 1604
rect 15740 1660 15804 1664
rect 15740 1604 15744 1660
rect 15744 1604 15800 1660
rect 15800 1604 15804 1660
rect 15740 1600 15804 1604
rect 15820 1660 15884 1664
rect 15820 1604 15824 1660
rect 15824 1604 15880 1660
rect 15880 1604 15884 1660
rect 15820 1600 15884 1604
rect 23170 1660 23234 1664
rect 23170 1604 23174 1660
rect 23174 1604 23230 1660
rect 23230 1604 23234 1660
rect 23170 1600 23234 1604
rect 23250 1660 23314 1664
rect 23250 1604 23254 1660
rect 23254 1604 23310 1660
rect 23310 1604 23314 1660
rect 23250 1600 23314 1604
rect 23330 1660 23394 1664
rect 23330 1604 23334 1660
rect 23334 1604 23390 1660
rect 23390 1604 23394 1660
rect 23330 1600 23394 1604
rect 23410 1660 23474 1664
rect 23410 1604 23414 1660
rect 23414 1604 23470 1660
rect 23470 1604 23474 1660
rect 23410 1600 23474 1604
rect 30760 1660 30824 1664
rect 30760 1604 30764 1660
rect 30764 1604 30820 1660
rect 30820 1604 30824 1660
rect 30760 1600 30824 1604
rect 30840 1660 30904 1664
rect 30840 1604 30844 1660
rect 30844 1604 30900 1660
rect 30900 1604 30904 1660
rect 30840 1600 30904 1604
rect 30920 1660 30984 1664
rect 30920 1604 30924 1660
rect 30924 1604 30980 1660
rect 30980 1604 30984 1660
rect 30920 1600 30984 1604
rect 31000 1660 31064 1664
rect 31000 1604 31004 1660
rect 31004 1604 31060 1660
rect 31060 1604 31064 1660
rect 31000 1600 31064 1604
rect 4195 1116 4259 1120
rect 4195 1060 4199 1116
rect 4199 1060 4255 1116
rect 4255 1060 4259 1116
rect 4195 1056 4259 1060
rect 4275 1116 4339 1120
rect 4275 1060 4279 1116
rect 4279 1060 4335 1116
rect 4335 1060 4339 1116
rect 4275 1056 4339 1060
rect 4355 1116 4419 1120
rect 4355 1060 4359 1116
rect 4359 1060 4415 1116
rect 4415 1060 4419 1116
rect 4355 1056 4419 1060
rect 4435 1116 4499 1120
rect 4435 1060 4439 1116
rect 4439 1060 4495 1116
rect 4495 1060 4499 1116
rect 4435 1056 4499 1060
rect 11785 1116 11849 1120
rect 11785 1060 11789 1116
rect 11789 1060 11845 1116
rect 11845 1060 11849 1116
rect 11785 1056 11849 1060
rect 11865 1116 11929 1120
rect 11865 1060 11869 1116
rect 11869 1060 11925 1116
rect 11925 1060 11929 1116
rect 11865 1056 11929 1060
rect 11945 1116 12009 1120
rect 11945 1060 11949 1116
rect 11949 1060 12005 1116
rect 12005 1060 12009 1116
rect 11945 1056 12009 1060
rect 12025 1116 12089 1120
rect 12025 1060 12029 1116
rect 12029 1060 12085 1116
rect 12085 1060 12089 1116
rect 12025 1056 12089 1060
rect 19375 1116 19439 1120
rect 19375 1060 19379 1116
rect 19379 1060 19435 1116
rect 19435 1060 19439 1116
rect 19375 1056 19439 1060
rect 19455 1116 19519 1120
rect 19455 1060 19459 1116
rect 19459 1060 19515 1116
rect 19515 1060 19519 1116
rect 19455 1056 19519 1060
rect 19535 1116 19599 1120
rect 19535 1060 19539 1116
rect 19539 1060 19595 1116
rect 19595 1060 19599 1116
rect 19535 1056 19599 1060
rect 19615 1116 19679 1120
rect 19615 1060 19619 1116
rect 19619 1060 19675 1116
rect 19675 1060 19679 1116
rect 19615 1056 19679 1060
rect 26965 1116 27029 1120
rect 26965 1060 26969 1116
rect 26969 1060 27025 1116
rect 27025 1060 27029 1116
rect 26965 1056 27029 1060
rect 27045 1116 27109 1120
rect 27045 1060 27049 1116
rect 27049 1060 27105 1116
rect 27105 1060 27109 1116
rect 27045 1056 27109 1060
rect 27125 1116 27189 1120
rect 27125 1060 27129 1116
rect 27129 1060 27185 1116
rect 27185 1060 27189 1116
rect 27125 1056 27189 1060
rect 27205 1116 27269 1120
rect 27205 1060 27209 1116
rect 27209 1060 27265 1116
rect 27265 1060 27269 1116
rect 27205 1056 27269 1060
rect 7990 572 8054 576
rect 7990 516 7994 572
rect 7994 516 8050 572
rect 8050 516 8054 572
rect 7990 512 8054 516
rect 8070 572 8134 576
rect 8070 516 8074 572
rect 8074 516 8130 572
rect 8130 516 8134 572
rect 8070 512 8134 516
rect 8150 572 8214 576
rect 8150 516 8154 572
rect 8154 516 8210 572
rect 8210 516 8214 572
rect 8150 512 8214 516
rect 8230 572 8294 576
rect 8230 516 8234 572
rect 8234 516 8290 572
rect 8290 516 8294 572
rect 8230 512 8294 516
rect 15580 572 15644 576
rect 15580 516 15584 572
rect 15584 516 15640 572
rect 15640 516 15644 572
rect 15580 512 15644 516
rect 15660 572 15724 576
rect 15660 516 15664 572
rect 15664 516 15720 572
rect 15720 516 15724 572
rect 15660 512 15724 516
rect 15740 572 15804 576
rect 15740 516 15744 572
rect 15744 516 15800 572
rect 15800 516 15804 572
rect 15740 512 15804 516
rect 15820 572 15884 576
rect 15820 516 15824 572
rect 15824 516 15880 572
rect 15880 516 15884 572
rect 15820 512 15884 516
rect 23170 572 23234 576
rect 23170 516 23174 572
rect 23174 516 23230 572
rect 23230 516 23234 572
rect 23170 512 23234 516
rect 23250 572 23314 576
rect 23250 516 23254 572
rect 23254 516 23310 572
rect 23310 516 23314 572
rect 23250 512 23314 516
rect 23330 572 23394 576
rect 23330 516 23334 572
rect 23334 516 23390 572
rect 23390 516 23394 572
rect 23330 512 23394 516
rect 23410 572 23474 576
rect 23410 516 23414 572
rect 23414 516 23470 572
rect 23470 516 23474 572
rect 23410 512 23474 516
rect 30760 572 30824 576
rect 30760 516 30764 572
rect 30764 516 30820 572
rect 30820 516 30824 572
rect 30760 512 30824 516
rect 30840 572 30904 576
rect 30840 516 30844 572
rect 30844 516 30900 572
rect 30900 516 30904 572
rect 30840 512 30904 516
rect 30920 572 30984 576
rect 30920 516 30924 572
rect 30924 516 30980 572
rect 30980 516 30984 572
rect 30920 512 30984 516
rect 31000 572 31064 576
rect 31000 516 31004 572
rect 31004 516 31060 572
rect 31060 516 31064 572
rect 31000 512 31064 516
<< metal4 >>
rect 2819 22132 2885 22133
rect 2819 22068 2820 22132
rect 2884 22068 2885 22132
rect 4294 22130 4354 22304
rect 4478 22174 4722 22234
rect 4478 22130 4538 22174
rect 4294 22070 4538 22130
rect 2819 22067 2885 22068
rect 2822 6901 2882 22067
rect 4187 21792 4507 21808
rect 4187 21728 4195 21792
rect 4259 21728 4275 21792
rect 4339 21728 4355 21792
rect 4419 21728 4435 21792
rect 4499 21728 4507 21792
rect 4187 20704 4507 21728
rect 4187 20640 4195 20704
rect 4259 20640 4275 20704
rect 4339 20640 4355 20704
rect 4419 20640 4435 20704
rect 4499 20640 4507 20704
rect 4187 19616 4507 20640
rect 4187 19552 4195 19616
rect 4259 19552 4275 19616
rect 4339 19552 4355 19616
rect 4419 19552 4435 19616
rect 4499 19552 4507 19616
rect 4187 18528 4507 19552
rect 4662 19277 4722 22174
rect 4659 19276 4725 19277
rect 4659 19212 4660 19276
rect 4724 19212 4725 19276
rect 4659 19211 4725 19212
rect 4187 18464 4195 18528
rect 4259 18464 4275 18528
rect 4339 18464 4355 18528
rect 4419 18464 4435 18528
rect 4499 18464 4507 18528
rect 4187 17440 4507 18464
rect 4187 17376 4195 17440
rect 4259 17376 4275 17440
rect 4339 17376 4355 17440
rect 4419 17376 4435 17440
rect 4499 17376 4507 17440
rect 4187 16352 4507 17376
rect 4187 16288 4195 16352
rect 4259 16288 4275 16352
rect 4339 16288 4355 16352
rect 4419 16288 4435 16352
rect 4499 16288 4507 16352
rect 4187 15264 4507 16288
rect 4187 15200 4195 15264
rect 4259 15200 4275 15264
rect 4339 15200 4355 15264
rect 4419 15200 4435 15264
rect 4499 15200 4507 15264
rect 4187 14176 4507 15200
rect 4187 14112 4195 14176
rect 4259 14112 4275 14176
rect 4339 14112 4355 14176
rect 4419 14112 4435 14176
rect 4499 14112 4507 14176
rect 4187 13088 4507 14112
rect 4846 13701 4906 22304
rect 5398 18053 5458 22304
rect 5950 18461 6010 22304
rect 5947 18460 6013 18461
rect 5947 18396 5948 18460
rect 6012 18396 6013 18460
rect 5947 18395 6013 18396
rect 6502 18053 6562 22304
rect 7054 18053 7114 22304
rect 7606 18461 7666 22304
rect 7790 22174 8034 22234
rect 7790 19005 7850 22174
rect 7974 22130 8034 22174
rect 8158 22130 8218 22304
rect 7974 22070 8218 22130
rect 7982 21248 8302 21808
rect 7982 21184 7990 21248
rect 8054 21184 8070 21248
rect 8134 21184 8150 21248
rect 8214 21184 8230 21248
rect 8294 21184 8302 21248
rect 7982 20160 8302 21184
rect 7982 20096 7990 20160
rect 8054 20096 8070 20160
rect 8134 20096 8150 20160
rect 8214 20096 8230 20160
rect 8294 20096 8302 20160
rect 7982 19072 8302 20096
rect 8523 19412 8589 19413
rect 8523 19348 8524 19412
rect 8588 19348 8589 19412
rect 8523 19347 8589 19348
rect 7982 19008 7990 19072
rect 8054 19008 8070 19072
rect 8134 19008 8150 19072
rect 8214 19008 8230 19072
rect 8294 19008 8302 19072
rect 7787 19004 7853 19005
rect 7787 18940 7788 19004
rect 7852 18940 7853 19004
rect 7787 18939 7853 18940
rect 7419 18460 7485 18461
rect 7419 18396 7420 18460
rect 7484 18396 7485 18460
rect 7419 18395 7485 18396
rect 7603 18460 7669 18461
rect 7603 18396 7604 18460
rect 7668 18396 7669 18460
rect 7603 18395 7669 18396
rect 5211 18052 5277 18053
rect 5211 17988 5212 18052
rect 5276 17988 5277 18052
rect 5211 17987 5277 17988
rect 5395 18052 5461 18053
rect 5395 17988 5396 18052
rect 5460 17988 5461 18052
rect 5395 17987 5461 17988
rect 6499 18052 6565 18053
rect 6499 17988 6500 18052
rect 6564 17988 6565 18052
rect 6499 17987 6565 17988
rect 7051 18052 7117 18053
rect 7051 17988 7052 18052
rect 7116 17988 7117 18052
rect 7051 17987 7117 17988
rect 4843 13700 4909 13701
rect 4843 13636 4844 13700
rect 4908 13636 4909 13700
rect 4843 13635 4909 13636
rect 5214 13157 5274 17987
rect 7422 14789 7482 18395
rect 7982 17984 8302 19008
rect 7982 17920 7990 17984
rect 8054 17920 8070 17984
rect 8134 17920 8150 17984
rect 8214 17920 8230 17984
rect 8294 17920 8302 17984
rect 7982 16896 8302 17920
rect 7982 16832 7990 16896
rect 8054 16832 8070 16896
rect 8134 16832 8150 16896
rect 8214 16832 8230 16896
rect 8294 16832 8302 16896
rect 7982 15808 8302 16832
rect 8526 16690 8586 19347
rect 8710 16965 8770 22304
rect 8891 20772 8957 20773
rect 8891 20708 8892 20772
rect 8956 20708 8957 20772
rect 8891 20707 8957 20708
rect 8707 16964 8773 16965
rect 8707 16900 8708 16964
rect 8772 16900 8773 16964
rect 8707 16899 8773 16900
rect 8526 16630 8770 16690
rect 8523 16420 8589 16421
rect 8523 16356 8524 16420
rect 8588 16356 8589 16420
rect 8523 16355 8589 16356
rect 7982 15744 7990 15808
rect 8054 15744 8070 15808
rect 8134 15744 8150 15808
rect 8214 15744 8230 15808
rect 8294 15744 8302 15808
rect 7419 14788 7485 14789
rect 7419 14724 7420 14788
rect 7484 14724 7485 14788
rect 7419 14723 7485 14724
rect 7982 14720 8302 15744
rect 7982 14656 7990 14720
rect 8054 14656 8070 14720
rect 8134 14656 8150 14720
rect 8214 14656 8230 14720
rect 8294 14656 8302 14720
rect 7982 13632 8302 14656
rect 7982 13568 7990 13632
rect 8054 13568 8070 13632
rect 8134 13568 8150 13632
rect 8214 13568 8230 13632
rect 8294 13568 8302 13632
rect 5211 13156 5277 13157
rect 5211 13092 5212 13156
rect 5276 13092 5277 13156
rect 5211 13091 5277 13092
rect 4187 13024 4195 13088
rect 4259 13024 4275 13088
rect 4339 13024 4355 13088
rect 4419 13024 4435 13088
rect 4499 13024 4507 13088
rect 3003 12476 3069 12477
rect 3003 12412 3004 12476
rect 3068 12412 3069 12476
rect 3003 12411 3069 12412
rect 2819 6900 2885 6901
rect 2819 6836 2820 6900
rect 2884 6836 2885 6900
rect 2819 6835 2885 6836
rect 3006 4045 3066 12411
rect 4187 12000 4507 13024
rect 7982 12544 8302 13568
rect 8526 13565 8586 16355
rect 8523 13564 8589 13565
rect 8523 13500 8524 13564
rect 8588 13500 8589 13564
rect 8523 13499 8589 13500
rect 8710 12885 8770 16630
rect 8707 12884 8773 12885
rect 8707 12820 8708 12884
rect 8772 12820 8773 12884
rect 8707 12819 8773 12820
rect 7982 12480 7990 12544
rect 8054 12480 8070 12544
rect 8134 12480 8150 12544
rect 8214 12480 8230 12544
rect 8294 12480 8302 12544
rect 5395 12340 5461 12341
rect 5395 12276 5396 12340
rect 5460 12276 5461 12340
rect 5395 12275 5461 12276
rect 4187 11936 4195 12000
rect 4259 11936 4275 12000
rect 4339 11936 4355 12000
rect 4419 11936 4435 12000
rect 4499 11936 4507 12000
rect 4187 10912 4507 11936
rect 5398 11661 5458 12275
rect 5395 11660 5461 11661
rect 5395 11596 5396 11660
rect 5460 11596 5461 11660
rect 5395 11595 5461 11596
rect 4187 10848 4195 10912
rect 4259 10848 4275 10912
rect 4339 10848 4355 10912
rect 4419 10848 4435 10912
rect 4499 10848 4507 10912
rect 4187 9824 4507 10848
rect 4187 9760 4195 9824
rect 4259 9760 4275 9824
rect 4339 9760 4355 9824
rect 4419 9760 4435 9824
rect 4499 9760 4507 9824
rect 4187 8736 4507 9760
rect 4187 8672 4195 8736
rect 4259 8672 4275 8736
rect 4339 8672 4355 8736
rect 4419 8672 4435 8736
rect 4499 8672 4507 8736
rect 4187 7648 4507 8672
rect 4187 7584 4195 7648
rect 4259 7584 4275 7648
rect 4339 7584 4355 7648
rect 4419 7584 4435 7648
rect 4499 7584 4507 7648
rect 4187 6560 4507 7584
rect 4187 6496 4195 6560
rect 4259 6496 4275 6560
rect 4339 6496 4355 6560
rect 4419 6496 4435 6560
rect 4499 6496 4507 6560
rect 4187 5472 4507 6496
rect 4187 5408 4195 5472
rect 4259 5408 4275 5472
rect 4339 5408 4355 5472
rect 4419 5408 4435 5472
rect 4499 5408 4507 5472
rect 4187 4384 4507 5408
rect 4187 4320 4195 4384
rect 4259 4320 4275 4384
rect 4339 4320 4355 4384
rect 4419 4320 4435 4384
rect 4499 4320 4507 4384
rect 3003 4044 3069 4045
rect 3003 3980 3004 4044
rect 3068 3980 3069 4044
rect 3003 3979 3069 3980
rect 4187 3296 4507 4320
rect 4187 3232 4195 3296
rect 4259 3232 4275 3296
rect 4339 3232 4355 3296
rect 4419 3232 4435 3296
rect 4499 3232 4507 3296
rect 4187 2208 4507 3232
rect 4187 2144 4195 2208
rect 4259 2144 4275 2208
rect 4339 2144 4355 2208
rect 4419 2144 4435 2208
rect 4499 2144 4507 2208
rect 4187 1120 4507 2144
rect 5398 1733 5458 11595
rect 7982 11456 8302 12480
rect 7982 11392 7990 11456
rect 8054 11392 8070 11456
rect 8134 11392 8150 11456
rect 8214 11392 8230 11456
rect 8294 11392 8302 11456
rect 6683 10980 6749 10981
rect 6683 10916 6684 10980
rect 6748 10916 6749 10980
rect 6683 10915 6749 10916
rect 5579 9756 5645 9757
rect 5579 9692 5580 9756
rect 5644 9692 5645 9756
rect 5579 9691 5645 9692
rect 5582 2685 5642 9691
rect 6686 2685 6746 10915
rect 7982 10368 8302 11392
rect 8894 10709 8954 20707
rect 9262 19821 9322 22304
rect 9814 20770 9874 22304
rect 10179 21316 10245 21317
rect 10179 21252 10180 21316
rect 10244 21252 10245 21316
rect 10179 21251 10245 21252
rect 9630 20710 9874 20770
rect 9630 20637 9690 20710
rect 9627 20636 9693 20637
rect 9627 20572 9628 20636
rect 9692 20572 9693 20636
rect 9627 20571 9693 20572
rect 9443 20092 9509 20093
rect 9443 20028 9444 20092
rect 9508 20028 9509 20092
rect 9443 20027 9509 20028
rect 9259 19820 9325 19821
rect 9259 19756 9260 19820
rect 9324 19756 9325 19820
rect 9259 19755 9325 19756
rect 9259 19412 9325 19413
rect 9259 19348 9260 19412
rect 9324 19348 9325 19412
rect 9259 19347 9325 19348
rect 9262 19005 9322 19347
rect 9259 19004 9325 19005
rect 9259 18940 9260 19004
rect 9324 18940 9325 19004
rect 9259 18939 9325 18940
rect 9446 18730 9506 20027
rect 9627 19820 9693 19821
rect 9627 19756 9628 19820
rect 9692 19756 9693 19820
rect 9627 19755 9693 19756
rect 9078 18670 9506 18730
rect 9078 13021 9138 18670
rect 9443 18188 9509 18189
rect 9443 18124 9444 18188
rect 9508 18124 9509 18188
rect 9443 18123 9509 18124
rect 9446 16421 9506 18123
rect 9443 16420 9509 16421
rect 9443 16356 9444 16420
rect 9508 16356 9509 16420
rect 9443 16355 9509 16356
rect 9630 16010 9690 19755
rect 9262 15950 9690 16010
rect 9075 13020 9141 13021
rect 9075 12956 9076 13020
rect 9140 12956 9141 13020
rect 9075 12955 9141 12956
rect 8891 10708 8957 10709
rect 8891 10644 8892 10708
rect 8956 10644 8957 10708
rect 8891 10643 8957 10644
rect 7982 10304 7990 10368
rect 8054 10304 8070 10368
rect 8134 10304 8150 10368
rect 8214 10304 8230 10368
rect 8294 10304 8302 10368
rect 6867 9484 6933 9485
rect 6867 9420 6868 9484
rect 6932 9420 6933 9484
rect 6867 9419 6933 9420
rect 6870 6493 6930 9419
rect 7982 9280 8302 10304
rect 9262 10029 9322 15950
rect 9443 15468 9509 15469
rect 9443 15404 9444 15468
rect 9508 15404 9509 15468
rect 9443 15403 9509 15404
rect 9627 15468 9693 15469
rect 9627 15404 9628 15468
rect 9692 15404 9693 15468
rect 9627 15403 9693 15404
rect 9446 13021 9506 15403
rect 9443 13020 9509 13021
rect 9443 12956 9444 13020
rect 9508 12956 9509 13020
rect 9443 12955 9509 12956
rect 9630 10981 9690 15403
rect 9811 12340 9877 12341
rect 9811 12276 9812 12340
rect 9876 12276 9877 12340
rect 9811 12275 9877 12276
rect 9814 10981 9874 12275
rect 10182 11661 10242 21251
rect 10366 20637 10426 22304
rect 10918 21997 10978 22304
rect 10915 21996 10981 21997
rect 10915 21932 10916 21996
rect 10980 21932 10981 21996
rect 10915 21931 10981 21932
rect 10363 20636 10429 20637
rect 10363 20572 10364 20636
rect 10428 20572 10429 20636
rect 10363 20571 10429 20572
rect 11470 19141 11530 22304
rect 12022 21963 12082 22304
rect 12019 21962 12085 21963
rect 12019 21898 12020 21962
rect 12084 21898 12085 21962
rect 12019 21897 12085 21898
rect 11777 21792 12097 21808
rect 11777 21728 11785 21792
rect 11849 21728 11865 21792
rect 11929 21728 11945 21792
rect 12009 21728 12025 21792
rect 12089 21728 12097 21792
rect 11777 20704 12097 21728
rect 11777 20640 11785 20704
rect 11849 20640 11865 20704
rect 11929 20640 11945 20704
rect 12009 20640 12025 20704
rect 12089 20640 12097 20704
rect 11777 19616 12097 20640
rect 11777 19552 11785 19616
rect 11849 19552 11865 19616
rect 11929 19552 11945 19616
rect 12009 19552 12025 19616
rect 12089 19552 12097 19616
rect 11467 19140 11533 19141
rect 11467 19076 11468 19140
rect 11532 19076 11533 19140
rect 11467 19075 11533 19076
rect 11777 18528 12097 19552
rect 12203 19140 12269 19141
rect 12203 19076 12204 19140
rect 12268 19076 12269 19140
rect 12203 19075 12269 19076
rect 11777 18464 11785 18528
rect 11849 18464 11865 18528
rect 11929 18464 11945 18528
rect 12009 18464 12025 18528
rect 12089 18464 12097 18528
rect 11777 17440 12097 18464
rect 11777 17376 11785 17440
rect 11849 17376 11865 17440
rect 11929 17376 11945 17440
rect 12009 17376 12025 17440
rect 12089 17376 12097 17440
rect 10731 16692 10797 16693
rect 10731 16628 10732 16692
rect 10796 16628 10797 16692
rect 10731 16627 10797 16628
rect 10734 12205 10794 16627
rect 11777 16352 12097 17376
rect 11777 16288 11785 16352
rect 11849 16288 11865 16352
rect 11929 16288 11945 16352
rect 12009 16288 12025 16352
rect 12089 16288 12097 16352
rect 11777 15264 12097 16288
rect 11777 15200 11785 15264
rect 11849 15200 11865 15264
rect 11929 15200 11945 15264
rect 12009 15200 12025 15264
rect 12089 15200 12097 15264
rect 11777 14176 12097 15200
rect 11777 14112 11785 14176
rect 11849 14112 11865 14176
rect 11929 14112 11945 14176
rect 12009 14112 12025 14176
rect 12089 14112 12097 14176
rect 11777 13088 12097 14112
rect 11777 13024 11785 13088
rect 11849 13024 11865 13088
rect 11929 13024 11945 13088
rect 12009 13024 12025 13088
rect 12089 13024 12097 13088
rect 10731 12204 10797 12205
rect 10731 12140 10732 12204
rect 10796 12140 10797 12204
rect 10731 12139 10797 12140
rect 11777 12000 12097 13024
rect 12206 12613 12266 19075
rect 12574 18733 12634 22304
rect 13126 21963 13186 22304
rect 13123 21962 13189 21963
rect 13123 21898 13124 21962
rect 13188 21898 13189 21962
rect 13123 21897 13189 21898
rect 12571 18732 12637 18733
rect 12571 18668 12572 18732
rect 12636 18668 12637 18732
rect 12571 18667 12637 18668
rect 13678 18325 13738 22304
rect 14230 20637 14290 22304
rect 14411 22268 14477 22269
rect 14411 22204 14412 22268
rect 14476 22234 14477 22268
rect 14476 22204 14658 22234
rect 14411 22203 14658 22204
rect 14414 22174 14658 22203
rect 14598 22130 14658 22174
rect 14782 22130 14842 22304
rect 14598 22070 14842 22130
rect 14227 20636 14293 20637
rect 14227 20572 14228 20636
rect 14292 20572 14293 20636
rect 14227 20571 14293 20572
rect 14043 19412 14109 19413
rect 14043 19348 14044 19412
rect 14108 19348 14109 19412
rect 14043 19347 14109 19348
rect 13675 18324 13741 18325
rect 13675 18260 13676 18324
rect 13740 18260 13741 18324
rect 13675 18259 13741 18260
rect 12203 12612 12269 12613
rect 12203 12548 12204 12612
rect 12268 12548 12269 12612
rect 12203 12547 12269 12548
rect 13491 12612 13557 12613
rect 13491 12548 13492 12612
rect 13556 12548 13557 12612
rect 13491 12547 13557 12548
rect 11777 11936 11785 12000
rect 11849 11936 11865 12000
rect 11929 11936 11945 12000
rect 12009 11936 12025 12000
rect 12089 11936 12097 12000
rect 10179 11660 10245 11661
rect 10179 11596 10180 11660
rect 10244 11596 10245 11660
rect 10179 11595 10245 11596
rect 9627 10980 9693 10981
rect 9627 10916 9628 10980
rect 9692 10916 9693 10980
rect 9627 10915 9693 10916
rect 9811 10980 9877 10981
rect 9811 10916 9812 10980
rect 9876 10916 9877 10980
rect 9811 10915 9877 10916
rect 11777 10912 12097 11936
rect 13494 11250 13554 12547
rect 14046 11797 14106 19347
rect 15147 19276 15213 19277
rect 15147 19212 15148 19276
rect 15212 19212 15213 19276
rect 15147 19211 15213 19212
rect 15150 18053 15210 19211
rect 15334 19005 15394 22304
rect 15886 21960 15946 22304
rect 15886 21900 16130 21960
rect 15572 21248 15892 21808
rect 15572 21184 15580 21248
rect 15644 21184 15660 21248
rect 15724 21184 15740 21248
rect 15804 21184 15820 21248
rect 15884 21184 15892 21248
rect 15572 20160 15892 21184
rect 15572 20096 15580 20160
rect 15644 20096 15660 20160
rect 15724 20096 15740 20160
rect 15804 20096 15820 20160
rect 15884 20096 15892 20160
rect 15572 19072 15892 20096
rect 15572 19008 15580 19072
rect 15644 19008 15660 19072
rect 15724 19008 15740 19072
rect 15804 19008 15820 19072
rect 15884 19008 15892 19072
rect 15331 19004 15397 19005
rect 15331 18940 15332 19004
rect 15396 18940 15397 19004
rect 15331 18939 15397 18940
rect 15147 18052 15213 18053
rect 15147 17988 15148 18052
rect 15212 17988 15213 18052
rect 15147 17987 15213 17988
rect 15150 15197 15210 17987
rect 15572 17984 15892 19008
rect 16070 18869 16130 21900
rect 16438 19141 16498 22304
rect 16990 19141 17050 22304
rect 17542 22104 17602 22304
rect 18094 22104 18154 22304
rect 18646 22104 18706 22304
rect 19198 22104 19258 22304
rect 19750 22104 19810 22304
rect 20302 22104 20362 22304
rect 20854 22104 20914 22304
rect 21406 22104 21466 22304
rect 21958 21861 22018 22304
rect 21955 21860 22021 21861
rect 19367 21792 19687 21808
rect 21955 21796 21956 21860
rect 22020 21796 22021 21860
rect 21955 21795 22021 21796
rect 19367 21728 19375 21792
rect 19439 21728 19455 21792
rect 19519 21728 19535 21792
rect 19599 21728 19615 21792
rect 19679 21728 19687 21792
rect 19367 20704 19687 21728
rect 19367 20640 19375 20704
rect 19439 20640 19455 20704
rect 19519 20640 19535 20704
rect 19599 20640 19615 20704
rect 19679 20640 19687 20704
rect 19367 19616 19687 20640
rect 19367 19552 19375 19616
rect 19439 19552 19455 19616
rect 19519 19552 19535 19616
rect 19599 19552 19615 19616
rect 19679 19552 19687 19616
rect 16435 19140 16501 19141
rect 16435 19076 16436 19140
rect 16500 19076 16501 19140
rect 16435 19075 16501 19076
rect 16987 19140 17053 19141
rect 16987 19076 16988 19140
rect 17052 19076 17053 19140
rect 16987 19075 17053 19076
rect 16067 18868 16133 18869
rect 16067 18804 16068 18868
rect 16132 18804 16133 18868
rect 16067 18803 16133 18804
rect 15572 17920 15580 17984
rect 15644 17920 15660 17984
rect 15724 17920 15740 17984
rect 15804 17920 15820 17984
rect 15884 17920 15892 17984
rect 15572 16896 15892 17920
rect 19367 18528 19687 19552
rect 22510 18597 22570 22304
rect 23062 22130 23122 22304
rect 22878 22070 23122 22130
rect 22878 19277 22938 22070
rect 23614 21861 23674 22304
rect 23611 21860 23677 21861
rect 23162 21248 23482 21808
rect 23611 21796 23612 21860
rect 23676 21796 23677 21860
rect 23611 21795 23677 21796
rect 23162 21184 23170 21248
rect 23234 21184 23250 21248
rect 23314 21184 23330 21248
rect 23394 21184 23410 21248
rect 23474 21184 23482 21248
rect 23162 20160 23482 21184
rect 23162 20096 23170 20160
rect 23234 20096 23250 20160
rect 23314 20096 23330 20160
rect 23394 20096 23410 20160
rect 23474 20096 23482 20160
rect 22875 19276 22941 19277
rect 22875 19212 22876 19276
rect 22940 19212 22941 19276
rect 22875 19211 22941 19212
rect 23162 19072 23482 20096
rect 23162 19008 23170 19072
rect 23234 19008 23250 19072
rect 23314 19008 23330 19072
rect 23394 19008 23410 19072
rect 23474 19008 23482 19072
rect 22507 18596 22573 18597
rect 22507 18532 22508 18596
rect 22572 18532 22573 18596
rect 22507 18531 22573 18532
rect 19367 18464 19375 18528
rect 19439 18464 19455 18528
rect 19519 18464 19535 18528
rect 19599 18464 19615 18528
rect 19679 18464 19687 18528
rect 16067 17916 16133 17917
rect 16067 17852 16068 17916
rect 16132 17852 16133 17916
rect 16067 17851 16133 17852
rect 15572 16832 15580 16896
rect 15644 16832 15660 16896
rect 15724 16832 15740 16896
rect 15804 16832 15820 16896
rect 15884 16832 15892 16896
rect 15572 15808 15892 16832
rect 15572 15744 15580 15808
rect 15644 15744 15660 15808
rect 15724 15744 15740 15808
rect 15804 15744 15820 15808
rect 15884 15744 15892 15808
rect 15147 15196 15213 15197
rect 15147 15132 15148 15196
rect 15212 15132 15213 15196
rect 15147 15131 15213 15132
rect 15572 14720 15892 15744
rect 15572 14656 15580 14720
rect 15644 14656 15660 14720
rect 15724 14656 15740 14720
rect 15804 14656 15820 14720
rect 15884 14656 15892 14720
rect 15572 13632 15892 14656
rect 15572 13568 15580 13632
rect 15644 13568 15660 13632
rect 15724 13568 15740 13632
rect 15804 13568 15820 13632
rect 15884 13568 15892 13632
rect 15572 12544 15892 13568
rect 15572 12480 15580 12544
rect 15644 12480 15660 12544
rect 15724 12480 15740 12544
rect 15804 12480 15820 12544
rect 15884 12480 15892 12544
rect 14043 11796 14109 11797
rect 14043 11732 14044 11796
rect 14108 11732 14109 11796
rect 14043 11731 14109 11732
rect 15572 11456 15892 12480
rect 16070 11661 16130 17851
rect 19367 17440 19687 18464
rect 19367 17376 19375 17440
rect 19439 17376 19455 17440
rect 19519 17376 19535 17440
rect 19599 17376 19615 17440
rect 19679 17376 19687 17440
rect 19367 16352 19687 17376
rect 19367 16288 19375 16352
rect 19439 16288 19455 16352
rect 19519 16288 19535 16352
rect 19599 16288 19615 16352
rect 19679 16288 19687 16352
rect 19367 15264 19687 16288
rect 19367 15200 19375 15264
rect 19439 15200 19455 15264
rect 19519 15200 19535 15264
rect 19599 15200 19615 15264
rect 19679 15200 19687 15264
rect 19367 14176 19687 15200
rect 19367 14112 19375 14176
rect 19439 14112 19455 14176
rect 19519 14112 19535 14176
rect 19599 14112 19615 14176
rect 19679 14112 19687 14176
rect 19367 13088 19687 14112
rect 23162 17984 23482 19008
rect 24166 18461 24226 22304
rect 24350 22174 24594 22234
rect 24350 20773 24410 22174
rect 24534 22130 24594 22174
rect 24718 22130 24778 22304
rect 24534 22070 24778 22130
rect 24347 20772 24413 20773
rect 24347 20708 24348 20772
rect 24412 20708 24413 20772
rect 24347 20707 24413 20708
rect 25270 19277 25330 22304
rect 25822 21450 25882 22304
rect 25638 21390 25882 21450
rect 25638 21045 25698 21390
rect 26374 21181 26434 22304
rect 26926 22104 26986 22304
rect 27478 22104 27538 22304
rect 26957 21792 27277 21808
rect 26957 21728 26965 21792
rect 27029 21728 27045 21792
rect 27109 21728 27125 21792
rect 27189 21728 27205 21792
rect 27269 21728 27277 21792
rect 26371 21180 26437 21181
rect 26371 21116 26372 21180
rect 26436 21116 26437 21180
rect 26371 21115 26437 21116
rect 25635 21044 25701 21045
rect 25635 20980 25636 21044
rect 25700 20980 25701 21044
rect 25635 20979 25701 20980
rect 26957 20704 27277 21728
rect 30752 21248 31072 21808
rect 30752 21184 30760 21248
rect 30824 21184 30840 21248
rect 30904 21184 30920 21248
rect 30984 21184 31000 21248
rect 31064 21184 31072 21248
rect 27659 20908 27725 20909
rect 27659 20844 27660 20908
rect 27724 20844 27725 20908
rect 27659 20843 27725 20844
rect 26957 20640 26965 20704
rect 27029 20640 27045 20704
rect 27109 20640 27125 20704
rect 27189 20640 27205 20704
rect 27269 20640 27277 20704
rect 26957 19616 27277 20640
rect 26957 19552 26965 19616
rect 27029 19552 27045 19616
rect 27109 19552 27125 19616
rect 27189 19552 27205 19616
rect 27269 19552 27277 19616
rect 25267 19276 25333 19277
rect 25267 19212 25268 19276
rect 25332 19212 25333 19276
rect 25267 19211 25333 19212
rect 26739 19140 26805 19141
rect 26739 19076 26740 19140
rect 26804 19076 26805 19140
rect 26739 19075 26805 19076
rect 24163 18460 24229 18461
rect 24163 18396 24164 18460
rect 24228 18396 24229 18460
rect 24163 18395 24229 18396
rect 24163 18052 24229 18053
rect 24163 17988 24164 18052
rect 24228 17988 24229 18052
rect 24163 17987 24229 17988
rect 23162 17920 23170 17984
rect 23234 17920 23250 17984
rect 23314 17920 23330 17984
rect 23394 17920 23410 17984
rect 23474 17920 23482 17984
rect 23162 16896 23482 17920
rect 23162 16832 23170 16896
rect 23234 16832 23250 16896
rect 23314 16832 23330 16896
rect 23394 16832 23410 16896
rect 23474 16832 23482 16896
rect 23162 15808 23482 16832
rect 24166 16285 24226 17987
rect 26187 16828 26253 16829
rect 26187 16764 26188 16828
rect 26252 16764 26253 16828
rect 26187 16763 26253 16764
rect 24163 16284 24229 16285
rect 24163 16220 24164 16284
rect 24228 16220 24229 16284
rect 24163 16219 24229 16220
rect 23162 15744 23170 15808
rect 23234 15744 23250 15808
rect 23314 15744 23330 15808
rect 23394 15744 23410 15808
rect 23474 15744 23482 15808
rect 23162 14720 23482 15744
rect 26190 15061 26250 16763
rect 26742 15061 26802 19075
rect 26957 18528 27277 19552
rect 26957 18464 26965 18528
rect 27029 18464 27045 18528
rect 27109 18464 27125 18528
rect 27189 18464 27205 18528
rect 27269 18464 27277 18528
rect 26957 17440 27277 18464
rect 26957 17376 26965 17440
rect 27029 17376 27045 17440
rect 27109 17376 27125 17440
rect 27189 17376 27205 17440
rect 27269 17376 27277 17440
rect 26957 16352 27277 17376
rect 27475 16964 27541 16965
rect 27475 16900 27476 16964
rect 27540 16900 27541 16964
rect 27475 16899 27541 16900
rect 26957 16288 26965 16352
rect 27029 16288 27045 16352
rect 27109 16288 27125 16352
rect 27189 16288 27205 16352
rect 27269 16288 27277 16352
rect 26957 15264 27277 16288
rect 26957 15200 26965 15264
rect 27029 15200 27045 15264
rect 27109 15200 27125 15264
rect 27189 15200 27205 15264
rect 27269 15200 27277 15264
rect 26187 15060 26253 15061
rect 26187 14996 26188 15060
rect 26252 14996 26253 15060
rect 26187 14995 26253 14996
rect 26739 15060 26805 15061
rect 26739 14996 26740 15060
rect 26804 14996 26805 15060
rect 26739 14995 26805 14996
rect 23162 14656 23170 14720
rect 23234 14656 23250 14720
rect 23314 14656 23330 14720
rect 23394 14656 23410 14720
rect 23474 14656 23482 14720
rect 20667 13836 20733 13837
rect 20667 13772 20668 13836
rect 20732 13772 20733 13836
rect 20667 13771 20733 13772
rect 19367 13024 19375 13088
rect 19439 13024 19455 13088
rect 19519 13024 19535 13088
rect 19599 13024 19615 13088
rect 19679 13024 19687 13088
rect 19367 12000 19687 13024
rect 19747 12884 19813 12885
rect 19747 12820 19748 12884
rect 19812 12820 19813 12884
rect 19747 12819 19813 12820
rect 19367 11936 19375 12000
rect 19439 11936 19455 12000
rect 19519 11936 19535 12000
rect 19599 11936 19615 12000
rect 19679 11936 19687 12000
rect 16067 11660 16133 11661
rect 16067 11596 16068 11660
rect 16132 11596 16133 11660
rect 16067 11595 16133 11596
rect 15572 11392 15580 11456
rect 15644 11392 15660 11456
rect 15724 11392 15740 11456
rect 15804 11392 15820 11456
rect 15884 11392 15892 11456
rect 13494 11190 14106 11250
rect 11777 10848 11785 10912
rect 11849 10848 11865 10912
rect 11929 10848 11945 10912
rect 12009 10848 12025 10912
rect 12089 10848 12097 10912
rect 9259 10028 9325 10029
rect 9259 9964 9260 10028
rect 9324 9964 9325 10028
rect 9259 9963 9325 9964
rect 7982 9216 7990 9280
rect 8054 9216 8070 9280
rect 8134 9216 8150 9280
rect 8214 9216 8230 9280
rect 8294 9216 8302 9280
rect 7982 8192 8302 9216
rect 7982 8128 7990 8192
rect 8054 8128 8070 8192
rect 8134 8128 8150 8192
rect 8214 8128 8230 8192
rect 8294 8128 8302 8192
rect 7982 7104 8302 8128
rect 7982 7040 7990 7104
rect 8054 7040 8070 7104
rect 8134 7040 8150 7104
rect 8214 7040 8230 7104
rect 8294 7040 8302 7104
rect 6867 6492 6933 6493
rect 6867 6428 6868 6492
rect 6932 6428 6933 6492
rect 6867 6427 6933 6428
rect 7982 6016 8302 7040
rect 7982 5952 7990 6016
rect 8054 5952 8070 6016
rect 8134 5952 8150 6016
rect 8214 5952 8230 6016
rect 8294 5952 8302 6016
rect 7982 4928 8302 5952
rect 7982 4864 7990 4928
rect 8054 4864 8070 4928
rect 8134 4864 8150 4928
rect 8214 4864 8230 4928
rect 8294 4864 8302 4928
rect 7982 3840 8302 4864
rect 7982 3776 7990 3840
rect 8054 3776 8070 3840
rect 8134 3776 8150 3840
rect 8214 3776 8230 3840
rect 8294 3776 8302 3840
rect 7982 2752 8302 3776
rect 7982 2688 7990 2752
rect 8054 2688 8070 2752
rect 8134 2688 8150 2752
rect 8214 2688 8230 2752
rect 8294 2688 8302 2752
rect 5579 2684 5645 2685
rect 5579 2620 5580 2684
rect 5644 2620 5645 2684
rect 5579 2619 5645 2620
rect 6683 2684 6749 2685
rect 6683 2620 6684 2684
rect 6748 2620 6749 2684
rect 6683 2619 6749 2620
rect 5395 1732 5461 1733
rect 5395 1668 5396 1732
rect 5460 1668 5461 1732
rect 5395 1667 5461 1668
rect 4187 1056 4195 1120
rect 4259 1056 4275 1120
rect 4339 1056 4355 1120
rect 4419 1056 4435 1120
rect 4499 1056 4507 1120
rect 4187 496 4507 1056
rect 7982 1664 8302 2688
rect 7982 1600 7990 1664
rect 8054 1600 8070 1664
rect 8134 1600 8150 1664
rect 8214 1600 8230 1664
rect 8294 1600 8302 1664
rect 7982 576 8302 1600
rect 7982 512 7990 576
rect 8054 512 8070 576
rect 8134 512 8150 576
rect 8214 512 8230 576
rect 8294 512 8302 576
rect 7982 496 8302 512
rect 11777 9824 12097 10848
rect 11777 9760 11785 9824
rect 11849 9760 11865 9824
rect 11929 9760 11945 9824
rect 12009 9760 12025 9824
rect 12089 9760 12097 9824
rect 11777 8736 12097 9760
rect 14046 8941 14106 11190
rect 15572 10368 15892 11392
rect 15572 10304 15580 10368
rect 15644 10304 15660 10368
rect 15724 10304 15740 10368
rect 15804 10304 15820 10368
rect 15884 10304 15892 10368
rect 15572 9280 15892 10304
rect 15572 9216 15580 9280
rect 15644 9216 15660 9280
rect 15724 9216 15740 9280
rect 15804 9216 15820 9280
rect 15884 9216 15892 9280
rect 14043 8940 14109 8941
rect 14043 8876 14044 8940
rect 14108 8876 14109 8940
rect 14043 8875 14109 8876
rect 11777 8672 11785 8736
rect 11849 8672 11865 8736
rect 11929 8672 11945 8736
rect 12009 8672 12025 8736
rect 12089 8672 12097 8736
rect 11777 7648 12097 8672
rect 11777 7584 11785 7648
rect 11849 7584 11865 7648
rect 11929 7584 11945 7648
rect 12009 7584 12025 7648
rect 12089 7584 12097 7648
rect 11777 6560 12097 7584
rect 11777 6496 11785 6560
rect 11849 6496 11865 6560
rect 11929 6496 11945 6560
rect 12009 6496 12025 6560
rect 12089 6496 12097 6560
rect 11777 5472 12097 6496
rect 11777 5408 11785 5472
rect 11849 5408 11865 5472
rect 11929 5408 11945 5472
rect 12009 5408 12025 5472
rect 12089 5408 12097 5472
rect 11777 4384 12097 5408
rect 11777 4320 11785 4384
rect 11849 4320 11865 4384
rect 11929 4320 11945 4384
rect 12009 4320 12025 4384
rect 12089 4320 12097 4384
rect 11777 3296 12097 4320
rect 11777 3232 11785 3296
rect 11849 3232 11865 3296
rect 11929 3232 11945 3296
rect 12009 3232 12025 3296
rect 12089 3232 12097 3296
rect 11777 2208 12097 3232
rect 11777 2144 11785 2208
rect 11849 2144 11865 2208
rect 11929 2144 11945 2208
rect 12009 2144 12025 2208
rect 12089 2144 12097 2208
rect 11777 1120 12097 2144
rect 11777 1056 11785 1120
rect 11849 1056 11865 1120
rect 11929 1056 11945 1120
rect 12009 1056 12025 1120
rect 12089 1056 12097 1120
rect 11777 496 12097 1056
rect 15572 8192 15892 9216
rect 15572 8128 15580 8192
rect 15644 8128 15660 8192
rect 15724 8128 15740 8192
rect 15804 8128 15820 8192
rect 15884 8128 15892 8192
rect 15572 7104 15892 8128
rect 15572 7040 15580 7104
rect 15644 7040 15660 7104
rect 15724 7040 15740 7104
rect 15804 7040 15820 7104
rect 15884 7040 15892 7104
rect 15572 6016 15892 7040
rect 15572 5952 15580 6016
rect 15644 5952 15660 6016
rect 15724 5952 15740 6016
rect 15804 5952 15820 6016
rect 15884 5952 15892 6016
rect 15572 4928 15892 5952
rect 15572 4864 15580 4928
rect 15644 4864 15660 4928
rect 15724 4864 15740 4928
rect 15804 4864 15820 4928
rect 15884 4864 15892 4928
rect 15572 3840 15892 4864
rect 15572 3776 15580 3840
rect 15644 3776 15660 3840
rect 15724 3776 15740 3840
rect 15804 3776 15820 3840
rect 15884 3776 15892 3840
rect 15572 2752 15892 3776
rect 15572 2688 15580 2752
rect 15644 2688 15660 2752
rect 15724 2688 15740 2752
rect 15804 2688 15820 2752
rect 15884 2688 15892 2752
rect 15572 1664 15892 2688
rect 15572 1600 15580 1664
rect 15644 1600 15660 1664
rect 15724 1600 15740 1664
rect 15804 1600 15820 1664
rect 15884 1600 15892 1664
rect 15572 576 15892 1600
rect 15572 512 15580 576
rect 15644 512 15660 576
rect 15724 512 15740 576
rect 15804 512 15820 576
rect 15884 512 15892 576
rect 15572 496 15892 512
rect 19367 10912 19687 11936
rect 19367 10848 19375 10912
rect 19439 10848 19455 10912
rect 19519 10848 19535 10912
rect 19599 10848 19615 10912
rect 19679 10848 19687 10912
rect 19367 9824 19687 10848
rect 19750 10165 19810 12819
rect 20670 11117 20730 13771
rect 23162 13632 23482 14656
rect 23162 13568 23170 13632
rect 23234 13568 23250 13632
rect 23314 13568 23330 13632
rect 23394 13568 23410 13632
rect 23474 13568 23482 13632
rect 23162 12544 23482 13568
rect 23162 12480 23170 12544
rect 23234 12480 23250 12544
rect 23314 12480 23330 12544
rect 23394 12480 23410 12544
rect 23474 12480 23482 12544
rect 23162 11456 23482 12480
rect 23162 11392 23170 11456
rect 23234 11392 23250 11456
rect 23314 11392 23330 11456
rect 23394 11392 23410 11456
rect 23474 11392 23482 11456
rect 20667 11116 20733 11117
rect 20667 11052 20668 11116
rect 20732 11052 20733 11116
rect 20667 11051 20733 11052
rect 23162 10368 23482 11392
rect 23162 10304 23170 10368
rect 23234 10304 23250 10368
rect 23314 10304 23330 10368
rect 23394 10304 23410 10368
rect 23474 10304 23482 10368
rect 19747 10164 19813 10165
rect 19747 10100 19748 10164
rect 19812 10100 19813 10164
rect 19747 10099 19813 10100
rect 19367 9760 19375 9824
rect 19439 9760 19455 9824
rect 19519 9760 19535 9824
rect 19599 9760 19615 9824
rect 19679 9760 19687 9824
rect 19367 8736 19687 9760
rect 19367 8672 19375 8736
rect 19439 8672 19455 8736
rect 19519 8672 19535 8736
rect 19599 8672 19615 8736
rect 19679 8672 19687 8736
rect 19367 7648 19687 8672
rect 19367 7584 19375 7648
rect 19439 7584 19455 7648
rect 19519 7584 19535 7648
rect 19599 7584 19615 7648
rect 19679 7584 19687 7648
rect 19367 6560 19687 7584
rect 19367 6496 19375 6560
rect 19439 6496 19455 6560
rect 19519 6496 19535 6560
rect 19599 6496 19615 6560
rect 19679 6496 19687 6560
rect 19367 5472 19687 6496
rect 19367 5408 19375 5472
rect 19439 5408 19455 5472
rect 19519 5408 19535 5472
rect 19599 5408 19615 5472
rect 19679 5408 19687 5472
rect 19367 4384 19687 5408
rect 19367 4320 19375 4384
rect 19439 4320 19455 4384
rect 19519 4320 19535 4384
rect 19599 4320 19615 4384
rect 19679 4320 19687 4384
rect 19367 3296 19687 4320
rect 19367 3232 19375 3296
rect 19439 3232 19455 3296
rect 19519 3232 19535 3296
rect 19599 3232 19615 3296
rect 19679 3232 19687 3296
rect 19367 2208 19687 3232
rect 19367 2144 19375 2208
rect 19439 2144 19455 2208
rect 19519 2144 19535 2208
rect 19599 2144 19615 2208
rect 19679 2144 19687 2208
rect 19367 1120 19687 2144
rect 19367 1056 19375 1120
rect 19439 1056 19455 1120
rect 19519 1056 19535 1120
rect 19599 1056 19615 1120
rect 19679 1056 19687 1120
rect 19367 496 19687 1056
rect 23162 9280 23482 10304
rect 23162 9216 23170 9280
rect 23234 9216 23250 9280
rect 23314 9216 23330 9280
rect 23394 9216 23410 9280
rect 23474 9216 23482 9280
rect 23162 8192 23482 9216
rect 23162 8128 23170 8192
rect 23234 8128 23250 8192
rect 23314 8128 23330 8192
rect 23394 8128 23410 8192
rect 23474 8128 23482 8192
rect 23162 7104 23482 8128
rect 23162 7040 23170 7104
rect 23234 7040 23250 7104
rect 23314 7040 23330 7104
rect 23394 7040 23410 7104
rect 23474 7040 23482 7104
rect 23162 6016 23482 7040
rect 23162 5952 23170 6016
rect 23234 5952 23250 6016
rect 23314 5952 23330 6016
rect 23394 5952 23410 6016
rect 23474 5952 23482 6016
rect 23162 4928 23482 5952
rect 23162 4864 23170 4928
rect 23234 4864 23250 4928
rect 23314 4864 23330 4928
rect 23394 4864 23410 4928
rect 23474 4864 23482 4928
rect 23162 3840 23482 4864
rect 23162 3776 23170 3840
rect 23234 3776 23250 3840
rect 23314 3776 23330 3840
rect 23394 3776 23410 3840
rect 23474 3776 23482 3840
rect 23162 2752 23482 3776
rect 23162 2688 23170 2752
rect 23234 2688 23250 2752
rect 23314 2688 23330 2752
rect 23394 2688 23410 2752
rect 23474 2688 23482 2752
rect 23162 1664 23482 2688
rect 23162 1600 23170 1664
rect 23234 1600 23250 1664
rect 23314 1600 23330 1664
rect 23394 1600 23410 1664
rect 23474 1600 23482 1664
rect 23162 576 23482 1600
rect 23162 512 23170 576
rect 23234 512 23250 576
rect 23314 512 23330 576
rect 23394 512 23410 576
rect 23474 512 23482 576
rect 23162 496 23482 512
rect 26957 14176 27277 15200
rect 27478 14381 27538 16899
rect 27662 14925 27722 20843
rect 30752 20160 31072 21184
rect 30752 20096 30760 20160
rect 30824 20096 30840 20160
rect 30904 20096 30920 20160
rect 30984 20096 31000 20160
rect 31064 20096 31072 20160
rect 29315 19140 29381 19141
rect 29315 19076 29316 19140
rect 29380 19076 29381 19140
rect 29315 19075 29381 19076
rect 28395 18460 28461 18461
rect 28395 18396 28396 18460
rect 28460 18396 28461 18460
rect 28395 18395 28461 18396
rect 27659 14924 27725 14925
rect 27659 14860 27660 14924
rect 27724 14860 27725 14924
rect 27659 14859 27725 14860
rect 27475 14380 27541 14381
rect 27475 14316 27476 14380
rect 27540 14316 27541 14380
rect 27475 14315 27541 14316
rect 26957 14112 26965 14176
rect 27029 14112 27045 14176
rect 27109 14112 27125 14176
rect 27189 14112 27205 14176
rect 27269 14112 27277 14176
rect 26957 13088 27277 14112
rect 28398 13837 28458 18395
rect 29318 15877 29378 19075
rect 30752 19072 31072 20096
rect 30752 19008 30760 19072
rect 30824 19008 30840 19072
rect 30904 19008 30920 19072
rect 30984 19008 31000 19072
rect 31064 19008 31072 19072
rect 30419 18052 30485 18053
rect 30419 17988 30420 18052
rect 30484 17988 30485 18052
rect 30419 17987 30485 17988
rect 29499 17644 29565 17645
rect 29499 17580 29500 17644
rect 29564 17580 29565 17644
rect 29499 17579 29565 17580
rect 29315 15876 29381 15877
rect 29315 15812 29316 15876
rect 29380 15812 29381 15876
rect 29315 15811 29381 15812
rect 29131 15468 29197 15469
rect 29131 15404 29132 15468
rect 29196 15404 29197 15468
rect 29131 15403 29197 15404
rect 28579 13972 28645 13973
rect 28579 13908 28580 13972
rect 28644 13908 28645 13972
rect 28579 13907 28645 13908
rect 28395 13836 28461 13837
rect 28395 13772 28396 13836
rect 28460 13772 28461 13836
rect 28395 13771 28461 13772
rect 26957 13024 26965 13088
rect 27029 13024 27045 13088
rect 27109 13024 27125 13088
rect 27189 13024 27205 13088
rect 27269 13024 27277 13088
rect 26957 12000 27277 13024
rect 26957 11936 26965 12000
rect 27029 11936 27045 12000
rect 27109 11936 27125 12000
rect 27189 11936 27205 12000
rect 27269 11936 27277 12000
rect 26957 10912 27277 11936
rect 26957 10848 26965 10912
rect 27029 10848 27045 10912
rect 27109 10848 27125 10912
rect 27189 10848 27205 10912
rect 27269 10848 27277 10912
rect 26957 9824 27277 10848
rect 26957 9760 26965 9824
rect 27029 9760 27045 9824
rect 27109 9760 27125 9824
rect 27189 9760 27205 9824
rect 27269 9760 27277 9824
rect 26957 8736 27277 9760
rect 26957 8672 26965 8736
rect 27029 8672 27045 8736
rect 27109 8672 27125 8736
rect 27189 8672 27205 8736
rect 27269 8672 27277 8736
rect 26957 7648 27277 8672
rect 26957 7584 26965 7648
rect 27029 7584 27045 7648
rect 27109 7584 27125 7648
rect 27189 7584 27205 7648
rect 27269 7584 27277 7648
rect 26957 6560 27277 7584
rect 28582 6901 28642 13907
rect 29134 12069 29194 15403
rect 29502 15333 29562 17579
rect 29683 16692 29749 16693
rect 29683 16628 29684 16692
rect 29748 16628 29749 16692
rect 29683 16627 29749 16628
rect 29686 15605 29746 16627
rect 30422 15605 30482 17987
rect 30752 17984 31072 19008
rect 30752 17920 30760 17984
rect 30824 17920 30840 17984
rect 30904 17920 30920 17984
rect 30984 17920 31000 17984
rect 31064 17920 31072 17984
rect 30752 16896 31072 17920
rect 30752 16832 30760 16896
rect 30824 16832 30840 16896
rect 30904 16832 30920 16896
rect 30984 16832 31000 16896
rect 31064 16832 31072 16896
rect 30752 15808 31072 16832
rect 30752 15744 30760 15808
rect 30824 15744 30840 15808
rect 30904 15744 30920 15808
rect 30984 15744 31000 15808
rect 31064 15744 31072 15808
rect 29683 15604 29749 15605
rect 29683 15540 29684 15604
rect 29748 15540 29749 15604
rect 29683 15539 29749 15540
rect 30419 15604 30485 15605
rect 30419 15540 30420 15604
rect 30484 15540 30485 15604
rect 30419 15539 30485 15540
rect 29499 15332 29565 15333
rect 29499 15268 29500 15332
rect 29564 15268 29565 15332
rect 29499 15267 29565 15268
rect 30752 14720 31072 15744
rect 30752 14656 30760 14720
rect 30824 14656 30840 14720
rect 30904 14656 30920 14720
rect 30984 14656 31000 14720
rect 31064 14656 31072 14720
rect 30752 13632 31072 14656
rect 30752 13568 30760 13632
rect 30824 13568 30840 13632
rect 30904 13568 30920 13632
rect 30984 13568 31000 13632
rect 31064 13568 31072 13632
rect 30752 12544 31072 13568
rect 30752 12480 30760 12544
rect 30824 12480 30840 12544
rect 30904 12480 30920 12544
rect 30984 12480 31000 12544
rect 31064 12480 31072 12544
rect 29131 12068 29197 12069
rect 29131 12004 29132 12068
rect 29196 12004 29197 12068
rect 29131 12003 29197 12004
rect 30752 11456 31072 12480
rect 30752 11392 30760 11456
rect 30824 11392 30840 11456
rect 30904 11392 30920 11456
rect 30984 11392 31000 11456
rect 31064 11392 31072 11456
rect 30752 10368 31072 11392
rect 30752 10304 30760 10368
rect 30824 10304 30840 10368
rect 30904 10304 30920 10368
rect 30984 10304 31000 10368
rect 31064 10304 31072 10368
rect 30752 9280 31072 10304
rect 30752 9216 30760 9280
rect 30824 9216 30840 9280
rect 30904 9216 30920 9280
rect 30984 9216 31000 9280
rect 31064 9216 31072 9280
rect 30752 8192 31072 9216
rect 30752 8128 30760 8192
rect 30824 8128 30840 8192
rect 30904 8128 30920 8192
rect 30984 8128 31000 8192
rect 31064 8128 31072 8192
rect 30752 7104 31072 8128
rect 30752 7040 30760 7104
rect 30824 7040 30840 7104
rect 30904 7040 30920 7104
rect 30984 7040 31000 7104
rect 31064 7040 31072 7104
rect 28579 6900 28645 6901
rect 28579 6836 28580 6900
rect 28644 6836 28645 6900
rect 28579 6835 28645 6836
rect 26957 6496 26965 6560
rect 27029 6496 27045 6560
rect 27109 6496 27125 6560
rect 27189 6496 27205 6560
rect 27269 6496 27277 6560
rect 26957 5472 27277 6496
rect 26957 5408 26965 5472
rect 27029 5408 27045 5472
rect 27109 5408 27125 5472
rect 27189 5408 27205 5472
rect 27269 5408 27277 5472
rect 26957 4384 27277 5408
rect 26957 4320 26965 4384
rect 27029 4320 27045 4384
rect 27109 4320 27125 4384
rect 27189 4320 27205 4384
rect 27269 4320 27277 4384
rect 26957 3296 27277 4320
rect 26957 3232 26965 3296
rect 27029 3232 27045 3296
rect 27109 3232 27125 3296
rect 27189 3232 27205 3296
rect 27269 3232 27277 3296
rect 26957 2208 27277 3232
rect 26957 2144 26965 2208
rect 27029 2144 27045 2208
rect 27109 2144 27125 2208
rect 27189 2144 27205 2208
rect 27269 2144 27277 2208
rect 26957 1120 27277 2144
rect 26957 1056 26965 1120
rect 27029 1056 27045 1120
rect 27109 1056 27125 1120
rect 27189 1056 27205 1120
rect 27269 1056 27277 1120
rect 26957 496 27277 1056
rect 30752 6016 31072 7040
rect 30752 5952 30760 6016
rect 30824 5952 30840 6016
rect 30904 5952 30920 6016
rect 30984 5952 31000 6016
rect 31064 5952 31072 6016
rect 30752 4928 31072 5952
rect 30752 4864 30760 4928
rect 30824 4864 30840 4928
rect 30904 4864 30920 4928
rect 30984 4864 31000 4928
rect 31064 4864 31072 4928
rect 30752 3840 31072 4864
rect 30752 3776 30760 3840
rect 30824 3776 30840 3840
rect 30904 3776 30920 3840
rect 30984 3776 31000 3840
rect 31064 3776 31072 3840
rect 30752 2752 31072 3776
rect 30752 2688 30760 2752
rect 30824 2688 30840 2752
rect 30904 2688 30920 2752
rect 30984 2688 31000 2752
rect 31064 2688 31072 2752
rect 30752 1664 31072 2688
rect 30752 1600 30760 1664
rect 30824 1600 30840 1664
rect 30904 1600 30920 1664
rect 30984 1600 31000 1664
rect 31064 1600 31072 1664
rect 30752 576 31072 1600
rect 30752 512 30760 576
rect 30824 512 30840 576
rect 30904 512 30920 576
rect 30984 512 31000 576
rect 31064 512 31072 576
rect 30752 496 31072 512
use sky130_fd_sc_hd__inv_2  _05_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 15732 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _06_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 21252 0 1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _07_
timestamp 1693170804
transform 1 0 23828 0 1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _08_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 23000 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _09_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 23184 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _10_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 18124 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _11_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 13156 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4600 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _21_
timestamp 1693170804
transform 1 0 11224 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _22_
timestamp 1693170804
transform 1 0 3496 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _23_
timestamp 1693170804
transform 1 0 20424 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _24_
timestamp 1693170804
transform 1 0 4048 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _25_
timestamp 1693170804
transform 1 0 4600 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _26_
timestamp 1693170804
transform 1 0 3496 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _27_
timestamp 1693170804
transform 1 0 8096 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 12328 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1693170804
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1693170804
transform 1 0 26036 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1693170804
transform 1 0 24012 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1693170804
transform 1 0 16284 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1693170804
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1693170804
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1693170804
transform 1 0 16560 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1693170804
transform 1 0 12696 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1693170804
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1693170804
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1693170804
transform 1 0 30360 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1693170804
transform 1 0 15732 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1693170804
transform 1 0 1288 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1693170804
transform 1 0 11868 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1693170804
transform 1 0 29992 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1693170804
transform 1 0 11500 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1693170804
transform 1 0 20976 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1693170804
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1693170804
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1693170804
transform 1 0 15364 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1693170804
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1693170804
transform 1 0 11132 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1693170804
transform 1 0 12236 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1693170804
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1693170804
transform 1 0 29992 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1693170804
transform 1 0 30360 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1693170804
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1693170804
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1693170804
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1693170804
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1693170804
transform 1 0 1288 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1693170804
transform 1 0 29624 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1693170804
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1693170804
transform 1 0 15364 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1693170804
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1693170804
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1693170804
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1693170804
transform 1 0 30360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1693170804
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1693170804
transform 1 0 30176 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_42
timestamp 1693170804
transform 1 0 13708 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_43
timestamp 1693170804
transform 1 0 20148 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_44
timestamp 1693170804
transform 1 0 4968 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_45
timestamp 1693170804
transform 1 0 30360 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_46
timestamp 1693170804
transform 1 0 1104 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_47
timestamp 1693170804
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_48
timestamp 1693170804
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_49
timestamp 1693170804
transform 1 0 6348 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_50
timestamp 1693170804
transform 1 0 30176 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_51
timestamp 1693170804
transform 1 0 30176 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_52
timestamp 1693170804
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_53
timestamp 1693170804
transform 1 0 29808 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_54
timestamp 1693170804
transform 1 0 29440 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_55
timestamp 1693170804
transform 1 0 4600 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_56
timestamp 1693170804
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2i_2  ct.cw.cc_test_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28980 0 1 20128
box -38 -48 1050 592
use sky130_ht_sc_tt05__mux2i_2  ct.cw.cc_test_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699029708
transform 1 0 28980 0 1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__maj3_2  ct.cw.cc_test_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28980 0 1 21216
box -38 -48 866 592
use sky130_ht_sc_tt05__maj3_2  ct.cw.cc_test_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699029708
transform 1 0 28980 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dlrtp_1  ct.cw.cc_test_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28980 0 1 19040
box -38 -48 1234 592
use sky130_ht_sc_tt05__dlrtp_1  ct.cw.cc_test_5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699029708
transform 1 0 28980 0 1 17952
box -38 -48 1418 592
use sky130_fd_sc_hd__dfrtp_1  ct.cw.cc_test_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28612 0 -1 17952
box -38 -48 1878 592
use sky130_ht_sc_tt05__dfrtp_1  ct.cw.cc_test_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699029708
transform 1 0 26404 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[0\].bits\[0\].cc_flop $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28612 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[0\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[0\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 14536 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[0\].cc_clkbuf
timestamp 1693170804
transform 1 0 28152 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[1\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[1\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[1\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 16836 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[1\].cc_clkbuf
timestamp 1693170804
transform 1 0 29808 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[2\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 26404 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[2\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[2\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 26772 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[2\].cc_clkbuf
timestamp 1693170804
transform 1 0 29992 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[3\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 6716 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[3\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[3\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[3\].cc_clkbuf
timestamp 1693170804
transform 1 0 26036 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[4\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 26404 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[4\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 24564 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[4\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 21988 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[4\].cc_clkbuf
timestamp 1693170804
transform 1 0 23552 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[5\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 828 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[5\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[5\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 16836 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[5\].cc_clkbuf
timestamp 1693170804
transform 1 0 23828 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[6\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 21988 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[6\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 16836 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[6\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[6\].cc_clkbuf
timestamp 1693170804
transform 1 0 23092 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[7\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 26864 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[7\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 26404 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[7\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[7\].cc_clkbuf
timestamp 1693170804
transform 1 0 23828 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[8\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 21252 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[8\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 19136 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[8\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 18676 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[8\].cc_clkbuf
timestamp 1693170804
transform 1 0 22540 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[9\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 18308 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[9\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 18676 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[9\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 24288 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[9\].cc_clkbuf
timestamp 1693170804
transform 1 0 18400 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[10\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 17940 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[10\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 16100 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[10\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 14260 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[10\].cc_clkbuf
timestamp 1693170804
transform 1 0 18676 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[11\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 18676 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[11\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 20424 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[11\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 16100 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[11\].cc_clkbuf
timestamp 1693170804
transform 1 0 10304 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[0\].cc_scanflop $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 13524 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 14904 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 7452 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 8464 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 20056 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8004 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 13800 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 12144 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[0\].cc_clkbuf
timestamp 1693170804
transform 1 0 17848 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[0\].rs_mbuf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8096 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 10764 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 17848 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 8464 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 10948 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[1\].bits\[6\].rs_cbuf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 5244 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[1\].cc_clkbuf
timestamp 1693170804
transform 1 0 5244 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[1\].rs_mbuf
timestamp 1693170804
transform 1 0 10672 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[2\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 10948 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[2\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 9200 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[2\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[2\].cc_clkbuf
timestamp 1693170804
transform 1 0 5152 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[2\].rs_mbuf
timestamp 1693170804
transform 1 0 5796 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 26036 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 24380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 5888 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 18032 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 11868 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 8648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 15732 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 8924 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11868 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 13432 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 12052 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[3\].cc_clkbuf
timestamp 1693170804
transform 1 0 2576 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[3\].rs_mbuf
timestamp 1693170804
transform 1 0 920 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5152 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 3772 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 5152 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[4\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 9844 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[4\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10396 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[4\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10120 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[4\].cc_clkbuf
timestamp 1693170804
transform 1 0 4048 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[4\].rs_mbuf
timestamp 1693170804
transform 1 0 3220 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 4324 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3772 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 4600 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3772 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 13248 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 1196 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 8924 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 6072 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[5\].cc_clkbuf
timestamp 1693170804
transform 1 0 3220 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[5\].rs_mbuf
timestamp 1693170804
transform 1 0 3220 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5980 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 6256 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 6532 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 9108 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 9384 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[6\].cc_clkbuf
timestamp 1693170804
transform 1 0 5796 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[6\].rs_mbuf
timestamp 1693170804
transform 1 0 8372 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 12696 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 11040 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 11316 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 11776 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 12972 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11500 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[7\].cc_clkbuf
timestamp 1693170804
transform 1 0 9936 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[7\].rs_mbuf
timestamp 1693170804
transform 1 0 11868 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 14168 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16836 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 14536 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 13616 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 13892 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 14628 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 13984 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[8\].cc_clkbuf
timestamp 1693170804
transform 1 0 11040 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[8\].rs_mbuf
timestamp 1693170804
transform 1 0 14720 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 17112 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 19136 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 19228 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 17112 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 19504 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 16652 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 19228 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 16560 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 16928 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 28152 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 16928 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[9\].cc_clkbuf
timestamp 1693170804
transform 1 0 16100 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[9\].rs_mbuf
timestamp 1693170804
transform 1 0 18676 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 21620 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 19412 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 19688 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 22172 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 19688 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 20332 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 20424 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 28612 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[10\].cc_clkbuf
timestamp 1693170804
transform 1 0 18676 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[10\].rs_mbuf
timestamp 1693170804
transform 1 0 22632 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 22724 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 23000 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 28612 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 23920 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24656 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[11\].cc_clkbuf
timestamp 1693170804
transform 1 0 23460 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[11\].rs_mbuf
timestamp 1693170804
transform 1 0 23184 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 26128 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 26036 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 26036 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 29992 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 28152 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 28612 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 24472 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 30176 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[12\].cc_clkbuf
timestamp 1693170804
transform 1 0 25668 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[12\].rs_mbuf
timestamp 1693170804
transform 1 0 26864 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 24472 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 26036 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 24104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 23184 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26036 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 28336 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 28428 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 29532 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 29808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[13\].cc_clkbuf
timestamp 1693170804
transform 1 0 28980 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[13\].rs_mbuf
timestamp 1693170804
transform 1 0 26680 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 22724 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 22448 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 21896 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 22172 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 29808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 27968 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 30084 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 27968 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 29900 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[14\].cc_clkbuf
timestamp 1693170804
transform 1 0 28980 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[14\].rs_mbuf
timestamp 1693170804
transform 1 0 23920 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 20700 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 19964 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 21528 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 19964 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 20240 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 21712 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 24472 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 27692 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 30268 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 27692 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[15\].cc_clkbuf
timestamp 1693170804
transform 1 0 28244 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[15\].rs_mbuf
timestamp 1693170804
transform 1 0 29532 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 18952 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 19228 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 19136 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 17940 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 23920 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 28520 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 28244 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[16\].cc_clkbuf
timestamp 1693170804
transform 1 0 25668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[16\].rs_mbuf
timestamp 1693170804
transform 1 0 17388 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 17112 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16836 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16744 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 17020 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 19504 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 19964 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 21712 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 24564 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 23184 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 26036 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 26036 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 25944 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[17\].cc_clkbuf
timestamp 1693170804
transform 1 0 18676 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[17\].rs_mbuf
timestamp 1693170804
transform 1 0 19320 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16560 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 19044 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 16836 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 16560 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 19320 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 25668 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 25392 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 22908 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 25116 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[18\].cc_clkbuf
timestamp 1693170804
transform 1 0 23828 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[18\].rs_mbuf
timestamp 1693170804
transform 1 0 20332 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 17756 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18032 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 17756 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 17756 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 18032 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 17480 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 20332 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 21988 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[19\].cc_clkbuf
timestamp 1693170804
transform 1 0 17940 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[19\].rs_mbuf
timestamp 1693170804
transform 1 0 18032 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 24288 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 27876 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 28520 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 27416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26312 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 25668 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 27968 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 27968 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 30084 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[20\].cc_clkbuf
timestamp 1693170804
transform 1 0 22356 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[20\].rs_mbuf
timestamp 1693170804
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3772 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 28612 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 27600 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[21\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[21\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__dlymetal6s2s_1  ct.oc.frame\[21\].bits\[6\].rs_cbuf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28980 0 1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[21\].cc_clkbuf
timestamp 1693170804
transform 1 0 27140 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[21\].rs_mbuf
timestamp 1693170804
transform 1 0 27324 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 27048 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18952 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26220 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 26680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26036 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 24472 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3588 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 27324 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 14168 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 27048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[22\].cc_clkbuf
timestamp 1693170804
transform 1 0 27232 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[22\].rs_mbuf
timestamp 1693170804
transform 1 0 26680 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[23\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 26680 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[23\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 25300 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 24472 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 24012 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 25944 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 24012 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 26220 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 25576 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[23\].cc_clkbuf
timestamp 1693170804
transform 1 0 26404 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[23\].rs_mbuf
timestamp 1693170804
transform 1 0 24748 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 23736 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 22264 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 23184 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 22080 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 23368 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 23092 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 22080 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 23092 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[24\].cc_clkbuf
timestamp 1693170804
transform 1 0 23184 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[24\].rs_mbuf
timestamp 1693170804
transform 1 0 22632 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 23092 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 23736 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 20332 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 20792 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 20608 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 23368 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[25\].cc_clkbuf
timestamp 1693170804
transform 1 0 20608 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[25\].rs_mbuf
timestamp 1693170804
transform 1 0 21252 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 20792 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 20608 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 18400 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 18400 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 20240 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 21804 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[26\].cc_clkbuf
timestamp 1693170804
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[26\].rs_mbuf
timestamp 1693170804
transform 1 0 19780 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 20516 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 16192 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 17204 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 16192 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 16192 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 18676 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 16192 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 13616 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[27\].cc_clkbuf
timestamp 1693170804
transform 1 0 19228 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[27\].rs_mbuf
timestamp 1693170804
transform 1 0 18676 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13892 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 12880 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 13708 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 14076 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 13984 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 13800 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 13984 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[28\].cc_clkbuf
timestamp 1693170804
transform 1 0 12880 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[28\].rs_mbuf
timestamp 1693170804
transform 1 0 11040 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5152 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 5888 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 11316 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 12788 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 13064 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 11040 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[29\].cc_clkbuf
timestamp 1693170804
transform 1 0 10304 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[29\].rs_mbuf
timestamp 1693170804
transform 1 0 11040 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 3588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[30\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 10212 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 10580 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 10120 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11500 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[30\].cc_clkbuf
timestamp 1693170804
transform 1 0 10948 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[30\].rs_mbuf
timestamp 1693170804
transform 1 0 9568 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 7728 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 6164 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 10212 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 8004 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8004 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 6716 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8096 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[31\].cc_clkbuf
timestamp 1693170804
transform 1 0 8464 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[31\].rs_mbuf
timestamp 1693170804
transform 1 0 8372 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[32\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16928 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[32\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 3588 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 5980 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 1196 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[32\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 5888 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[32\].cc_clkbuf
timestamp 1693170804
transform 1 0 7728 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[32\].rs_mbuf
timestamp 1693170804
transform 1 0 8372 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 2392 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 21528 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 17112 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 12880 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 17480 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 4876 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[33\].cc_clkbuf
timestamp 1693170804
transform 1 0 8372 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[33\].rs_mbuf
timestamp 1693170804
transform 1 0 4232 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 21804 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 17204 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 5980 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 5152 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10488 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 17388 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 16376 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[34\].cc_clkbuf
timestamp 1693170804
transform 1 0 8924 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[34\].rs_mbuf
timestamp 1693170804
transform 1 0 1472 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 3864 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 4140 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 2392 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 2024 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 828 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[35\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 12604 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[35\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[35\].cc_clkbuf
timestamp 1693170804
transform 1 0 3220 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[35\].rs_mbuf
timestamp 1693170804
transform 1 0 1656 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8188 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 5152 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 6440 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 6164 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 8832 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 8280 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 9108 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10396 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[36\].cc_clkbuf
timestamp 1693170804
transform 1 0 4600 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[36\].rs_mbuf
timestamp 1693170804
transform 1 0 7728 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 14352 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 14076 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 15732 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 17572 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 14352 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 15732 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11316 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11408 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11132 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10672 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[37\].cc_clkbuf
timestamp 1693170804
transform 1 0 9752 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[37\].rs_mbuf
timestamp 1693170804
transform 1 0 13524 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 14628 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 15732 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 10948 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 10948 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 10764 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10304 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[38\].cc_clkbuf
timestamp 1693170804
transform 1 0 11684 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[38\].rs_mbuf
timestamp 1693170804
transform 1 0 15732 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 12420 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 12420 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 12880 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 12420 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 12788 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 12144 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 12604 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 9476 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 9384 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[39\].cc_clkbuf
timestamp 1693170804
transform 1 0 11868 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[39\].rs_mbuf
timestamp 1693170804
transform 1 0 14628 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 9660 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 11500 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 9660 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 10212 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 9660 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 9660 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 7544 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 7268 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[40\].cc_clkbuf
timestamp 1693170804
transform 1 0 9476 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[40\].rs_mbuf
timestamp 1693170804
transform 1 0 8832 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 6532 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6808 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 7728 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6808 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6808 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 8740 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 9016 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[41\].cc_clkbuf
timestamp 1693170804
transform 1 0 6256 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[41\].rs_mbuf
timestamp 1693170804
transform 1 0 5888 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 6072 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 3588 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 3312 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 4232 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 4600 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3588 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 5152 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[42\].cc_clkbuf
timestamp 1693170804
transform 1 0 4600 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[42\].rs_mbuf
timestamp 1693170804
transform 1 0 3680 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 1472 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 3588 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 1472 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 1104 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[43\].cc_clkbuf
timestamp 1693170804
transform 1 0 920 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[43\].rs_mbuf
timestamp 1693170804
transform 1 0 1656 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dlclkp_4  ct.ro.cc_clock_gate $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 22172 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_4  ct.ro.cc_clock_inv $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 30176 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  ct.ro.cc_ring_osc_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 21252 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  ct.ro.cc_ring_osc_1
timestamp 1693170804
transform 1 0 25760 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  ct.ro.cc_ring_osc_2
timestamp 1693170804
transform 1 0 23092 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[1\].cc_div_flop $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 18952 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[2\].cc_div_flop
timestamp 1693170804
transform 1 0 19228 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[3\].cc_div_flop
timestamp 1693170804
transform 1 0 21252 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[4\].cc_div_flop
timestamp 1693170804
transform 1 0 23460 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[5\].cc_div_flop
timestamp 1693170804
transform 1 0 22080 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[6\].cc_div_flop
timestamp 1693170804
transform 1 0 21528 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[7\].cc_div_flop
timestamp 1693170804
transform 1 0 23828 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2i_2  cw.cc_test_0
timestamp 1693170804
transform 1 0 19688 0 -1 20128
box -38 -48 1050 592
use sky130_ht_sc_tt05__mux2i_2  cw.cc_test_1
timestamp 1699029708
transform 1 0 20056 0 -1 19040
box -38 -48 1050 592
use sky130_fd_sc_hd__maj3_2  cw.cc_test_2
timestamp 1693170804
transform 1 0 16100 0 -1 17952
box -38 -48 866 592
use sky130_ht_sc_tt05__maj3_2  cw.cc_test_3
timestamp 1699029708
transform 1 0 13524 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dlrtp_1  cw.cc_test_4
timestamp 1693170804
transform 1 0 4048 0 1 19040
box -38 -48 1234 592
use sky130_ht_sc_tt05__dlrtp_1  cw.cc_test_5
timestamp 1699029708
transform 1 0 18676 0 1 17952
box -38 -48 1418 592
use sky130_fd_sc_hd__dfrtp_1  cw.cc_test_6
timestamp 1693170804
transform 1 0 16100 0 -1 20128
box -38 -48 1878 592
use sky130_ht_sc_tt05__dfrtp_1  cw.cc_test_7
timestamp 1699029708
transform 1 0 16100 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  fanout5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 7912 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 12236 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout7
timestamp 1693170804
transform 1 0 10948 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout8
timestamp 1693170804
transform 1 0 28980 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout9
timestamp 1693170804
transform 1 0 30084 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout10
timestamp 1693170804
transform 1 0 9016 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout11
timestamp 1693170804
transform 1 0 13156 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout12
timestamp 1693170804
transform 1 0 10672 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 1693170804
transform 1 0 29532 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1693170804
transform 1 0 29532 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout15
timestamp 1693170804
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 1693170804
transform 1 0 12972 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout17
timestamp 1693170804
transform 1 0 10948 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 1693170804
transform 1 0 30084 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout19
timestamp 1693170804
transform 1 0 29532 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout20
timestamp 1693170804
transform 1 0 30084 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout21
timestamp 1693170804
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout22
timestamp 1693170804
transform 1 0 13064 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1693170804
transform 1 0 13616 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 1693170804
transform 1 0 30084 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout25
timestamp 1693170804
transform 1 0 28336 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp 1693170804
transform 1 0 17204 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1693170804
transform 1 0 16100 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout28
timestamp 1693170804
transform 1 0 15732 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1693170804
transform 1 0 28612 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout30
timestamp 1693170804
transform 1 0 27232 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout31
timestamp 1693170804
transform 1 0 29992 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout32
timestamp 1693170804
transform 1 0 16652 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 1693170804
transform 1 0 5796 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp 1693170804
transform 1 0 10856 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout35
timestamp 1693170804
transform 1 0 28980 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1693170804
transform 1 0 26496 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout37
timestamp 1693170804
transform 1 0 16100 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 1693170804
transform 1 0 15272 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout39
timestamp 1693170804
transform 1 0 14168 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout40
timestamp 1693170804
transform 1 0 29532 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 1693170804
transform 1 0 28244 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 1693170804
transform 1 0 30176 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp 1693170804
transform 1 0 16560 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 1693170804
transform 1 0 16468 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout45
timestamp 1693170804
transform 1 0 14076 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1693170804
transform 1 0 26404 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 1693170804
transform 1 0 26312 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp 1693170804
transform 1 0 27600 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1693170804
transform 1 0 12328 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp 1693170804
transform 1 0 13156 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 1693170804
transform 1 0 7728 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout52
timestamp 1693170804
transform 1 0 28980 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout53
timestamp 1693170804
transform 1 0 25668 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 1693170804
transform 1 0 23368 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 828 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_32
timestamp 1693170804
transform 1 0 3496 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4416 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_46
timestamp 1693170804
transform 1 0 4784 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1693170804
transform 1 0 10948 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_117
timestamp 1693170804
transform 1 0 11316 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_121
timestamp 1693170804
transform 1 0 11684 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_125
timestamp 1693170804
transform 1 0 12052 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_129 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 12420 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_312
timestamp 1693170804
transform 1 0 29256 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_316
timestamp 1693170804
transform 1 0 29624 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_320
timestamp 1693170804
transform 1 0 29992 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_324
timestamp 1693170804
transform 1 0 30360 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 1693170804
transform 1 0 828 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1693170804
transform 1 0 5796 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_119
timestamp 1693170804
transform 1 0 11500 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1693170804
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_255
timestamp 1693170804
transform 1 0 24012 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_287
timestamp 1693170804
transform 1 0 26956 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_318
timestamp 1693170804
transform 1 0 29808 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_322
timestamp 1693170804
transform 1 0 30176 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_326
timestamp 1693170804
transform 1 0 30544 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 1693170804
transform 1 0 828 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_32
timestamp 1693170804
transform 1 0 3496 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_91
timestamp 1693170804
transform 1 0 8924 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 1693170804
transform 1 0 13524 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1693170804
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_277
timestamp 1693170804
transform 1 0 26036 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_303
timestamp 1693170804
transform 1 0 28428 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_312 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 29256 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_318
timestamp 1693170804
transform 1 0 29808 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_322
timestamp 1693170804
transform 1 0 30176 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_326
timestamp 1693170804
transform 1 0 30544 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_3
timestamp 1693170804
transform 1 0 828 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_7
timestamp 1693170804
transform 1 0 1196 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_57
timestamp 1693170804
transform 1 0 5796 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_113
timestamp 1693170804
transform 1 0 10948 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_217
timestamp 1693170804
transform 1 0 20516 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_255
timestamp 1693170804
transform 1 0 24012 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_287
timestamp 1693170804
transform 1 0 26956 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_296
timestamp 1693170804
transform 1 0 27784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_322
timestamp 1693170804
transform 1 0 30176 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_326
timestamp 1693170804
transform 1 0 30544 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_3
timestamp 1693170804
transform 1 0 828 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_32
timestamp 1693170804
transform 1 0 3496 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1693170804
transform 1 0 8372 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_144
timestamp 1693170804
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1693170804
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_245
timestamp 1693170804
transform 1 0 23092 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1693170804
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_319
timestamp 1693170804
transform 1 0 29900 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_324
timestamp 1693170804
transform 1 0 30360 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_3
timestamp 1693170804
transform 1 0 828 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_57
timestamp 1693170804
transform 1 0 5796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_83
timestamp 1693170804
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp 1693170804
transform 1 0 10948 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1693170804
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_234
timestamp 1693170804
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_260
timestamp 1693170804
transform 1 0 24472 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_275
timestamp 1693170804
transform 1 0 25852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1693170804
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_290
timestamp 1693170804
transform 1 0 27232 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_297
timestamp 1693170804
transform 1 0 27876 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_322
timestamp 1693170804
transform 1 0 30176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_326
timestamp 1693170804
transform 1 0 30544 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1693170804
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 1693170804
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_33
timestamp 1693170804
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1693170804
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_97
timestamp 1693170804
transform 1 0 9476 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_141
timestamp 1693170804
transform 1 0 13524 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_146
timestamp 1693170804
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_239
timestamp 1693170804
transform 1 0 22540 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1693170804
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_257
timestamp 1693170804
transform 1 0 24196 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_312 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 29256 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_320
timestamp 1693170804
transform 1 0 29992 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_324
timestamp 1693170804
transform 1 0 30360 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_3
timestamp 1693170804
transform 1 0 828 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_108
timestamp 1693170804
transform 1 0 10488 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1693170804
transform 1 0 10948 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_169
timestamp 1693170804
transform 1 0 16100 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_258
timestamp 1693170804
transform 1 0 24288 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_263 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 24748 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_275
timestamp 1693170804
transform 1 0 25852 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1693170804
transform 1 0 26220 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_287
timestamp 1693170804
transform 1 0 26956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_291
timestamp 1693170804
transform 1 0 27324 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_321
timestamp 1693170804
transform 1 0 30084 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1693170804
transform 1 0 828 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_35
timestamp 1693170804
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_91
timestamp 1693170804
transform 1 0 8924 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_141
timestamp 1693170804
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_194
timestamp 1693170804
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1693170804
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_253
timestamp 1693170804
transform 1 0 23828 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_282
timestamp 1693170804
transform 1 0 26496 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_315
timestamp 1693170804
transform 1 0 29532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_3
timestamp 1693170804
transform 1 0 828 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_7
timestamp 1693170804
transform 1 0 1196 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_108
timestamp 1693170804
transform 1 0 10488 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_119
timestamp 1693170804
transform 1 0 11500 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_169
timestamp 1693170804
transform 1 0 16100 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1693170804
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_315
timestamp 1693170804
transform 1 0 29532 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 1693170804
transform 1 0 828 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_53
timestamp 1693170804
transform 1 0 5428 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1693170804
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_174
timestamp 1693170804
transform 1 0 16560 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_248
timestamp 1693170804
transform 1 0 23368 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_253
timestamp 1693170804
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_279
timestamp 1693170804
transform 1 0 26220 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1693170804
transform 1 0 28980 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_321
timestamp 1693170804
transform 1 0 30084 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_3
timestamp 1693170804
transform 1 0 828 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_46
timestamp 1693170804
transform 1 0 4784 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_81
timestamp 1693170804
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1693170804
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 1693170804
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_142
timestamp 1693170804
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1693170804
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_225
timestamp 1693170804
transform 1 0 21252 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_233
timestamp 1693170804
transform 1 0 21988 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_287
timestamp 1693170804
transform 1 0 26956 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_319
timestamp 1693170804
transform 1 0 29900 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 1693170804
transform 1 0 828 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_53
timestamp 1693170804
transform 1 0 5428 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_109
timestamp 1693170804
transform 1 0 10580 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_186
timestamp 1693170804
transform 1 0 17664 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_221
timestamp 1693170804
transform 1 0 20884 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_253
timestamp 1693170804
transform 1 0 23828 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1693170804
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_315
timestamp 1693170804
transform 1 0 29532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_6
timestamp 1693170804
transform 1 0 1104 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_10
timestamp 1693170804
transform 1 0 1472 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_18
timestamp 1693170804
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1693170804
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_116
timestamp 1693170804
transform 1 0 11224 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_188
timestamp 1693170804
transform 1 0 17848 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_214
timestamp 1693170804
transform 1 0 20240 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_218
timestamp 1693170804
transform 1 0 20608 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1693170804
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_281
timestamp 1693170804
transform 1 0 26404 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_289
timestamp 1693170804
transform 1 0 27140 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_319
timestamp 1693170804
transform 1 0 29900 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 1693170804
transform 1 0 828 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_53
timestamp 1693170804
transform 1 0 5428 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_88
timestamp 1693170804
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_96
timestamp 1693170804
transform 1 0 9384 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1693170804
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_221
timestamp 1693170804
transform 1 0 20884 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_227
timestamp 1693170804
transform 1 0 21436 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_280
timestamp 1693170804
transform 1 0 26312 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_325
timestamp 1693170804
transform 1 0 30452 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_3
timestamp 1693170804
transform 1 0 828 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_10
timestamp 1693170804
transform 1 0 1472 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_18
timestamp 1693170804
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_60
timestamp 1693170804
transform 1 0 6072 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1693170804
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_173
timestamp 1693170804
transform 1 0 16468 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_207
timestamp 1693170804
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_211
timestamp 1693170804
transform 1 0 19964 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_221
timestamp 1693170804
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_228
timestamp 1693170804
transform 1 0 21528 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_232
timestamp 1693170804
transform 1 0 21896 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_236
timestamp 1693170804
transform 1 0 22264 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1693170804
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 1693170804
transform 1 0 828 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_29
timestamp 1693170804
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 1693170804
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1693170804
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_171
timestamp 1693170804
transform 1 0 16284 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_245
timestamp 1693170804
transform 1 0 23092 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1693170804
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_312
timestamp 1693170804
transform 1 0 29256 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_326
timestamp 1693170804
transform 1 0 30544 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1693170804
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1693170804
transform 1 0 5796 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_172
timestamp 1693170804
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_210
timestamp 1693170804
transform 1 0 19872 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_214
timestamp 1693170804
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_218
timestamp 1693170804
transform 1 0 20608 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_252
timestamp 1693170804
transform 1 0 23736 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_3
timestamp 1693170804
transform 1 0 828 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_53
timestamp 1693170804
transform 1 0 5428 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_78
timestamp 1693170804
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_89
timestamp 1693170804
transform 1 0 8740 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_132
timestamp 1693170804
transform 1 0 12696 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_136
timestamp 1693170804
transform 1 0 13064 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_165
timestamp 1693170804
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_169
timestamp 1693170804
transform 1 0 16100 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_259
timestamp 1693170804
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_304
timestamp 1693170804
transform 1 0 28520 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_325
timestamp 1693170804
transform 1 0 30452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 1693170804
transform 1 0 828 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_7
timestamp 1693170804
transform 1 0 1196 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_43
timestamp 1693170804
transform 1 0 4508 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_60
timestamp 1693170804
transform 1 0 6072 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_96
timestamp 1693170804
transform 1 0 9384 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_103
timestamp 1693170804
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1693170804
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_125
timestamp 1693170804
transform 1 0 12052 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_159
timestamp 1693170804
transform 1 0 15180 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_163
timestamp 1693170804
transform 1 0 15548 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1693170804
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_169
timestamp 1693170804
transform 1 0 16100 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_173
timestamp 1693170804
transform 1 0 16468 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_228
timestamp 1693170804
transform 1 0 21528 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_278
timestamp 1693170804
transform 1 0 26128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_3
timestamp 1693170804
transform 1 0 828 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_29
timestamp 1693170804
transform 1 0 3220 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_97
timestamp 1693170804
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_126
timestamp 1693170804
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_130
timestamp 1693170804
transform 1 0 12512 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_165
timestamp 1693170804
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_221
timestamp 1693170804
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_225
timestamp 1693170804
transform 1 0 21252 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_253
timestamp 1693170804
transform 1 0 23828 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1693170804
transform 1 0 828 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_63
timestamp 1693170804
transform 1 0 6348 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_125
timestamp 1693170804
transform 1 0 12052 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_159
timestamp 1693170804
transform 1 0 15180 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_163
timestamp 1693170804
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1693170804
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_169
timestamp 1693170804
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_173
timestamp 1693170804
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_177
timestamp 1693170804
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_182
timestamp 1693170804
transform 1 0 17296 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_213
timestamp 1693170804
transform 1 0 20148 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_217
timestamp 1693170804
transform 1 0 20516 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 1693170804
transform 1 0 20976 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1693170804
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_3
timestamp 1693170804
transform 1 0 828 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_32
timestamp 1693170804
transform 1 0 3496 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_98
timestamp 1693170804
transform 1 0 9568 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_129
timestamp 1693170804
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_165
timestamp 1693170804
transform 1 0 15732 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_169
timestamp 1693170804
transform 1 0 16100 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_197
timestamp 1693170804
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_238
timestamp 1693170804
transform 1 0 22448 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_244
timestamp 1693170804
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1693170804
transform 1 0 28796 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_322
timestamp 1693170804
transform 1 0 30176 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp 1693170804
transform 1 0 828 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_63
timestamp 1693170804
transform 1 0 6348 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1693170804
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_128
timestamp 1693170804
transform 1 0 12328 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_153
timestamp 1693170804
transform 1 0 14628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 1693170804
transform 1 0 15824 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_172
timestamp 1693170804
transform 1 0 16376 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_177
timestamp 1693170804
transform 1 0 16836 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_204
timestamp 1693170804
transform 1 0 19320 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_231
timestamp 1693170804
transform 1 0 21804 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_3
timestamp 1693170804
transform 1 0 828 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_29
timestamp 1693170804
transform 1 0 3220 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_97
timestamp 1693170804
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1693170804
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1693170804
transform 1 0 13524 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_209
timestamp 1693170804
transform 1 0 19780 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_247
timestamp 1693170804
transform 1 0 23276 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_259
timestamp 1693170804
transform 1 0 24380 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_3
timestamp 1693170804
transform 1 0 828 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_34
timestamp 1693170804
transform 1 0 3680 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_57
timestamp 1693170804
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_92
timestamp 1693170804
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1693170804
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_113
timestamp 1693170804
transform 1 0 10948 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_173
timestamp 1693170804
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_199
timestamp 1693170804
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_203
timestamp 1693170804
transform 1 0 19228 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_225
timestamp 1693170804
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_296
timestamp 1693170804
transform 1 0 27784 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_325
timestamp 1693170804
transform 1 0 30452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_3
timestamp 1693170804
transform 1 0 828 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_59
timestamp 1693170804
transform 1 0 5980 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_112
timestamp 1693170804
transform 1 0 10856 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_151
timestamp 1693170804
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_206
timestamp 1693170804
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_232
timestamp 1693170804
transform 1 0 21896 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_325
timestamp 1693170804
transform 1 0 30452 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_6
timestamp 1693170804
transform 1 0 1104 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_63
timestamp 1693170804
transform 1 0 6348 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_113
timestamp 1693170804
transform 1 0 10948 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_175
timestamp 1693170804
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_204
timestamp 1693170804
transform 1 0 19320 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1693170804
transform 1 0 26220 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_281
timestamp 1693170804
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_292
timestamp 1693170804
transform 1 0 27416 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_326
timestamp 1693170804
transform 1 0 30544 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_3
timestamp 1693170804
transform 1 0 828 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_59
timestamp 1693170804
transform 1 0 5980 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_112
timestamp 1693170804
transform 1 0 10856 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1693170804
transform 1 0 13524 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_176
timestamp 1693170804
transform 1 0 16744 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1693170804
transform 1 0 23552 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_3
timestamp 1693170804
transform 1 0 828 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_31
timestamp 1693170804
transform 1 0 3404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_81
timestamp 1693170804
transform 1 0 8004 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_119
timestamp 1693170804
transform 1 0 11500 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_172
timestamp 1693170804
transform 1 0 16376 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_255
timestamp 1693170804
transform 1 0 24012 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_3
timestamp 1693170804
transform 1 0 828 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_29
timestamp 1693170804
transform 1 0 3220 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_54
timestamp 1693170804
transform 1 0 5520 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_150
timestamp 1693170804
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_171
timestamp 1693170804
transform 1 0 16284 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_253
timestamp 1693170804
transform 1 0 23828 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_3
timestamp 1693170804
transform 1 0 828 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_7
timestamp 1693170804
transform 1 0 1196 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_63
timestamp 1693170804
transform 1 0 6348 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_143
timestamp 1693170804
transform 1 0 13708 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_249
timestamp 1693170804
transform 1 0 23460 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_325
timestamp 1693170804
transform 1 0 30452 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_3
timestamp 1693170804
transform 1 0 828 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_35
timestamp 1693170804
transform 1 0 3772 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 1693170804
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_135
timestamp 1693170804
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_141
timestamp 1693170804
transform 1 0 13524 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_168
timestamp 1693170804
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_172
timestamp 1693170804
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1693170804
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_3
timestamp 1693170804
transform 1 0 828 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_57
timestamp 1693170804
transform 1 0 5796 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_137
timestamp 1693170804
transform 1 0 13156 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1693170804
transform 1 0 21068 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_326
timestamp 1693170804
transform 1 0 30544 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_109
timestamp 1693170804
transform 1 0 10580 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_141
timestamp 1693170804
transform 1 0 13524 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_145
timestamp 1693170804
transform 1 0 13892 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_149
timestamp 1693170804
transform 1 0 14260 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_152
timestamp 1693170804
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_159
timestamp 1693170804
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_163
timestamp 1693170804
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_259
timestamp 1693170804
transform 1 0 24380 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_3
timestamp 1693170804
transform 1 0 828 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_61
timestamp 1693170804
transform 1 0 6164 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_65
timestamp 1693170804
transform 1 0 6532 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_110
timestamp 1693170804
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_219
timestamp 1693170804
transform 1 0 20700 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_3
timestamp 1693170804
transform 1 0 828 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_29
timestamp 1693170804
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_33
timestamp 1693170804
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_37
timestamp 1693170804
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_50
timestamp 1693170804
transform 1 0 5152 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_85
timestamp 1693170804
transform 1 0 8372 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_189
timestamp 1693170804
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_227
timestamp 1693170804
transform 1 0 21436 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_283
timestamp 1693170804
transform 1 0 26588 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_326
timestamp 1693170804
transform 1 0 30544 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_3
timestamp 1693170804
transform 1 0 828 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_105
timestamp 1693170804
transform 1 0 10212 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_164
timestamp 1693170804
transform 1 0 15640 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_193
timestamp 1693170804
transform 1 0 18308 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1693170804
transform 1 0 26220 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_3
timestamp 1693170804
transform 1 0 828 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 1693170804
transform 1 0 18400 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_222
timestamp 1693170804
transform 1 0 20976 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_279
timestamp 1693170804
transform 1 0 26220 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 1693170804
transform 1 0 28704 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1693170804
transform 1 0 30360 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1693170804
transform 1 0 30360 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1693170804
transform 1 0 30084 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1693170804
transform 1 0 15732 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_39
timestamp 1693170804
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1693170804
transform -1 0 30912 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_40
timestamp 1693170804
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1693170804
transform -1 0 30912 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_41
timestamp 1693170804
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1693170804
transform -1 0 30912 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_42
timestamp 1693170804
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1693170804
transform -1 0 30912 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_43
timestamp 1693170804
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1693170804
transform -1 0 30912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_44
timestamp 1693170804
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1693170804
transform -1 0 30912 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_45
timestamp 1693170804
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1693170804
transform -1 0 30912 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_46
timestamp 1693170804
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1693170804
transform -1 0 30912 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_47
timestamp 1693170804
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1693170804
transform -1 0 30912 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_48
timestamp 1693170804
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1693170804
transform -1 0 30912 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_49
timestamp 1693170804
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1693170804
transform -1 0 30912 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_50
timestamp 1693170804
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1693170804
transform -1 0 30912 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_51
timestamp 1693170804
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1693170804
transform -1 0 30912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_52
timestamp 1693170804
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1693170804
transform -1 0 30912 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_53
timestamp 1693170804
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1693170804
transform -1 0 30912 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_54
timestamp 1693170804
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1693170804
transform -1 0 30912 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_55
timestamp 1693170804
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1693170804
transform -1 0 30912 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_56
timestamp 1693170804
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1693170804
transform -1 0 30912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_57
timestamp 1693170804
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1693170804
transform -1 0 30912 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_58
timestamp 1693170804
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1693170804
transform -1 0 30912 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_59
timestamp 1693170804
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1693170804
transform -1 0 30912 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_60
timestamp 1693170804
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1693170804
transform -1 0 30912 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_61
timestamp 1693170804
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1693170804
transform -1 0 30912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_62
timestamp 1693170804
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1693170804
transform -1 0 30912 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_63
timestamp 1693170804
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1693170804
transform -1 0 30912 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_64
timestamp 1693170804
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1693170804
transform -1 0 30912 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_65
timestamp 1693170804
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1693170804
transform -1 0 30912 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_66
timestamp 1693170804
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1693170804
transform -1 0 30912 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_67
timestamp 1693170804
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1693170804
transform -1 0 30912 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_68
timestamp 1693170804
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1693170804
transform -1 0 30912 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_69
timestamp 1693170804
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1693170804
transform -1 0 30912 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_70
timestamp 1693170804
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1693170804
transform -1 0 30912 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_71
timestamp 1693170804
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1693170804
transform -1 0 30912 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_72
timestamp 1693170804
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1693170804
transform -1 0 30912 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_73
timestamp 1693170804
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1693170804
transform -1 0 30912 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_74
timestamp 1693170804
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1693170804
transform -1 0 30912 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_75
timestamp 1693170804
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1693170804
transform -1 0 30912 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_76
timestamp 1693170804
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1693170804
transform -1 0 30912 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_77
timestamp 1693170804
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1693170804
transform -1 0 30912 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp 1693170804
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp 1693170804
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_81
timestamp 1693170804
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82
timestamp 1693170804
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_83
timestamp 1693170804
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 1693170804
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1693170804
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1693170804
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1693170804
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1693170804
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_89
timestamp 1693170804
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_90
timestamp 1693170804
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_91
timestamp 1693170804
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1693170804
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1693170804
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_94
timestamp 1693170804
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_95
timestamp 1693170804
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1693170804
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1693170804
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1693170804
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1693170804
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1693170804
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1693170804
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1693170804
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1693170804
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_104
timestamp 1693170804
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1693170804
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1693170804
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1693170804
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_108
timestamp 1693170804
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_109
timestamp 1693170804
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_110
timestamp 1693170804
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1693170804
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_112
timestamp 1693170804
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_113
timestamp 1693170804
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_114
timestamp 1693170804
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_115
timestamp 1693170804
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_116
timestamp 1693170804
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_117
timestamp 1693170804
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_118
timestamp 1693170804
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_119
timestamp 1693170804
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_120
timestamp 1693170804
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_121
timestamp 1693170804
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_122
timestamp 1693170804
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_123
timestamp 1693170804
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_124
timestamp 1693170804
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_125
timestamp 1693170804
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_126
timestamp 1693170804
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_127
timestamp 1693170804
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_128
timestamp 1693170804
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_129
timestamp 1693170804
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_130
timestamp 1693170804
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_131
timestamp 1693170804
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_132
timestamp 1693170804
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_133
timestamp 1693170804
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_134
timestamp 1693170804
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_135
timestamp 1693170804
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_136
timestamp 1693170804
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_137
timestamp 1693170804
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_138
timestamp 1693170804
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_139
timestamp 1693170804
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_140
timestamp 1693170804
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 1693170804
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_142
timestamp 1693170804
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 1693170804
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp 1693170804
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp 1693170804
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp 1693170804
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp 1693170804
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp 1693170804
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_149
timestamp 1693170804
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_150
timestamp 1693170804
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_151
timestamp 1693170804
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_152
timestamp 1693170804
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_153
timestamp 1693170804
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_154
timestamp 1693170804
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_155
timestamp 1693170804
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_156
timestamp 1693170804
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_157
timestamp 1693170804
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_158
timestamp 1693170804
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_159
timestamp 1693170804
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_160
timestamp 1693170804
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_161
timestamp 1693170804
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_162
timestamp 1693170804
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp 1693170804
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_164
timestamp 1693170804
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_165
timestamp 1693170804
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_166
timestamp 1693170804
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_167
timestamp 1693170804
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_168
timestamp 1693170804
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_169
timestamp 1693170804
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_170
timestamp 1693170804
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_171
timestamp 1693170804
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_172
timestamp 1693170804
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_173
timestamp 1693170804
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_174
timestamp 1693170804
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_175
timestamp 1693170804
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_176
timestamp 1693170804
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_177
timestamp 1693170804
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_178
timestamp 1693170804
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_179
timestamp 1693170804
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_180
timestamp 1693170804
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_181
timestamp 1693170804
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_182
timestamp 1693170804
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_183
timestamp 1693170804
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_184
timestamp 1693170804
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 1693170804
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_186
timestamp 1693170804
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_187
timestamp 1693170804
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_188
timestamp 1693170804
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_189
timestamp 1693170804
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_190
timestamp 1693170804
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_191
timestamp 1693170804
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_192
timestamp 1693170804
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_193
timestamp 1693170804
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_194
timestamp 1693170804
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_195
timestamp 1693170804
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_196
timestamp 1693170804
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_197
timestamp 1693170804
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_198
timestamp 1693170804
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_199
timestamp 1693170804
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_200
timestamp 1693170804
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_201
timestamp 1693170804
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_202
timestamp 1693170804
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_203
timestamp 1693170804
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_204
timestamp 1693170804
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_205
timestamp 1693170804
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_206
timestamp 1693170804
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_207
timestamp 1693170804
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_208
timestamp 1693170804
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp 1693170804
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_210
timestamp 1693170804
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_211
timestamp 1693170804
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_212
timestamp 1693170804
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_213
timestamp 1693170804
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp 1693170804
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_215
timestamp 1693170804
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_216
timestamp 1693170804
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_217
timestamp 1693170804
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_218
timestamp 1693170804
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp 1693170804
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp 1693170804
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_221
timestamp 1693170804
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_222
timestamp 1693170804
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_223
timestamp 1693170804
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp 1693170804
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp 1693170804
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_226
timestamp 1693170804
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_227
timestamp 1693170804
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_228
timestamp 1693170804
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp 1693170804
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp 1693170804
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp 1693170804
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_232
timestamp 1693170804
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_233
timestamp 1693170804
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp 1693170804
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp 1693170804
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp 1693170804
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_237
timestamp 1693170804
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_238
timestamp 1693170804
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp 1693170804
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp 1693170804
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp 1693170804
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp 1693170804
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_243
timestamp 1693170804
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp 1693170804
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp 1693170804
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp 1693170804
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp 1693170804
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_248
timestamp 1693170804
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp 1693170804
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp 1693170804
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp 1693170804
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp 1693170804
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 1693170804
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp 1693170804
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp 1693170804
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp 1693170804
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp 1693170804
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 1693170804
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp 1693170804
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp 1693170804
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp 1693170804
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp 1693170804
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 1693170804
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 1693170804
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1693170804
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp 1693170804
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp 1693170804
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 1693170804
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 1693170804
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp 1693170804
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp 1693170804
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp 1693170804
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 1693170804
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 1693170804
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1693170804
transform 1 0 28888 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp 1693170804
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp 1693170804
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 1693170804
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 1693170804
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1693170804
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp 1693170804
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp 1693170804
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 1693170804
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 1693170804
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1693170804
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 1693170804
transform 1 0 28888 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp 1693170804
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 1693170804
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 1693170804
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1693170804
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 1693170804
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp 1693170804
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 1693170804
transform 1 0 5704 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 1693170804
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1693170804
transform 1 0 10856 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 1693170804
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 1693170804
transform 1 0 16008 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_298
timestamp 1693170804
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp 1693170804
transform 1 0 21160 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_300
timestamp 1693170804
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp 1693170804
transform 1 0 26312 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_302
timestamp 1693170804
transform 1 0 28888 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 13524 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_56
timestamp 1693170804
transform 1 0 9200 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_57
timestamp 1693170804
transform 1 0 9016 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_58
timestamp 1693170804
transform 1 0 9568 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_59
timestamp 1693170804
transform 1 0 9292 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_60
timestamp 1693170804
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_61
timestamp 1693170804
transform 1 0 11224 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_62
timestamp 1693170804
transform 1 0 11500 0 -1 13600
box -38 -48 314 592
<< labels >>
flabel metal4 s 7982 496 8302 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15572 496 15892 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 23162 496 23482 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 30752 496 31072 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4187 496 4507 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11777 496 12097 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19367 496 19687 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26957 496 27277 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26926 22104 26986 22304 0 FreeSans 480 90 0 0 clk
port 2 nsew signal input
flabel metal4 s 27478 22104 27538 22304 0 FreeSans 480 90 0 0 ena
port 3 nsew signal input
flabel metal4 s 26374 22104 26434 22304 0 FreeSans 480 90 0 0 rst_n
port 4 nsew signal input
flabel metal4 s 25822 22104 25882 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 5 nsew signal input
flabel metal4 s 25270 22104 25330 22304 0 FreeSans 480 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal4 s 24718 22104 24778 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal4 s 24166 22104 24226 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal4 s 23614 22104 23674 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal4 s 23062 22104 23122 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal4 s 22510 22104 22570 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal4 s 21958 22104 22018 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal4 s 21406 22104 21466 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal4 s 20854 22104 20914 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal4 s 20302 22104 20362 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal4 s 19750 22104 19810 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal4 s 19198 22104 19258 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal4 s 18646 22104 18706 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal4 s 18094 22104 18154 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal4 s 17542 22104 17602 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal4 s 8158 22104 8218 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 21 nsew signal tristate
flabel metal4 s 7606 22104 7666 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 22 nsew signal tristate
flabel metal4 s 7054 22104 7114 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 23 nsew signal tristate
flabel metal4 s 6502 22104 6562 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 24 nsew signal tristate
flabel metal4 s 5950 22104 6010 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 25 nsew signal tristate
flabel metal4 s 5398 22104 5458 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 26 nsew signal tristate
flabel metal4 s 4846 22104 4906 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 27 nsew signal tristate
flabel metal4 s 4294 22104 4354 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 28 nsew signal tristate
flabel metal4 s 12574 22104 12634 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 29 nsew signal tristate
flabel metal4 s 12022 22104 12082 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 30 nsew signal tristate
flabel metal4 s 11470 22104 11530 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 31 nsew signal tristate
flabel metal4 s 10918 22104 10978 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 32 nsew signal tristate
flabel metal4 s 10366 22104 10426 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 33 nsew signal tristate
flabel metal4 s 9814 22104 9874 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 34 nsew signal tristate
flabel metal4 s 9262 22104 9322 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 35 nsew signal tristate
flabel metal4 s 8710 22104 8770 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 36 nsew signal tristate
flabel metal4 s 16990 22104 17050 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 37 nsew signal tristate
flabel metal4 s 16438 22104 16498 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 38 nsew signal tristate
flabel metal4 s 15886 22104 15946 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 39 nsew signal tristate
flabel metal4 s 15334 22104 15394 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 40 nsew signal tristate
flabel metal4 s 14782 22104 14842 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 41 nsew signal tristate
flabel metal4 s 14230 22104 14290 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 42 nsew signal tristate
flabel metal4 s 13678 22104 13738 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 43 nsew signal tristate
flabel metal4 s 13126 22104 13186 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 44 nsew signal tristate
rlabel via1 15812 21216 15812 21216 0 VGND
rlabel metal1 15732 21760 15732 21760 0 VPWR
rlabel metal1 18998 20808 18998 20808 0 _00_
rlabel metal1 23230 18938 23230 18938 0 _01_
rlabel metal1 24610 18938 24610 18938 0 _02_
rlabel metal1 23000 18666 23000 18666 0 _03_
rlabel metal2 18538 20672 18538 20672 0 _04_
rlabel metal1 29440 20366 29440 20366 0 ct.cw.source\[0\]
rlabel metal1 29716 19346 29716 19346 0 ct.cw.source\[1\]
rlabel metal1 17112 17306 17112 17306 0 ct.cw.source\[2\]
rlabel metal2 1978 11169 1978 11169 0 ct.cw.target\[0\]
rlabel via2 2254 13277 2254 13277 0 ct.cw.target\[1\]
rlabel metal2 1978 14433 1978 14433 0 ct.cw.target\[2\]
rlabel metal1 1840 8058 1840 8058 0 ct.cw.target\[3\]
rlabel metal3 14904 19652 14904 19652 0 ct.cw.target\[4\]
rlabel metal2 14260 18700 14260 18700 0 ct.cw.target\[5\]
rlabel metal1 15042 19346 15042 19346 0 ct.cw.target\[6\]
rlabel metal2 20332 13396 20332 13396 0 ct.cw.target\[7\]
rlabel metal1 29486 13158 29486 13158 0 ct.ic.data_chain\[10\]
rlabel metal2 21022 13702 21022 13702 0 ct.ic.data_chain\[11\]
rlabel metal2 7038 20655 7038 20655 0 ct.ic.data_chain\[12\]
rlabel metal1 27324 13158 27324 13158 0 ct.ic.data_chain\[13\]
rlabel metal1 20562 15538 20562 15538 0 ct.ic.data_chain\[14\]
rlabel metal2 2530 20621 2530 20621 0 ct.ic.data_chain\[15\]
rlabel metal1 21620 13294 21620 13294 0 ct.ic.data_chain\[16\]
rlabel metal1 18446 15096 18446 15096 0 ct.ic.data_chain\[17\]
rlabel metal1 828 19210 828 19210 0 ct.ic.data_chain\[18\]
rlabel metal1 19826 13294 19826 13294 0 ct.ic.data_chain\[19\]
rlabel via2 17158 15011 17158 15011 0 ct.ic.data_chain\[20\]
rlabel metal1 29302 18394 29302 18394 0 ct.ic.data_chain\[21\]
rlabel metal1 22034 21624 22034 21624 0 ct.ic.data_chain\[22\]
rlabel via2 21114 16643 21114 16643 0 ct.ic.data_chain\[23\]
rlabel metal1 26634 18258 26634 18258 0 ct.ic.data_chain\[24\]
rlabel metal1 21160 17510 21160 17510 0 ct.ic.data_chain\[25\]
rlabel metal1 19918 16626 19918 16626 0 ct.ic.data_chain\[26\]
rlabel metal1 21114 18802 21114 18802 0 ct.ic.data_chain\[27\]
rlabel metal1 19780 17714 19780 17714 0 ct.ic.data_chain\[28\]
rlabel metal2 22172 19380 22172 19380 0 ct.ic.data_chain\[29\]
rlabel metal1 18814 18802 18814 18802 0 ct.ic.data_chain\[30\]
rlabel metal1 18906 19278 18906 19278 0 ct.ic.data_chain\[31\]
rlabel metal2 18906 19975 18906 19975 0 ct.ic.data_chain\[32\]
rlabel metal1 19182 19822 19182 19822 0 ct.ic.data_chain\[33\]
rlabel metal2 19366 19295 19366 19295 0 ct.ic.data_chain\[34\]
rlabel metal1 15042 19890 15042 19890 0 ct.ic.data_chain\[35\]
rlabel metal1 29486 9010 29486 9010 0 ct.ic.data_chain\[3\]
rlabel metal3 20217 13804 20217 13804 0 ct.ic.data_chain\[4\]
rlabel metal1 14904 17102 14904 17102 0 ct.ic.data_chain\[5\]
rlabel metal2 30130 18564 30130 18564 0 ct.ic.data_chain\[6\]
rlabel metal2 28934 11084 28934 11084 0 ct.ic.data_chain\[7\]
rlabel metal1 17342 16014 17342 16014 0 ct.ic.data_chain\[8\]
rlabel metal2 26358 20927 26358 20927 0 ct.ic.data_chain\[9\]
rlabel metal1 28290 21488 28290 21488 0 ct.ic.trig_chain\[0\]
rlabel metal1 18998 20298 18998 20298 0 ct.ic.trig_chain\[10\]
rlabel metal1 14306 19788 14306 19788 0 ct.ic.trig_chain\[11\]
rlabel metal2 19366 21250 19366 21250 0 ct.ic.trig_chain\[12\]
rlabel metal1 19458 14348 19458 14348 0 ct.ic.trig_chain\[1\]
rlabel metal2 16882 15793 16882 15793 0 ct.ic.trig_chain\[2\]
rlabel metal1 27140 19822 27140 19822 0 ct.ic.trig_chain\[3\]
rlabel metal2 19274 15912 19274 15912 0 ct.ic.trig_chain\[4\]
rlabel metal1 25116 20774 25116 20774 0 ct.ic.trig_chain\[5\]
rlabel metal2 874 18785 874 18785 0 ct.ic.trig_chain\[6\]
rlabel metal3 20516 18360 20516 18360 0 ct.ic.trig_chain\[7\]
rlabel metal2 21206 16592 21206 16592 0 ct.ic.trig_chain\[8\]
rlabel metal1 18998 17714 18998 17714 0 ct.ic.trig_chain\[9\]
rlabel metal1 14628 18802 14628 18802 0 ct.oc.capture_buffer\[0\]
rlabel metal1 29716 20910 29716 20910 0 ct.oc.capture_buffer\[100\]
rlabel metal1 29946 20026 29946 20026 0 ct.oc.capture_buffer\[101\]
rlabel metal1 30130 14314 30130 14314 0 ct.oc.capture_buffer\[102\]
rlabel metal1 29946 18598 29946 18598 0 ct.oc.capture_buffer\[103\]
rlabel metal1 25668 13906 25668 13906 0 ct.oc.capture_buffer\[104\]
rlabel metal1 27094 13362 27094 13362 0 ct.oc.capture_buffer\[105\]
rlabel metal1 23046 12614 23046 12614 0 ct.oc.capture_buffer\[106\]
rlabel metal1 26772 12818 26772 12818 0 ct.oc.capture_buffer\[107\]
rlabel metal1 28290 14042 28290 14042 0 ct.oc.capture_buffer\[108\]
rlabel metal1 29210 14042 29210 14042 0 ct.oc.capture_buffer\[109\]
rlabel metal1 20930 19992 20930 19992 0 ct.oc.capture_buffer\[10\]
rlabel metal1 29394 19822 29394 19822 0 ct.oc.capture_buffer\[110\]
rlabel metal2 29854 15215 29854 15215 0 ct.oc.capture_buffer\[111\]
rlabel metal1 24288 12750 24288 12750 0 ct.oc.capture_buffer\[112\]
rlabel metal2 24886 13702 24886 13702 0 ct.oc.capture_buffer\[113\]
rlabel metal1 22448 12954 22448 12954 0 ct.oc.capture_buffer\[114\]
rlabel metal1 23828 12614 23828 12614 0 ct.oc.capture_buffer\[115\]
rlabel metal2 27186 12359 27186 12359 0 ct.oc.capture_buffer\[116\]
rlabel metal1 27968 11730 27968 11730 0 ct.oc.capture_buffer\[117\]
rlabel metal2 28750 13600 28750 13600 0 ct.oc.capture_buffer\[118\]
rlabel metal2 29946 13668 29946 13668 0 ct.oc.capture_buffer\[119\]
rlabel metal1 11270 21114 11270 21114 0 ct.oc.capture_buffer\[11\]
rlabel metal1 21712 12274 21712 12274 0 ct.oc.capture_buffer\[120\]
rlabel metal1 21160 13498 21160 13498 0 ct.oc.capture_buffer\[121\]
rlabel metal1 20516 12750 20516 12750 0 ct.oc.capture_buffer\[122\]
rlabel metal2 22310 11220 22310 11220 0 ct.oc.capture_buffer\[123\]
rlabel metal1 23690 9622 23690 9622 0 ct.oc.capture_buffer\[124\]
rlabel metal1 28198 8398 28198 8398 0 ct.oc.capture_buffer\[125\]
rlabel metal1 29394 6834 29394 6834 0 ct.oc.capture_buffer\[126\]
rlabel metal2 28474 9520 28474 9520 0 ct.oc.capture_buffer\[127\]
rlabel metal2 19274 10982 19274 10982 0 ct.oc.capture_buffer\[128\]
rlabel metal1 19274 12614 19274 12614 0 ct.oc.capture_buffer\[129\]
rlabel metal1 9522 14280 9522 14280 0 ct.oc.capture_buffer\[12\]
rlabel metal2 18906 12517 18906 12517 0 ct.oc.capture_buffer\[130\]
rlabel metal2 22034 10251 22034 10251 0 ct.oc.capture_buffer\[131\]
rlabel metal1 24288 10234 24288 10234 0 ct.oc.capture_buffer\[132\]
rlabel metal1 28060 9622 28060 9622 0 ct.oc.capture_buffer\[133\]
rlabel metal1 27646 8942 27646 8942 0 ct.oc.capture_buffer\[134\]
rlabel metal2 28290 9860 28290 9860 0 ct.oc.capture_buffer\[135\]
rlabel metal1 17572 10098 17572 10098 0 ct.oc.capture_buffer\[136\]
rlabel metal1 16836 11186 16836 11186 0 ct.oc.capture_buffer\[137\]
rlabel metal1 17112 11730 17112 11730 0 ct.oc.capture_buffer\[138\]
rlabel metal1 20148 10234 20148 10234 0 ct.oc.capture_buffer\[139\]
rlabel metal2 9522 21471 9522 21471 0 ct.oc.capture_buffer\[13\]
rlabel metal1 23552 10234 23552 10234 0 ct.oc.capture_buffer\[140\]
rlabel metal1 23184 9622 23184 9622 0 ct.oc.capture_buffer\[141\]
rlabel metal1 26266 8602 26266 8602 0 ct.oc.capture_buffer\[142\]
rlabel metal1 25990 9112 25990 9112 0 ct.oc.capture_buffer\[143\]
rlabel metal1 16882 9146 16882 9146 0 ct.oc.capture_buffer\[144\]
rlabel metal1 19274 9146 19274 9146 0 ct.oc.capture_buffer\[145\]
rlabel metal1 17296 9010 17296 9010 0 ct.oc.capture_buffer\[146\]
rlabel metal1 19412 8466 19412 8466 0 ct.oc.capture_buffer\[147\]
rlabel metal1 21482 9146 21482 9146 0 ct.oc.capture_buffer\[148\]
rlabel metal2 25714 9316 25714 9316 0 ct.oc.capture_buffer\[149\]
rlabel metal2 4554 20910 4554 20910 0 ct.oc.capture_buffer\[14\]
rlabel metal1 25024 8466 25024 8466 0 ct.oc.capture_buffer\[150\]
rlabel metal1 24426 8942 24426 8942 0 ct.oc.capture_buffer\[151\]
rlabel metal1 19136 6222 19136 6222 0 ct.oc.capture_buffer\[152\]
rlabel metal2 17802 7599 17802 7599 0 ct.oc.capture_buffer\[153\]
rlabel metal2 17802 7072 17802 7072 0 ct.oc.capture_buffer\[154\]
rlabel metal1 18446 6834 18446 6834 0 ct.oc.capture_buffer\[155\]
rlabel metal1 21620 7922 21620 7922 0 ct.oc.capture_buffer\[156\]
rlabel metal1 23138 7480 23138 7480 0 ct.oc.capture_buffer\[157\]
rlabel metal1 22264 8466 22264 8466 0 ct.oc.capture_buffer\[158\]
rlabel metal1 22264 7378 22264 7378 0 ct.oc.capture_buffer\[159\]
rlabel metal1 5934 11322 5934 11322 0 ct.oc.capture_buffer\[15\]
rlabel metal1 24610 6630 24610 6630 0 ct.oc.capture_buffer\[160\]
rlabel metal1 28612 4658 28612 4658 0 ct.oc.capture_buffer\[161\]
rlabel metal2 27462 7004 27462 7004 0 ct.oc.capture_buffer\[162\]
rlabel metal2 25714 6562 25714 6562 0 ct.oc.capture_buffer\[163\]
rlabel metal1 27508 5202 27508 5202 0 ct.oc.capture_buffer\[164\]
rlabel metal1 29256 2482 29256 2482 0 ct.oc.capture_buffer\[165\]
rlabel metal1 28796 3570 28796 3570 0 ct.oc.capture_buffer\[166\]
rlabel metal1 28934 4114 28934 4114 0 ct.oc.capture_buffer\[167\]
rlabel metal1 17480 12750 17480 12750 0 ct.oc.capture_buffer\[168\]
rlabel metal1 12144 986 12144 986 0 ct.oc.capture_buffer\[169\]
rlabel metal1 1909 19686 1909 19686 0 ct.oc.capture_buffer\[16\]
rlabel metal2 19182 10132 19182 10132 0 ct.oc.capture_buffer\[170\]
rlabel metal2 21666 4896 21666 4896 0 ct.oc.capture_buffer\[171\]
rlabel metal1 28704 5610 28704 5610 0 ct.oc.capture_buffer\[172\]
rlabel metal1 28382 850 28382 850 0 ct.oc.capture_buffer\[173\]
rlabel metal2 2162 3553 2162 3553 0 ct.oc.capture_buffer\[174\]
rlabel metal1 18216 1734 18216 1734 0 ct.oc.capture_buffer\[175\]
rlabel metal1 27278 1496 27278 1496 0 ct.oc.capture_buffer\[176\]
rlabel metal2 4600 1700 4600 1700 0 ct.oc.capture_buffer\[177\]
rlabel metal2 19826 3060 19826 3060 0 ct.oc.capture_buffer\[178\]
rlabel metal1 26956 1938 26956 1938 0 ct.oc.capture_buffer\[179\]
rlabel metal2 9338 18547 9338 18547 0 ct.oc.capture_buffer\[17\]
rlabel metal1 26726 3026 26726 3026 0 ct.oc.capture_buffer\[180\]
rlabel metal1 25852 4046 25852 4046 0 ct.oc.capture_buffer\[181\]
rlabel via2 4370 1955 4370 1955 0 ct.oc.capture_buffer\[182\]
rlabel metal1 15594 4182 15594 4182 0 ct.oc.capture_buffer\[183\]
rlabel metal2 24886 799 24886 799 0 ct.oc.capture_buffer\[184\]
rlabel via2 4278 1309 4278 1309 0 ct.oc.capture_buffer\[185\]
rlabel metal1 25116 2482 25116 2482 0 ct.oc.capture_buffer\[186\]
rlabel metal1 25300 4794 25300 4794 0 ct.oc.capture_buffer\[187\]
rlabel metal1 25392 5134 25392 5134 0 ct.oc.capture_buffer\[188\]
rlabel metal1 25898 5270 25898 5270 0 ct.oc.capture_buffer\[189\]
rlabel metal3 8832 12988 8832 12988 0 ct.oc.capture_buffer\[18\]
rlabel metal2 14582 612 14582 612 0 ct.oc.capture_buffer\[190\]
rlabel metal1 25254 1326 25254 1326 0 ct.oc.capture_buffer\[191\]
rlabel metal1 24564 1938 24564 1938 0 ct.oc.capture_buffer\[192\]
rlabel metal1 22908 850 22908 850 0 ct.oc.capture_buffer\[193\]
rlabel metal2 23046 3740 23046 3740 0 ct.oc.capture_buffer\[194\]
rlabel metal1 23230 5338 23230 5338 0 ct.oc.capture_buffer\[195\]
rlabel metal2 23138 5406 23138 5406 0 ct.oc.capture_buffer\[196\]
rlabel metal2 22862 5372 22862 5372 0 ct.oc.capture_buffer\[197\]
rlabel metal1 24610 816 24610 816 0 ct.oc.capture_buffer\[198\]
rlabel metal1 23782 2618 23782 2618 0 ct.oc.capture_buffer\[199\]
rlabel metal1 9476 17714 9476 17714 0 ct.oc.capture_buffer\[19\]
rlabel metal1 11684 19278 11684 19278 0 ct.oc.capture_buffer\[1\]
rlabel metal1 22310 1972 22310 1972 0 ct.oc.capture_buffer\[200\]
rlabel metal1 23736 1530 23736 1530 0 ct.oc.capture_buffer\[201\]
rlabel metal1 21068 4114 21068 4114 0 ct.oc.capture_buffer\[202\]
rlabel metal1 21620 6222 21620 6222 0 ct.oc.capture_buffer\[203\]
rlabel metal1 21942 5746 21942 5746 0 ct.oc.capture_buffer\[204\]
rlabel metal1 21574 5202 21574 5202 0 ct.oc.capture_buffer\[205\]
rlabel metal2 22770 1530 22770 1530 0 ct.oc.capture_buffer\[206\]
rlabel metal1 21574 3026 21574 3026 0 ct.oc.capture_buffer\[207\]
rlabel metal1 20148 1530 20148 1530 0 ct.oc.capture_buffer\[208\]
rlabel metal1 23506 1496 23506 1496 0 ct.oc.capture_buffer\[209\]
rlabel metal1 5244 11322 5244 11322 0 ct.oc.capture_buffer\[20\]
rlabel metal2 19090 4012 19090 4012 0 ct.oc.capture_buffer\[210\]
rlabel metal1 19090 4658 19090 4658 0 ct.oc.capture_buffer\[211\]
rlabel metal1 19780 5746 19780 5746 0 ct.oc.capture_buffer\[212\]
rlabel metal1 19872 5202 19872 5202 0 ct.oc.capture_buffer\[213\]
rlabel metal1 21114 986 21114 986 0 ct.oc.capture_buffer\[214\]
rlabel metal1 20056 3026 20056 3026 0 ct.oc.capture_buffer\[215\]
rlabel metal1 16422 986 16422 986 0 ct.oc.capture_buffer\[216\]
rlabel metal2 20562 1768 20562 1768 0 ct.oc.capture_buffer\[217\]
rlabel metal1 18170 2074 18170 2074 0 ct.oc.capture_buffer\[218\]
rlabel metal1 17112 4658 17112 4658 0 ct.oc.capture_buffer\[219\]
rlabel metal2 1886 16116 1886 16116 0 ct.oc.capture_buffer\[21\]
rlabel metal1 16928 5746 16928 5746 0 ct.oc.capture_buffer\[220\]
rlabel metal2 16974 5644 16974 5644 0 ct.oc.capture_buffer\[221\]
rlabel metal1 17802 986 17802 986 0 ct.oc.capture_buffer\[222\]
rlabel metal1 14398 2074 14398 2074 0 ct.oc.capture_buffer\[223\]
rlabel metal1 13340 918 13340 918 0 ct.oc.capture_buffer\[224\]
rlabel metal1 14536 2482 14536 2482 0 ct.oc.capture_buffer\[225\]
rlabel metal1 13892 986 13892 986 0 ct.oc.capture_buffer\[226\]
rlabel metal1 14168 4658 14168 4658 0 ct.oc.capture_buffer\[227\]
rlabel metal1 14536 5746 14536 5746 0 ct.oc.capture_buffer\[228\]
rlabel metal1 14674 5202 14674 5202 0 ct.oc.capture_buffer\[229\]
rlabel metal1 9545 11866 9545 11866 0 ct.oc.capture_buffer\[22\]
rlabel metal2 14398 884 14398 884 0 ct.oc.capture_buffer\[230\]
rlabel metal1 13662 2890 13662 2890 0 ct.oc.capture_buffer\[231\]
rlabel metal2 5198 1071 5198 1071 0 ct.oc.capture_buffer\[232\]
rlabel via2 5934 1547 5934 1547 0 ct.oc.capture_buffer\[233\]
rlabel metal1 12282 3570 12282 3570 0 ct.oc.capture_buffer\[234\]
rlabel metal1 13570 5780 13570 5780 0 ct.oc.capture_buffer\[235\]
rlabel metal2 12834 5644 12834 5644 0 ct.oc.capture_buffer\[236\]
rlabel metal2 13110 5372 13110 5372 0 ct.oc.capture_buffer\[237\]
rlabel via1 10810 629 10810 629 0 ct.oc.capture_buffer\[238\]
rlabel metal1 11776 2958 11776 2958 0 ct.oc.capture_buffer\[239\]
rlabel metal2 2070 18173 2070 18173 0 ct.oc.capture_buffer\[23\]
rlabel metal1 9476 1870 9476 1870 0 ct.oc.capture_buffer\[240\]
rlabel metal2 12650 10353 12650 10353 0 ct.oc.capture_buffer\[241\]
rlabel metal1 9476 3570 9476 3570 0 ct.oc.capture_buffer\[242\]
rlabel metal1 10994 5610 10994 5610 0 ct.oc.capture_buffer\[243\]
rlabel metal1 10810 4114 10810 4114 0 ct.oc.capture_buffer\[244\]
rlabel metal1 10212 4794 10212 4794 0 ct.oc.capture_buffer\[245\]
rlabel metal1 9798 1326 9798 1326 0 ct.oc.capture_buffer\[246\]
rlabel metal1 7958 2074 7958 2074 0 ct.oc.capture_buffer\[247\]
rlabel metal1 6808 850 6808 850 0 ct.oc.capture_buffer\[248\]
rlabel metal1 2116 1870 2116 1870 0 ct.oc.capture_buffer\[249\]
rlabel metal2 20654 17816 20654 17816 0 ct.oc.capture_buffer\[24\]
rlabel metal1 6210 1292 6210 1292 0 ct.oc.capture_buffer\[250\]
rlabel metal1 7176 5134 7176 5134 0 ct.oc.capture_buffer\[251\]
rlabel metal1 8510 3706 8510 3706 0 ct.oc.capture_buffer\[252\]
rlabel metal1 8556 986 8556 986 0 ct.oc.capture_buffer\[253\]
rlabel metal2 2070 1717 2070 1717 0 ct.oc.capture_buffer\[254\]
rlabel metal1 9614 2482 9614 2482 0 ct.oc.capture_buffer\[255\]
rlabel metal1 17296 18734 17296 18734 0 ct.oc.capture_buffer\[256\]
rlabel metal2 1702 1020 1702 1020 0 ct.oc.capture_buffer\[257\]
rlabel metal1 4140 986 4140 986 0 ct.oc.capture_buffer\[258\]
rlabel metal1 6486 5746 6486 5746 0 ct.oc.capture_buffer\[259\]
rlabel metal2 20746 18020 20746 18020 0 ct.oc.capture_buffer\[25\]
rlabel metal1 6486 4590 6486 4590 0 ct.oc.capture_buffer\[260\]
rlabel metal1 2346 6392 2346 6392 0 ct.oc.capture_buffer\[261\]
rlabel metal1 14490 20366 14490 20366 0 ct.oc.capture_buffer\[262\]
rlabel via3 6693 2652 6693 2652 0 ct.oc.capture_buffer\[263\]
rlabel metal2 21758 5066 21758 5066 0 ct.oc.capture_buffer\[264\]
rlabel metal1 9246 8296 9246 8296 0 ct.oc.capture_buffer\[265\]
rlabel metal2 2438 5865 2438 5865 0 ct.oc.capture_buffer\[266\]
rlabel metal2 3818 4386 3818 4386 0 ct.oc.capture_buffer\[267\]
rlabel metal1 1334 4488 1334 4488 0 ct.oc.capture_buffer\[268\]
rlabel metal2 966 3247 966 3247 0 ct.oc.capture_buffer\[269\]
rlabel metal2 18078 20825 18078 20825 0 ct.oc.capture_buffer\[26\]
rlabel metal2 1702 11322 1702 11322 0 ct.oc.capture_buffer\[270\]
rlabel metal1 4600 3502 4600 3502 0 ct.oc.capture_buffer\[271\]
rlabel metal1 21942 4794 21942 4794 0 ct.oc.capture_buffer\[272\]
rlabel metal1 2162 13838 2162 13838 0 ct.oc.capture_buffer\[273\]
rlabel metal1 18170 6086 18170 6086 0 ct.oc.capture_buffer\[274\]
rlabel metal1 3450 2074 3450 2074 0 ct.oc.capture_buffer\[275\]
rlabel metal1 3450 5712 3450 5712 0 ct.oc.capture_buffer\[276\]
rlabel metal2 1702 5389 1702 5389 0 ct.oc.capture_buffer\[277\]
rlabel metal2 2484 14484 2484 14484 0 ct.oc.capture_buffer\[278\]
rlabel metal2 16698 5542 16698 5542 0 ct.oc.capture_buffer\[279\]
rlabel metal2 8878 11866 8878 11866 0 ct.oc.capture_buffer\[27\]
rlabel metal1 2622 952 2622 952 0 ct.oc.capture_buffer\[280\]
rlabel metal2 1702 8602 1702 8602 0 ct.oc.capture_buffer\[281\]
rlabel metal1 1536 7310 1536 7310 0 ct.oc.capture_buffer\[282\]
rlabel metal1 1150 1530 1150 1530 0 ct.oc.capture_buffer\[283\]
rlabel metal2 3266 4964 3266 4964 0 ct.oc.capture_buffer\[284\]
rlabel metal1 3312 986 3312 986 0 ct.oc.capture_buffer\[285\]
rlabel metal2 1610 4947 1610 4947 0 ct.oc.capture_buffer\[286\]
rlabel metal2 2070 4845 2070 4845 0 ct.oc.capture_buffer\[287\]
rlabel metal2 8970 7242 8970 7242 0 ct.oc.capture_buffer\[288\]
rlabel metal1 6164 7922 6164 7922 0 ct.oc.capture_buffer\[289\]
rlabel metal2 1702 21658 1702 21658 0 ct.oc.capture_buffer\[28\]
rlabel metal1 5152 6970 5152 6970 0 ct.oc.capture_buffer\[290\]
rlabel metal1 6394 6290 6394 6290 0 ct.oc.capture_buffer\[291\]
rlabel metal2 6578 7837 6578 7837 0 ct.oc.capture_buffer\[292\]
rlabel metal2 9154 7582 9154 7582 0 ct.oc.capture_buffer\[293\]
rlabel metal1 9108 7922 9108 7922 0 ct.oc.capture_buffer\[294\]
rlabel metal1 9798 6222 9798 6222 0 ct.oc.capture_buffer\[295\]
rlabel metal1 15364 6766 15364 6766 0 ct.oc.capture_buffer\[296\]
rlabel metal1 14904 7310 14904 7310 0 ct.oc.capture_buffer\[297\]
rlabel metal1 14260 7922 14260 7922 0 ct.oc.capture_buffer\[298\]
rlabel metal2 17618 8228 17618 8228 0 ct.oc.capture_buffer\[299\]
rlabel metal2 16146 19261 16146 19261 0 ct.oc.capture_buffer\[29\]
rlabel metal1 8556 20570 8556 20570 0 ct.oc.capture_buffer\[2\]
rlabel metal1 15318 6222 15318 6222 0 ct.oc.capture_buffer\[300\]
rlabel metal1 11132 7446 11132 7446 0 ct.oc.capture_buffer\[301\]
rlabel metal1 11822 6834 11822 6834 0 ct.oc.capture_buffer\[302\]
rlabel metal1 11684 7310 11684 7310 0 ct.oc.capture_buffer\[303\]
rlabel metal1 14490 9554 14490 9554 0 ct.oc.capture_buffer\[304\]
rlabel metal1 13984 10574 13984 10574 0 ct.oc.capture_buffer\[305\]
rlabel metal1 15042 10030 15042 10030 0 ct.oc.capture_buffer\[306\]
rlabel metal1 14628 9010 14628 9010 0 ct.oc.capture_buffer\[307\]
rlabel metal1 14996 8398 14996 8398 0 ct.oc.capture_buffer\[308\]
rlabel metal2 10626 9486 10626 9486 0 ct.oc.capture_buffer\[309\]
rlabel metal1 12880 19686 12880 19686 0 ct.oc.capture_buffer\[30\]
rlabel metal1 11684 9010 11684 9010 0 ct.oc.capture_buffer\[310\]
rlabel metal1 10948 9146 10948 9146 0 ct.oc.capture_buffer\[311\]
rlabel metal1 13294 12274 13294 12274 0 ct.oc.capture_buffer\[312\]
rlabel metal1 13156 11186 13156 11186 0 ct.oc.capture_buffer\[313\]
rlabel metal1 12926 11866 12926 11866 0 ct.oc.capture_buffer\[314\]
rlabel metal2 14306 11968 14306 11968 0 ct.oc.capture_buffer\[315\]
rlabel metal1 14122 12750 14122 12750 0 ct.oc.capture_buffer\[316\]
rlabel metal1 9936 9486 9936 9486 0 ct.oc.capture_buffer\[317\]
rlabel metal1 10626 8466 10626 8466 0 ct.oc.capture_buffer\[318\]
rlabel metal2 9430 10268 9430 10268 0 ct.oc.capture_buffer\[319\]
rlabel metal2 13386 16541 13386 16541 0 ct.oc.capture_buffer\[31\]
rlabel metal1 10534 11730 10534 11730 0 ct.oc.capture_buffer\[320\]
rlabel metal1 10488 12206 10488 12206 0 ct.oc.capture_buffer\[321\]
rlabel metal1 10350 11322 10350 11322 0 ct.oc.capture_buffer\[322\]
rlabel metal1 10856 12750 10856 12750 0 ct.oc.capture_buffer\[323\]
rlabel metal1 10764 10642 10764 10642 0 ct.oc.capture_buffer\[324\]
rlabel metal1 8188 8602 8188 8602 0 ct.oc.capture_buffer\[325\]
rlabel metal2 8418 9044 8418 9044 0 ct.oc.capture_buffer\[326\]
rlabel metal1 7268 9146 7268 9146 0 ct.oc.capture_buffer\[327\]
rlabel metal1 6854 13158 6854 13158 0 ct.oc.capture_buffer\[328\]
rlabel metal2 7590 11356 7590 11356 0 ct.oc.capture_buffer\[329\]
rlabel metal1 4968 14586 4968 14586 0 ct.oc.capture_buffer\[32\]
rlabel metal1 7820 11866 7820 11866 0 ct.oc.capture_buffer\[330\]
rlabel metal2 8786 13124 8786 13124 0 ct.oc.capture_buffer\[331\]
rlabel metal1 7958 12818 7958 12818 0 ct.oc.capture_buffer\[332\]
rlabel metal1 6072 9690 6072 9690 0 ct.oc.capture_buffer\[333\]
rlabel metal1 5474 11220 5474 11220 0 ct.oc.capture_buffer\[334\]
rlabel metal1 6072 8398 6072 8398 0 ct.oc.capture_buffer\[335\]
rlabel metal1 4600 11730 4600 11730 0 ct.oc.capture_buffer\[336\]
rlabel metal1 4692 13294 4692 13294 0 ct.oc.capture_buffer\[337\]
rlabel metal2 5842 13668 5842 13668 0 ct.oc.capture_buffer\[338\]
rlabel metal1 4416 12750 4416 12750 0 ct.oc.capture_buffer\[339\]
rlabel metal2 16146 16643 16146 16643 0 ct.oc.capture_buffer\[33\]
rlabel metal1 4186 12206 4186 12206 0 ct.oc.capture_buffer\[340\]
rlabel metal1 4324 10098 4324 10098 0 ct.oc.capture_buffer\[341\]
rlabel metal2 4646 9860 4646 9860 0 ct.oc.capture_buffer\[342\]
rlabel metal2 5198 8772 5198 8772 0 ct.oc.capture_buffer\[343\]
rlabel metal1 3680 13702 3680 13702 0 ct.oc.capture_buffer\[344\]
rlabel metal1 1886 13362 1886 13362 0 ct.oc.capture_buffer\[345\]
rlabel metal1 1932 14450 1932 14450 0 ct.oc.capture_buffer\[346\]
rlabel metal1 1656 12818 1656 12818 0 ct.oc.capture_buffer\[347\]
rlabel metal1 2024 12206 2024 12206 0 ct.oc.capture_buffer\[348\]
rlabel metal1 2208 10030 2208 10030 0 ct.oc.capture_buffer\[349\]
rlabel metal1 4324 14314 4324 14314 0 ct.oc.capture_buffer\[34\]
rlabel metal1 966 4794 966 4794 0 ct.oc.capture_buffer\[350\]
rlabel metal1 1012 5882 1012 5882 0 ct.oc.capture_buffer\[351\]
rlabel metal1 10994 16082 10994 16082 0 ct.oc.capture_buffer\[35\]
rlabel metal1 2668 17646 2668 17646 0 ct.oc.capture_buffer\[36\]
rlabel metal2 2530 17085 2530 17085 0 ct.oc.capture_buffer\[37\]
rlabel metal2 1702 18105 1702 18105 0 ct.oc.capture_buffer\[38\]
rlabel metal2 9154 13362 9154 13362 0 ct.oc.capture_buffer\[39\]
rlabel metal1 11684 20366 11684 20366 0 ct.oc.capture_buffer\[3\]
rlabel metal1 4508 14246 4508 14246 0 ct.oc.capture_buffer\[40\]
rlabel metal1 4600 14586 4600 14586 0 ct.oc.capture_buffer\[41\]
rlabel metal1 4278 14586 4278 14586 0 ct.oc.capture_buffer\[42\]
rlabel metal2 4922 15164 4922 15164 0 ct.oc.capture_buffer\[43\]
rlabel metal2 2070 15521 2070 15521 0 ct.oc.capture_buffer\[44\]
rlabel metal1 1518 14926 1518 14926 0 ct.oc.capture_buffer\[45\]
rlabel metal1 9062 13974 9062 13974 0 ct.oc.capture_buffer\[46\]
rlabel metal2 6118 14688 6118 14688 0 ct.oc.capture_buffer\[47\]
rlabel metal1 6578 13838 6578 13838 0 ct.oc.capture_buffer\[48\]
rlabel metal1 6256 14586 6256 14586 0 ct.oc.capture_buffer\[49\]
rlabel metal1 20010 18326 20010 18326 0 ct.oc.capture_buffer\[4\]
rlabel metal1 6716 14586 6716 14586 0 ct.oc.capture_buffer\[50\]
rlabel metal2 5474 14943 5474 14943 0 ct.oc.capture_buffer\[51\]
rlabel metal1 9246 14586 9246 14586 0 ct.oc.capture_buffer\[52\]
rlabel metal2 9430 15606 9430 15606 0 ct.oc.capture_buffer\[53\]
rlabel metal1 9108 14926 9108 14926 0 ct.oc.capture_buffer\[54\]
rlabel metal1 9179 16014 9179 16014 0 ct.oc.capture_buffer\[55\]
rlabel metal2 12742 14722 12742 14722 0 ct.oc.capture_buffer\[56\]
rlabel metal1 11178 14586 11178 14586 0 ct.oc.capture_buffer\[57\]
rlabel metal1 11684 14586 11684 14586 0 ct.oc.capture_buffer\[58\]
rlabel metal2 12374 14212 12374 14212 0 ct.oc.capture_buffer\[59\]
rlabel metal1 8694 20978 8694 20978 0 ct.oc.capture_buffer\[5\]
rlabel metal1 12788 14042 12788 14042 0 ct.oc.capture_buffer\[60\]
rlabel metal2 10994 16048 10994 16048 0 ct.oc.capture_buffer\[61\]
rlabel metal2 5842 17408 5842 17408 0 ct.oc.capture_buffer\[62\]
rlabel metal1 9384 16218 9384 16218 0 ct.oc.capture_buffer\[63\]
rlabel metal1 15410 13906 15410 13906 0 ct.oc.capture_buffer\[64\]
rlabel metal1 13846 13974 13846 13974 0 ct.oc.capture_buffer\[65\]
rlabel metal1 14260 14042 14260 14042 0 ct.oc.capture_buffer\[66\]
rlabel metal1 15778 13498 15778 13498 0 ct.oc.capture_buffer\[67\]
rlabel metal1 13892 17714 13892 17714 0 ct.oc.capture_buffer\[68\]
rlabel metal1 14260 19686 14260 19686 0 ct.oc.capture_buffer\[69\]
rlabel metal2 13846 14569 13846 14569 0 ct.oc.capture_buffer\[6\]
rlabel metal1 15272 15538 15272 15538 0 ct.oc.capture_buffer\[70\]
rlabel metal1 14260 18190 14260 18190 0 ct.oc.capture_buffer\[71\]
rlabel metal1 18538 15538 18538 15538 0 ct.oc.capture_buffer\[72\]
rlabel metal1 18216 13838 18216 13838 0 ct.oc.capture_buffer\[73\]
rlabel metal1 18308 13362 18308 13362 0 ct.oc.capture_buffer\[74\]
rlabel metal1 18354 14450 18354 14450 0 ct.oc.capture_buffer\[75\]
rlabel metal1 19136 16014 19136 16014 0 ct.oc.capture_buffer\[76\]
rlabel metal2 17158 17612 17158 17612 0 ct.oc.capture_buffer\[77\]
rlabel metal3 19964 19448 19964 19448 0 ct.oc.capture_buffer\[78\]
rlabel metal1 18446 16626 18446 16626 0 ct.oc.capture_buffer\[79\]
rlabel metal1 12282 12954 12282 12954 0 ct.oc.capture_buffer\[7\]
rlabel metal1 21666 13192 21666 13192 0 ct.oc.capture_buffer\[80\]
rlabel metal1 19642 12614 19642 12614 0 ct.oc.capture_buffer\[81\]
rlabel metal2 21482 14450 21482 14450 0 ct.oc.capture_buffer\[82\]
rlabel metal2 19734 13022 19734 13022 0 ct.oc.capture_buffer\[83\]
rlabel metal2 21758 20196 21758 20196 0 ct.oc.capture_buffer\[84\]
rlabel metal2 21390 19278 21390 19278 0 ct.oc.capture_buffer\[85\]
rlabel metal1 22954 17680 22954 17680 0 ct.oc.capture_buffer\[86\]
rlabel via2 21206 17187 21206 17187 0 ct.oc.capture_buffer\[87\]
rlabel metal1 23874 13770 23874 13770 0 ct.oc.capture_buffer\[88\]
rlabel metal1 23644 13974 23644 13974 0 ct.oc.capture_buffer\[89\]
rlabel metal1 7314 18802 7314 18802 0 ct.oc.capture_buffer\[8\]
rlabel metal2 23046 14280 23046 14280 0 ct.oc.capture_buffer\[90\]
rlabel metal1 24564 15538 24564 15538 0 ct.oc.capture_buffer\[91\]
rlabel metal1 30360 13226 30360 13226 0 ct.oc.capture_buffer\[92\]
rlabel metal1 28750 18088 28750 18088 0 ct.oc.capture_buffer\[93\]
rlabel metal2 21942 20451 21942 20451 0 ct.oc.capture_buffer\[94\]
rlabel metal1 18768 20502 18768 20502 0 ct.oc.capture_buffer\[95\]
rlabel metal1 28658 17170 28658 17170 0 ct.oc.capture_buffer\[96\]
rlabel metal1 27899 16082 27899 16082 0 ct.oc.capture_buffer\[97\]
rlabel metal2 26082 15878 26082 15878 0 ct.oc.capture_buffer\[98\]
rlabel metal1 30360 9622 30360 9622 0 ct.oc.capture_buffer\[99\]
rlabel metal1 13846 18360 13846 18360 0 ct.oc.capture_buffer\[9\]
rlabel metal1 5934 20400 5934 20400 0 ct.oc.data_chain\[0\]
rlabel metal1 24725 17646 24725 17646 0 ct.oc.data_chain\[100\]
rlabel viali 24611 16576 24611 16576 0 ct.oc.data_chain\[101\]
rlabel metal1 25415 17170 25415 17170 0 ct.oc.data_chain\[102\]
rlabel metal1 25415 18258 25415 18258 0 ct.oc.data_chain\[103\]
rlabel metal1 26589 17170 26589 17170 0 ct.oc.data_chain\[104\]
rlabel viali 26543 16080 26543 16080 0 ct.oc.data_chain\[105\]
rlabel viali 26913 16559 26913 16559 0 ct.oc.data_chain\[106\]
rlabel via1 26911 17646 26911 17646 0 ct.oc.data_chain\[107\]
rlabel via1 28659 20910 28659 20910 0 ct.oc.data_chain\[108\]
rlabel metal1 28727 20434 28727 20434 0 ct.oc.data_chain\[109\]
rlabel metal1 10718 20570 10718 20570 0 ct.oc.data_chain\[10\]
rlabel metal1 25875 19346 25875 19346 0 ct.oc.data_chain\[110\]
rlabel metal1 24725 18734 24725 18734 0 ct.oc.data_chain\[111\]
rlabel metal1 25093 13906 25093 13906 0 ct.oc.data_chain\[112\]
rlabel metal1 26913 13329 26913 13329 0 ct.oc.data_chain\[113\]
rlabel metal1 27095 13906 27095 13906 0 ct.oc.data_chain\[114\]
rlabel metal1 26083 12818 26083 12818 0 ct.oc.data_chain\[115\]
rlabel metal1 27416 14246 27416 14246 0 ct.oc.data_chain\[116\]
rlabel metal1 28796 11866 28796 11866 0 ct.oc.data_chain\[117\]
rlabel viali 28935 19824 28935 19824 0 ct.oc.data_chain\[118\]
rlabel metal3 28106 19380 28106 19380 0 ct.oc.data_chain\[119\]
rlabel metal2 12834 20876 12834 20876 0 ct.oc.data_chain\[11\]
rlabel metal1 24197 12818 24197 12818 0 ct.oc.data_chain\[120\]
rlabel metal1 24613 13331 24613 13331 0 ct.oc.data_chain\[121\]
rlabel metal2 22402 13090 22402 13090 0 ct.oc.data_chain\[122\]
rlabel metal1 23782 11866 23782 11866 0 ct.oc.data_chain\[123\]
rlabel metal1 26726 11866 26726 11866 0 ct.oc.data_chain\[124\]
rlabel metal1 27301 11730 27301 11730 0 ct.oc.data_chain\[125\]
rlabel metal3 29095 6868 29095 6868 0 ct.oc.data_chain\[126\]
rlabel metal1 28429 14382 28429 14382 0 ct.oc.data_chain\[127\]
rlabel metal1 21436 11322 21436 11322 0 ct.oc.data_chain\[128\]
rlabel via1 20562 13905 20562 13905 0 ct.oc.data_chain\[129\]
rlabel metal1 8516 19244 8516 19244 0 ct.oc.data_chain\[12\]
rlabel metal1 20333 12818 20333 12818 0 ct.oc.data_chain\[130\]
rlabel metal1 22517 11730 22517 11730 0 ct.oc.data_chain\[131\]
rlabel metal1 25277 11730 25277 11730 0 ct.oc.data_chain\[132\]
rlabel metal1 27669 8466 27669 8466 0 ct.oc.data_chain\[133\]
rlabel via1 28267 6766 28267 6766 0 ct.oc.data_chain\[134\]
rlabel metal1 28244 9894 28244 9894 0 ct.oc.data_chain\[135\]
rlabel metal1 19136 10234 19136 10234 0 ct.oc.data_chain\[136\]
rlabel metal1 18999 11730 18999 11730 0 ct.oc.data_chain\[137\]
rlabel metal2 18446 12036 18446 12036 0 ct.oc.data_chain\[138\]
rlabel metal1 21621 10030 21621 10030 0 ct.oc.data_chain\[139\]
rlabel metal1 8465 20910 8465 20910 0 ct.oc.data_chain\[13\]
rlabel metal1 24335 11118 24335 11118 0 ct.oc.data_chain\[140\]
rlabel metal1 26726 10778 26726 10778 0 ct.oc.data_chain\[141\]
rlabel metal1 27025 8942 27025 8942 0 ct.oc.data_chain\[142\]
rlabel viali 26911 10030 26911 10030 0 ct.oc.data_chain\[143\]
rlabel metal1 17733 10030 17733 10030 0 ct.oc.data_chain\[144\]
rlabel metal1 18101 11118 18101 11118 0 ct.oc.data_chain\[145\]
rlabel metal2 17894 10404 17894 10404 0 ct.oc.data_chain\[146\]
rlabel metal1 20401 10642 20401 10642 0 ct.oc.data_chain\[147\]
rlabel metal1 22333 11118 22333 11118 0 ct.oc.data_chain\[148\]
rlabel metal1 25415 10642 25415 10642 0 ct.oc.data_chain\[149\]
rlabel metal1 6211 20928 6211 20928 0 ct.oc.data_chain\[14\]
rlabel metal1 26221 9554 26221 9554 0 ct.oc.data_chain\[150\]
rlabel viali 24621 10030 24621 10030 0 ct.oc.data_chain\[151\]
rlabel metal1 17757 9554 17757 9554 0 ct.oc.data_chain\[152\]
rlabel metal1 19573 9554 19573 9554 0 ct.oc.data_chain\[153\]
rlabel metal1 18423 8942 18423 8942 0 ct.oc.data_chain\[154\]
rlabel via1 19183 8466 19183 8466 0 ct.oc.data_chain\[155\]
rlabel metal1 21345 9552 21345 9552 0 ct.oc.data_chain\[156\]
rlabel metal1 24863 9554 24863 9554 0 ct.oc.data_chain\[157\]
rlabel metal1 24013 8466 24013 8466 0 ct.oc.data_chain\[158\]
rlabel metal1 23529 8942 23529 8942 0 ct.oc.data_chain\[159\]
rlabel viali 4005 21521 4005 21521 0 ct.oc.data_chain\[15\]
rlabel metal2 19274 6511 19274 6511 0 ct.oc.data_chain\[160\]
rlabel metal1 29670 6154 29670 6154 0 ct.oc.data_chain\[161\]
rlabel metal2 21758 6800 21758 6800 0 ct.oc.data_chain\[162\]
rlabel metal2 18630 6817 18630 6817 0 ct.oc.data_chain\[163\]
rlabel metal1 22862 7786 22862 7786 0 ct.oc.data_chain\[164\]
rlabel metal1 26864 6970 26864 6970 0 ct.oc.data_chain\[165\]
rlabel via2 22034 8483 22034 8483 0 ct.oc.data_chain\[166\]
rlabel metal2 22034 6987 22034 6987 0 ct.oc.data_chain\[167\]
rlabel metal1 18446 12920 18446 12920 0 ct.oc.data_chain\[168\]
rlabel metal2 5934 4403 5934 4403 0 ct.oc.data_chain\[169\]
rlabel metal2 8924 18734 8924 18734 0 ct.oc.data_chain\[16\]
rlabel metal1 20378 9928 20378 9928 0 ct.oc.data_chain\[170\]
rlabel metal1 18538 4148 18538 4148 0 ct.oc.data_chain\[171\]
rlabel metal1 29256 1530 29256 1530 0 ct.oc.data_chain\[172\]
rlabel viali 28475 2416 28475 2416 0 ct.oc.data_chain\[173\]
rlabel via2 3082 2907 3082 2907 0 ct.oc.data_chain\[174\]
rlabel viali 27222 4113 27222 4113 0 ct.oc.data_chain\[175\]
rlabel metal1 12558 12920 12558 12920 0 ct.oc.data_chain\[176\]
rlabel viali 4279 4112 4279 4112 0 ct.oc.data_chain\[177\]
rlabel metal2 20838 1873 20838 1873 0 ct.oc.data_chain\[178\]
rlabel metal2 17894 3859 17894 3859 0 ct.oc.data_chain\[179\]
rlabel metal1 10995 18258 10995 18258 0 ct.oc.data_chain\[17\]
rlabel via1 28107 1326 28107 1326 0 ct.oc.data_chain\[180\]
rlabel metal1 26726 884 26726 884 0 ct.oc.data_chain\[181\]
rlabel metal1 5014 2074 5014 2074 0 ct.oc.data_chain\[182\]
rlabel metal2 16376 1836 16376 1836 0 ct.oc.data_chain\[183\]
rlabel metal1 10534 2482 10534 2482 0 ct.oc.data_chain\[184\]
rlabel metal2 5566 2023 5566 2023 0 ct.oc.data_chain\[185\]
rlabel metal1 19573 850 19573 850 0 ct.oc.data_chain\[186\]
rlabel viali 26769 1920 26769 1920 0 ct.oc.data_chain\[187\]
rlabel metal1 26451 3026 26451 3026 0 ct.oc.data_chain\[188\]
rlabel metal1 25461 4114 25461 4114 0 ct.oc.data_chain\[189\]
rlabel metal2 10258 19958 10258 19958 0 ct.oc.data_chain\[18\]
rlabel metal2 15318 357 15318 357 0 ct.oc.data_chain\[190\]
rlabel metal1 14306 4114 14306 4114 0 ct.oc.data_chain\[191\]
rlabel metal2 9246 595 9246 595 0 ct.oc.data_chain\[192\]
rlabel metal2 4094 1105 4094 1105 0 ct.oc.data_chain\[193\]
rlabel via1 24611 2414 24611 2414 0 ct.oc.data_chain\[194\]
rlabel metal1 26865 5678 26865 5678 0 ct.oc.data_chain\[195\]
rlabel metal1 24771 5202 24771 5202 0 ct.oc.data_chain\[196\]
rlabel metal1 24427 6290 24427 6290 0 ct.oc.data_chain\[197\]
rlabel metal2 14306 578 14306 578 0 ct.oc.data_chain\[198\]
rlabel metal1 24656 1326 24656 1326 0 ct.oc.data_chain\[199\]
rlabel metal1 11133 21522 11133 21522 0 ct.oc.data_chain\[19\]
rlabel metal1 12880 19482 12880 19482 0 ct.oc.data_chain\[1\]
rlabel metal1 24337 1901 24337 1901 0 ct.oc.data_chain\[200\]
rlabel metal1 22149 850 22149 850 0 ct.oc.data_chain\[201\]
rlabel viali 22773 3503 22773 3503 0 ct.oc.data_chain\[202\]
rlabel metal1 22701 6766 22701 6766 0 ct.oc.data_chain\[203\]
rlabel viali 23967 5678 23967 5678 0 ct.oc.data_chain\[204\]
rlabel metal1 22701 4590 22701 4590 0 ct.oc.data_chain\[205\]
rlabel via1 24335 850 24335 850 0 ct.oc.data_chain\[206\]
rlabel metal1 24197 3026 24197 3026 0 ct.oc.data_chain\[207\]
rlabel metal1 21445 1936 21445 1936 0 ct.oc.data_chain\[208\]
rlabel metal1 21713 2414 21713 2414 0 ct.oc.data_chain\[209\]
rlabel metal1 5981 19346 5981 19346 0 ct.oc.data_chain\[20\]
rlabel via1 20839 4114 20839 4114 0 ct.oc.data_chain\[210\]
rlabel metal1 20977 6290 20977 6290 0 ct.oc.data_chain\[211\]
rlabel metal1 21161 5678 21161 5678 0 ct.oc.data_chain\[212\]
rlabel metal1 21115 5202 21115 5202 0 ct.oc.data_chain\[213\]
rlabel metal1 21433 1326 21433 1326 0 ct.oc.data_chain\[214\]
rlabel metal1 21115 3026 21115 3026 0 ct.oc.data_chain\[215\]
rlabel metal1 18723 1938 18723 1938 0 ct.oc.data_chain\[216\]
rlabel viali 18815 2414 18815 2414 0 ct.oc.data_chain\[217\]
rlabel metal1 18817 3537 18817 3537 0 ct.oc.data_chain\[218\]
rlabel viali 18907 4590 18907 4590 0 ct.oc.data_chain\[219\]
rlabel metal1 6165 21522 6165 21522 0 ct.oc.data_chain\[21\]
rlabel viali 18907 5678 18907 5678 0 ct.oc.data_chain\[220\]
rlabel metal1 18769 5202 18769 5202 0 ct.oc.data_chain\[221\]
rlabel viali 18815 1326 18815 1326 0 ct.oc.data_chain\[222\]
rlabel metal1 18769 3026 18769 3026 0 ct.oc.data_chain\[223\]
rlabel metal1 16423 1938 16423 1938 0 ct.oc.data_chain\[224\]
rlabel viali 16607 2414 16607 2414 0 ct.oc.data_chain\[225\]
rlabel metal1 16609 3537 16609 3537 0 ct.oc.data_chain\[226\]
rlabel viali 16699 4590 16699 4590 0 ct.oc.data_chain\[227\]
rlabel viali 16699 5678 16699 5678 0 ct.oc.data_chain\[228\]
rlabel metal1 16423 5202 16423 5202 0 ct.oc.data_chain\[229\]
rlabel metal1 12788 18666 12788 18666 0 ct.oc.data_chain\[22\]
rlabel viali 16607 1326 16607 1326 0 ct.oc.data_chain\[230\]
rlabel metal1 16423 3026 16423 3026 0 ct.oc.data_chain\[231\]
rlabel metal1 13893 1938 13893 1938 0 ct.oc.data_chain\[232\]
rlabel viali 14307 2414 14307 2414 0 ct.oc.data_chain\[233\]
rlabel metal1 14309 3537 14309 3537 0 ct.oc.data_chain\[234\]
rlabel via1 14307 4590 14307 4590 0 ct.oc.data_chain\[235\]
rlabel metal1 13524 5338 13524 5338 0 ct.oc.data_chain\[236\]
rlabel metal1 14307 5202 14307 5202 0 ct.oc.data_chain\[237\]
rlabel viali 14307 1326 14307 1326 0 ct.oc.data_chain\[238\]
rlabel metal1 13939 3026 13939 3026 0 ct.oc.data_chain\[239\]
rlabel metal1 4555 20434 4555 20434 0 ct.oc.data_chain\[23\]
rlabel metal1 11455 1938 11455 1938 0 ct.oc.data_chain\[240\]
rlabel metal1 9936 1530 9936 1530 0 ct.oc.data_chain\[241\]
rlabel metal1 11915 3502 11915 3502 0 ct.oc.data_chain\[242\]
rlabel metal1 12213 5678 12213 5678 0 ct.oc.data_chain\[243\]
rlabel via1 11731 5202 11731 5202 0 ct.oc.data_chain\[244\]
rlabel via1 12099 4592 12099 4592 0 ct.oc.data_chain\[245\]
rlabel viali 12099 1344 12099 1344 0 ct.oc.data_chain\[246\]
rlabel metal1 11455 3026 11455 3026 0 ct.oc.data_chain\[247\]
rlabel metal1 9201 1938 9201 1938 0 ct.oc.data_chain\[248\]
rlabel viali 6973 1344 6973 1344 0 ct.oc.data_chain\[249\]
rlabel metal1 8971 17170 8971 17170 0 ct.oc.data_chain\[24\]
rlabel metal1 8694 3162 8694 3162 0 ct.oc.data_chain\[250\]
rlabel via1 11087 6290 11087 6290 0 ct.oc.data_chain\[251\]
rlabel metal1 10351 4114 10351 4114 0 ct.oc.data_chain\[252\]
rlabel viali 9523 5200 9523 5200 0 ct.oc.data_chain\[253\]
rlabel via1 9155 1326 9155 1326 0 ct.oc.data_chain\[254\]
rlabel metal1 9798 2618 9798 2618 0 ct.oc.data_chain\[255\]
rlabel metal2 18170 15509 18170 15509 0 ct.oc.data_chain\[256\]
rlabel metal2 2806 1462 2806 1462 0 ct.oc.data_chain\[257\]
rlabel viali 6624 3025 6624 3025 0 ct.oc.data_chain\[258\]
rlabel metal1 6831 5202 6831 5202 0 ct.oc.data_chain\[259\]
rlabel metal3 9016 17884 9016 17884 0 ct.oc.data_chain\[25\]
rlabel metal1 8327 4590 8327 4590 0 ct.oc.data_chain\[260\]
rlabel metal1 8326 3638 8326 3638 0 ct.oc.data_chain\[261\]
rlabel metal2 2254 1394 2254 1394 0 ct.oc.data_chain\[262\]
rlabel metal1 8419 2414 8419 2414 0 ct.oc.data_chain\[263\]
rlabel metal1 4646 9078 4646 9078 0 ct.oc.data_chain\[264\]
rlabel metal1 1610 816 1610 816 0 ct.oc.data_chain\[265\]
rlabel metal1 6165 1938 6165 1938 0 ct.oc.data_chain\[266\]
rlabel metal1 6118 5338 6118 5338 0 ct.oc.data_chain\[267\]
rlabel metal1 6305 4627 6305 4627 0 ct.oc.data_chain\[268\]
rlabel via1 6487 3502 6487 3502 0 ct.oc.data_chain\[269\]
rlabel metal1 8741 19346 8741 19346 0 ct.oc.data_chain\[26\]
rlabel via3 14053 19380 14053 19380 0 ct.oc.data_chain\[270\]
rlabel via1 6486 2415 6486 2415 0 ct.oc.data_chain\[271\]
rlabel metal3 9729 20740 9729 20740 0 ct.oc.data_chain\[272\]
rlabel metal1 3405 8466 3405 8466 0 ct.oc.data_chain\[273\]
rlabel metal1 1840 3536 1840 3536 0 ct.oc.data_chain\[274\]
rlabel metal1 4761 5202 4761 5202 0 ct.oc.data_chain\[275\]
rlabel via1 4003 4590 4003 4590 0 ct.oc.data_chain\[276\]
rlabel metal1 3542 5338 3542 5338 0 ct.oc.data_chain\[277\]
rlabel metal2 2116 14076 2116 14076 0 ct.oc.data_chain\[278\]
rlabel metal1 3450 2618 3450 2618 0 ct.oc.data_chain\[279\]
rlabel metal1 9017 17646 9017 17646 0 ct.oc.data_chain\[27\]
rlabel via1 9155 21522 9155 21522 0 ct.oc.data_chain\[280\]
rlabel metal1 2139 13906 2139 13906 0 ct.oc.data_chain\[281\]
rlabel metal1 6489 4079 6489 4079 0 ct.oc.data_chain\[282\]
rlabel metal1 3933 6290 3933 6290 0 ct.oc.data_chain\[283\]
rlabel metal1 1978 5712 1978 5712 0 ct.oc.data_chain\[284\]
rlabel viali 1462 5193 1462 5193 0 ct.oc.data_chain\[285\]
rlabel metal2 1518 16677 1518 16677 0 ct.oc.data_chain\[286\]
rlabel metal1 1909 2414 1909 2414 0 ct.oc.data_chain\[287\]
rlabel via2 2162 6307 2162 6307 0 ct.oc.data_chain\[288\]
rlabel metal1 2093 8466 2093 8466 0 ct.oc.data_chain\[289\]
rlabel metal1 4005 18769 4005 18769 0 ct.oc.data_chain\[28\]
rlabel metal1 2116 7378 2116 7378 0 ct.oc.data_chain\[290\]
rlabel metal1 4255 7854 4255 7854 0 ct.oc.data_chain\[291\]
rlabel metal1 2548 6784 2548 6784 0 ct.oc.data_chain\[292\]
rlabel metal2 7682 7344 7682 7344 0 ct.oc.data_chain\[293\]
rlabel metal2 1334 4063 1334 4063 0 ct.oc.data_chain\[294\]
rlabel metal2 8970 5661 8970 5661 0 ct.oc.data_chain\[295\]
rlabel via2 15686 6715 15686 6715 0 ct.oc.data_chain\[296\]
rlabel metal2 16238 7667 16238 7667 0 ct.oc.data_chain\[297\]
rlabel metal2 15686 7565 15686 7565 0 ct.oc.data_chain\[298\]
rlabel metal2 17618 9027 17618 9027 0 ct.oc.data_chain\[299\]
rlabel metal1 17204 20230 17204 20230 0 ct.oc.data_chain\[29\]
rlabel metal1 12926 22032 12926 22032 0 ct.oc.data_chain\[2\]
rlabel metal2 13754 6749 13754 6749 0 ct.oc.data_chain\[300\]
rlabel metal2 13202 7616 13202 7616 0 ct.oc.data_chain\[301\]
rlabel metal2 13294 6528 13294 6528 0 ct.oc.data_chain\[302\]
rlabel metal2 13110 6732 13110 6732 0 ct.oc.data_chain\[303\]
rlabel metal1 14421 6766 14421 6766 0 ct.oc.data_chain\[304\]
rlabel metal1 15111 7378 15111 7378 0 ct.oc.data_chain\[305\]
rlabel metal1 14881 7854 14881 7854 0 ct.oc.data_chain\[306\]
rlabel metal1 15917 8466 15917 8466 0 ct.oc.data_chain\[307\]
rlabel metal1 15065 6290 15065 6290 0 ct.oc.data_chain\[308\]
rlabel metal1 12512 9894 12512 9894 0 ct.oc.data_chain\[309\]
rlabel metal2 14030 17901 14030 17901 0 ct.oc.data_chain\[30\]
rlabel metal2 12374 7786 12374 7786 0 ct.oc.data_chain\[310\]
rlabel metal2 12650 8364 12650 8364 0 ct.oc.data_chain\[311\]
rlabel viali 14033 9553 14033 9553 0 ct.oc.data_chain\[312\]
rlabel metal1 14145 10642 14145 10642 0 ct.oc.data_chain\[313\]
rlabel via1 14042 10032 14042 10032 0 ct.oc.data_chain\[314\]
rlabel metal1 14651 8942 14651 8942 0 ct.oc.data_chain\[315\]
rlabel metal1 15870 12682 15870 12682 0 ct.oc.data_chain\[316\]
rlabel metal1 10856 9554 10856 9554 0 ct.oc.data_chain\[317\]
rlabel viali 11455 8944 11455 8944 0 ct.oc.data_chain\[318\]
rlabel metal1 10948 9894 10948 9894 0 ct.oc.data_chain\[319\]
rlabel metal2 1978 20910 1978 20910 0 ct.oc.data_chain\[31\]
rlabel metal2 11546 12036 11546 12036 0 ct.oc.data_chain\[320\]
rlabel metal1 12929 11155 12929 11155 0 ct.oc.data_chain\[321\]
rlabel metal1 12929 13331 12929 13331 0 ct.oc.data_chain\[322\]
rlabel metal1 14145 11730 14145 11730 0 ct.oc.data_chain\[323\]
rlabel viali 14076 12817 14076 12817 0 ct.oc.data_chain\[324\]
rlabel metal1 9177 9554 9177 9554 0 ct.oc.data_chain\[325\]
rlabel metal2 9062 8466 9062 8466 0 ct.oc.data_chain\[326\]
rlabel viali 9155 10030 9155 10030 0 ct.oc.data_chain\[327\]
rlabel metal1 9339 11730 9339 11730 0 ct.oc.data_chain\[328\]
rlabel metal1 9016 11322 9016 11322 0 ct.oc.data_chain\[329\]
rlabel metal1 6027 17170 6027 17170 0 ct.oc.data_chain\[32\]
rlabel metal1 9430 13872 9430 13872 0 ct.oc.data_chain\[330\]
rlabel via1 9522 13243 9522 13243 0 ct.oc.data_chain\[331\]
rlabel metal1 8947 12682 8947 12682 0 ct.oc.data_chain\[332\]
rlabel viali 8053 8951 8053 8951 0 ct.oc.data_chain\[333\]
rlabel metal1 6831 9554 6831 9554 0 ct.oc.data_chain\[334\]
rlabel metal1 7061 10030 7061 10030 0 ct.oc.data_chain\[335\]
rlabel metal1 5704 11730 5704 11730 0 ct.oc.data_chain\[336\]
rlabel via1 7315 11120 7315 11120 0 ct.oc.data_chain\[337\]
rlabel metal1 6624 14042 6624 14042 0 ct.oc.data_chain\[338\]
rlabel metal1 6624 12954 6624 12954 0 ct.oc.data_chain\[339\]
rlabel viali 6949 17647 6949 17647 0 ct.oc.data_chain\[33\]
rlabel metal1 6119 12818 6119 12818 0 ct.oc.data_chain\[340\]
rlabel metal1 5935 10642 5935 10642 0 ct.oc.data_chain\[341\]
rlabel viali 6027 11728 6027 11728 0 ct.oc.data_chain\[342\]
rlabel metal1 5981 8466 5981 8466 0 ct.oc.data_chain\[343\]
rlabel metal1 3727 11730 3727 11730 0 ct.oc.data_chain\[344\]
rlabel via1 4003 13294 4003 13294 0 ct.oc.data_chain\[345\]
rlabel metal1 4279 13906 4279 13906 0 ct.oc.data_chain\[346\]
rlabel metal1 4325 12818 4325 12818 0 ct.oc.data_chain\[347\]
rlabel viali 4003 12206 4003 12206 0 ct.oc.data_chain\[348\]
rlabel viali 3819 10030 3819 10030 0 ct.oc.data_chain\[349\]
rlabel metal1 6164 18394 6164 18394 0 ct.oc.data_chain\[34\]
rlabel metal1 3405 10642 3405 10642 0 ct.oc.data_chain\[350\]
rlabel metal1 3589 9554 3589 9554 0 ct.oc.data_chain\[351\]
rlabel metal1 6119 18258 6119 18258 0 ct.oc.data_chain\[35\]
rlabel metal2 3174 19686 3174 19686 0 ct.oc.data_chain\[36\]
rlabel via2 15226 20451 15226 20451 0 ct.oc.data_chain\[37\]
rlabel metal1 14123 21522 14123 21522 0 ct.oc.data_chain\[38\]
rlabel metal1 10856 21386 10856 21386 0 ct.oc.data_chain\[39\]
rlabel metal1 19642 21352 19642 21352 0 ct.oc.data_chain\[3\]
rlabel metal1 4255 17170 4255 17170 0 ct.oc.data_chain\[40\]
rlabel metal1 5888 15130 5888 15130 0 ct.oc.data_chain\[41\]
rlabel metal1 4991 18258 4991 18258 0 ct.oc.data_chain\[42\]
rlabel viali 4029 17664 4029 17664 0 ct.oc.data_chain\[43\]
rlabel metal1 1978 17680 1978 17680 0 ct.oc.data_chain\[44\]
rlabel metal1 1978 18768 1978 18768 0 ct.oc.data_chain\[45\]
rlabel metal2 3082 17510 3082 17510 0 ct.oc.data_chain\[46\]
rlabel metal1 1610 17136 1610 17136 0 ct.oc.data_chain\[47\]
rlabel via1 4003 15470 4003 15470 0 ct.oc.data_chain\[48\]
rlabel metal1 5221 14994 5221 14994 0 ct.oc.data_chain\[49\]
rlabel metal1 4186 19992 4186 19992 0 ct.oc.data_chain\[4\]
rlabel viali 4048 16559 4048 16559 0 ct.oc.data_chain\[50\]
rlabel metal1 5221 16082 5221 16082 0 ct.oc.data_chain\[51\]
rlabel metal1 5750 15606 5750 15606 0 ct.oc.data_chain\[52\]
rlabel metal2 10534 16932 10534 16932 0 ct.oc.data_chain\[53\]
rlabel metal2 1794 15725 1794 15725 0 ct.oc.data_chain\[54\]
rlabel metal1 3818 16150 3818 16150 0 ct.oc.data_chain\[55\]
rlabel metal1 8234 13974 8234 13974 0 ct.oc.data_chain\[56\]
rlabel metal2 13110 15776 13110 15776 0 ct.oc.data_chain\[57\]
rlabel metal1 8694 15062 8694 15062 0 ct.oc.data_chain\[58\]
rlabel metal2 13018 15215 13018 15215 0 ct.oc.data_chain\[59\]
rlabel metal2 4738 20366 4738 20366 0 ct.oc.data_chain\[5\]
rlabel via1 9155 15470 9155 15470 0 ct.oc.data_chain\[60\]
rlabel metal2 11914 16864 11914 16864 0 ct.oc.data_chain\[61\]
rlabel metal2 10810 15742 10810 15742 0 ct.oc.data_chain\[62\]
rlabel metal2 13478 16320 13478 16320 0 ct.oc.data_chain\[63\]
rlabel metal1 12213 15470 12213 15470 0 ct.oc.data_chain\[64\]
rlabel metal1 12926 16082 12926 16082 0 ct.oc.data_chain\[65\]
rlabel metal1 13478 14960 13478 14960 0 ct.oc.data_chain\[66\]
rlabel metal1 12213 14382 12213 14382 0 ct.oc.data_chain\[67\]
rlabel metal1 15502 17850 15502 17850 0 ct.oc.data_chain\[68\]
rlabel metal2 12834 16966 12834 16966 0 ct.oc.data_chain\[69\]
rlabel metal1 4784 19210 4784 19210 0 ct.oc.data_chain\[6\]
rlabel metal1 13754 17578 13754 17578 0 ct.oc.data_chain\[70\]
rlabel metal1 12949 16558 12949 16558 0 ct.oc.data_chain\[71\]
rlabel viali 14675 13904 14675 13904 0 ct.oc.data_chain\[72\]
rlabel metal1 14951 16082 14951 16082 0 ct.oc.data_chain\[73\]
rlabel metal1 14421 14382 14421 14382 0 ct.oc.data_chain\[74\]
rlabel metal1 15985 14994 15985 14994 0 ct.oc.data_chain\[75\]
rlabel metal1 15249 17646 15249 17646 0 ct.oc.data_chain\[76\]
rlabel metal2 17066 16864 17066 16864 0 ct.oc.data_chain\[77\]
rlabel metal1 14421 15470 14421 15470 0 ct.oc.data_chain\[78\]
rlabel metal1 15295 18258 15295 18258 0 ct.oc.data_chain\[79\]
rlabel metal1 7774 16694 7774 16694 0 ct.oc.data_chain\[7\]
rlabel metal1 19366 15572 19366 15572 0 ct.oc.data_chain\[80\]
rlabel metal2 21942 13991 21942 13991 0 ct.oc.data_chain\[81\]
rlabel metal1 18515 13294 18515 13294 0 ct.oc.data_chain\[82\]
rlabel metal1 19366 14416 19366 14416 0 ct.oc.data_chain\[83\]
rlabel metal1 20654 16150 20654 16150 0 ct.oc.data_chain\[84\]
rlabel metal2 20010 16983 20010 16983 0 ct.oc.data_chain\[85\]
rlabel metal1 18446 17782 18446 17782 0 ct.oc.data_chain\[86\]
rlabel metal1 20194 17000 20194 17000 0 ct.oc.data_chain\[87\]
rlabel metal1 22181 14382 22181 14382 0 ct.oc.data_chain\[88\]
rlabel viali 21804 15471 21804 15471 0 ct.oc.data_chain\[89\]
rlabel metal1 14033 18769 14033 18769 0 ct.oc.data_chain\[8\]
rlabel metal1 20585 14994 20585 14994 0 ct.oc.data_chain\[90\]
rlabel metal1 23690 15980 23690 15980 0 ct.oc.data_chain\[91\]
rlabel metal2 24058 18054 24058 18054 0 ct.oc.data_chain\[92\]
rlabel metal1 24058 16490 24058 16490 0 ct.oc.data_chain\[93\]
rlabel metal1 22862 17612 22862 17612 0 ct.oc.data_chain\[94\]
rlabel metal2 21114 17459 21114 17459 0 ct.oc.data_chain\[95\]
rlabel metal1 25185 16082 25185 16082 0 ct.oc.data_chain\[96\]
rlabel metal2 24334 15130 24334 15130 0 ct.oc.data_chain\[97\]
rlabel metal1 24587 14994 24587 14994 0 ct.oc.data_chain\[98\]
rlabel metal2 28290 17153 28290 17153 0 ct.oc.data_chain\[99\]
rlabel metal1 13018 19244 13018 19244 0 ct.oc.data_chain\[9\]
rlabel metal1 6121 21114 6121 21114 0 ct.oc.mode_buffer\[0\]
rlabel metal1 21485 14586 21485 14586 0 ct.oc.mode_buffer\[10\]
rlabel metal1 24727 17714 24727 17714 0 ct.oc.mode_buffer\[11\]
rlabel metal1 27281 20230 27281 20230 0 ct.oc.mode_buffer\[12\]
rlabel via1 28845 18938 28845 18938 0 ct.oc.mode_buffer\[13\]
rlabel metal1 28385 14586 28385 14586 0 ct.oc.mode_buffer\[14\]
rlabel metal1 21255 12614 21255 12614 0 ct.oc.mode_buffer\[15\]
rlabel metal2 21666 10540 21666 10540 0 ct.oc.mode_buffer\[16\]
rlabel metal1 18222 10234 18222 10234 0 ct.oc.mode_buffer\[17\]
rlabel metal1 17299 9146 17299 9146 0 ct.oc.mode_buffer\[18\]
rlabel metal2 21942 8160 21942 8160 0 ct.oc.mode_buffer\[19\]
rlabel metal1 5661 20230 5661 20230 0 ct.oc.mode_buffer\[1\]
rlabel metal1 28060 2618 28060 2618 0 ct.oc.mode_buffer\[20\]
rlabel metal1 17391 646 17391 646 0 ct.oc.mode_buffer\[21\]
rlabel metal2 19274 1139 19274 1139 0 ct.oc.mode_buffer\[22\]
rlabel via1 9041 782 9041 782 0 ct.oc.mode_buffer\[23\]
rlabel metal1 22543 4794 22543 4794 0 ct.oc.mode_buffer\[24\]
rlabel metal1 21669 5882 21669 5882 0 ct.oc.mode_buffer\[25\]
rlabel metal1 19001 4998 19001 4998 0 ct.oc.mode_buffer\[26\]
rlabel metal1 16747 3706 16747 3706 0 ct.oc.mode_buffer\[27\]
rlabel metal1 14401 2618 14401 2618 0 ct.oc.mode_buffer\[28\]
rlabel metal1 11500 2550 11500 2550 0 ct.oc.mode_buffer\[29\]
rlabel metal1 1705 20026 1705 20026 0 ct.oc.mode_buffer\[2\]
rlabel metal1 10951 3910 10951 3910 0 ct.oc.mode_buffer\[30\]
rlabel metal1 1613 1734 1613 1734 0 ct.oc.mode_buffer\[31\]
rlabel metal1 14217 20230 14217 20230 0 ct.oc.mode_buffer\[32\]
rlabel metal1 2165 11526 2165 11526 0 ct.oc.mode_buffer\[33\]
rlabel via1 1797 21114 1797 21114 0 ct.oc.mode_buffer\[34\]
rlabel metal1 1589 4590 1589 4590 0 ct.oc.mode_buffer\[35\]
rlabel metal1 6051 6834 6051 6834 0 ct.oc.mode_buffer\[36\]
rlabel metal1 15183 8058 15183 8058 0 ct.oc.mode_buffer\[37\]
rlabel via1 13917 10030 13917 10030 0 ct.oc.mode_buffer\[38\]
rlabel metal1 9341 9350 9341 9350 0 ct.oc.mode_buffer\[39\]
rlabel metal1 1889 21318 1889 21318 0 ct.oc.mode_buffer\[3\]
rlabel metal1 9246 10506 9246 10506 0 ct.oc.mode_buffer\[40\]
rlabel via1 6029 8262 6029 8262 0 ct.oc.mode_buffer\[41\]
rlabel metal1 4465 12614 4465 12614 0 ct.oc.mode_buffer\[42\]
rlabel metal1 1751 13498 1751 13498 0 ct.oc.mode_buffer\[43\]
rlabel metal1 4143 18054 4143 18054 0 ct.oc.mode_buffer\[4\]
rlabel via1 1681 15470 1681 15470 0 ct.oc.mode_buffer\[5\]
rlabel via1 6465 14926 6465 14926 0 ct.oc.mode_buffer\[6\]
rlabel via1 12169 19822 12169 19822 0 ct.oc.mode_buffer\[7\]
rlabel via1 14193 17646 14193 17646 0 ct.oc.mode_buffer\[8\]
rlabel metal1 17183 16626 17183 16626 0 ct.oc.mode_buffer\[9\]
rlabel metal2 17158 13498 17158 13498 0 ct.oc.trig_chain\[10\]
rlabel metal1 19090 14858 19090 14858 0 ct.oc.trig_chain\[11\]
rlabel metal1 24196 17714 24196 17714 0 ct.oc.trig_chain\[12\]
rlabel metal1 27002 15470 27002 15470 0 ct.oc.trig_chain\[13\]
rlabel metal1 28382 19822 28382 19822 0 ct.oc.trig_chain\[14\]
rlabel metal2 28014 14960 28014 14960 0 ct.oc.trig_chain\[15\]
rlabel metal1 27048 8398 27048 8398 0 ct.oc.trig_chain\[16\]
rlabel metal1 26404 9010 26404 9010 0 ct.oc.trig_chain\[17\]
rlabel metal1 16882 11118 16882 11118 0 ct.oc.trig_chain\[18\]
rlabel metal1 20930 9418 20930 9418 0 ct.oc.trig_chain\[19\]
rlabel metal1 5842 21012 5842 21012 0 ct.oc.trig_chain\[1\]
rlabel metal2 21942 8636 21942 8636 0 ct.oc.trig_chain\[20\]
rlabel metal1 23414 7378 23414 7378 0 ct.oc.trig_chain\[21\]
rlabel metal2 16422 408 16422 408 0 ct.oc.trig_chain\[22\]
rlabel metal1 19044 782 19044 782 0 ct.oc.trig_chain\[23\]
rlabel metal1 13846 816 13846 816 0 ct.oc.trig_chain\[24\]
rlabel metal1 22172 4658 22172 4658 0 ct.oc.trig_chain\[25\]
rlabel metal1 21252 5746 21252 5746 0 ct.oc.trig_chain\[26\]
rlabel metal1 18722 1836 18722 1836 0 ct.oc.trig_chain\[27\]
rlabel metal1 16100 2414 16100 2414 0 ct.oc.trig_chain\[28\]
rlabel metal2 13892 2414 13892 2414 0 ct.oc.trig_chain\[29\]
rlabel metal1 5704 19414 5704 19414 0 ct.oc.trig_chain\[2\]
rlabel metal1 11546 2414 11546 2414 0 ct.oc.trig_chain\[30\]
rlabel metal1 10718 1292 10718 1292 0 ct.oc.trig_chain\[31\]
rlabel metal1 1150 1870 1150 1870 0 ct.oc.trig_chain\[32\]
rlabel metal1 13248 20366 13248 20366 0 ct.oc.trig_chain\[33\]
rlabel metal1 8970 3978 8970 3978 0 ct.oc.trig_chain\[34\]
rlabel metal1 1058 2414 1058 2414 0 ct.oc.trig_chain\[35\]
rlabel metal1 1104 4590 1104 4590 0 ct.oc.trig_chain\[36\]
rlabel metal1 8372 7922 8372 7922 0 ct.oc.trig_chain\[37\]
rlabel metal1 14444 7310 14444 7310 0 ct.oc.trig_chain\[38\]
rlabel metal2 13570 10336 13570 10336 0 ct.oc.trig_chain\[39\]
rlabel metal2 1334 20128 1334 20128 0 ct.oc.trig_chain\[3\]
rlabel metal1 9568 11186 9568 11186 0 ct.oc.trig_chain\[40\]
rlabel metal1 6394 11220 6394 11220 0 ct.oc.trig_chain\[41\]
rlabel metal2 6854 13872 6854 13872 0 ct.oc.trig_chain\[42\]
rlabel metal2 1978 9214 1978 9214 0 ct.oc.trig_chain\[43\]
rlabel via1 1334 13379 1334 13379 0 ct.oc.trig_chain\[44\]
rlabel metal2 1242 20468 1242 20468 0 ct.oc.trig_chain\[4\]
rlabel metal1 1334 17578 1334 17578 0 ct.oc.trig_chain\[5\]
rlabel metal1 1334 15402 1334 15402 0 ct.oc.trig_chain\[6\]
rlabel metal1 6486 15402 6486 15402 0 ct.oc.trig_chain\[7\]
rlabel metal1 11592 17714 11592 17714 0 ct.oc.trig_chain\[8\]
rlabel metal1 13662 15538 13662 15538 0 ct.oc.trig_chain\[9\]
rlabel metal2 21482 21692 21482 21692 0 ct.ro.counter\[0\]
rlabel metal1 21068 21454 21068 21454 0 ct.ro.counter\[1\]
rlabel metal1 21666 20230 21666 20230 0 ct.ro.counter\[2\]
rlabel metal2 22218 21284 22218 21284 0 ct.ro.counter\[3\]
rlabel metal1 24012 21454 24012 21454 0 ct.ro.counter\[4\]
rlabel metal2 23874 20740 23874 20740 0 ct.ro.counter\[5\]
rlabel metal1 23414 20298 23414 20298 0 ct.ro.counter\[6\]
rlabel metal1 25254 20230 25254 20230 0 ct.ro.counter\[7\]
rlabel metal1 18998 22236 18998 22236 0 ct.ro.counter_n\[0\]
rlabel metal1 20148 20910 20148 20910 0 ct.ro.counter_n\[1\]
rlabel metal1 20422 20434 20422 20434 0 ct.ro.counter_n\[2\]
rlabel metal1 23322 20944 23322 20944 0 ct.ro.counter_n\[3\]
rlabel metal1 23690 20910 23690 20910 0 ct.ro.counter_n\[4\]
rlabel metal1 21850 19822 21850 19822 0 ct.ro.counter_n\[5\]
rlabel metal1 23598 20400 23598 20400 0 ct.ro.counter_n\[6\]
rlabel metal1 25898 20400 25898 20400 0 ct.ro.counter_n\[7\]
rlabel metal2 13202 21896 13202 21896 0 ct.ro.gate
rlabel metal2 22034 19312 22034 19312 0 ct.ro.ring\[0\]
rlabel metal1 21666 19754 21666 19754 0 ct.ro.ring\[1\]
rlabel metal1 23046 16014 23046 16014 0 ct.ro.ring\[2\]
rlabel metal2 30406 13311 30406 13311 0 net1
rlabel metal1 9200 11050 9200 11050 0 net10
rlabel metal1 6026 884 6026 884 0 net11
rlabel metal1 12972 9010 12972 9010 0 net12
rlabel metal1 21482 748 21482 748 0 net13
rlabel metal2 20746 19839 20746 19839 0 net14
rlabel metal1 1426 2482 1426 2482 0 net15
rlabel metal1 9062 8432 9062 8432 0 net16
rlabel metal1 3128 21454 3128 21454 0 net17
rlabel metal1 21482 7242 21482 7242 0 net18
rlabel metal1 30130 10608 30130 10608 0 net19
rlabel metal1 31142 21556 31142 21556 0 net2
rlabel metal1 16790 18224 16790 18224 0 net20
rlabel metal1 3496 2958 3496 2958 0 net21
rlabel metal1 15732 9010 15732 9010 0 net22
rlabel metal1 19826 18292 19826 18292 0 net23
rlabel metal1 16882 6324 16882 6324 0 net24
rlabel metal2 16468 12852 16468 12852 0 net25
rlabel metal1 17618 7786 17618 7786 0 net26
rlabel metal1 8878 12750 8878 12750 0 net27
rlabel metal2 1242 18598 1242 18598 0 net28
rlabel metal1 20194 10132 20194 10132 0 net29
rlabel metal1 31234 22032 31234 22032 0 net3
rlabel metal1 27692 5746 27692 5746 0 net30
rlabel metal1 16790 7990 16790 7990 0 net31
rlabel metal1 5336 6834 5336 6834 0 net32
rlabel metal1 6256 19686 6256 19686 0 net33
rlabel metal2 21114 19839 21114 19839 0 net34
rlabel metal2 18538 2315 18538 2315 0 net35
rlabel metal1 14720 13838 14720 13838 0 net36
rlabel metal2 12374 10353 12374 10353 0 net37
rlabel metal2 24610 17629 24610 17629 0 net38
rlabel metal1 9200 20910 9200 20910 0 net39
rlabel metal2 22034 21233 22034 21233 0 net4
rlabel metal1 17986 7276 17986 7276 0 net40
rlabel metal2 19274 13022 19274 13022 0 net41
rlabel metal2 14306 16184 14306 16184 0 net42
rlabel metal1 12788 782 12788 782 0 net43
rlabel metal1 1932 19346 1932 19346 0 net44
rlabel metal1 14398 15130 14398 15130 0 net45
rlabel metal1 17066 1190 17066 1190 0 net46
rlabel metal2 17066 10268 17066 10268 0 net47
rlabel metal1 16560 13362 16560 13362 0 net48
rlabel metal1 5796 10098 5796 10098 0 net49
rlabel metal1 12098 11186 12098 11186 0 net5
rlabel metal2 13386 10472 13386 10472 0 net50
rlabel metal1 13110 10098 13110 10098 0 net51
rlabel metal1 20378 8976 20378 8976 0 net52
rlabel metal1 18400 19278 18400 19278 0 net53
rlabel metal1 18768 14926 18768 14926 0 net54
rlabel via2 13570 15011 13570 15011 0 net55
rlabel metal1 8556 13770 8556 13770 0 net56
rlabel metal1 8464 13498 8464 13498 0 net57
rlabel via2 9614 13413 9614 13413 0 net58
rlabel metal1 8510 12614 8510 12614 0 net59
rlabel metal2 8142 2074 8142 2074 0 net6
rlabel metal4 5428 20097 5428 20097 0 net60
rlabel metal2 11270 13124 11270 13124 0 net61
rlabel metal1 11454 13294 11454 13294 0 net62
rlabel metal1 6302 13396 6302 13396 0 net7
rlabel metal1 18722 2040 18722 2040 0 net8
rlabel metal2 18630 18836 18630 18836 0 net9
rlabel metal2 20286 20672 20286 20672 0 rst_n
rlabel metal1 20516 18802 20516 18802 0 ui_in[0]
rlabel metal1 20378 19822 20378 19822 0 ui_in[1]
rlabel metal2 19826 20281 19826 20281 0 ui_in[2]
rlabel metal4 24196 20301 24196 20301 0 ui_in[3]
rlabel metal2 17986 21488 17986 21488 0 ui_in[4]
rlabel metal4 23092 22137 23092 22137 0 ui_in[5]
rlabel metal4 22540 20369 22540 20369 0 ui_in[6]
rlabel metal4 21988 22001 21988 22001 0 ui_in[7]
rlabel metal4 12604 20437 12604 20437 0 uio_out[0]
rlabel metal1 11684 19958 11684 19958 0 uio_out[1]
rlabel metal1 4002 19686 4002 19686 0 uio_out[2]
rlabel metal2 20746 21726 20746 21726 0 uio_out[3]
rlabel metal2 4554 20213 4554 20213 0 uio_out[4]
rlabel metal2 5106 20281 5106 20281 0 uio_out[5]
rlabel metal1 6072 19482 6072 19482 0 uio_out[6]
rlabel metal1 8602 16762 8602 16762 0 uio_out[7]
rlabel metal2 20654 19312 20654 19312 0 uo_out[0]
rlabel metal1 19642 18598 19642 18598 0 uo_out[1]
rlabel metal1 16744 17850 16744 17850 0 uo_out[2]
rlabel metal1 14628 17306 14628 17306 0 uo_out[3]
rlabel metal4 14812 22137 14812 22137 0 uo_out[4]
rlabel metal2 20010 19261 20010 19261 0 uo_out[5]
rlabel metal1 17342 19686 17342 19686 0 uo_out[6]
rlabel metal1 17342 21114 17342 21114 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 31464 22304
<< end >>
