VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ht_sc_tt05__mux2i_2
  CLASS CORE ;
  FOREIGN sky130_ht_sc_tt05__mux2i_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.055 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.014 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.075 3.535 1.275 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.170 ;
    ANTENNAGATEAREA 0.852 ;
    PORT
      LAYER li1 ;
        RECT 4.255 0.995 4.425 1.105 ;
        RECT 4.255 1.105 4.475 1.325 ;
        RECT 4.285 1.325 4.475 1.615 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.308 ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.765 0.785 0.995 ;
        RECT 0.445 0.995 0.785 1.275 ;
        RECT 0.445 1.275 0.615 1.325 ;
    END
  END S
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.170 ;
    PORT
      LAYER li1 ;
        RECT 2.715 0.295 4.965 0.465 ;
        RECT 4.795 0.465 4.965 1.785 ;
        RECT 4.735 1.785 4.965 2.255 ;
        RECT 2.715 2.255 4.965 2.425 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 2.275 2.175 2.445 2.255 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.355 2.255 1.685 2.635 ;
        RECT 2.275 2.255 2.445 2.635 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 1.855 1.835 2.965 1.915 ;
        RECT 1.855 1.915 4.355 2.005 ;
        RECT 1.855 2.005 2.025 2.085 ;
        RECT 2.795 2.005 4.355 2.085 ;
        RECT 1.855 2.085 2.025 2.465 ;
        RECT 0.095 0.255 0.345 0.585 ;
        RECT 0.095 0.585 0.265 1.075 ;
        RECT 0.095 1.075 0.265 1.155 ;
        RECT 1.435 1.075 1.955 1.155 ;
        RECT 0.095 1.155 0.265 1.245 ;
        RECT 1.015 1.155 1.955 1.245 ;
        RECT 0.095 1.245 0.265 1.325 ;
        RECT 1.015 1.245 1.605 1.325 ;
        RECT 0.095 1.325 0.265 1.495 ;
        RECT 1.015 1.325 1.185 1.495 ;
        RECT 0.095 1.495 1.185 1.665 ;
        RECT 0.095 1.665 0.265 2.135 ;
        RECT 0.095 2.135 0.345 2.465 ;
        RECT 1.435 1.495 3.465 1.665 ;
        RECT 1.435 1.665 1.605 1.745 ;
        RECT 3.135 1.665 3.465 1.745 ;
        RECT 1.435 1.745 1.605 1.835 ;
        RECT 0.935 1.835 1.605 2.005 ;
        RECT 1.015 0.555 1.245 0.965 ;
        RECT 3.815 0.635 4.355 0.805 ;
        RECT 3.815 0.805 4.005 0.935 ;
        RECT 1.855 0.255 2.025 0.635 ;
        RECT 1.855 0.635 2.025 0.715 ;
        RECT 3.135 0.635 3.465 0.715 ;
        RECT 1.855 0.715 3.465 0.885 ;
        RECT 0.000 -0.085 5.060 0.085 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 1.435 0.085 1.605 0.545 ;
        RECT 2.275 0.085 2.445 0.545 ;
        RECT 1.435 0.545 1.605 0.885 ;
      LAYER mcon ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 3.825 0.765 3.995 0.935 ;
        RECT 1.065 0.765 1.235 0.935 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
      LAYER met1 ;
        RECT 1.005 0.735 1.295 0.780 ;
        RECT 3.765 0.735 4.055 0.780 ;
        RECT 1.005 0.780 4.055 0.920 ;
        RECT 1.005 0.920 1.295 0.965 ;
        RECT 3.765 0.920 4.055 0.965 ;
  END
END sky130_ht_sc_tt05__mux2i_2
MACRO sky130_ht_sc_tt05__maj3_2
  CLASS CORE ;
  FOREIGN sky130_ht_sc_tt05__maj3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.135 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.842 ;
    PORT
      LAYER li1 ;
        RECT 1.055 0.995 1.225 1.105 ;
        RECT 1.055 1.105 1.695 1.275 ;
        RECT 1.055 1.275 1.225 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.842 ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.995 2.065 1.105 ;
        RECT 1.895 1.105 2.155 1.275 ;
        RECT 1.895 1.275 2.065 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.850 ;
    ANTENNAGATEAREA 0.416 ;
    PORT
      LAYER li1 ;
        RECT 0.435 0.995 0.745 1.105 ;
        RECT 2.535 0.995 2.705 1.105 ;
        RECT 0.435 1.105 0.775 1.325 ;
        RECT 2.445 1.105 2.705 1.325 ;
        RECT 0.605 1.325 0.775 1.575 ;
        RECT 2.445 1.325 2.615 1.575 ;
        RECT 0.605 1.575 2.615 1.745 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.502 ;
    PORT
      LAYER li1 ;
        RECT 3.285 0.295 3.615 0.805 ;
        RECT 3.445 0.805 3.615 1.575 ;
        RECT 3.285 1.575 3.615 2.425 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 3.785 1.495 3.955 1.915 ;
        RECT 2.705 1.915 3.035 2.255 ;
        RECT 3.785 1.915 3.955 2.255 ;
        RECT 0.985 2.255 1.315 2.635 ;
        RECT 2.705 2.255 3.035 2.635 ;
        RECT 3.785 2.255 3.955 2.635 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 0.295 0.435 0.635 ;
        RECT 1.825 0.295 2.155 0.635 ;
        RECT 0.085 0.635 3.115 0.805 ;
        RECT 0.085 0.805 0.255 0.995 ;
        RECT 2.945 0.805 3.115 0.995 ;
        RECT 0.085 0.995 0.255 1.245 ;
        RECT 2.945 0.995 3.225 1.245 ;
        RECT 0.085 1.245 0.255 1.325 ;
        RECT 3.055 1.245 3.225 1.325 ;
        RECT 0.085 1.325 0.255 1.915 ;
        RECT 0.085 1.915 2.155 2.085 ;
        RECT 0.085 2.085 0.435 2.425 ;
        RECT 1.825 2.085 2.155 2.425 ;
        RECT 0.000 -0.085 4.140 0.085 ;
        RECT 0.985 0.085 1.315 0.465 ;
        RECT 2.705 0.085 3.035 0.465 ;
        RECT 3.785 0.085 3.955 0.465 ;
        RECT 3.785 0.465 3.955 0.885 ;
      LAYER mcon ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
      LAYER met1 ;
  END
END sky130_ht_sc_tt05__maj3_2
MACRO sky130_ht_sc_tt05__dlrtp_1
  CLASS CORE ;
  FOREIGN sky130_ht_sc_tt05__dlrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.895 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.090 ;
    ANTENNAGATEAREA 0.476 ;
    PORT
      LAYER li1 ;
        RECT 0.145 0.995 0.315 1.105 ;
        RECT 0.135 1.105 0.325 1.615 ;
    END
  END GATE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.449 ;
    PORT
      LAYER li1 ;
        RECT 1.505 1.075 1.835 1.275 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.059 ;
    ANTENNAGATEAREA 0.416 ;
    PORT
      LAYER li1 ;
        RECT 5.655 0.425 5.845 1.075 ;
        RECT 5.655 1.075 5.995 1.245 ;
        RECT 5.655 1.245 5.845 1.275 ;
    END
  END RESET_B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.355 0.295 6.805 0.595 ;
        RECT 6.635 0.595 6.805 1.785 ;
        RECT 6.355 1.785 6.805 2.425 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 2.015 1.835 2.185 2.175 ;
        RECT 2.015 2.175 2.185 2.255 ;
        RECT 4.535 2.175 5.225 2.255 ;
        RECT 6.015 2.175 6.185 2.255 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 2.015 2.255 2.185 2.635 ;
        RECT 4.535 2.255 5.225 2.635 ;
        RECT 6.015 2.255 6.185 2.635 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 1.015 1.755 1.245 2.465 ;
        RECT 0.095 0.635 0.765 0.805 ;
        RECT 0.595 0.805 0.765 0.995 ;
        RECT 0.595 0.995 0.975 1.325 ;
        RECT 0.595 1.325 0.785 1.615 ;
        RECT 0.595 1.615 0.765 1.875 ;
        RECT 0.095 1.875 0.765 2.045 ;
        RECT 0.175 2.045 0.345 2.465 ;
        RECT 1.535 0.255 1.705 0.715 ;
        RECT 1.535 0.715 2.185 0.885 ;
        RECT 2.015 0.885 2.185 0.995 ;
        RECT 2.015 0.995 2.395 1.325 ;
        RECT 2.015 1.325 2.185 1.445 ;
        RECT 1.535 1.445 2.185 1.615 ;
        RECT 1.535 1.615 1.705 2.465 ;
        RECT 3.015 0.635 3.345 0.715 ;
        RECT 3.015 0.715 4.445 0.885 ;
        RECT 4.275 0.885 4.445 1.445 ;
        RECT 4.275 1.445 4.465 1.615 ;
        RECT 4.275 1.615 4.445 1.785 ;
        RECT 4.195 1.785 4.445 1.955 ;
        RECT 4.195 1.955 4.365 2.255 ;
        RECT 3.555 2.255 4.365 2.425 ;
        RECT 2.475 2.255 3.345 2.425 ;
        RECT 5.455 2.255 5.785 2.425 ;
        RECT 4.875 0.295 5.305 0.465 ;
        RECT 4.875 0.465 5.045 0.715 ;
        RECT 4.655 0.715 5.045 0.885 ;
        RECT 4.655 0.885 4.825 0.995 ;
        RECT 4.645 0.995 4.825 1.075 ;
        RECT 6.285 0.995 6.455 1.075 ;
        RECT 4.645 1.075 4.825 1.325 ;
        RECT 6.275 1.075 6.455 1.325 ;
        RECT 4.655 1.325 4.825 1.445 ;
        RECT 6.275 1.325 6.445 1.445 ;
        RECT 4.655 1.445 4.825 1.615 ;
        RECT 5.655 1.445 6.445 1.615 ;
        RECT 4.655 1.615 4.825 1.785 ;
        RECT 5.655 1.615 5.825 1.785 ;
        RECT 4.655 1.785 5.825 1.955 ;
        RECT 2.435 0.425 2.745 0.595 ;
        RECT 2.575 0.595 2.745 1.075 ;
        RECT 2.575 1.075 3.015 1.245 ;
        RECT 3.765 1.075 4.095 1.245 ;
        RECT 2.575 1.245 2.745 1.785 ;
        RECT 3.855 1.245 4.025 1.785 ;
        RECT 2.435 1.785 4.025 1.955 ;
        RECT 5.125 1.075 5.455 1.245 ;
        RECT 5.195 1.245 5.365 1.445 ;
        RECT 5.195 1.445 5.385 1.615 ;
        RECT 3.225 1.075 3.555 1.275 ;
        RECT 3.355 1.275 3.545 1.615 ;
        RECT 1.015 0.255 1.245 0.625 ;
        RECT 0.000 -0.085 6.900 0.085 ;
        RECT 0.515 0.085 0.845 0.465 ;
        RECT 1.935 0.085 2.265 0.465 ;
        RECT 4.535 0.085 4.705 0.465 ;
        RECT 6.015 0.085 6.185 0.465 ;
        RECT 4.535 0.465 4.705 0.545 ;
        RECT 6.015 0.465 6.185 0.545 ;
        RECT 3.555 0.295 4.365 0.465 ;
      LAYER mcon ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 1.065 1.785 1.235 1.955 ;
        RECT 2.445 1.785 2.615 1.955 ;
        RECT 3.365 1.445 3.535 1.615 ;
        RECT 4.285 1.445 4.455 1.615 ;
        RECT 5.205 1.445 5.375 1.615 ;
        RECT 0.605 1.445 0.775 1.615 ;
        RECT 2.445 0.425 2.615 0.595 ;
        RECT 1.065 0.425 1.235 0.595 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
      LAYER met1 ;
        RECT 1.005 1.755 1.295 1.800 ;
        RECT 2.385 1.755 2.675 1.800 ;
        RECT 1.005 1.800 2.675 1.940 ;
        RECT 1.005 1.940 1.295 1.985 ;
        RECT 2.385 1.940 2.675 1.985 ;
        RECT 0.545 1.415 0.835 1.460 ;
        RECT 3.305 1.415 3.595 1.460 ;
        RECT 0.545 1.460 3.595 1.600 ;
        RECT 0.545 1.600 0.835 1.645 ;
        RECT 3.305 1.600 3.595 1.645 ;
        RECT 4.225 1.415 4.515 1.460 ;
        RECT 5.145 1.415 5.435 1.460 ;
        RECT 4.225 1.460 5.435 1.600 ;
        RECT 4.225 1.600 4.515 1.645 ;
        RECT 5.145 1.600 5.435 1.645 ;
        RECT 1.005 0.395 1.295 0.440 ;
        RECT 2.385 0.395 2.675 0.440 ;
        RECT 1.005 0.440 2.675 0.580 ;
        RECT 1.005 0.580 1.295 0.625 ;
        RECT 2.385 0.580 2.675 0.625 ;
  END
END sky130_ht_sc_tt05__dlrtp_1
MACRO sky130_ht_sc_tt05__dfrtp_1
  CLASS CORE ;
  FOREIGN sky130_ht_sc_tt05__dfrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 10.580 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 10.580 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 10.575 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 10.770 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 10.580 2.960 ;
    END
  END VPWR
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.740 ;
    PORT
      LAYER li1 ;
        RECT 1.495 0.295 1.825 0.425 ;
        RECT 1.495 0.425 2.165 0.635 ;
        RECT 1.495 0.635 1.825 2.255 ;
        RECT 0.575 2.255 2.745 2.425 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.740 ;
    PORT
      LAYER li1 ;
        RECT 3.335 0.295 4.125 0.425 ;
        RECT 3.335 0.425 4.465 0.635 ;
        RECT 2.875 0.635 4.585 0.805 ;
        RECT 2.875 0.805 3.205 1.915 ;
        RECT 4.255 0.805 4.585 1.915 ;
        RECT 2.875 1.915 4.585 2.085 ;
        RECT 3.335 2.085 4.125 2.425 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.740 ;
    PORT
      LAYER li1 ;
        RECT 5.175 0.295 6.425 0.425 ;
        RECT 5.175 0.425 6.765 0.465 ;
        RECT 5.175 0.465 5.505 0.635 ;
        RECT 6.095 0.465 6.765 0.635 ;
        RECT 5.175 0.635 5.505 0.805 ;
        RECT 6.095 0.635 6.885 0.805 ;
        RECT 5.175 0.805 5.505 1.915 ;
        RECT 6.555 0.805 6.885 1.915 ;
        RECT 5.175 1.915 5.505 2.085 ;
        RECT 6.095 1.915 6.885 2.085 ;
        RECT 5.175 2.085 5.505 2.255 ;
        RECT 6.095 2.085 6.425 2.255 ;
        RECT 5.175 2.255 6.425 2.425 ;
    END
  END RESET_B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.740 ;
    PORT
      LAYER li1 ;
        RECT 7.935 0.295 8.725 0.425 ;
        RECT 7.935 0.425 9.065 0.635 ;
        RECT 7.475 0.635 9.185 0.805 ;
        RECT 7.475 0.805 7.805 1.915 ;
        RECT 8.855 0.805 9.185 1.915 ;
        RECT 7.475 1.915 9.185 2.085 ;
        RECT 7.935 2.085 8.725 2.425 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 0.000 2.635 10.580 2.805 ;
        RECT 0.000 -0.085 10.580 0.085 ;
      LAYER mcon ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 9.805 2.635 9.975 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 10.265 2.635 10.435 2.805 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 9.805 -0.085 9.975 0.085 ;
        RECT 10.265 -0.085 10.435 0.085 ;
      LAYER met1 ;
        RECT 5.220 0.440 6.280 0.580 ;
        RECT 5.220 0.580 5.360 0.780 ;
        RECT 6.140 0.580 6.280 0.780 ;
        RECT 5.220 0.780 5.360 0.920 ;
        RECT 6.140 0.780 6.740 0.920 ;
        RECT 5.220 0.920 5.360 1.800 ;
        RECT 6.600 0.920 6.740 1.800 ;
        RECT 5.220 1.800 5.360 1.940 ;
        RECT 6.140 1.800 6.740 1.940 ;
        RECT 5.220 1.940 5.360 2.140 ;
        RECT 6.140 1.940 6.280 2.140 ;
        RECT 5.220 2.140 6.280 2.280 ;
        RECT 1.540 0.440 1.680 2.140 ;
        RECT 0.620 2.140 2.600 2.280 ;
        RECT 3.380 0.440 3.980 0.580 ;
        RECT 3.380 0.580 3.520 0.780 ;
        RECT 3.840 0.580 3.980 0.780 ;
        RECT 2.920 0.780 3.520 0.920 ;
        RECT 3.840 0.780 4.440 0.920 ;
        RECT 2.920 0.920 3.060 1.800 ;
        RECT 4.300 0.920 4.440 1.800 ;
        RECT 2.920 1.800 3.520 1.940 ;
        RECT 3.840 1.800 4.440 1.940 ;
        RECT 3.380 1.940 3.520 2.140 ;
        RECT 3.840 1.940 3.980 2.140 ;
        RECT 3.380 2.140 3.980 2.280 ;
        RECT 7.980 0.440 8.580 0.580 ;
        RECT 7.980 0.580 8.120 0.780 ;
        RECT 8.440 0.580 8.580 0.780 ;
        RECT 7.520 0.780 8.120 0.920 ;
        RECT 8.440 0.780 9.040 0.920 ;
        RECT 7.520 0.920 7.660 1.800 ;
        RECT 8.900 0.920 9.040 1.800 ;
        RECT 7.520 1.800 8.120 1.940 ;
        RECT 8.440 1.800 9.040 1.940 ;
        RECT 7.980 1.940 8.120 2.140 ;
        RECT 8.440 1.940 8.580 2.140 ;
        RECT 7.980 2.140 8.580 2.280 ;
  END
END sky130_ht_sc_tt05__dfrtp_1
