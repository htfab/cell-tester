magic
tech sky130A
magscale 1 2
timestamp 1698685089
<< nwell >>
rect -38 261 2154 582
<< pwell >>
rect 1 21 2115 203
rect 29 -17 63 21
<< scnmos >>
rect 87 47 117 177
rect 179 47 209 177
rect 271 47 301 177
rect 363 47 393 177
rect 455 47 485 177
rect 547 47 577 177
rect 639 47 669 177
rect 731 47 761 177
rect 823 47 853 177
rect 915 47 945 177
rect 1007 47 1037 177
rect 1099 47 1129 177
rect 1191 47 1221 177
rect 1283 47 1313 177
rect 1375 47 1405 177
rect 1467 47 1497 177
rect 1559 47 1589 177
rect 1651 47 1681 177
rect 1743 47 1773 177
rect 1835 47 1865 177
rect 1927 47 1957 177
<< scpmoshvt >>
rect 87 297 117 497
rect 179 297 209 497
rect 271 297 301 497
rect 363 297 393 497
rect 455 297 485 497
rect 547 297 577 497
rect 639 297 669 497
rect 731 297 761 497
rect 823 297 853 497
rect 915 297 945 497
rect 1007 297 1037 497
rect 1099 297 1129 497
rect 1191 297 1221 497
rect 1283 297 1313 497
rect 1375 297 1405 497
rect 1467 297 1497 497
rect 1559 297 1589 497
rect 1651 297 1681 497
rect 1743 297 1773 497
rect 1835 297 1865 497
rect 1927 297 1957 497
<< ndiff >>
rect 1865 47 1927 177
rect 1037 47 1099 59
rect 1037 59 1051 93
rect 1085 59 1099 93
rect 1037 93 1099 127
rect 1037 127 1051 161
rect 1085 127 1099 161
rect 1037 161 1099 177
rect 117 47 179 177
rect 209 47 271 177
rect 301 47 363 59
rect 301 59 315 93
rect 349 59 363 93
rect 301 93 363 127
rect 301 127 315 161
rect 349 127 363 161
rect 301 161 363 177
rect 393 47 455 177
rect 485 47 547 177
rect 577 47 639 127
rect 577 127 591 161
rect 625 127 639 161
rect 577 161 639 177
rect 669 47 731 59
rect 669 59 683 93
rect 717 59 731 93
rect 669 93 731 127
rect 669 127 683 161
rect 717 127 731 161
rect 669 161 731 177
rect 761 47 823 59
rect 761 59 775 93
rect 809 59 823 93
rect 761 93 823 127
rect 761 127 775 161
rect 809 127 823 161
rect 761 161 823 177
rect 853 47 915 127
rect 853 127 867 161
rect 901 127 915 161
rect 853 161 915 177
rect 945 47 1007 177
rect 31 47 87 177
rect 1129 47 1191 59
rect 1129 59 1143 93
rect 1177 59 1191 93
rect 1129 93 1191 177
rect 1221 47 1283 59
rect 1221 59 1235 93
rect 1269 59 1283 93
rect 1221 93 1283 127
rect 1221 127 1235 161
rect 1269 127 1283 161
rect 1221 161 1283 177
rect 1313 47 1375 127
rect 1313 127 1327 161
rect 1361 127 1375 161
rect 1313 161 1375 177
rect 1405 47 1467 177
rect 1497 47 1559 127
rect 1497 127 1511 161
rect 1545 127 1559 161
rect 1497 161 1559 177
rect 1589 47 1651 59
rect 1589 59 1603 93
rect 1637 59 1651 93
rect 1589 93 1651 127
rect 1589 127 1603 161
rect 1637 127 1651 161
rect 1589 161 1651 177
rect 1681 47 1743 59
rect 1681 59 1695 93
rect 1729 59 1743 93
rect 1681 93 1743 127
rect 1681 127 1695 161
rect 1729 127 1743 161
rect 1681 161 1743 177
rect 1773 47 1835 127
rect 1773 127 1787 161
rect 1821 127 1835 161
rect 1773 161 1835 177
rect 1957 47 2013 177
<< pdiff >>
rect 1865 297 1927 497
rect 1957 297 2013 497
rect 31 297 87 497
rect 117 297 179 451
rect 117 451 131 485
rect 165 451 179 485
rect 117 485 179 497
rect 209 297 271 451
rect 209 451 223 485
rect 257 451 271 485
rect 209 485 271 497
rect 301 297 363 315
rect 301 315 315 349
rect 349 315 363 349
rect 301 349 363 383
rect 301 383 315 417
rect 349 383 363 417
rect 301 417 363 451
rect 301 451 315 485
rect 349 451 363 485
rect 301 485 363 497
rect 393 297 455 451
rect 393 451 407 485
rect 441 451 455 485
rect 393 485 455 497
rect 485 297 547 451
rect 485 451 499 485
rect 533 451 547 485
rect 485 485 547 497
rect 577 297 639 315
rect 577 315 591 349
rect 625 315 639 349
rect 577 349 639 383
rect 577 383 591 417
rect 625 383 639 417
rect 577 417 639 497
rect 669 297 731 383
rect 669 383 683 417
rect 717 383 731 417
rect 669 417 731 451
rect 669 451 683 485
rect 717 451 731 485
rect 669 485 731 497
rect 761 297 823 383
rect 761 383 775 417
rect 809 383 823 417
rect 761 417 823 451
rect 761 451 775 485
rect 809 451 823 485
rect 761 485 823 497
rect 853 297 915 315
rect 853 315 867 349
rect 901 315 915 349
rect 853 349 915 383
rect 853 383 867 417
rect 901 383 915 417
rect 853 417 915 497
rect 1037 297 1099 315
rect 1037 315 1051 349
rect 1085 315 1099 349
rect 1037 349 1099 383
rect 1037 383 1051 417
rect 1085 383 1099 417
rect 1037 417 1099 451
rect 1037 451 1051 485
rect 1085 451 1099 485
rect 1037 485 1099 497
rect 1129 297 1191 451
rect 1129 451 1143 485
rect 1177 451 1191 485
rect 1129 485 1191 497
rect 1221 297 1283 383
rect 1221 383 1235 417
rect 1269 383 1283 417
rect 1221 417 1283 451
rect 1221 451 1235 485
rect 1269 451 1283 485
rect 1221 485 1283 497
rect 1313 297 1375 315
rect 1313 315 1327 349
rect 1361 315 1375 349
rect 1313 349 1375 383
rect 1313 383 1327 417
rect 1361 383 1375 417
rect 1313 417 1375 497
rect 1405 297 1467 497
rect 1497 297 1559 315
rect 1497 315 1511 349
rect 1545 315 1559 349
rect 1497 349 1559 383
rect 1497 383 1511 417
rect 1545 383 1559 417
rect 1497 417 1559 497
rect 1589 297 1651 383
rect 1589 383 1603 417
rect 1637 383 1651 417
rect 1589 417 1651 451
rect 1589 451 1603 485
rect 1637 451 1651 485
rect 1589 485 1651 497
rect 1681 297 1743 383
rect 1681 383 1695 417
rect 1729 383 1743 417
rect 1681 417 1743 451
rect 1681 451 1695 485
rect 1729 451 1743 485
rect 1681 485 1743 497
rect 1773 297 1835 315
rect 1773 315 1787 349
rect 1821 315 1835 349
rect 1773 349 1835 383
rect 1773 383 1787 417
rect 1821 383 1835 417
rect 1773 417 1835 497
rect 945 297 1007 497
<< ndiffc >>
rect 591 127 625 161
rect 1511 127 1545 161
rect 1787 127 1821 161
rect 1695 127 1729 161
rect 1327 127 1361 161
rect 867 127 901 161
rect 1235 127 1269 161
rect 683 127 717 161
rect 1603 127 1637 161
rect 1051 127 1085 161
rect 775 127 809 161
rect 315 127 349 161
rect 1235 59 1269 93
rect 1603 59 1637 93
rect 1143 59 1177 93
rect 775 59 809 93
rect 683 59 717 93
rect 1695 59 1729 93
rect 1051 59 1085 93
rect 315 59 349 93
<< pdiffc >>
rect 1051 451 1085 485
rect 223 451 257 485
rect 1603 451 1637 485
rect 1143 451 1177 485
rect 775 451 809 485
rect 499 451 533 485
rect 131 451 165 485
rect 407 451 441 485
rect 683 451 717 485
rect 1235 451 1269 485
rect 315 451 349 485
rect 1695 451 1729 485
rect 1787 383 1821 417
rect 867 383 901 417
rect 1603 383 1637 417
rect 1051 383 1085 417
rect 683 383 717 417
rect 1695 383 1729 417
rect 315 383 349 417
rect 591 383 625 417
rect 1511 383 1545 417
rect 775 383 809 417
rect 1235 383 1269 417
rect 1327 383 1361 417
rect 1787 315 1821 349
rect 1051 315 1085 349
rect 1511 315 1545 349
rect 315 315 349 349
rect 1327 315 1361 349
rect 867 315 901 349
rect 591 315 625 349
<< poly >>
rect 1099 497 1129 523
rect 271 497 301 523
rect 363 497 393 523
rect 455 497 485 523
rect 547 497 577 523
rect 639 497 669 523
rect 731 497 761 523
rect 915 497 945 523
rect 1007 497 1037 523
rect 179 497 209 523
rect 1191 497 1221 523
rect 1283 497 1313 523
rect 1375 497 1405 523
rect 1467 497 1497 523
rect 1559 497 1589 523
rect 1651 497 1681 523
rect 1743 497 1773 523
rect 87 497 117 523
rect 1835 497 1865 523
rect 1927 497 1957 523
rect 823 497 853 523
rect 87 177 117 199
rect 179 177 209 199
rect 271 177 301 199
rect 363 177 393 199
rect 455 177 485 199
rect 547 177 577 199
rect 639 177 669 199
rect 731 177 761 199
rect 823 177 853 199
rect 915 177 945 199
rect 1007 177 1037 199
rect 1099 177 1129 199
rect 1191 177 1221 199
rect 1283 177 1313 199
rect 1375 177 1405 199
rect 1467 177 1497 199
rect 1559 177 1589 199
rect 1651 177 1681 199
rect 1743 177 1773 199
rect 1835 177 1865 199
rect 1927 177 1957 199
rect 75 199 1969 215
rect 75 215 315 249
rect 349 215 591 249
rect 625 215 867 249
rect 901 215 1051 249
rect 1085 215 1327 249
rect 1361 215 1511 249
rect 1545 215 1787 249
rect 1821 215 1969 249
rect 75 249 1969 265
rect 87 265 117 297
rect 179 265 209 297
rect 271 265 301 297
rect 363 265 393 297
rect 455 265 485 297
rect 547 265 577 297
rect 639 265 669 297
rect 731 265 761 297
rect 823 265 853 297
rect 915 265 945 297
rect 1007 265 1037 297
rect 1099 265 1129 297
rect 1191 265 1221 297
rect 1283 265 1313 297
rect 1375 265 1405 297
rect 1467 265 1497 297
rect 1559 265 1589 297
rect 1651 265 1681 297
rect 1743 265 1773 297
rect 1835 265 1865 297
rect 1927 265 1957 297
rect 1099 21 1129 47
rect 1927 21 1957 47
rect 1191 21 1221 47
rect 1283 21 1313 47
rect 1375 21 1405 47
rect 1467 21 1497 47
rect 1559 21 1589 47
rect 1651 21 1681 47
rect 1743 21 1773 47
rect 1835 21 1865 47
rect 1007 21 1037 47
rect 915 21 945 47
rect 87 21 117 47
rect 179 21 209 47
rect 271 21 301 47
rect 363 21 393 47
rect 455 21 485 47
rect 547 21 577 47
rect 639 21 669 47
rect 731 21 761 47
rect 823 21 853 47
<< polycont >>
rect 591 215 625 249
rect 1511 215 1545 249
rect 1327 215 1361 249
rect 1051 215 1085 249
rect 315 215 349 249
rect 867 215 901 249
rect 1787 215 1821 249
<< locali >>
rect 2087 527 2116 561
rect 1177 59 1235 85
rect 1269 59 1285 85
rect 1177 85 1235 93
rect 1269 85 1353 93
rect 1219 93 1353 127
rect 1219 127 1235 161
rect 1269 127 1327 161
rect 1361 127 1377 161
rect 1311 161 1377 215
rect 1311 215 1327 249
rect 1361 215 1377 249
rect 1311 249 1377 315
rect 1311 315 1327 349
rect 1361 315 1377 349
rect 1311 349 1377 383
rect 1219 383 1235 417
rect 1269 383 1327 417
rect 1361 383 1377 417
rect 1219 417 1285 451
rect 1177 451 1235 485
rect 1269 451 1285 485
rect 1035 59 1051 93
rect 1085 59 1143 93
rect 1035 93 1101 127
rect 1035 127 1051 161
rect 1085 127 1101 161
rect 1035 161 1101 215
rect 1035 215 1051 249
rect 1085 215 1101 249
rect 1035 249 1101 315
rect 1035 315 1051 349
rect 1085 315 1101 349
rect 1035 349 1101 383
rect 1035 383 1051 417
rect 1085 383 1101 417
rect 1035 417 1101 451
rect 1035 451 1051 485
rect 1085 451 1143 485
rect 299 59 315 85
rect 349 59 365 85
rect 299 85 315 93
rect 349 85 433 93
rect 299 93 433 127
rect 299 127 315 161
rect 349 127 365 161
rect 299 161 365 215
rect 299 215 315 249
rect 349 215 365 249
rect 299 249 365 315
rect 299 315 315 349
rect 349 315 365 349
rect 299 349 365 383
rect 299 383 315 417
rect 349 383 365 417
rect 299 417 365 451
rect 257 451 315 485
rect 349 451 407 485
rect 441 451 499 485
rect 533 451 549 485
rect 165 451 223 485
rect 115 451 131 485
rect 2087 -17 2116 17
rect 1995 527 2053 561
rect 1903 527 1961 561
rect 1811 527 1869 561
rect 1719 527 1777 561
rect 1627 527 1685 561
rect 1535 527 1593 561
rect 1443 527 1501 561
rect 1351 527 1409 561
rect 1259 527 1317 561
rect 1167 527 1225 561
rect 1075 527 1133 561
rect 983 527 1041 561
rect 891 527 949 561
rect 799 527 857 561
rect 707 527 765 561
rect 615 527 673 561
rect 523 527 581 561
rect 431 527 489 561
rect 339 527 397 561
rect 247 527 305 561
rect 155 527 213 561
rect 63 527 121 561
rect 0 527 29 561
rect 1587 59 1603 85
rect 1637 59 1695 85
rect 1729 59 1745 85
rect 1587 85 1603 93
rect 1637 85 1695 93
rect 1729 85 1813 93
rect 1587 93 1813 127
rect 1495 127 1511 161
rect 1545 127 1603 161
rect 1637 127 1695 161
rect 1729 127 1787 161
rect 1821 127 1837 161
rect 1495 161 1561 215
rect 1771 161 1837 215
rect 1495 215 1511 249
rect 1545 215 1561 249
rect 1771 215 1787 249
rect 1821 215 1837 249
rect 1495 249 1561 315
rect 1771 249 1837 315
rect 1495 315 1511 349
rect 1545 315 1561 349
rect 1771 315 1787 349
rect 1821 315 1837 349
rect 1495 349 1561 383
rect 1771 349 1837 383
rect 1495 383 1511 417
rect 1545 383 1603 417
rect 1637 383 1695 417
rect 1729 383 1787 417
rect 1821 383 1837 417
rect 1587 417 1745 451
rect 1587 451 1603 485
rect 1637 451 1695 485
rect 1729 451 1745 485
rect 667 59 683 85
rect 717 59 775 85
rect 809 59 825 85
rect 667 85 683 93
rect 717 85 775 93
rect 809 85 893 93
rect 667 93 893 127
rect 575 127 591 161
rect 625 127 683 161
rect 717 127 775 161
rect 809 127 867 161
rect 901 127 917 161
rect 575 161 641 215
rect 851 161 917 215
rect 575 215 591 249
rect 625 215 641 249
rect 851 215 867 249
rect 901 215 917 249
rect 575 249 641 315
rect 851 249 917 315
rect 575 315 591 349
rect 625 315 641 349
rect 851 315 867 349
rect 901 315 917 349
rect 575 349 641 383
rect 851 349 917 383
rect 575 383 591 417
rect 625 383 683 417
rect 717 383 775 417
rect 809 383 867 417
rect 901 383 917 417
rect 667 417 825 451
rect 667 451 683 485
rect 717 451 775 485
rect 809 451 825 485
rect 1995 -17 2053 17
rect 1903 -17 1961 17
rect 1811 -17 1869 17
rect 1719 -17 1777 17
rect 1627 -17 1685 17
rect 1535 -17 1593 17
rect 1443 -17 1501 17
rect 1351 -17 1409 17
rect 1259 -17 1317 17
rect 1167 -17 1225 17
rect 1075 -17 1133 17
rect 983 -17 1041 17
rect 891 -17 949 17
rect 799 -17 857 17
rect 707 -17 765 17
rect 615 -17 673 17
rect 523 -17 581 17
rect 431 -17 489 17
rect 339 -17 397 17
rect 247 -17 305 17
rect 155 -17 213 17
rect 63 -17 121 17
rect 0 -17 29 17
<< viali >>
rect 765 527 799 561
rect 213 527 247 561
rect 1685 527 1719 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1593 527 1627 561
rect 121 527 155 561
rect 1869 527 1903 561
rect 305 527 339 561
rect 857 527 891 561
rect 489 527 523 561
rect 949 527 983 561
rect 397 527 431 561
rect 1961 527 1995 561
rect 1409 527 1443 561
rect 1317 527 1351 561
rect 581 527 615 561
rect 29 527 63 561
rect 1777 527 1811 561
rect 1041 527 1075 561
rect 1501 527 1535 561
rect 673 527 707 561
rect 2053 527 2087 561
rect 1041 -17 1075 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 29 -17 63 17
rect 857 -17 891 17
rect 121 -17 155 17
rect 949 -17 983 17
rect 213 -17 247 17
rect 1501 -17 1535 17
rect 305 -17 339 17
rect 1593 -17 1627 17
rect 1133 -17 1167 17
rect 1685 -17 1719 17
rect 1225 -17 1259 17
rect 1777 -17 1811 17
rect 1317 -17 1351 17
rect 1869 -17 1903 17
rect 1409 -17 1443 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
<< metal1 >>
rect 0 496 2116 527
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 561 2116 592
rect 308 88 336 428
rect 124 428 520 456
rect 1044 88 1256 116
rect 1044 116 1072 156
rect 1228 116 1256 156
rect 1044 156 1072 184
rect 1228 156 1348 184
rect 1044 184 1072 360
rect 1320 184 1348 360
rect 1044 360 1072 388
rect 1228 360 1348 388
rect 1044 388 1072 428
rect 1228 388 1256 428
rect 1044 428 1256 456
rect 0 -48 2116 -17
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 17 2116 48
rect 676 88 796 116
rect 676 116 704 156
rect 768 116 796 156
rect 584 156 704 184
rect 768 156 888 184
rect 584 184 612 360
rect 860 184 888 360
rect 584 360 704 388
rect 768 360 888 388
rect 676 388 704 428
rect 768 388 796 428
rect 676 428 796 456
rect 1596 88 1716 116
rect 1596 116 1624 156
rect 1688 116 1716 156
rect 1504 156 1624 184
rect 1688 156 1808 184
rect 1504 184 1532 360
rect 1780 184 1808 360
rect 1504 360 1624 388
rect 1688 360 1808 388
rect 1596 388 1624 428
rect 1688 388 1716 428
rect 1596 428 1716 456
<< labels >>
flabel locali s 397 85 431 119 0 FreeSans 200 0 0 0 CLK
port 5 nsew signal input
flabel locali s 857 85 891 119 0 FreeSans 200 0 0 0 D
port 6 nsew signal input
flabel locali s 1317 85 1351 119 0 FreeSans 200 0 0 0 RESET_B
port 7 nsew signal input
flabel locali s 1777 85 1811 119 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 -48 2116 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2116 592 1 VPWR
port 4 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 dfrtp_1
<< properties >>
string FIXED_BBOX 0 0 2116 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ht_sc_tt05.gds
string GDS_START 24132
string GDS_END 35028
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
