magic
tech sky130A
magscale 1 2
timestamp 1698676621
<< nwell >>
rect -38 261 1050 582
<< pwell >>
rect 1 21 1011 203
rect 29 -17 63 21
<< scnmos >>
rect 603 47 633 177
rect 687 47 717 177
rect 775 47 805 177
rect 865 47 895 177
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
<< scpmoshvt >>
rect 603 297 633 497
rect 687 297 717 497
rect 775 297 805 497
rect 865 297 895 497
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
<< ndiff >>
rect 361 47 415 67
rect 361 67 371 101
rect 405 67 415 101
rect 361 101 415 177
rect 445 47 497 59
rect 445 59 455 93
rect 489 59 497 93
rect 445 93 497 177
rect 277 47 331 59
rect 277 59 287 93
rect 321 59 331 93
rect 277 93 331 127
rect 277 127 287 161
rect 321 127 331 161
rect 277 161 331 177
rect 193 47 247 127
rect 193 127 203 161
rect 237 127 247 161
rect 193 161 247 177
rect 109 47 163 59
rect 109 59 119 93
rect 153 59 163 93
rect 109 93 163 177
rect 895 47 985 59
rect 895 59 943 93
rect 977 59 985 93
rect 895 93 985 177
rect 805 47 865 127
rect 805 127 821 161
rect 855 127 865 161
rect 805 161 865 177
rect 717 47 775 59
rect 717 59 731 93
rect 765 59 775 93
rect 717 93 775 177
rect 633 47 687 127
rect 633 127 643 161
rect 677 127 687 161
rect 633 161 687 177
rect 551 47 603 59
rect 551 59 559 93
rect 593 59 603 93
rect 551 93 603 177
rect 27 47 79 67
rect 27 67 35 101
rect 69 67 79 101
rect 27 101 79 177
<< pdiff >>
rect 361 297 415 443
rect 361 443 371 477
rect 405 443 415 477
rect 361 477 415 497
rect 445 297 497 451
rect 445 451 455 485
rect 489 451 497 485
rect 445 485 497 497
rect 27 297 79 443
rect 27 443 35 477
rect 69 443 79 477
rect 27 477 79 497
rect 551 297 603 451
rect 551 451 559 485
rect 593 451 603 485
rect 551 485 603 497
rect 633 297 687 315
rect 633 315 643 349
rect 677 315 687 349
rect 633 349 687 497
rect 717 297 775 451
rect 717 451 731 485
rect 765 451 775 485
rect 717 485 775 497
rect 805 297 865 383
rect 805 383 821 417
rect 855 383 865 417
rect 805 417 865 497
rect 895 297 985 451
rect 895 451 943 485
rect 977 451 985 485
rect 895 485 985 497
rect 109 297 163 451
rect 109 451 119 485
rect 153 451 163 485
rect 109 485 163 497
rect 193 297 247 367
rect 193 367 203 401
rect 237 367 247 401
rect 193 401 247 497
rect 277 297 331 451
rect 277 451 287 485
rect 321 451 331 485
rect 277 485 331 497
<< ndiffc >>
rect 821 127 855 161
rect 643 127 677 161
rect 203 127 237 161
rect 287 127 321 161
rect 371 67 405 101
rect 35 67 69 101
rect 287 59 321 93
rect 943 59 977 93
rect 559 59 593 93
rect 455 59 489 93
rect 731 59 765 93
rect 119 59 153 93
<< pdiffc >>
rect 943 451 977 485
rect 455 451 489 485
rect 731 451 765 485
rect 287 451 321 485
rect 559 451 593 485
rect 119 451 153 485
rect 371 443 405 477
rect 35 443 69 477
rect 821 383 855 417
rect 203 367 237 401
rect 643 315 677 349
<< poly >>
rect 865 497 895 523
rect 603 497 633 523
rect 687 497 717 523
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 775 497 805 523
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 79 199 277 215
rect 79 215 89 249
rect 123 215 277 249
rect 79 249 277 265
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 177 361 199
rect 415 177 445 199
rect 331 199 445 215
rect 331 215 341 249
rect 375 215 445 249
rect 331 249 445 265
rect 331 265 361 297
rect 415 265 445 297
rect 603 177 633 199
rect 687 177 717 199
rect 499 199 717 215
rect 499 215 509 249
rect 543 215 577 249
rect 611 215 645 249
rect 679 215 717 249
rect 499 249 717 265
rect 603 265 633 297
rect 687 265 717 297
rect 775 177 805 199
rect 865 177 895 199
rect 775 199 895 215
rect 775 215 851 249
rect 885 215 895 249
rect 775 249 895 265
rect 775 265 805 297
rect 865 265 895 297
rect 775 21 805 47
rect 687 21 717 47
rect 603 21 633 47
rect 865 21 895 47
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
<< polycont >>
rect 645 215 679 249
rect 509 215 543 249
rect 89 215 123 249
rect 577 215 611 249
rect 851 215 885 249
rect 341 215 375 249
<< locali >>
rect 103 451 119 485
rect 153 451 169 485
rect 103 485 169 527
rect 63 527 121 561
rect 155 527 213 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 19 51 69 67
rect 19 67 35 101
rect 19 101 69 117
rect 19 117 53 215
rect 19 215 53 231
rect 287 215 341 231
rect 19 231 53 249
rect 203 231 341 249
rect 19 249 53 265
rect 203 249 321 265
rect 19 265 53 299
rect 203 265 237 299
rect 19 299 237 333
rect 19 333 53 427
rect 19 427 69 443
rect 19 443 35 477
rect 19 477 69 493
rect 371 477 405 493
rect 543 451 559 485
rect 977 59 993 93
rect 959 93 993 357
rect 947 357 993 451
rect 977 451 993 485
rect 765 451 943 485
rect 593 451 731 485
rect 455 435 489 451
rect 371 367 593 383
rect 371 383 821 401
rect 371 401 405 417
rect 559 401 821 417
rect 371 417 405 443
rect 855 383 871 417
rect 187 367 203 401
rect 287 299 693 315
rect 287 315 643 333
rect 677 315 693 333
rect 287 333 321 349
rect 627 333 643 349
rect 677 333 693 349
rect 287 349 321 367
rect 237 367 321 401
rect 885 221 895 249
rect 851 249 895 265
rect 857 265 895 323
rect 119 153 157 199
rect 89 199 157 215
rect 123 215 157 249
rect 89 249 157 255
rect 89 255 123 265
rect 489 215 509 249
rect 543 215 577 249
rect 611 215 645 249
rect 679 215 707 249
rect 489 249 707 255
rect 375 215 391 249
rect 851 199 885 215
rect 203 111 249 127
rect 237 127 249 153
rect 247 153 249 161
rect 203 161 213 187
rect 247 161 249 187
rect 203 187 249 193
rect 763 127 821 153
rect 763 153 765 161
rect 799 153 821 161
rect 763 161 765 187
rect 799 161 801 187
rect 371 101 405 127
rect 371 127 405 143
rect 627 127 643 143
rect 677 127 693 143
rect 371 143 643 161
rect 677 143 693 161
rect 371 161 693 177
rect 287 161 321 177
rect 855 127 871 161
rect 287 93 321 127
rect 119 93 153 109
rect 455 93 489 109
rect 543 59 559 93
rect 765 59 943 93
rect 593 59 731 93
rect 371 51 405 67
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 527 29 561
rect 271 451 287 485
rect 321 451 337 485
rect 271 485 337 527
rect 247 527 305 561
rect 455 485 489 527
rect 431 527 489 561
rect 339 527 397 561
rect 523 -17 581 17
rect 431 -17 489 17
rect 455 17 489 59
rect 339 -17 397 17
rect 247 -17 305 17
rect 287 17 321 59
rect 63 -17 121 17
rect 155 -17 213 17
rect 119 17 153 59
rect 0 -17 29 17
<< viali >>
rect 949 527 983 561
rect 857 527 891 561
rect 765 527 799 561
rect 673 527 707 561
rect 581 527 615 561
rect 489 527 523 561
rect 397 527 431 561
rect 305 527 339 561
rect 213 527 247 561
rect 121 527 155 561
rect 29 527 63 561
rect 765 153 799 187
rect 213 153 247 187
rect 305 -17 339 17
rect 949 -17 983 17
rect 581 -17 615 17
rect 213 -17 247 17
rect 857 -17 891 17
rect 489 -17 523 17
rect 121 -17 155 17
rect 765 -17 799 17
rect 397 -17 431 17
rect 29 -17 63 17
rect 673 -17 707 17
<< metal1 >>
rect 0 496 1012 527
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1012 561
rect 0 561 1012 592
rect 201 147 259 153
rect 753 147 811 153
rect 201 153 213 156
rect 247 153 259 156
rect 753 153 765 156
rect 799 153 811 156
rect 201 156 213 184
rect 247 156 765 184
rect 799 156 811 184
rect 201 184 213 187
rect 247 184 259 187
rect 753 184 765 187
rect 799 184 811 187
rect 201 187 259 193
rect 753 187 811 193
rect 0 -48 1012 -17
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1012 17
rect 0 17 1012 48
<< labels >>
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 A0
port 5 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 A0
port 5 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 200 0 0 0 A0
port 5 nsew signal input
flabel locali s 857 221 891 255 0 FreeSans 200 0 0 0 A1
port 6 nsew signal input
flabel locali s 857 289 891 323 0 FreeSans 200 0 0 0 A1
port 6 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 S
port 7 nsew signal input
flabel locali s 949 357 983 391 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 949 425 983 459 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 -48 1012 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1012 592 1 VPWR
port 4 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 mux2i_2
<< properties >>
string FIXED_BBOX 0 0 1012 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ht_sc_tt05.gds
string GDS_START 134
string GDS_END 7254
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
