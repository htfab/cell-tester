magic
tech sky130A
magscale 1 2
timestamp 1699069689
<< viali >>
rect 12817 21641 12851 21675
rect 18429 21641 18463 21675
rect 23213 21641 23247 21675
rect 5089 21573 5123 21607
rect 18981 21573 19015 21607
rect 21925 21573 21959 21607
rect 26065 21573 26099 21607
rect 949 21505 983 21539
rect 1455 21505 1489 21539
rect 3712 21505 3746 21539
rect 6288 21505 6322 21539
rect 6561 21505 6595 21539
rect 8864 21503 8898 21537
rect 9137 21505 9171 21539
rect 11440 21505 11474 21539
rect 14289 21505 14323 21539
rect 16129 21505 16163 21539
rect 16773 21505 16807 21539
rect 22318 21505 22352 21539
rect 22477 21505 22511 21539
rect 23857 21505 23891 21539
rect 24041 21505 24075 21539
rect 24501 21505 24535 21539
rect 24777 21505 24811 21539
rect 26709 21505 26743 21539
rect 27215 21505 27249 21539
rect 1685 21437 1719 21471
rect 3249 21437 3283 21471
rect 3985 21437 4019 21471
rect 5641 21437 5675 21471
rect 5825 21437 5859 21471
rect 8217 21437 8251 21471
rect 8401 21437 8435 21471
rect 8728 21437 8762 21471
rect 10793 21437 10827 21471
rect 10977 21437 11011 21471
rect 11304 21437 11338 21471
rect 11713 21437 11747 21471
rect 13369 21437 13403 21471
rect 14565 21437 14599 21471
rect 16681 21437 16715 21471
rect 16865 21437 16899 21471
rect 17141 21437 17175 21471
rect 18705 21437 18739 21471
rect 19349 21437 19383 21471
rect 19441 21437 19475 21471
rect 19717 21437 19751 21471
rect 21281 21437 21315 21471
rect 21465 21437 21499 21471
rect 22201 21437 22235 21471
rect 23121 21437 23155 21471
rect 23397 21437 23431 21471
rect 23581 21437 23615 21471
rect 23673 21437 23707 21471
rect 24915 21437 24949 21471
rect 25053 21437 25087 21471
rect 25881 21437 25915 21471
rect 26617 21437 26651 21471
rect 27036 21437 27070 21471
rect 27445 21437 27479 21471
rect 29101 21437 29135 21471
rect 30113 21437 30147 21471
rect 3065 21369 3099 21403
rect 13645 21369 13679 21403
rect 15945 21369 15979 21403
rect 29469 21369 29503 21403
rect 29653 21369 29687 21403
rect 1415 21301 1449 21335
rect 3715 21301 3749 21335
rect 5457 21301 5491 21335
rect 6291 21301 6325 21335
rect 7665 21301 7699 21335
rect 8033 21301 8067 21335
rect 10241 21301 10275 21335
rect 10609 21301 10643 21335
rect 13185 21301 13219 21335
rect 13737 21301 13771 21335
rect 19165 21301 19199 21335
rect 21005 21301 21039 21335
rect 25697 21301 25731 21335
rect 26433 21301 26467 21335
rect 28549 21301 28583 21335
rect 29929 21301 29963 21335
rect 30297 21301 30331 21335
rect 10149 21097 10183 21131
rect 11719 21097 11753 21131
rect 13645 21097 13679 21131
rect 15945 21097 15979 21131
rect 18797 21097 18831 21131
rect 20821 21097 20855 21131
rect 23121 21097 23155 21131
rect 25329 21097 25363 21131
rect 30481 21097 30515 21131
rect 1593 21029 1627 21063
rect 1961 21029 1995 21063
rect 2145 21029 2179 21063
rect 5273 21029 5307 21063
rect 28089 21029 28123 21063
rect 949 20961 983 20995
rect 1225 20961 1259 20995
rect 2932 20961 2966 20995
rect 4813 20961 4847 20995
rect 6009 20961 6043 20995
rect 6193 20961 6227 20995
rect 6474 20961 6508 20995
rect 8125 20961 8159 20995
rect 10701 20961 10735 20995
rect 11161 20961 11195 20995
rect 11253 20961 11287 20995
rect 11989 20961 12023 20995
rect 13553 20961 13587 20995
rect 14105 20961 14139 20995
rect 14381 20961 14415 20995
rect 16129 20961 16163 20995
rect 17969 20961 18003 20995
rect 18429 20961 18463 20995
rect 18705 20961 18739 20995
rect 21005 20961 21039 20995
rect 23305 20961 23339 20995
rect 25513 20961 25547 20995
rect 25697 20961 25731 20995
rect 28365 20961 28399 20995
rect 2605 20893 2639 20927
rect 3101 20911 3135 20945
rect 3341 20893 3375 20927
rect 5549 20893 5583 20927
rect 8309 20893 8343 20927
rect 8636 20893 8670 20927
rect 8772 20893 8806 20927
rect 9045 20893 9079 20927
rect 11716 20893 11750 20927
rect 16405 20893 16439 20927
rect 18981 20893 19015 20927
rect 19257 20893 19291 20927
rect 21281 20893 21315 20927
rect 21557 20893 21591 20927
rect 23489 20893 23523 20927
rect 23765 20893 23799 20927
rect 25973 20893 26007 20927
rect 26433 20893 26467 20927
rect 26709 20893 26743 20927
rect 28457 20893 28491 20927
rect 28784 20893 28818 20927
rect 28963 20893 28997 20927
rect 29193 20893 29227 20927
rect 15669 20825 15703 20859
rect 28181 20825 28215 20859
rect 2421 20757 2455 20791
rect 4445 20757 4479 20791
rect 4997 20757 5031 20791
rect 5825 20757 5859 20791
rect 7573 20757 7607 20791
rect 7941 20757 7975 20791
rect 10517 20757 10551 20791
rect 10977 20757 11011 20791
rect 13093 20757 13127 20791
rect 17509 20757 17543 20791
rect 3709 20553 3743 20587
rect 5917 20553 5951 20587
rect 7941 20553 7975 20587
rect 10517 20553 10551 20587
rect 13093 20553 13127 20587
rect 16037 20553 16071 20587
rect 19073 20553 19107 20587
rect 28549 20553 28583 20587
rect 26341 20485 26375 20519
rect 1363 20417 1397 20451
rect 4399 20417 4433 20451
rect 4629 20417 4663 20451
rect 6607 20415 6641 20449
rect 6837 20417 6871 20451
rect 8999 20417 9033 20451
rect 11164 20417 11198 20451
rect 14105 20417 14139 20451
rect 16405 20417 16439 20451
rect 18705 20417 18739 20451
rect 19349 20417 19383 20451
rect 21833 20417 21867 20451
rect 24133 20417 24167 20451
rect 27215 20417 27249 20451
rect 30389 20417 30423 20451
rect 857 20349 891 20383
rect 1593 20349 1627 20383
rect 3893 20349 3927 20383
rect 6101 20349 6135 20383
rect 8493 20349 8527 20383
rect 9229 20349 9263 20383
rect 10701 20349 10735 20383
rect 11437 20349 11471 20383
rect 14289 20349 14323 20383
rect 16129 20349 16163 20383
rect 18889 20349 18923 20383
rect 21373 20349 21407 20383
rect 21557 20349 21591 20383
rect 23581 20349 23615 20383
rect 23857 20349 23891 20383
rect 25881 20349 25915 20383
rect 26157 20349 26191 20383
rect 26709 20349 26743 20383
rect 27445 20349 27479 20383
rect 29469 20349 29503 20383
rect 29837 20349 29871 20383
rect 3433 20281 3467 20315
rect 13001 20281 13035 20315
rect 13829 20281 13863 20315
rect 14565 20281 14599 20315
rect 17969 20281 18003 20315
rect 19625 20281 19659 20315
rect 29101 20281 29135 20315
rect 30113 20281 30147 20315
rect 1323 20213 1357 20247
rect 2881 20213 2915 20247
rect 4359 20213 4393 20247
rect 6567 20213 6601 20247
rect 8959 20213 8993 20247
rect 11167 20213 11201 20247
rect 12541 20213 12575 20247
rect 17509 20213 17543 20247
rect 18061 20213 18095 20247
rect 21189 20213 21223 20247
rect 23397 20213 23431 20247
rect 25697 20213 25731 20247
rect 27175 20213 27209 20247
rect 29929 20213 29963 20247
rect 8959 20009 8993 20043
rect 11897 20009 11931 20043
rect 12639 20009 12673 20043
rect 14013 20009 14047 20043
rect 15485 20009 15519 20043
rect 16773 20009 16807 20043
rect 20085 20009 20119 20043
rect 20545 20009 20579 20043
rect 21097 20009 21131 20043
rect 24041 20009 24075 20043
rect 28831 20009 28865 20043
rect 2973 19941 3007 19975
rect 8033 19941 8067 19975
rect 1184 19873 1218 19907
rect 5641 19873 5675 19907
rect 8125 19873 8159 19907
rect 8493 19873 8527 19907
rect 10977 19873 11011 19907
rect 11253 19873 11287 19907
rect 12909 19873 12943 19907
rect 14657 19873 14691 19907
rect 15945 19873 15979 19907
rect 16313 19873 16347 19907
rect 16497 19873 16531 19907
rect 18613 19873 18647 19907
rect 18981 19873 19015 19907
rect 20637 19873 20671 19907
rect 20913 19873 20947 19907
rect 21557 19873 21591 19907
rect 21833 19873 21867 19907
rect 22201 19873 22235 19907
rect 24225 19873 24259 19907
rect 26065 19873 26099 19907
rect 26709 19873 26743 19907
rect 28365 19873 28399 19907
rect 30481 19873 30515 19907
rect 857 19805 891 19839
rect 1363 19805 1397 19839
rect 1593 19805 1627 19839
rect 3065 19805 3099 19839
rect 3392 19805 3426 19839
rect 3571 19807 3605 19841
rect 3801 19805 3835 19839
rect 5917 19805 5951 19839
rect 6244 19805 6278 19839
rect 6380 19805 6414 19839
rect 6653 19805 6687 19839
rect 8972 19823 9006 19857
rect 9229 19805 9263 19839
rect 12173 19805 12207 19839
rect 12636 19805 12670 19839
rect 14381 19805 14415 19839
rect 16221 19805 16255 19839
rect 16957 19805 16991 19839
rect 17233 19805 17267 19839
rect 18705 19805 18739 19839
rect 22477 19805 22511 19839
rect 24409 19805 24443 19839
rect 24685 19805 24719 19839
rect 26433 19805 26467 19839
rect 28871 19805 28905 19839
rect 29101 19805 29135 19839
rect 5089 19669 5123 19703
rect 5457 19669 5491 19703
rect 8309 19669 8343 19703
rect 10333 19669 10367 19703
rect 12081 19669 12115 19703
rect 15669 19669 15703 19703
rect 15761 19669 15795 19703
rect 21373 19669 21407 19703
rect 27997 19669 28031 19703
rect 10241 19465 10275 19499
rect 11069 19465 11103 19499
rect 13093 19465 13127 19499
rect 18061 19465 18095 19499
rect 949 19329 983 19363
rect 1445 19311 1479 19345
rect 3249 19329 3283 19363
rect 3755 19329 3789 19363
rect 5920 19329 5954 19363
rect 8864 19329 8898 19363
rect 11759 19329 11793 19363
rect 14016 19329 14050 19363
rect 15945 19329 15979 19363
rect 18705 19329 18739 19363
rect 22063 19329 22097 19363
rect 24501 19329 24535 19363
rect 25191 19329 25225 19363
rect 1685 19261 1719 19295
rect 3576 19261 3610 19295
rect 3985 19261 4019 19295
rect 5365 19261 5399 19295
rect 5457 19261 5491 19295
rect 6193 19261 6227 19295
rect 7573 19261 7607 19295
rect 7757 19261 7791 19295
rect 8401 19261 8435 19295
rect 9137 19261 9171 19295
rect 11253 19261 11287 19295
rect 11989 19261 12023 19295
rect 13553 19261 13587 19295
rect 14289 19261 14323 19295
rect 16221 19261 16255 19295
rect 17601 19261 17635 19295
rect 18245 19261 18279 19295
rect 18521 19261 18555 19295
rect 18981 19261 19015 19295
rect 20545 19261 20579 19295
rect 21557 19261 21591 19295
rect 22293 19261 22327 19295
rect 24225 19261 24259 19295
rect 24317 19261 24351 19295
rect 24685 19261 24719 19295
rect 25421 19261 25455 19295
rect 26893 19261 26927 19295
rect 27169 19261 27203 19295
rect 28641 19261 28675 19295
rect 28733 19261 28767 19295
rect 29009 19261 29043 19295
rect 29285 19261 29319 19295
rect 30573 19261 30607 19295
rect 8033 19193 8067 19227
rect 10793 19193 10827 19227
rect 17785 19193 17819 19227
rect 20729 19193 20763 19227
rect 29929 19193 29963 19227
rect 1415 19125 1449 19159
rect 2973 19125 3007 19159
rect 5923 19125 5957 19159
rect 8867 19125 8901 19159
rect 11719 19125 11753 19159
rect 14019 19125 14053 19159
rect 15393 19125 15427 19159
rect 17877 19125 17911 19159
rect 18337 19125 18371 19159
rect 20085 19125 20119 19159
rect 20821 19125 20855 19159
rect 21097 19125 21131 19159
rect 22023 19125 22057 19159
rect 23581 19125 23615 19159
rect 23857 19125 23891 19159
rect 25151 19125 25185 19159
rect 26525 19125 26559 19159
rect 28273 19125 28307 19159
rect 30113 19125 30147 19159
rect 30389 19125 30423 19159
rect 857 18921 891 18955
rect 4261 18921 4295 18955
rect 9143 18921 9177 18955
rect 10701 18921 10735 18955
rect 15853 18921 15887 18955
rect 21465 18921 21499 18955
rect 22391 18921 22425 18955
rect 24599 18921 24633 18955
rect 25973 18921 26007 18955
rect 26899 18921 26933 18955
rect 30481 18921 30515 18955
rect 1409 18853 1443 18887
rect 4721 18853 4755 18887
rect 5457 18853 5491 18887
rect 8033 18853 8067 18887
rect 20545 18853 20579 18887
rect 1041 18785 1075 18819
rect 1133 18785 1167 18819
rect 1777 18785 1811 18819
rect 2748 18785 2782 18819
rect 5181 18785 5215 18819
rect 6653 18785 6687 18819
rect 8217 18785 8251 18819
rect 8585 18785 8619 18819
rect 11161 18785 11195 18819
rect 11345 18785 11379 18819
rect 14197 18785 14231 18819
rect 14289 18785 14323 18819
rect 16405 18785 16439 18819
rect 16497 18785 16531 18819
rect 17233 18785 17267 18819
rect 18613 18785 18647 18819
rect 18981 18785 19015 18819
rect 21373 18785 21407 18819
rect 21925 18785 21959 18819
rect 24869 18785 24903 18819
rect 28641 18785 28675 18819
rect 28917 18785 28951 18819
rect 2421 18717 2455 18751
rect 2884 18719 2918 18753
rect 3157 18717 3191 18751
rect 5917 18717 5951 18751
rect 6244 18717 6278 18751
rect 6380 18717 6414 18751
rect 8677 18717 8711 18751
rect 9183 18717 9217 18751
rect 9413 18717 9447 18751
rect 11805 18717 11839 18751
rect 12132 18717 12166 18751
rect 12311 18717 12345 18751
rect 12541 18717 12575 18751
rect 14565 18717 14599 18751
rect 16221 18717 16255 18751
rect 16957 18717 16991 18751
rect 18705 18717 18739 18751
rect 20821 18717 20855 18751
rect 22388 18719 22422 18753
rect 22661 18717 22695 18751
rect 24133 18717 24167 18751
rect 24639 18717 24673 18751
rect 26433 18717 26467 18751
rect 26939 18717 26973 18751
rect 27169 18717 27203 18751
rect 1961 18649 1995 18683
rect 16773 18649 16807 18683
rect 30205 18649 30239 18683
rect 4813 18581 4847 18615
rect 10977 18581 11011 18615
rect 11437 18581 11471 18615
rect 13645 18581 13679 18615
rect 14013 18581 14047 18615
rect 20085 18581 20119 18615
rect 23949 18581 23983 18615
rect 28273 18581 28307 18615
rect 2973 18377 3007 18411
rect 5917 18377 5951 18411
rect 12633 18377 12667 18411
rect 17233 18377 17267 18411
rect 22201 18377 22235 18411
rect 22937 18377 22971 18411
rect 28273 18377 28307 18411
rect 30389 18377 30423 18411
rect 23305 18309 23339 18343
rect 28641 18309 28675 18343
rect 949 18241 983 18275
rect 1455 18241 1489 18275
rect 4220 18241 4254 18275
rect 4356 18241 4390 18275
rect 4629 18241 4663 18275
rect 6564 18241 6598 18275
rect 8585 18241 8619 18275
rect 9048 18241 9082 18275
rect 10701 18241 10735 18275
rect 11256 18241 11290 18275
rect 11529 18241 11563 18275
rect 14049 18223 14083 18257
rect 15853 18241 15887 18275
rect 16129 18241 16163 18275
rect 18521 18241 18555 18275
rect 20177 18241 20211 18275
rect 20867 18241 20901 18275
rect 24685 18241 24719 18275
rect 25148 18241 25182 18275
rect 26893 18241 26927 18275
rect 1685 18173 1719 18207
rect 3341 18173 3375 18207
rect 3893 18173 3927 18207
rect 6101 18173 6135 18207
rect 6837 18173 6871 18207
rect 9321 18173 9355 18207
rect 10793 18173 10827 18207
rect 13369 18173 13403 18207
rect 13553 18173 13587 18207
rect 14289 18173 14323 18207
rect 18061 18173 18095 18207
rect 18429 18173 18463 18207
rect 20361 18173 20395 18207
rect 21097 18173 21131 18207
rect 23121 18173 23155 18207
rect 23673 18173 23707 18207
rect 24317 18173 24351 18207
rect 24593 18173 24627 18207
rect 25421 18173 25455 18207
rect 27169 18173 27203 18207
rect 28825 18173 28859 18207
rect 29009 18173 29043 18207
rect 29285 18173 29319 18207
rect 30113 18173 30147 18207
rect 30573 18173 30607 18207
rect 8217 18105 8251 18139
rect 17693 18105 17727 18139
rect 19073 18105 19107 18139
rect 22661 18105 22695 18139
rect 23949 18105 23983 18139
rect 1415 18037 1449 18071
rect 3617 18037 3651 18071
rect 6567 18037 6601 18071
rect 9051 18037 9085 18071
rect 11259 18037 11293 18071
rect 13185 18037 13219 18071
rect 14019 18037 14053 18071
rect 15577 18037 15611 18071
rect 20827 18037 20861 18071
rect 23489 18037 23523 18071
rect 24409 18037 24443 18071
rect 25151 18037 25185 18071
rect 26525 18037 26559 18071
rect 30297 18037 30331 18071
rect 1415 17833 1449 17867
rect 2789 17833 2823 17867
rect 3157 17833 3191 17867
rect 3991 17833 4025 17867
rect 6193 17833 6227 17867
rect 10977 17833 11011 17867
rect 11621 17833 11655 17867
rect 16589 17833 16623 17867
rect 23581 17833 23615 17867
rect 23857 17833 23891 17867
rect 24599 17833 24633 17867
rect 5641 17765 5675 17799
rect 8585 17765 8619 17799
rect 16313 17765 16347 17799
rect 28917 17765 28951 17799
rect 949 17697 983 17731
rect 3341 17697 3375 17731
rect 6101 17697 6135 17731
rect 6377 17697 6411 17731
rect 10793 17697 10827 17731
rect 11161 17697 11195 17731
rect 11345 17697 11379 17731
rect 12541 17697 12575 17731
rect 14197 17697 14231 17731
rect 17693 17697 17727 17731
rect 19165 17697 19199 17731
rect 19441 17697 19475 17731
rect 21097 17697 21131 17731
rect 21281 17697 21315 17731
rect 21608 17697 21642 17731
rect 22017 17697 22051 17731
rect 23765 17697 23799 17731
rect 24041 17697 24075 17731
rect 24869 17697 24903 17731
rect 26433 17697 26467 17731
rect 26760 17697 26794 17731
rect 27169 17697 27203 17731
rect 1445 17647 1479 17681
rect 1685 17629 1719 17663
rect 3525 17629 3559 17663
rect 3988 17647 4022 17681
rect 4261 17629 4295 17663
rect 6469 17629 6503 17663
rect 6796 17629 6830 17663
rect 6932 17631 6966 17665
rect 7205 17629 7239 17663
rect 8677 17629 8711 17663
rect 9004 17629 9038 17663
rect 9140 17631 9174 17665
rect 9413 17629 9447 17663
rect 11805 17629 11839 17663
rect 12132 17629 12166 17663
rect 12311 17629 12345 17663
rect 14289 17629 14323 17663
rect 14565 17629 14599 17663
rect 16957 17629 16991 17663
rect 17284 17629 17318 17663
rect 17463 17631 17497 17665
rect 21744 17629 21778 17663
rect 24133 17629 24167 17663
rect 24639 17631 24673 17665
rect 26896 17631 26930 17665
rect 28641 17629 28675 17663
rect 5917 17561 5951 17595
rect 15853 17561 15887 17595
rect 13645 17493 13679 17527
rect 14013 17493 14047 17527
rect 18797 17493 18831 17527
rect 20729 17493 20763 17527
rect 20913 17493 20947 17527
rect 23121 17493 23155 17527
rect 25973 17493 26007 17527
rect 28273 17493 28307 17527
rect 30389 17493 30423 17527
rect 2789 17289 2823 17323
rect 10517 17289 10551 17323
rect 10885 17289 10919 17323
rect 16037 17289 16071 17323
rect 18981 17289 19015 17323
rect 19257 17289 19291 17323
rect 25605 17289 25639 17323
rect 30389 17289 30423 17323
rect 8401 17221 8435 17255
rect 14013 17221 14047 17255
rect 19533 17221 19567 17255
rect 1455 17153 1489 17187
rect 3893 17153 3927 17187
rect 4399 17153 4433 17187
rect 6009 17153 6043 17187
rect 6564 17153 6598 17187
rect 8677 17153 8711 17187
rect 9140 17151 9174 17185
rect 9413 17153 9447 17187
rect 11253 17153 11287 17187
rect 11759 17153 11793 17187
rect 14703 17153 14737 17187
rect 16911 17153 16945 17187
rect 18705 17153 18739 17187
rect 20867 17153 20901 17187
rect 23489 17153 23523 17187
rect 24133 17153 24167 17187
rect 25513 17153 25547 17187
rect 26387 17153 26421 17187
rect 28181 17153 28215 17187
rect 29837 17153 29871 17187
rect 949 17085 983 17119
rect 1685 17085 1719 17119
rect 3249 17085 3283 17119
rect 4629 17085 4663 17119
rect 6101 17085 6135 17119
rect 6428 17085 6462 17119
rect 6837 17085 6871 17119
rect 8585 17085 8619 17119
rect 11069 17085 11103 17119
rect 11989 17085 12023 17119
rect 14197 17085 14231 17119
rect 14933 17085 14967 17119
rect 16405 17085 16439 17119
rect 16732 17085 16766 17119
rect 17141 17085 17175 17119
rect 19165 17085 19199 17119
rect 19441 17085 19475 17119
rect 19717 17085 19751 17119
rect 19809 17085 19843 17119
rect 20361 17085 20395 17119
rect 20688 17085 20722 17119
rect 21097 17085 21131 17119
rect 23213 17085 23247 17119
rect 23857 17085 23891 17119
rect 25789 17085 25823 17119
rect 25881 17085 25915 17119
rect 26617 17085 26651 17119
rect 28365 17085 28399 17119
rect 28457 17085 28491 17119
rect 29101 17085 29135 17119
rect 29653 17085 29687 17119
rect 3525 17017 3559 17051
rect 8217 17017 8251 17051
rect 13737 17017 13771 17051
rect 20085 17017 20119 17051
rect 22661 17017 22695 17051
rect 30113 17017 30147 17051
rect 1415 16949 1449 16983
rect 4359 16949 4393 16983
rect 9143 16949 9177 16983
rect 11719 16949 11753 16983
rect 13093 16949 13127 16983
rect 14663 16949 14697 16983
rect 18245 16949 18279 16983
rect 22201 16949 22235 16983
rect 22937 16949 22971 16983
rect 26347 16949 26381 16983
rect 27721 16949 27755 16983
rect 28733 16949 28767 16983
rect 29929 16949 29963 16983
rect 1415 16745 1449 16779
rect 3157 16745 3191 16779
rect 5365 16745 5399 16779
rect 7665 16745 7699 16779
rect 8401 16745 8435 16779
rect 13461 16745 13495 16779
rect 15669 16745 15703 16779
rect 16405 16745 16439 16779
rect 16681 16745 16715 16779
rect 17423 16745 17457 16779
rect 19165 16745 19199 16779
rect 23121 16745 23155 16779
rect 23765 16745 23799 16779
rect 29193 16745 29227 16779
rect 30389 16745 30423 16779
rect 8125 16677 8159 16711
rect 19073 16677 19107 16711
rect 26525 16677 26559 16711
rect 949 16609 983 16643
rect 3341 16609 3375 16643
rect 4261 16609 4295 16643
rect 6561 16609 6595 16643
rect 8585 16609 8619 16643
rect 9321 16609 9355 16643
rect 11069 16609 11103 16643
rect 11621 16609 11655 16643
rect 14565 16609 14599 16643
rect 16313 16609 16347 16643
rect 16589 16609 16623 16643
rect 16865 16609 16899 16643
rect 17693 16609 17727 16643
rect 19349 16609 19383 16643
rect 19717 16609 19751 16643
rect 23673 16609 23707 16643
rect 23949 16609 23983 16643
rect 24133 16609 24167 16643
rect 24869 16609 24903 16643
rect 26985 16609 27019 16643
rect 27353 16609 27387 16643
rect 27680 16609 27714 16643
rect 28089 16609 28123 16643
rect 29837 16609 29871 16643
rect 29929 16609 29963 16643
rect 30573 16609 30607 16643
rect 1445 16559 1479 16593
rect 1685 16541 1719 16575
rect 3525 16541 3559 16575
rect 3852 16541 3886 16575
rect 3988 16543 4022 16577
rect 5825 16541 5859 16575
rect 6152 16541 6186 16575
rect 6288 16543 6322 16577
rect 8912 16541 8946 16575
rect 9081 16559 9115 16593
rect 11345 16541 11379 16575
rect 11948 16541 11982 16575
rect 12127 16541 12161 16575
rect 12357 16541 12391 16575
rect 13829 16541 13863 16575
rect 14156 16541 14190 16575
rect 14292 16543 14326 16577
rect 16957 16541 16991 16575
rect 17463 16543 17497 16577
rect 19441 16541 19475 16575
rect 21281 16541 21315 16575
rect 21608 16541 21642 16575
rect 21787 16543 21821 16577
rect 22017 16541 22051 16575
rect 24460 16541 24494 16575
rect 24596 16543 24630 16577
rect 27859 16543 27893 16577
rect 29653 16541 29687 16575
rect 25973 16473 26007 16507
rect 2789 16405 2823 16439
rect 10425 16405 10459 16439
rect 16129 16405 16163 16439
rect 21005 16405 21039 16439
rect 23489 16405 23523 16439
rect 26801 16405 26835 16439
rect 27169 16405 27203 16439
rect 30205 16405 30239 16439
rect 2789 16201 2823 16235
rect 5641 16201 5675 16235
rect 7941 16201 7975 16235
rect 23397 16201 23431 16235
rect 10977 16133 11011 16167
rect 25697 16133 25731 16167
rect 1445 16047 1479 16081
rect 4307 16065 4341 16099
rect 6607 16063 6641 16097
rect 9183 16065 9217 16099
rect 11253 16065 11287 16099
rect 11716 16063 11750 16097
rect 14703 16065 14737 16099
rect 16911 16065 16945 16099
rect 19625 16065 19659 16099
rect 19952 16065 19986 16099
rect 20121 16047 20155 16081
rect 22109 16065 22143 16099
rect 24320 16063 24354 16097
rect 26571 16065 26605 16099
rect 30113 16065 30147 16099
rect 949 15997 983 16031
rect 1685 15997 1719 16031
rect 3341 15997 3375 16031
rect 3801 15997 3835 16031
rect 4537 15997 4571 16031
rect 6101 15997 6135 16031
rect 6837 15997 6871 16031
rect 8585 15997 8619 16031
rect 8677 15997 8711 16031
rect 9413 15997 9447 16031
rect 11161 15997 11195 16031
rect 11989 15997 12023 16031
rect 13645 15997 13679 16031
rect 14197 15997 14231 16031
rect 14933 15997 14967 16031
rect 16405 15997 16439 16031
rect 17141 15997 17175 16031
rect 18797 15997 18831 16031
rect 19165 15997 19199 16031
rect 19441 15997 19475 16031
rect 20361 15997 20395 16031
rect 21833 15997 21867 16031
rect 23857 15997 23891 16031
rect 24593 15997 24627 16031
rect 26065 15997 26099 16031
rect 26392 15997 26426 16031
rect 26801 15997 26835 16031
rect 28365 15997 28399 16031
rect 29837 15997 29871 16031
rect 30297 15997 30331 16031
rect 29285 15929 29319 15963
rect 1415 15861 1449 15895
rect 3617 15861 3651 15895
rect 4267 15861 4301 15895
rect 6567 15861 6601 15895
rect 8401 15861 8435 15895
rect 9143 15861 9177 15895
rect 10517 15861 10551 15895
rect 11719 15861 11753 15895
rect 13093 15861 13127 15895
rect 13921 15861 13955 15895
rect 14663 15861 14697 15895
rect 16037 15861 16071 15895
rect 16871 15861 16905 15895
rect 18245 15861 18279 15895
rect 19257 15861 19291 15895
rect 21465 15861 21499 15895
rect 24323 15861 24357 15895
rect 27905 15861 27939 15895
rect 28641 15861 28675 15895
rect 29561 15861 29595 15895
rect 30481 15861 30515 15895
rect 1783 15657 1817 15691
rect 3157 15657 3191 15691
rect 15669 15657 15703 15691
rect 23121 15657 23155 15691
rect 25697 15657 25731 15691
rect 27721 15657 27755 15691
rect 30389 15657 30423 15691
rect 5641 15589 5675 15623
rect 11437 15589 11471 15623
rect 1133 15521 1167 15555
rect 3525 15521 3559 15555
rect 4261 15521 4295 15555
rect 5917 15521 5951 15555
rect 6796 15521 6830 15555
rect 9413 15521 9447 15555
rect 11069 15521 11103 15555
rect 11856 15521 11890 15555
rect 14565 15521 14599 15555
rect 16313 15521 16347 15555
rect 16589 15521 16623 15555
rect 16865 15521 16899 15555
rect 17376 15521 17410 15555
rect 21097 15521 21131 15555
rect 24225 15521 24259 15555
rect 25881 15521 25915 15555
rect 25973 15521 26007 15555
rect 26709 15521 26743 15555
rect 27169 15521 27203 15555
rect 27881 15521 27915 15555
rect 27997 15521 28031 15555
rect 28324 15521 28358 15555
rect 30297 15521 30331 15555
rect 1317 15453 1351 15487
rect 1813 15471 1847 15505
rect 2053 15453 2087 15487
rect 3852 15453 3886 15487
rect 4031 15453 4065 15487
rect 6469 15453 6503 15487
rect 6965 15471 6999 15505
rect 7205 15453 7239 15487
rect 8677 15453 8711 15487
rect 9004 15453 9038 15487
rect 9183 15455 9217 15489
rect 11529 15453 11563 15487
rect 12035 15453 12069 15487
rect 12265 15453 12299 15487
rect 13829 15453 13863 15487
rect 14156 15453 14190 15487
rect 14335 15453 14369 15487
rect 17049 15453 17083 15487
rect 17555 15453 17589 15487
rect 17785 15453 17819 15487
rect 19441 15453 19475 15487
rect 19717 15453 19751 15487
rect 21281 15453 21315 15487
rect 21608 15453 21642 15487
rect 21777 15471 21811 15505
rect 22017 15453 22051 15487
rect 23489 15453 23523 15487
rect 23816 15453 23850 15487
rect 23995 15453 24029 15487
rect 27353 15453 27387 15487
rect 28503 15453 28537 15487
rect 28733 15453 28767 15487
rect 6193 15385 6227 15419
rect 16129 15385 16163 15419
rect 26157 15385 26191 15419
rect 949 15317 983 15351
rect 8309 15317 8343 15351
rect 10517 15317 10551 15351
rect 13369 15317 13403 15351
rect 16405 15317 16439 15351
rect 16681 15317 16715 15351
rect 18889 15317 18923 15351
rect 25329 15317 25363 15351
rect 26985 15317 27019 15351
rect 29837 15317 29871 15351
rect 2973 15113 3007 15147
rect 10517 15113 10551 15147
rect 10977 15113 11011 15147
rect 19349 15113 19383 15147
rect 25697 15113 25731 15147
rect 26065 15113 26099 15147
rect 28733 15113 28767 15147
rect 30205 15113 30239 15147
rect 13093 15045 13127 15079
rect 13921 15045 13955 15079
rect 14197 15045 14231 15079
rect 29285 15045 29319 15079
rect 29929 15045 29963 15079
rect 949 14977 983 15011
rect 1455 14977 1489 15011
rect 3893 14977 3927 15011
rect 4399 14977 4433 15011
rect 6607 14977 6641 15011
rect 9004 14977 9038 15011
rect 9183 14977 9217 15011
rect 11759 14977 11793 15011
rect 15071 14977 15105 15011
rect 17141 14977 17175 15011
rect 18521 14977 18555 15011
rect 20121 14959 20155 14993
rect 22293 14977 22327 15011
rect 24184 14977 24218 15011
rect 24363 14977 24397 15011
rect 27172 14975 27206 15009
rect 1685 14909 1719 14943
rect 3249 14909 3283 14943
rect 4629 14909 4663 14943
rect 6101 14909 6135 14943
rect 6837 14909 6871 14943
rect 8585 14909 8619 14943
rect 8677 14909 8711 14943
rect 9413 14909 9447 14943
rect 11161 14909 11195 14943
rect 11253 14909 11287 14943
rect 11989 14909 12023 14943
rect 14105 14909 14139 14943
rect 14381 14909 14415 14943
rect 14565 14909 14599 14943
rect 15301 14909 15335 14943
rect 16865 14909 16899 14943
rect 18705 14909 18739 14943
rect 19533 14909 19567 14943
rect 19625 14909 19659 14943
rect 20361 14909 20395 14943
rect 22017 14909 22051 14943
rect 23857 14909 23891 14943
rect 24593 14909 24627 14943
rect 26249 14909 26283 14943
rect 26341 14909 26375 14943
rect 26709 14909 26743 14943
rect 27445 14909 27479 14943
rect 29653 14909 29687 14943
rect 30389 14909 30423 14943
rect 3525 14841 3559 14875
rect 6009 14841 6043 14875
rect 13645 14841 13679 14875
rect 13829 14841 13863 14875
rect 18981 14841 19015 14875
rect 29101 14841 29135 14875
rect 1415 14773 1449 14807
rect 4359 14773 4393 14807
rect 6567 14773 6601 14807
rect 7941 14773 7975 14807
rect 8401 14773 8435 14807
rect 11719 14773 11753 14807
rect 15031 14773 15065 14807
rect 16405 14773 16439 14807
rect 20091 14773 20125 14807
rect 21465 14773 21499 14807
rect 23581 14773 23615 14807
rect 26525 14773 26559 14807
rect 27175 14773 27209 14807
rect 1225 14569 1259 14603
rect 4077 14569 4111 14603
rect 4353 14569 4387 14603
rect 4905 14569 4939 14603
rect 5181 14569 5215 14603
rect 5457 14569 5491 14603
rect 6285 14569 6319 14603
rect 9965 14569 9999 14603
rect 10609 14569 10643 14603
rect 11161 14569 11195 14603
rect 16497 14569 16531 14603
rect 16681 14569 16715 14603
rect 17423 14569 17457 14603
rect 18797 14569 18831 14603
rect 21005 14569 21039 14603
rect 21747 14569 21781 14603
rect 25329 14569 25363 14603
rect 28273 14569 28307 14603
rect 30389 14569 30423 14603
rect 9321 14501 9355 14535
rect 15945 14501 15979 14535
rect 1133 14433 1167 14467
rect 1409 14433 1443 14467
rect 1828 14433 1862 14467
rect 3893 14433 3927 14467
rect 4261 14433 4295 14467
rect 4537 14433 4571 14467
rect 4813 14433 4847 14467
rect 5089 14433 5123 14467
rect 5365 14437 5399 14471
rect 5641 14433 5675 14467
rect 6009 14433 6043 14467
rect 6469 14433 6503 14467
rect 6745 14433 6779 14467
rect 9045 14433 9079 14467
rect 9781 14433 9815 14467
rect 10517 14433 10551 14467
rect 10793 14433 10827 14467
rect 11069 14433 11103 14467
rect 12357 14433 12391 14467
rect 14565 14433 14599 14467
rect 16221 14433 16255 14467
rect 16865 14433 16899 14467
rect 19349 14433 19383 14467
rect 19441 14433 19475 14467
rect 19717 14433 19751 14467
rect 21281 14433 21315 14467
rect 23816 14433 23850 14467
rect 24225 14433 24259 14467
rect 25789 14433 25823 14467
rect 26433 14433 26467 14467
rect 26760 14433 26794 14467
rect 28917 14433 28951 14467
rect 30573 14433 30607 14467
rect 1501 14365 1535 14399
rect 2007 14367 2041 14401
rect 2237 14365 2271 14399
rect 6837 14365 6871 14399
rect 7164 14365 7198 14399
rect 7300 14365 7334 14399
rect 7573 14365 7607 14399
rect 10057 14365 10091 14399
rect 11621 14365 11655 14399
rect 11948 14365 11982 14399
rect 12127 14365 12161 14399
rect 13829 14365 13863 14399
rect 14156 14365 14190 14399
rect 14335 14367 14369 14401
rect 16957 14365 16991 14399
rect 17463 14367 17497 14401
rect 17693 14365 17727 14399
rect 21777 14383 21811 14417
rect 22017 14365 22051 14399
rect 23489 14365 23523 14399
rect 23995 14365 24029 14399
rect 26065 14365 26099 14399
rect 26939 14365 26973 14399
rect 27169 14365 27203 14399
rect 28641 14365 28675 14399
rect 8861 14297 8895 14331
rect 10333 14297 10367 14331
rect 19165 14297 19199 14331
rect 949 14229 983 14263
rect 3525 14229 3559 14263
rect 3709 14229 3743 14263
rect 4629 14229 4663 14263
rect 5825 14229 5859 14263
rect 6561 14229 6595 14263
rect 13461 14229 13495 14263
rect 23121 14229 23155 14263
rect 30021 14229 30055 14263
rect 2789 14025 2823 14059
rect 7941 14025 7975 14059
rect 8493 14025 8527 14059
rect 9229 14025 9263 14059
rect 9413 14025 9447 14059
rect 12449 14025 12483 14059
rect 13001 14025 13035 14059
rect 13921 14025 13955 14059
rect 18981 14025 19015 14059
rect 19625 14025 19659 14059
rect 22753 14025 22787 14059
rect 23029 14025 23063 14059
rect 24225 14025 24259 14059
rect 26525 14025 26559 14059
rect 29009 14025 29043 14059
rect 29285 14025 29319 14059
rect 29561 14025 29595 14059
rect 3341 13957 3375 13991
rect 5917 13957 5951 13991
rect 8769 13957 8803 13991
rect 12725 13957 12759 13991
rect 13645 13957 13679 13991
rect 19257 13957 19291 13991
rect 22201 13957 22235 13991
rect 23949 13957 23983 13991
rect 28549 13957 28583 13991
rect 1445 13871 1479 13905
rect 4389 13871 4423 13905
rect 4629 13889 4663 13923
rect 6428 13889 6462 13923
rect 6607 13889 6641 13923
rect 10152 13889 10186 13923
rect 14703 13889 14737 13923
rect 16911 13889 16945 13923
rect 17141 13889 17175 13923
rect 20364 13889 20398 13923
rect 24828 13889 24862 13923
rect 25007 13889 25041 13923
rect 27172 13889 27206 13923
rect 949 13821 983 13855
rect 1685 13821 1719 13855
rect 3525 13821 3559 13855
rect 3801 13821 3835 13855
rect 3893 13821 3927 13855
rect 6101 13821 6135 13855
rect 6837 13821 6871 13855
rect 8677 13821 8711 13855
rect 8953 13821 8987 13855
rect 9045 13821 9079 13855
rect 9597 13821 9631 13855
rect 9689 13821 9723 13855
rect 10425 13821 10459 13855
rect 11805 13821 11839 13855
rect 11897 13821 11931 13855
rect 12173 13821 12207 13855
rect 12633 13821 12667 13855
rect 12909 13821 12943 13855
rect 13185 13821 13219 13855
rect 13829 13821 13863 13855
rect 14105 13821 14139 13855
rect 14197 13821 14231 13855
rect 14933 13821 14967 13855
rect 16313 13821 16347 13855
rect 16405 13821 16439 13855
rect 18889 13821 18923 13855
rect 19165 13821 19199 13855
rect 19441 13821 19475 13855
rect 19809 13821 19843 13855
rect 19901 13821 19935 13855
rect 20637 13821 20671 13855
rect 22017 13821 22051 13855
rect 22385 13821 22419 13855
rect 22937 13821 22971 13855
rect 23213 13821 23247 13855
rect 23673 13821 23707 13855
rect 24133 13821 24167 13855
rect 24409 13821 24443 13855
rect 24501 13821 24535 13855
rect 25237 13821 25271 13855
rect 26709 13821 26743 13855
rect 27445 13821 27479 13855
rect 29193 13821 29227 13855
rect 29469 13821 29503 13855
rect 29745 13821 29779 13855
rect 1415 13685 1449 13719
rect 3617 13685 3651 13719
rect 4359 13685 4393 13719
rect 10155 13685 10189 13719
rect 14663 13685 14697 13719
rect 16871 13685 16905 13719
rect 18245 13685 18279 13719
rect 18705 13685 18739 13719
rect 20367 13685 20401 13719
rect 23489 13685 23523 13719
rect 27175 13685 27209 13719
rect 1783 13481 1817 13515
rect 3991 13481 4025 13515
rect 6561 13481 6595 13515
rect 9781 13481 9815 13515
rect 11437 13481 11471 13515
rect 12915 13481 12949 13515
rect 16313 13481 16347 13515
rect 16681 13481 16715 13515
rect 17515 13481 17549 13515
rect 18889 13481 18923 13515
rect 21649 13481 21683 13515
rect 22391 13481 22425 13515
rect 24599 13481 24633 13515
rect 26899 13481 26933 13515
rect 28273 13481 28307 13515
rect 5641 13413 5675 13447
rect 9321 13413 9355 13447
rect 24041 13413 24075 13447
rect 1225 13345 1259 13379
rect 3433 13345 3467 13379
rect 3525 13345 3559 13379
rect 6193 13345 6227 13379
rect 6469 13345 6503 13379
rect 6837 13345 6871 13379
rect 9229 13345 9263 13379
rect 9597 13345 9631 13379
rect 9873 13345 9907 13379
rect 10149 13345 10183 13379
rect 10425 13345 10459 13379
rect 10977 13345 11011 13379
rect 11253 13345 11287 13379
rect 11713 13345 11747 13379
rect 11989 13345 12023 13379
rect 12265 13345 12299 13379
rect 14841 13345 14875 13379
rect 15393 13345 15427 13379
rect 15945 13345 15979 13379
rect 16129 13345 16163 13379
rect 16497 13345 16531 13379
rect 17049 13345 17083 13379
rect 17785 13345 17819 13379
rect 19809 13345 19843 13379
rect 20361 13345 20395 13379
rect 20637 13345 20671 13379
rect 21833 13345 21867 13379
rect 22661 13345 22695 13379
rect 24869 13345 24903 13379
rect 26433 13345 26467 13379
rect 27169 13345 27203 13379
rect 28917 13345 28951 13379
rect 1317 13277 1351 13311
rect 1823 13279 1857 13313
rect 2053 13277 2087 13311
rect 3988 13277 4022 13311
rect 4261 13277 4295 13311
rect 7164 13277 7198 13311
rect 7300 13277 7334 13311
rect 7573 13277 7607 13311
rect 12449 13277 12483 13311
rect 12912 13277 12946 13311
rect 13185 13277 13219 13311
rect 15025 13277 15059 13311
rect 17545 13295 17579 13329
rect 21925 13277 21959 13311
rect 22388 13277 22422 13311
rect 24133 13277 24167 13311
rect 24596 13279 24630 13313
rect 26896 13277 26930 13311
rect 28641 13277 28675 13311
rect 6009 13209 6043 13243
rect 9045 13209 9079 13243
rect 10609 13209 10643 13243
rect 11529 13209 11563 13243
rect 12081 13209 12115 13243
rect 15577 13209 15611 13243
rect 19533 13209 19567 13243
rect 20177 13209 20211 13243
rect 26157 13209 26191 13243
rect 1041 13141 1075 13175
rect 6285 13141 6319 13175
rect 8861 13141 8895 13175
rect 10057 13141 10091 13175
rect 10333 13141 10367 13175
rect 11161 13141 11195 13175
rect 11805 13141 11839 13175
rect 14289 13141 14323 13175
rect 15761 13141 15795 13175
rect 20453 13141 20487 13175
rect 30021 13141 30055 13175
rect 5917 12937 5951 12971
rect 12173 12937 12207 12971
rect 16773 12937 16807 12971
rect 20085 12937 20119 12971
rect 25697 12937 25731 12971
rect 28733 12937 28767 12971
rect 29193 12937 29227 12971
rect 29837 12937 29871 12971
rect 9045 12869 9079 12903
rect 11897 12869 11931 12903
rect 12909 12869 12943 12903
rect 22845 12869 22879 12903
rect 23213 12869 23247 12903
rect 949 12801 983 12835
rect 1455 12801 1489 12835
rect 3065 12801 3099 12835
rect 3883 12801 3917 12835
rect 4356 12801 4390 12835
rect 6564 12801 6598 12835
rect 6837 12801 6871 12835
rect 10152 12801 10186 12835
rect 10425 12801 10459 12835
rect 13737 12801 13771 12835
rect 14565 12801 14599 12835
rect 14892 12801 14926 12835
rect 15071 12801 15105 12835
rect 15301 12801 15335 12835
rect 20824 12801 20858 12835
rect 23857 12801 23891 12835
rect 24320 12783 24354 12817
rect 24593 12801 24627 12835
rect 26709 12801 26743 12835
rect 27205 12783 27239 12817
rect 1685 12733 1719 12767
rect 3525 12733 3559 12767
rect 3801 12733 3835 12767
rect 4629 12733 4663 12767
rect 6101 12733 6135 12767
rect 6428 12733 6462 12767
rect 9229 12733 9263 12767
rect 9321 12733 9355 12767
rect 9689 12733 9723 12767
rect 12081 12733 12115 12767
rect 12365 12733 12399 12767
rect 12817 12733 12851 12767
rect 13093 12733 13127 12767
rect 13369 12733 13403 12767
rect 13553 12733 13587 12767
rect 16957 12733 16991 12767
rect 18889 12733 18923 12767
rect 19165 12733 19199 12767
rect 19993 12733 20027 12767
rect 20269 12733 20303 12767
rect 20361 12733 20395 12767
rect 20688 12733 20722 12767
rect 21097 12733 21131 12767
rect 23029 12733 23063 12767
rect 23397 12733 23431 12767
rect 23673 12733 23707 12767
rect 26157 12733 26191 12767
rect 27445 12733 27479 12767
rect 29745 12733 29779 12767
rect 30013 12733 30047 12767
rect 8217 12665 8251 12699
rect 8493 12665 8527 12699
rect 14197 12665 14231 12699
rect 17969 12665 18003 12699
rect 18337 12665 18371 12699
rect 22477 12665 22511 12699
rect 29101 12665 29135 12699
rect 1415 12597 1449 12631
rect 3617 12597 3651 12631
rect 4359 12597 4393 12631
rect 8585 12597 8619 12631
rect 10155 12597 10189 12631
rect 11713 12597 11747 12631
rect 12633 12597 12667 12631
rect 13185 12597 13219 12631
rect 14289 12597 14323 12631
rect 16405 12597 16439 12631
rect 17233 12597 17267 12631
rect 17601 12597 17635 12631
rect 18705 12597 18739 12631
rect 18981 12597 19015 12631
rect 19809 12597 19843 12631
rect 23489 12597 23523 12631
rect 24323 12597 24357 12631
rect 26433 12597 26467 12631
rect 27175 12597 27209 12631
rect 29561 12597 29595 12631
rect 3991 12393 4025 12427
rect 5549 12393 5583 12427
rect 10701 12393 10735 12427
rect 12265 12393 12299 12427
rect 13007 12393 13041 12427
rect 15301 12393 15335 12427
rect 15761 12393 15795 12427
rect 16405 12393 16439 12427
rect 16957 12393 16991 12427
rect 18527 12393 18561 12427
rect 20085 12393 20119 12427
rect 20821 12393 20855 12427
rect 21747 12393 21781 12427
rect 23305 12393 23339 12427
rect 23955 12393 23989 12427
rect 25513 12393 25547 12427
rect 26899 12393 26933 12427
rect 28273 12393 28307 12427
rect 30389 12393 30423 12427
rect 17785 12325 17819 12359
rect 1225 12257 1259 12291
rect 3433 12257 3467 12291
rect 4261 12257 4295 12291
rect 6009 12257 6043 12291
rect 6285 12257 6319 12291
rect 6469 12257 6503 12291
rect 7205 12257 7239 12291
rect 8585 12257 8619 12291
rect 11161 12257 11195 12291
rect 11437 12257 11471 12291
rect 11713 12257 11747 12291
rect 11989 12257 12023 12291
rect 12449 12257 12483 12291
rect 12541 12257 12575 12291
rect 13277 12257 13311 12291
rect 14933 12257 14967 12291
rect 15209 12257 15243 12291
rect 15485 12257 15519 12291
rect 15945 12257 15979 12291
rect 16313 12257 16347 12291
rect 16589 12257 16623 12291
rect 17233 12257 17267 12291
rect 17509 12257 17543 12291
rect 18797 12257 18831 12291
rect 21005 12257 21039 12291
rect 22017 12257 22051 12291
rect 23489 12257 23523 12291
rect 24225 12257 24259 12291
rect 25697 12257 25731 12291
rect 26433 12257 26467 12291
rect 28641 12257 28675 12291
rect 30573 12257 30607 12291
rect 1317 12189 1351 12223
rect 1644 12189 1678 12223
rect 1823 12189 1857 12223
rect 2053 12189 2087 12223
rect 3525 12189 3559 12223
rect 4004 12191 4038 12225
rect 6796 12189 6830 12223
rect 6932 12189 6966 12223
rect 8677 12189 8711 12223
rect 9004 12189 9038 12223
rect 9140 12191 9174 12225
rect 9413 12189 9447 12223
rect 13004 12189 13038 12223
rect 18061 12189 18095 12223
rect 18524 12189 18558 12223
rect 21281 12189 21315 12223
rect 21744 12189 21778 12223
rect 23952 12189 23986 12223
rect 25881 12189 25915 12223
rect 26896 12189 26930 12223
rect 27169 12189 27203 12223
rect 28917 12189 28951 12223
rect 5825 12121 5859 12155
rect 10977 12121 11011 12155
rect 11805 12121 11839 12155
rect 16129 12121 16163 12155
rect 1041 12053 1075 12087
rect 6101 12053 6135 12087
rect 11253 12053 11287 12087
rect 11529 12053 11563 12087
rect 14381 12053 14415 12087
rect 14749 12053 14783 12087
rect 15025 12053 15059 12087
rect 17049 12053 17083 12087
rect 30021 12053 30055 12087
rect 5365 11849 5399 11883
rect 8033 11849 8067 11883
rect 15945 11849 15979 11883
rect 18429 11849 18463 11883
rect 20729 11849 20763 11883
rect 23581 11849 23615 11883
rect 26709 11849 26743 11883
rect 28641 11849 28675 11883
rect 23857 11781 23891 11815
rect 1455 11713 1489 11747
rect 1685 11713 1719 11747
rect 3847 11713 3881 11747
rect 4077 11713 4111 11747
rect 6012 11713 6046 11747
rect 9508 11713 9542 11747
rect 9781 11713 9815 11747
rect 11161 11713 11195 11747
rect 11716 11695 11750 11729
rect 11989 11713 12023 11747
rect 14059 11711 14093 11745
rect 14289 11713 14323 11747
rect 16911 11711 16945 11745
rect 17141 11713 17175 11747
rect 19168 11713 19202 11747
rect 19441 11713 19475 11747
rect 21557 11713 21591 11747
rect 22063 11713 22097 11747
rect 25191 11713 25225 11747
rect 26893 11713 26927 11747
rect 27169 11713 27203 11747
rect 29745 11713 29779 11747
rect 949 11645 983 11679
rect 3341 11645 3375 11679
rect 5549 11645 5583 11679
rect 6285 11645 6319 11679
rect 7941 11645 7975 11679
rect 8217 11645 8251 11679
rect 8585 11645 8619 11679
rect 8677 11645 8711 11679
rect 9045 11645 9079 11679
rect 11253 11645 11287 11679
rect 13553 11645 13587 11679
rect 13880 11645 13914 11679
rect 16313 11645 16347 11679
rect 16405 11645 16439 11679
rect 18705 11645 18739 11679
rect 22293 11645 22327 11679
rect 24041 11645 24075 11679
rect 24225 11645 24259 11679
rect 24685 11645 24719 11679
rect 25421 11645 25455 11679
rect 28825 11645 28859 11679
rect 29469 11645 29503 11679
rect 29561 11645 29595 11679
rect 3065 11577 3099 11611
rect 13369 11577 13403 11611
rect 24593 11577 24627 11611
rect 29101 11577 29135 11611
rect 1415 11509 1449 11543
rect 3807 11509 3841 11543
rect 6015 11509 6049 11543
rect 7389 11509 7423 11543
rect 7757 11509 7791 11543
rect 8401 11509 8435 11543
rect 8861 11509 8895 11543
rect 9511 11509 9545 11543
rect 11719 11509 11753 11543
rect 15393 11509 15427 11543
rect 16129 11509 16163 11543
rect 16871 11509 16905 11543
rect 19171 11509 19205 11543
rect 22023 11509 22057 11543
rect 25151 11509 25185 11543
rect 28273 11509 28307 11543
rect 3525 11305 3559 11339
rect 4813 11305 4847 11339
rect 9689 11305 9723 11339
rect 11805 11305 11839 11339
rect 12081 11305 12115 11339
rect 12915 11305 12949 11339
rect 16681 11305 16715 11339
rect 17331 11305 17365 11339
rect 18889 11305 18923 11339
rect 21649 11305 21683 11339
rect 24599 11305 24633 11339
rect 25973 11305 26007 11339
rect 26899 11305 26933 11339
rect 30389 11305 30423 11339
rect 4721 11237 4755 11271
rect 5457 11237 5491 11271
rect 5917 11237 5951 11271
rect 19349 11237 19383 11271
rect 1225 11169 1259 11203
rect 2237 11169 2271 11203
rect 3709 11169 3743 11203
rect 4537 11169 4571 11203
rect 5181 11169 5215 11203
rect 6561 11169 6595 11203
rect 6745 11169 6779 11203
rect 7481 11169 7515 11203
rect 8953 11169 8987 11203
rect 9597 11169 9631 11203
rect 10425 11169 10459 11203
rect 10701 11169 10735 11203
rect 11161 11169 11195 11203
rect 11253 11169 11287 11203
rect 11529 11169 11563 11203
rect 11989 11169 12023 11203
rect 12265 11169 12299 11203
rect 13185 11169 13219 11203
rect 14841 11169 14875 11203
rect 15117 11169 15151 11203
rect 15485 11169 15519 11203
rect 15761 11169 15795 11203
rect 17601 11169 17635 11203
rect 19073 11169 19107 11203
rect 19809 11169 19843 11203
rect 21465 11169 21499 11203
rect 21833 11169 21867 11203
rect 22252 11169 22286 11203
rect 24041 11169 24075 11203
rect 27169 11169 27203 11203
rect 28917 11169 28951 11203
rect 30573 11169 30607 11203
rect 1501 11101 1535 11135
rect 1828 11101 1862 11135
rect 2007 11101 2041 11135
rect 3985 11101 4019 11135
rect 7072 11101 7106 11135
rect 7208 11103 7242 11137
rect 8861 11101 8895 11135
rect 12449 11101 12483 11135
rect 12912 11101 12946 11135
rect 16865 11101 16899 11135
rect 17371 11101 17405 11135
rect 21925 11101 21959 11135
rect 22431 11101 22465 11135
rect 22661 11101 22695 11135
rect 24133 11101 24167 11135
rect 24596 11103 24630 11137
rect 24869 11101 24903 11135
rect 26433 11101 26467 11135
rect 26896 11101 26930 11135
rect 28641 11101 28675 11135
rect 6101 11033 6135 11067
rect 6377 11033 6411 11067
rect 10241 11033 10275 11067
rect 10517 11033 10551 11067
rect 10977 11033 11011 11067
rect 14289 11033 14323 11067
rect 14933 11033 14967 11067
rect 28273 11033 28307 11067
rect 30021 11033 30055 11067
rect 4353 10965 4387 10999
rect 9137 10965 9171 10999
rect 11437 10965 11471 10999
rect 11713 10965 11747 10999
rect 14657 10965 14691 10999
rect 16313 10965 16347 10999
rect 19625 10965 19659 10999
rect 21281 10965 21315 10999
rect 11713 10761 11747 10795
rect 16313 10761 16347 10795
rect 20729 10761 20763 10795
rect 23121 10761 23155 10795
rect 23857 10761 23891 10795
rect 8033 10693 8067 10727
rect 12265 10693 12299 10727
rect 12449 10693 12483 10727
rect 18429 10693 18463 10727
rect 22753 10693 22787 10727
rect 30297 10693 30331 10727
rect 949 10625 983 10659
rect 1455 10625 1489 10659
rect 3755 10623 3789 10657
rect 5549 10625 5583 10659
rect 6012 10625 6046 10659
rect 7665 10625 7699 10659
rect 10152 10625 10186 10659
rect 10425 10625 10459 10659
rect 14016 10625 14050 10659
rect 14289 10625 14323 10659
rect 16868 10625 16902 10659
rect 18705 10625 18739 10659
rect 19184 10607 19218 10641
rect 20913 10625 20947 10659
rect 21409 10607 21443 10641
rect 25099 10625 25133 10659
rect 27077 10625 27111 10659
rect 1685 10557 1719 10591
rect 3249 10557 3283 10591
rect 3985 10557 4019 10591
rect 6285 10557 6319 10591
rect 8401 10557 8435 10591
rect 8953 10557 8987 10591
rect 9689 10557 9723 10591
rect 10016 10557 10050 10591
rect 12633 10557 12667 10591
rect 12725 10557 12759 10591
rect 13369 10557 13403 10591
rect 13553 10557 13587 10591
rect 16405 10557 16439 10591
rect 17141 10557 17175 10591
rect 19441 10557 19475 10591
rect 21649 10557 21683 10591
rect 23305 10557 23339 10591
rect 24041 10557 24075 10591
rect 24593 10557 24627 10591
rect 25329 10557 25363 10591
rect 26801 10557 26835 10591
rect 29101 10557 29135 10591
rect 30113 10557 30147 10591
rect 5365 10489 5399 10523
rect 7849 10489 7883 10523
rect 9229 10489 9263 10523
rect 11989 10489 12023 10523
rect 26709 10489 26743 10523
rect 29653 10489 29687 10523
rect 1415 10421 1449 10455
rect 2973 10421 3007 10455
rect 3715 10421 3749 10455
rect 6015 10421 6049 10455
rect 8585 10421 8619 10455
rect 12909 10421 12943 10455
rect 13185 10421 13219 10455
rect 14019 10421 14053 10455
rect 15393 10421 15427 10455
rect 16871 10421 16905 10455
rect 19171 10421 19205 10455
rect 21379 10421 21413 10455
rect 25059 10421 25093 10455
rect 28181 10421 28215 10455
rect 29193 10421 29227 10455
rect 29745 10421 29779 10455
rect 1507 10217 1541 10251
rect 3715 10217 3749 10251
rect 6935 10217 6969 10251
rect 17699 10217 17733 10251
rect 19257 10217 19291 10251
rect 21747 10217 21781 10251
rect 23121 10217 23155 10251
rect 26899 10217 26933 10251
rect 13277 10149 13311 10183
rect 20729 10149 20763 10183
rect 1041 10081 1075 10115
rect 5641 10081 5675 10115
rect 5917 10081 5951 10115
rect 6469 10081 6503 10115
rect 8585 10081 8619 10115
rect 9413 10081 9447 10115
rect 13553 10081 13587 10115
rect 15945 10081 15979 10115
rect 16313 10081 16347 10115
rect 16865 10081 16899 10115
rect 17141 10081 17175 10115
rect 20177 10081 20211 10115
rect 22017 10081 22051 10115
rect 24041 10081 24075 10115
rect 24460 10081 24494 10115
rect 26249 10081 26283 10115
rect 28641 10081 28675 10115
rect 30573 10081 30607 10115
rect 1537 10031 1571 10065
rect 1777 10013 1811 10047
rect 3249 10013 3283 10047
rect 3712 10013 3746 10047
rect 3985 10013 4019 10047
rect 5365 10013 5399 10047
rect 6101 10013 6135 10047
rect 6975 10013 7009 10047
rect 7205 10013 7239 10047
rect 8677 10013 8711 10047
rect 9004 10013 9038 10047
rect 9140 10015 9174 10049
rect 10977 10013 11011 10047
rect 11304 10013 11338 10047
rect 11440 10013 11474 10047
rect 11713 10013 11747 10047
rect 13880 10013 13914 10047
rect 14059 10013 14093 10047
rect 14289 10013 14323 10047
rect 17233 10013 17267 10047
rect 17739 10013 17773 10047
rect 17969 10013 18003 10047
rect 21281 10013 21315 10047
rect 21744 10013 21778 10047
rect 24133 10013 24167 10047
rect 24596 10013 24630 10047
rect 24869 10013 24903 10047
rect 26433 10013 26467 10047
rect 26896 10013 26930 10047
rect 27169 10013 27203 10047
rect 28917 10013 28951 10047
rect 15761 9945 15795 9979
rect 16681 9945 16715 9979
rect 19993 9945 20027 9979
rect 3065 9877 3099 9911
rect 5457 9877 5491 9911
rect 10701 9877 10735 9911
rect 12817 9877 12851 9911
rect 13369 9877 13403 9911
rect 15393 9877 15427 9911
rect 16129 9877 16163 9911
rect 16957 9877 16991 9911
rect 21005 9877 21039 9911
rect 23857 9877 23891 9911
rect 28457 9877 28491 9911
rect 30021 9877 30055 9911
rect 30389 9877 30423 9911
rect 18245 9673 18279 9707
rect 25697 9673 25731 9707
rect 28273 9673 28307 9707
rect 5365 9605 5399 9639
rect 10609 9605 10643 9639
rect 13185 9605 13219 9639
rect 22753 9605 22787 9639
rect 949 9537 983 9571
rect 1445 9519 1479 9553
rect 3804 9537 3838 9571
rect 6101 9537 6135 9571
rect 6564 9537 6598 9571
rect 8585 9537 8619 9571
rect 9091 9537 9125 9571
rect 10793 9537 10827 9571
rect 11120 9537 11154 9571
rect 11256 9537 11290 9571
rect 13553 9537 13587 9571
rect 14059 9537 14093 9571
rect 16911 9535 16945 9569
rect 19211 9535 19245 9569
rect 19441 9537 19475 9571
rect 20821 9537 20855 9571
rect 21409 9519 21443 9553
rect 24320 9537 24354 9571
rect 26065 9537 26099 9571
rect 26392 9537 26426 9571
rect 26528 9535 26562 9569
rect 1685 9469 1719 9503
rect 3341 9469 3375 9503
rect 4077 9469 4111 9503
rect 5733 9469 5767 9503
rect 6009 9469 6043 9503
rect 6837 9469 6871 9503
rect 9321 9469 9355 9503
rect 11529 9469 11563 9503
rect 13001 9469 13035 9503
rect 14289 9469 14323 9503
rect 16313 9469 16347 9503
rect 16405 9469 16439 9503
rect 16732 9469 16766 9503
rect 17141 9469 17175 9503
rect 18705 9469 18739 9503
rect 20913 9469 20947 9503
rect 21649 9469 21683 9503
rect 23581 9469 23615 9503
rect 23857 9469 23891 9503
rect 24593 9469 24627 9503
rect 26801 9469 26835 9503
rect 28457 9469 28491 9503
rect 28733 9469 28767 9503
rect 30481 9469 30515 9503
rect 16037 9401 16071 9435
rect 1415 9333 1449 9367
rect 2973 9333 3007 9367
rect 3807 9333 3841 9367
rect 5549 9333 5583 9367
rect 5825 9333 5859 9367
rect 6567 9333 6601 9367
rect 8125 9333 8159 9367
rect 9051 9333 9085 9367
rect 12633 9333 12667 9367
rect 14019 9333 14053 9367
rect 15393 9333 15427 9367
rect 16129 9333 16163 9367
rect 19171 9333 19205 9367
rect 21379 9333 21413 9367
rect 23397 9333 23431 9367
rect 24323 9333 24357 9367
rect 27905 9333 27939 9367
rect 28549 9333 28583 9367
rect 30297 9333 30331 9367
rect 3715 9129 3749 9163
rect 7297 9129 7331 9163
rect 9413 9129 9447 9163
rect 9781 9129 9815 9163
rect 10333 9129 10367 9163
rect 10609 9129 10643 9163
rect 15761 9129 15795 9163
rect 16589 9129 16623 9163
rect 21281 9129 21315 9163
rect 25697 9129 25731 9163
rect 25973 9129 26007 9163
rect 26899 9129 26933 9163
rect 30205 9129 30239 9163
rect 5365 9061 5399 9095
rect 13277 9061 13311 9095
rect 20545 9061 20579 9095
rect 25237 9061 25271 9095
rect 5641 8993 5675 9027
rect 6009 8993 6043 9027
rect 6377 8993 6411 9027
rect 6653 8993 6687 9027
rect 6745 8993 6779 9027
rect 7481 8993 7515 9027
rect 8309 8993 8343 9027
rect 9965 8993 9999 9027
rect 10241 8993 10275 9027
rect 10517 8993 10551 9027
rect 10793 8993 10827 9027
rect 11304 8993 11338 9027
rect 11713 8993 11747 9027
rect 13880 8993 13914 9027
rect 14289 8993 14323 9027
rect 15945 8993 15979 9027
rect 16313 8993 16347 9027
rect 16773 8993 16807 9027
rect 16865 8993 16899 9027
rect 19257 8993 19291 9027
rect 20269 8993 20303 9027
rect 21465 8993 21499 9027
rect 22201 8993 22235 9027
rect 22845 8993 22879 9027
rect 22937 8993 22971 9027
rect 23264 8993 23298 9027
rect 23673 8993 23707 9027
rect 25881 8993 25915 9027
rect 26157 8993 26191 9027
rect 26433 8993 26467 9027
rect 28641 8993 28675 9027
rect 28917 8993 28951 9027
rect 1041 8925 1075 8959
rect 1368 8925 1402 8959
rect 1537 8943 1571 8977
rect 1777 8925 1811 8959
rect 3157 8925 3191 8959
rect 3249 8925 3283 8959
rect 3712 8943 3746 8977
rect 3985 8925 4019 8959
rect 6929 8925 6963 8959
rect 7573 8925 7607 8959
rect 7900 8925 7934 8959
rect 8036 8925 8070 8959
rect 10977 8925 11011 8959
rect 11440 8927 11474 8961
rect 13553 8925 13587 8959
rect 14049 8943 14083 8977
rect 17192 8925 17226 8959
rect 17371 8925 17405 8959
rect 17601 8925 17635 8959
rect 23443 8925 23477 8959
rect 25513 8925 25547 8959
rect 26939 8925 26973 8959
rect 27169 8925 27203 8959
rect 5825 8857 5859 8891
rect 5457 8789 5491 8823
rect 6193 8789 6227 8823
rect 6469 8789 6503 8823
rect 10057 8789 10091 8823
rect 12817 8789 12851 8823
rect 13369 8789 13403 8823
rect 15393 8789 15427 8823
rect 16129 8789 16163 8823
rect 18705 8789 18739 8823
rect 19073 8789 19107 8823
rect 22017 8789 22051 8823
rect 22661 8789 22695 8823
rect 24961 8789 24995 8823
rect 28273 8789 28307 8823
rect 2789 8585 2823 8619
rect 7389 8585 7423 8619
rect 7757 8585 7791 8619
rect 11529 8585 11563 8619
rect 18245 8585 18279 8619
rect 20729 8585 20763 8619
rect 22753 8585 22787 8619
rect 26065 8585 26099 8619
rect 26341 8585 26375 8619
rect 28549 8585 28583 8619
rect 29193 8585 29227 8619
rect 30297 8585 30331 8619
rect 5181 8517 5215 8551
rect 9137 8517 9171 8551
rect 12817 8517 12851 8551
rect 25881 8517 25915 8551
rect 1455 8449 1489 8483
rect 3341 8449 3375 8483
rect 3847 8449 3881 8483
rect 4077 8449 4111 8483
rect 5549 8449 5583 8483
rect 6012 8449 6046 8483
rect 9968 8449 10002 8483
rect 10241 8449 10275 8483
rect 12081 8449 12115 8483
rect 13553 8449 13587 8483
rect 14059 8449 14093 8483
rect 14289 8449 14323 8483
rect 16732 8449 16766 8483
rect 16901 8431 16935 8465
rect 18705 8449 18739 8483
rect 19032 8449 19066 8483
rect 19211 8449 19245 8483
rect 21240 8449 21274 8483
rect 21419 8449 21453 8483
rect 24320 8449 24354 8483
rect 24593 8449 24627 8483
rect 26709 8449 26743 8483
rect 27036 8449 27070 8483
rect 27215 8449 27249 8483
rect 949 8381 983 8415
rect 1685 8381 1719 8415
rect 3668 8381 3702 8415
rect 6285 8381 6319 8415
rect 7941 8381 7975 8415
rect 8217 8381 8251 8415
rect 8861 8381 8895 8415
rect 9321 8381 9355 8415
rect 9505 8381 9539 8415
rect 9832 8381 9866 8415
rect 12541 8381 12575 8415
rect 12633 8381 12667 8415
rect 12909 8381 12943 8415
rect 13185 8381 13219 8415
rect 13880 8381 13914 8415
rect 15853 8381 15887 8415
rect 16405 8381 16439 8415
rect 17141 8381 17175 8415
rect 19441 8381 19475 8415
rect 20913 8381 20947 8415
rect 21649 8381 21683 8415
rect 23213 8381 23247 8415
rect 23857 8381 23891 8415
rect 24184 8381 24218 8415
rect 26249 8381 26283 8415
rect 26525 8381 26559 8415
rect 27445 8381 27479 8415
rect 29101 8381 29135 8415
rect 30205 8381 30239 8415
rect 8493 8313 8527 8347
rect 11805 8313 11839 8347
rect 12321 8313 12355 8347
rect 23581 8313 23615 8347
rect 29653 8313 29687 8347
rect 1415 8245 1449 8279
rect 6015 8245 6049 8279
rect 8033 8245 8067 8279
rect 15393 8245 15427 8279
rect 16129 8245 16163 8279
rect 29745 8245 29779 8279
rect 5457 8041 5491 8075
rect 5825 8041 5859 8075
rect 8033 8041 8067 8075
rect 13461 8041 13495 8075
rect 14295 8041 14329 8075
rect 18527 8041 18561 8075
rect 19901 8041 19935 8075
rect 20453 8041 20487 8075
rect 21281 8041 21315 8075
rect 23581 8041 23615 8075
rect 25973 8041 26007 8075
rect 29653 8041 29687 8075
rect 11069 7973 11103 8007
rect 16957 7973 16991 8007
rect 17509 7973 17543 8007
rect 3249 7905 3283 7939
rect 3985 7905 4019 7939
rect 5641 7905 5675 7939
rect 6009 7905 6043 7939
rect 8401 7905 8435 7939
rect 10793 7905 10827 7939
rect 11948 7905 11982 7939
rect 14565 7905 14599 7939
rect 16405 7905 16439 7939
rect 18061 7905 18095 7939
rect 20637 7905 20671 7939
rect 21097 7905 21131 7939
rect 21441 7905 21475 7939
rect 22293 7905 22327 7939
rect 26433 7905 26467 7939
rect 27721 7905 27755 7939
rect 28140 7905 28174 7939
rect 28549 7905 28583 7939
rect 30297 7905 30331 7939
rect 30573 7905 30607 7939
rect 1041 7837 1075 7871
rect 1368 7837 1402 7871
rect 1547 7837 1581 7871
rect 1777 7837 1811 7871
rect 3576 7837 3610 7871
rect 3728 7855 3762 7889
rect 6193 7837 6227 7871
rect 6520 7837 6554 7871
rect 6699 7839 6733 7873
rect 6929 7837 6963 7871
rect 8728 7837 8762 7871
rect 8907 7837 8941 7871
rect 9137 7837 9171 7871
rect 11345 7837 11379 7871
rect 11621 7837 11655 7871
rect 12127 7837 12161 7871
rect 12357 7837 12391 7871
rect 13829 7837 13863 7871
rect 14335 7837 14369 7871
rect 18567 7839 18601 7873
rect 18797 7837 18831 7871
rect 21557 7837 21591 7871
rect 21884 7837 21918 7871
rect 22063 7837 22097 7871
rect 24133 7837 24167 7871
rect 24460 7837 24494 7871
rect 24596 7839 24630 7873
rect 24869 7837 24903 7871
rect 26709 7837 26743 7871
rect 27813 7837 27847 7871
rect 28319 7837 28353 7871
rect 10609 7769 10643 7803
rect 17693 7769 17727 7803
rect 30389 7769 30423 7803
rect 2881 7701 2915 7735
rect 5089 7701 5123 7735
rect 10241 7701 10275 7735
rect 15669 7701 15703 7735
rect 16681 7701 16715 7735
rect 17049 7701 17083 7735
rect 20913 7701 20947 7735
rect 27537 7701 27571 7735
rect 30113 7701 30147 7735
rect 7941 7497 7975 7531
rect 13093 7497 13127 7531
rect 17877 7497 17911 7531
rect 20545 7497 20579 7531
rect 23581 7497 23615 7531
rect 28457 7497 28491 7531
rect 5365 7429 5399 7463
rect 10333 7429 10367 7463
rect 10977 7429 11011 7463
rect 14105 7429 14139 7463
rect 25881 7429 25915 7463
rect 28089 7429 28123 7463
rect 29285 7429 29319 7463
rect 1455 7361 1489 7395
rect 3525 7361 3559 7395
rect 4031 7361 4065 7395
rect 4261 7361 4295 7395
rect 6239 7359 6273 7393
rect 8493 7361 8527 7395
rect 8999 7361 9033 7395
rect 11759 7361 11793 7395
rect 14887 7361 14921 7395
rect 19211 7361 19245 7395
rect 22063 7359 22097 7393
rect 22293 7361 22327 7395
rect 24504 7361 24538 7395
rect 26712 7361 26746 7395
rect 949 7293 983 7327
rect 1685 7293 1719 7327
rect 3433 7293 3467 7327
rect 5733 7293 5767 7327
rect 6469 7293 6503 7327
rect 8125 7293 8159 7327
rect 8820 7293 8854 7327
rect 9229 7293 9263 7327
rect 10885 7293 10919 7327
rect 11161 7293 11195 7327
rect 11253 7293 11287 7327
rect 11989 7293 12023 7327
rect 13553 7293 13587 7327
rect 14289 7293 14323 7327
rect 14381 7293 14415 7327
rect 15117 7293 15151 7327
rect 16773 7293 16807 7327
rect 16865 7293 16899 7327
rect 17417 7293 17451 7327
rect 17601 7293 17635 7327
rect 18061 7293 18095 7327
rect 18337 7293 18371 7327
rect 18705 7293 18739 7327
rect 19441 7293 19475 7327
rect 21557 7293 21591 7327
rect 24041 7293 24075 7327
rect 24777 7293 24811 7327
rect 26249 7293 26283 7327
rect 26576 7293 26610 7327
rect 26985 7293 27019 7327
rect 28641 7293 28675 7327
rect 29193 7293 29227 7327
rect 29469 7293 29503 7327
rect 13829 7225 13863 7259
rect 21097 7225 21131 7259
rect 1415 7157 1449 7191
rect 2789 7157 2823 7191
rect 3249 7157 3283 7191
rect 3991 7157 4025 7191
rect 6199 7157 6233 7191
rect 7573 7157 7607 7191
rect 10701 7157 10735 7191
rect 11719 7157 11753 7191
rect 14847 7157 14881 7191
rect 16221 7157 16255 7191
rect 16589 7157 16623 7191
rect 17049 7157 17083 7191
rect 17233 7157 17267 7191
rect 19171 7157 19205 7191
rect 22023 7157 22057 7191
rect 24507 7157 24541 7191
rect 29009 7157 29043 7191
rect 13185 6953 13219 6987
rect 14295 6953 14329 6987
rect 16129 6953 16163 6987
rect 17509 6953 17543 6987
rect 18527 6953 18561 6987
rect 26433 6953 26467 6987
rect 28279 6953 28313 6987
rect 27353 6885 27387 6919
rect 5641 6817 5675 6851
rect 8217 6817 8251 6851
rect 10793 6817 10827 6851
rect 11253 6817 11287 6851
rect 11672 6817 11706 6851
rect 13553 6817 13587 6851
rect 15945 6817 15979 6851
rect 16313 6817 16347 6851
rect 16405 6817 16439 6851
rect 16681 6817 16715 6851
rect 16957 6817 16991 6851
rect 17417 6817 17451 6851
rect 17693 6817 17727 6851
rect 17785 6817 17819 6851
rect 18061 6817 18095 6851
rect 20453 6817 20487 6851
rect 20729 6817 20763 6851
rect 21005 6817 21039 6851
rect 21465 6817 21499 6851
rect 22477 6817 22511 6851
rect 23857 6817 23891 6851
rect 24368 6817 24402 6851
rect 26617 6817 26651 6851
rect 28549 6817 28583 6851
rect 1041 6749 1075 6783
rect 1368 6749 1402 6783
rect 1547 6749 1581 6783
rect 1777 6749 1811 6783
rect 3249 6749 3283 6783
rect 3576 6749 3610 6783
rect 3755 6749 3789 6783
rect 3985 6749 4019 6783
rect 5825 6749 5859 6783
rect 6152 6749 6186 6783
rect 6331 6749 6365 6783
rect 6561 6749 6595 6783
rect 8401 6749 8435 6783
rect 8728 6749 8762 6783
rect 8907 6751 8941 6785
rect 9137 6749 9171 6783
rect 11345 6749 11379 6783
rect 11851 6749 11885 6783
rect 12081 6749 12115 6783
rect 13829 6749 13863 6783
rect 14335 6749 14369 6783
rect 14565 6749 14599 6783
rect 18567 6751 18601 6785
rect 18797 6749 18831 6783
rect 21741 6749 21775 6783
rect 22068 6749 22102 6783
rect 22247 6749 22281 6783
rect 24049 6749 24083 6783
rect 24504 6749 24538 6783
rect 24777 6749 24811 6783
rect 27813 6749 27847 6783
rect 28276 6749 28310 6783
rect 19901 6681 19935 6715
rect 29653 6681 29687 6715
rect 2881 6613 2915 6647
rect 5089 6613 5123 6647
rect 5457 6613 5491 6647
rect 7665 6613 7699 6647
rect 8033 6613 8067 6647
rect 10241 6613 10275 6647
rect 10609 6613 10643 6647
rect 11069 6613 11103 6647
rect 13737 6613 13771 6647
rect 16589 6613 16623 6647
rect 16865 6613 16899 6647
rect 17141 6613 17175 6647
rect 17233 6613 17267 6647
rect 17969 6613 18003 6647
rect 20269 6613 20303 6647
rect 20545 6613 20579 6647
rect 20821 6613 20855 6647
rect 21281 6613 21315 6647
rect 26065 6613 26099 6647
rect 27445 6613 27479 6647
rect 10609 6409 10643 6443
rect 13093 6409 13127 6443
rect 13829 6409 13863 6443
rect 16221 6409 16255 6443
rect 18061 6409 18095 6443
rect 23489 6409 23523 6443
rect 28549 6409 28583 6443
rect 7389 6341 7423 6375
rect 8125 6341 8159 6375
rect 10885 6341 10919 6375
rect 17785 6341 17819 6375
rect 1455 6273 1489 6307
rect 3576 6273 3610 6307
rect 3755 6273 3789 6307
rect 5876 6273 5910 6307
rect 6055 6273 6089 6307
rect 6285 6273 6319 6307
rect 8864 6273 8898 6307
rect 11580 6273 11614 6307
rect 11759 6273 11793 6307
rect 14381 6273 14415 6307
rect 14708 6273 14742 6307
rect 14887 6273 14921 6307
rect 15117 6273 15151 6307
rect 19168 6273 19202 6307
rect 19441 6273 19475 6307
rect 20821 6273 20855 6307
rect 21376 6273 21410 6307
rect 21649 6273 21683 6307
rect 24547 6273 24581 6307
rect 27172 6273 27206 6307
rect 27445 6273 27479 6307
rect 949 6205 983 6239
rect 1685 6205 1719 6239
rect 3249 6205 3283 6239
rect 3985 6205 4019 6239
rect 5549 6205 5583 6239
rect 8401 6205 8435 6239
rect 9137 6205 9171 6239
rect 10793 6205 10827 6239
rect 11069 6205 11103 6239
rect 11253 6205 11287 6239
rect 11989 6205 12023 6239
rect 13737 6205 13771 6239
rect 14013 6205 14047 6239
rect 14289 6205 14323 6239
rect 16865 6205 16899 6239
rect 17141 6205 17175 6239
rect 17417 6205 17451 6239
rect 17509 6205 17543 6239
rect 17969 6205 18003 6239
rect 18245 6205 18279 6239
rect 18337 6205 18371 6239
rect 18705 6205 18739 6239
rect 20913 6205 20947 6239
rect 23305 6205 23339 6239
rect 23673 6205 23707 6239
rect 24041 6205 24075 6239
rect 24777 6205 24811 6239
rect 26617 6205 26651 6239
rect 26709 6205 26743 6239
rect 27036 6205 27070 6239
rect 29193 6205 29227 6239
rect 7849 6137 7883 6171
rect 23029 6137 23063 6171
rect 26157 6137 26191 6171
rect 1415 6069 1449 6103
rect 2789 6069 2823 6103
rect 5089 6069 5123 6103
rect 8867 6069 8901 6103
rect 10241 6069 10275 6103
rect 13553 6069 13587 6103
rect 14105 6069 14139 6103
rect 16681 6069 16715 6103
rect 16957 6069 16991 6103
rect 17233 6069 17267 6103
rect 17693 6069 17727 6103
rect 18521 6069 18555 6103
rect 19171 6069 19205 6103
rect 21379 6069 21413 6103
rect 23121 6069 23155 6103
rect 24507 6069 24541 6103
rect 26433 6069 26467 6103
rect 29009 6069 29043 6103
rect 1783 5865 1817 5899
rect 3991 5865 4025 5899
rect 8499 5865 8533 5899
rect 11069 5865 11103 5899
rect 21747 5865 21781 5899
rect 23955 5865 23989 5899
rect 25329 5865 25363 5899
rect 25973 5865 26007 5899
rect 26899 5865 26933 5899
rect 3433 5797 3467 5831
rect 1225 5729 1259 5763
rect 1317 5729 1351 5763
rect 4261 5729 4295 5763
rect 6561 5729 6595 5763
rect 10433 5729 10467 5763
rect 10793 5729 10827 5763
rect 11253 5729 11287 5763
rect 11529 5729 11563 5763
rect 12357 5729 12391 5763
rect 14565 5729 14599 5763
rect 15945 5729 15979 5763
rect 16957 5729 16991 5763
rect 18337 5729 18371 5763
rect 20821 5729 20855 5763
rect 21097 5729 21131 5763
rect 22017 5729 22051 5763
rect 23397 5729 23431 5763
rect 25881 5729 25915 5763
rect 26157 5729 26191 5763
rect 27169 5729 27203 5763
rect 28641 5729 28675 5763
rect 29009 5729 29043 5763
rect 29285 5729 29319 5763
rect 1813 5679 1847 5713
rect 2053 5661 2087 5695
rect 3525 5661 3559 5695
rect 4031 5661 4065 5695
rect 5825 5661 5859 5695
rect 6152 5661 6186 5695
rect 6288 5661 6322 5695
rect 8033 5661 8067 5695
rect 8496 5679 8530 5713
rect 8769 5661 8803 5695
rect 10149 5661 10183 5695
rect 11621 5661 11655 5695
rect 11948 5661 11982 5695
rect 12127 5661 12161 5695
rect 13829 5661 13863 5695
rect 14156 5661 14190 5695
rect 14292 5661 14326 5695
rect 16221 5661 16255 5695
rect 16548 5661 16582 5695
rect 16684 5663 16718 5697
rect 18429 5661 18463 5695
rect 18756 5661 18790 5695
rect 18892 5663 18926 5697
rect 19165 5661 19199 5695
rect 21281 5661 21315 5695
rect 21744 5661 21778 5695
rect 23489 5661 23523 5695
rect 23952 5661 23986 5695
rect 24225 5661 24259 5695
rect 26433 5661 26467 5695
rect 26896 5661 26930 5695
rect 20637 5593 20671 5627
rect 20913 5593 20947 5627
rect 25697 5593 25731 5627
rect 28825 5593 28859 5627
rect 1041 5525 1075 5559
rect 5549 5525 5583 5559
rect 7665 5525 7699 5559
rect 10241 5525 10275 5559
rect 10609 5525 10643 5559
rect 11345 5525 11379 5559
rect 13645 5525 13679 5559
rect 20453 5525 20487 5559
rect 28273 5525 28307 5559
rect 29193 5525 29227 5559
rect 29469 5525 29503 5559
rect 2973 5321 3007 5355
rect 5917 5321 5951 5355
rect 8401 5321 8435 5355
rect 13277 5321 13311 5355
rect 25881 5321 25915 5355
rect 28549 5321 28583 5355
rect 3617 5253 3651 5287
rect 8677 5253 8711 5287
rect 23397 5253 23431 5287
rect 949 5185 983 5219
rect 1455 5185 1489 5219
rect 3893 5185 3927 5219
rect 4399 5185 4433 5219
rect 6607 5185 6641 5219
rect 9551 5185 9585 5219
rect 9781 5185 9815 5219
rect 11716 5185 11750 5219
rect 14340 5185 14374 5219
rect 14476 5183 14510 5217
rect 14749 5185 14783 5219
rect 16129 5185 16163 5219
rect 16684 5185 16718 5219
rect 16957 5185 16991 5219
rect 18337 5185 18371 5219
rect 19168 5185 19202 5219
rect 19441 5185 19475 5219
rect 20821 5185 20855 5219
rect 21376 5185 21410 5219
rect 24320 5185 24354 5219
rect 27172 5185 27206 5219
rect 27445 5185 27479 5219
rect 1276 5117 1310 5151
rect 1685 5117 1719 5151
rect 4220 5117 4254 5151
rect 4629 5117 4663 5151
rect 6101 5117 6135 5151
rect 6837 5117 6871 5151
rect 8585 5117 8619 5151
rect 8861 5117 8895 5151
rect 9045 5117 9079 5151
rect 11253 5117 11287 5151
rect 11989 5117 12023 5151
rect 13921 5117 13955 5151
rect 14013 5117 14047 5151
rect 16221 5117 16255 5151
rect 16548 5117 16582 5151
rect 18705 5117 18739 5151
rect 20913 5117 20947 5151
rect 21649 5117 21683 5151
rect 23305 5117 23339 5151
rect 23581 5117 23615 5151
rect 23857 5117 23891 5151
rect 24593 5117 24627 5151
rect 26525 5117 26559 5151
rect 26709 5117 26743 5151
rect 3341 5049 3375 5083
rect 8217 5049 8251 5083
rect 6567 4981 6601 5015
rect 9511 4981 9545 5015
rect 11069 4981 11103 5015
rect 11719 4981 11753 5015
rect 13737 4981 13771 5015
rect 19171 4981 19205 5015
rect 21379 4981 21413 5015
rect 22753 4981 22787 5015
rect 23121 4981 23155 5015
rect 24323 4981 24357 5015
rect 26341 4981 26375 5015
rect 27175 4981 27209 5015
rect 2697 4777 2731 4811
rect 3991 4777 4025 4811
rect 7849 4777 7883 4811
rect 10977 4777 11011 4811
rect 12087 4777 12121 4811
rect 13645 4777 13679 4811
rect 14295 4777 14329 4811
rect 16687 4777 16721 4811
rect 19447 4777 19481 4811
rect 24225 4777 24259 4811
rect 24593 4777 24627 4811
rect 18337 4709 18371 4743
rect 857 4641 891 4675
rect 3433 4641 3467 4675
rect 4261 4641 4295 4675
rect 5641 4641 5675 4675
rect 8585 4641 8619 4675
rect 11161 4641 11195 4675
rect 11437 4641 11471 4675
rect 11621 4641 11655 4675
rect 12357 4641 12391 4675
rect 14565 4641 14599 4675
rect 15945 4641 15979 4675
rect 16957 4641 16991 4675
rect 18429 4641 18463 4675
rect 21465 4641 21499 4675
rect 21741 4641 21775 4675
rect 22017 4641 22051 4675
rect 22201 4641 22235 4675
rect 22937 4641 22971 4675
rect 24777 4641 24811 4675
rect 27077 4641 27111 4675
rect 27997 4641 28031 4675
rect 28733 4641 28767 4675
rect 1184 4573 1218 4607
rect 1363 4573 1397 4607
rect 1593 4573 1627 4607
rect 3525 4573 3559 4607
rect 3988 4573 4022 4607
rect 6009 4573 6043 4607
rect 6336 4573 6370 4607
rect 6472 4575 6506 4609
rect 6745 4573 6779 4607
rect 8677 4573 8711 4607
rect 9004 4573 9038 4607
rect 9140 4575 9174 4609
rect 9413 4573 9447 4607
rect 12084 4591 12118 4625
rect 13829 4573 13863 4607
rect 14292 4573 14326 4607
rect 16221 4573 16255 4607
rect 16684 4575 16718 4609
rect 18705 4573 18739 4607
rect 18981 4573 19015 4607
rect 19487 4573 19521 4607
rect 19717 4573 19751 4607
rect 22528 4573 22562 4607
rect 22664 4575 22698 4609
rect 28324 4573 28358 4607
rect 28503 4573 28537 4607
rect 8401 4505 8435 4539
rect 11253 4505 11287 4539
rect 29837 4505 29871 4539
rect 3249 4437 3283 4471
rect 10701 4437 10735 4471
rect 21005 4437 21039 4471
rect 21281 4437 21315 4471
rect 21557 4437 21591 4471
rect 21833 4437 21867 4471
rect 25053 4437 25087 4471
rect 26893 4437 26927 4471
rect 8953 4233 8987 4267
rect 11989 4233 12023 4267
rect 9873 4165 9907 4199
rect 949 4097 983 4131
rect 1445 4079 1479 4113
rect 3525 4097 3559 4131
rect 4307 4095 4341 4129
rect 4537 4097 4571 4131
rect 6472 4097 6506 4131
rect 8125 4097 8159 4131
rect 8677 4097 8711 4131
rect 10149 4097 10183 4131
rect 10612 4097 10646 4131
rect 10885 4097 10919 4131
rect 12541 4097 12575 4131
rect 14476 4097 14510 4131
rect 16129 4097 16163 4131
rect 16684 4097 16718 4131
rect 18337 4097 18371 4131
rect 19168 4097 19202 4131
rect 19441 4097 19475 4131
rect 20821 4097 20855 4131
rect 21376 4097 21410 4131
rect 21649 4097 21683 4131
rect 25145 4097 25179 4131
rect 26436 4097 26470 4131
rect 26709 4097 26743 4131
rect 1685 4029 1719 4063
rect 3249 4029 3283 4063
rect 3801 4029 3835 4063
rect 6009 4029 6043 4063
rect 6745 4029 6779 4063
rect 8401 4029 8435 4063
rect 9137 4029 9171 4063
rect 9505 4029 9539 4063
rect 9781 4029 9815 4063
rect 10057 4029 10091 4063
rect 12357 4029 12391 4063
rect 13921 4029 13955 4063
rect 14013 4029 14047 4063
rect 14749 4029 14783 4063
rect 16221 4029 16255 4063
rect 16957 4029 16991 4063
rect 18705 4029 18739 4063
rect 20913 4029 20947 4063
rect 21240 4029 21274 4063
rect 23121 4029 23155 4063
rect 24041 4029 24075 4063
rect 24317 4029 24351 4063
rect 24593 4029 24627 4063
rect 24869 4029 24903 4063
rect 25973 4029 26007 4063
rect 28181 4029 28215 4063
rect 29009 4029 29043 4063
rect 5917 3961 5951 3995
rect 13001 3961 13035 3995
rect 23397 3961 23431 3995
rect 1415 3893 1449 3927
rect 2789 3893 2823 3927
rect 4267 3893 4301 3927
rect 6475 3893 6509 3927
rect 9321 3893 9355 3927
rect 9597 3893 9631 3927
rect 10615 3893 10649 3927
rect 13093 3893 13127 3927
rect 13737 3893 13771 3927
rect 14479 3893 14513 3927
rect 16687 3893 16721 3927
rect 19171 3893 19205 3927
rect 22753 3893 22787 3927
rect 23857 3893 23891 3927
rect 24133 3893 24167 3927
rect 24409 3893 24443 3927
rect 24685 3893 24719 3927
rect 25513 3893 25547 3927
rect 26439 3893 26473 3927
rect 27813 3893 27847 3927
rect 28365 3893 28399 3927
rect 29193 3893 29227 3927
rect 1041 3689 1075 3723
rect 6935 3689 6969 3723
rect 11529 3689 11563 3723
rect 14105 3689 14139 3723
rect 15853 3689 15887 3723
rect 27077 3689 27111 3723
rect 29745 3689 29779 3723
rect 3433 3621 3467 3655
rect 11253 3621 11287 3655
rect 15025 3621 15059 3655
rect 15577 3621 15611 3655
rect 16497 3621 16531 3655
rect 21373 3621 21407 3655
rect 1225 3553 1259 3587
rect 6009 3553 6043 3587
rect 6469 3553 6503 3587
rect 7205 3553 7239 3587
rect 8585 3553 8619 3587
rect 9413 3553 9447 3587
rect 10977 3553 11011 3587
rect 11713 3553 11747 3587
rect 11989 3553 12023 3587
rect 12081 3553 12115 3587
rect 12817 3553 12851 3587
rect 14473 3553 14507 3587
rect 16221 3553 16255 3587
rect 17509 3553 17543 3587
rect 19308 3553 19342 3587
rect 21097 3553 21131 3587
rect 22017 3553 22051 3587
rect 22528 3553 22562 3587
rect 22937 3553 22971 3587
rect 24593 3537 24627 3571
rect 24685 3553 24719 3587
rect 25421 3577 25455 3611
rect 25697 3553 25731 3587
rect 25973 3553 26007 3587
rect 26709 3553 26743 3587
rect 27261 3553 27295 3587
rect 27353 3553 27387 3587
rect 27905 3553 27939 3587
rect 28232 3553 28266 3587
rect 28641 3553 28675 3587
rect 1317 3485 1351 3519
rect 1644 3485 1678 3519
rect 1813 3503 1847 3537
rect 2053 3485 2087 3519
rect 3525 3485 3559 3519
rect 3852 3485 3886 3519
rect 3988 3503 4022 3537
rect 4261 3485 4295 3519
rect 5641 3485 5675 3519
rect 6975 3485 7009 3519
rect 8677 3485 8711 3519
rect 9004 3485 9038 3519
rect 9140 3487 9174 3521
rect 12408 3485 12442 3519
rect 12544 3485 12578 3519
rect 16773 3485 16807 3519
rect 17100 3485 17134 3519
rect 17279 3485 17313 3519
rect 18981 3485 19015 3519
rect 19487 3485 19521 3519
rect 19717 3485 19751 3519
rect 22201 3485 22235 3519
rect 22664 3487 22698 3521
rect 24961 3485 24995 3519
rect 27537 3485 27571 3519
rect 28368 3485 28402 3519
rect 6193 3417 6227 3451
rect 10517 3417 10551 3451
rect 15209 3417 15243 3451
rect 25789 3417 25823 3451
rect 11805 3349 11839 3383
rect 14565 3349 14599 3383
rect 18613 3349 18647 3383
rect 21465 3349 21499 3383
rect 21833 3349 21867 3383
rect 24225 3349 24259 3383
rect 24409 3349 24443 3383
rect 25237 3349 25271 3383
rect 25513 3349 25547 3383
rect 26525 3349 26559 3383
rect 2973 3145 3007 3179
rect 949 3009 983 3043
rect 1445 2991 1479 3025
rect 4356 3009 4390 3043
rect 4629 3009 4663 3043
rect 6009 3009 6043 3043
rect 6564 3009 6598 3043
rect 6837 3009 6871 3043
rect 8217 3009 8251 3043
rect 9508 3009 9542 3043
rect 11161 3009 11195 3043
rect 11716 3009 11750 3043
rect 13369 3009 13403 3043
rect 14568 3009 14602 3043
rect 16221 3009 16255 3043
rect 16776 3009 16810 3043
rect 18429 3009 18463 3043
rect 19168 3009 19202 3043
rect 19441 3009 19475 3043
rect 20821 3009 20855 3043
rect 21376 3009 21410 3043
rect 21649 3009 21683 3043
rect 23029 3009 23063 3043
rect 24320 3009 24354 3043
rect 24593 3009 24627 3043
rect 26065 3009 26099 3043
rect 26392 3009 26426 3043
rect 26528 3009 26562 3043
rect 26801 3009 26835 3043
rect 29009 3009 29043 3043
rect 1685 2941 1719 2975
rect 3341 2941 3375 2975
rect 3617 2941 3651 2975
rect 3893 2941 3927 2975
rect 6101 2941 6135 2975
rect 8585 2941 8619 2975
rect 9045 2941 9079 2975
rect 9781 2941 9815 2975
rect 11253 2941 11287 2975
rect 11989 2941 12023 2975
rect 13553 2941 13587 2975
rect 14105 2941 14139 2975
rect 14432 2941 14466 2975
rect 14841 2941 14875 2975
rect 16313 2941 16347 2975
rect 16640 2941 16674 2975
rect 17049 2941 17083 2975
rect 18705 2941 18739 2975
rect 20913 2941 20947 2975
rect 21240 2941 21274 2975
rect 23213 2941 23247 2975
rect 23857 2941 23891 2975
rect 29285 2941 29319 2975
rect 13829 2873 13863 2907
rect 25973 2873 26007 2907
rect 1415 2805 1449 2839
rect 4359 2805 4393 2839
rect 6567 2805 6601 2839
rect 8677 2805 8711 2839
rect 9511 2805 9545 2839
rect 11719 2805 11753 2839
rect 19171 2805 19205 2839
rect 23305 2805 23339 2839
rect 24323 2805 24357 2839
rect 27905 2805 27939 2839
rect 1507 2601 1541 2635
rect 3065 2601 3099 2635
rect 5089 2601 5123 2635
rect 6291 2601 6325 2635
rect 7665 2601 7699 2635
rect 9143 2601 9177 2635
rect 11161 2601 11195 2635
rect 16687 2601 16721 2635
rect 21747 2601 21781 2635
rect 23857 2601 23891 2635
rect 27629 2601 27663 2635
rect 28463 2601 28497 2635
rect 29837 2601 29871 2635
rect 8309 2533 8343 2567
rect 10793 2533 10827 2567
rect 20545 2533 20579 2567
rect 1041 2465 1075 2499
rect 3576 2465 3610 2499
rect 5641 2465 5675 2499
rect 8033 2465 8067 2499
rect 9413 2465 9447 2499
rect 11069 2465 11103 2499
rect 11621 2465 11655 2499
rect 13737 2465 13771 2499
rect 16221 2465 16255 2499
rect 18429 2465 18463 2499
rect 18756 2465 18790 2499
rect 20637 2465 20671 2499
rect 21281 2465 21315 2499
rect 23581 2465 23615 2499
rect 24133 2465 24167 2499
rect 24869 2465 24903 2499
rect 26617 2465 26651 2499
rect 26709 2465 26743 2499
rect 27353 2465 27387 2499
rect 27997 2465 28031 2499
rect 28733 2465 28767 2499
rect 1547 2397 1581 2431
rect 1777 2397 1811 2431
rect 3249 2397 3283 2431
rect 3755 2397 3789 2431
rect 3985 2397 4019 2431
rect 5825 2397 5859 2431
rect 6288 2397 6322 2431
rect 6561 2397 6595 2431
rect 8677 2397 8711 2431
rect 9140 2397 9174 2431
rect 11948 2397 11982 2431
rect 12084 2399 12118 2433
rect 12357 2397 12391 2431
rect 13829 2397 13863 2431
rect 14156 2397 14190 2431
rect 14292 2397 14326 2431
rect 14565 2397 14599 2431
rect 15945 2397 15979 2431
rect 16684 2397 16718 2431
rect 16957 2397 16991 2431
rect 18337 2397 18371 2431
rect 18892 2415 18926 2449
rect 19165 2397 19199 2431
rect 20821 2397 20855 2431
rect 21744 2399 21778 2433
rect 22017 2397 22051 2431
rect 24460 2397 24494 2431
rect 24629 2399 24663 2433
rect 26893 2397 26927 2431
rect 28460 2397 28494 2431
rect 26433 2329 26467 2363
rect 5457 2261 5491 2295
rect 23305 2261 23339 2295
rect 25973 2261 26007 2295
rect 3249 2057 3283 2091
rect 13645 2057 13679 2091
rect 18337 2057 18371 2091
rect 23121 2057 23155 2091
rect 25881 2057 25915 2091
rect 28181 2057 28215 2091
rect 29193 2057 29227 2091
rect 29469 2057 29503 2091
rect 1455 1921 1489 1955
rect 3852 1921 3886 1955
rect 3988 1919 4022 1953
rect 4261 1921 4295 1955
rect 6101 1921 6135 1955
rect 6564 1921 6598 1955
rect 6837 1921 6871 1955
rect 8217 1921 8251 1955
rect 9508 1921 9542 1955
rect 9781 1921 9815 1955
rect 11161 1921 11195 1955
rect 11716 1921 11750 1955
rect 13369 1921 13403 1955
rect 14384 1921 14418 1955
rect 16129 1921 16163 1955
rect 16592 1903 16626 1937
rect 18245 1921 18279 1955
rect 19168 1921 19202 1955
rect 20821 1921 20855 1955
rect 21376 1921 21410 1955
rect 21649 1921 21683 1955
rect 24320 1903 24354 1937
rect 24593 1921 24627 1955
rect 26341 1921 26375 1955
rect 26847 1921 26881 1955
rect 949 1853 983 1887
rect 1685 1853 1719 1887
rect 3433 1853 3467 1887
rect 3525 1853 3559 1887
rect 8401 1853 8435 1887
rect 9045 1853 9079 1887
rect 11253 1853 11287 1887
rect 11989 1853 12023 1887
rect 13829 1853 13863 1887
rect 13921 1853 13955 1887
rect 14657 1853 14691 1887
rect 16037 1853 16071 1887
rect 16865 1853 16899 1887
rect 18521 1853 18555 1887
rect 18705 1853 18739 1887
rect 19032 1853 19066 1887
rect 19441 1853 19475 1887
rect 20913 1853 20947 1887
rect 21240 1853 21274 1887
rect 23305 1853 23339 1887
rect 23581 1853 23615 1887
rect 23857 1853 23891 1887
rect 26241 1853 26275 1887
rect 26668 1853 26702 1887
rect 27077 1853 27111 1887
rect 28549 1853 28583 1887
rect 29018 1853 29052 1887
rect 29285 1853 29319 1887
rect 3065 1785 3099 1819
rect 8677 1785 8711 1819
rect 23029 1785 23063 1819
rect 1415 1717 1449 1751
rect 5365 1717 5399 1751
rect 6009 1717 6043 1751
rect 6567 1717 6601 1751
rect 9511 1717 9545 1751
rect 11719 1717 11753 1751
rect 14387 1717 14421 1751
rect 16595 1717 16629 1751
rect 23397 1717 23431 1751
rect 24323 1717 24357 1751
rect 26065 1717 26099 1751
rect 28733 1717 28767 1751
rect 857 1513 891 1547
rect 3157 1513 3191 1547
rect 6935 1513 6969 1547
rect 8493 1513 8527 1547
rect 12087 1513 12121 1547
rect 16687 1513 16721 1547
rect 18895 1513 18929 1547
rect 20913 1513 20947 1547
rect 21747 1513 21781 1547
rect 28273 1513 28307 1547
rect 29101 1513 29135 1547
rect 29653 1513 29687 1547
rect 5917 1445 5951 1479
rect 10793 1445 10827 1479
rect 20545 1445 20579 1479
rect 25789 1445 25823 1479
rect 1041 1377 1075 1411
rect 1317 1377 1351 1411
rect 2605 1377 2639 1411
rect 2881 1377 2915 1411
rect 3065 1377 3099 1411
rect 5641 1377 5675 1411
rect 6469 1377 6503 1411
rect 11161 1377 11195 1411
rect 11529 1377 11563 1411
rect 11621 1377 11655 1411
rect 13737 1377 13771 1411
rect 16221 1377 16255 1411
rect 18337 1377 18371 1411
rect 20821 1377 20855 1411
rect 21097 1377 21131 1411
rect 23397 1377 23431 1411
rect 23816 1377 23850 1411
rect 28825 1361 28859 1395
rect 28917 1377 28951 1411
rect 29193 1377 29227 1411
rect 29469 1377 29503 1411
rect 2329 1309 2363 1343
rect 3525 1309 3559 1343
rect 3852 1309 3886 1343
rect 3988 1309 4022 1343
rect 4261 1309 4295 1343
rect 6193 1309 6227 1343
rect 6932 1309 6966 1343
rect 7205 1309 7239 1343
rect 8677 1309 8711 1343
rect 9004 1309 9038 1343
rect 9183 1309 9217 1343
rect 9413 1309 9447 1343
rect 12084 1309 12118 1343
rect 12357 1309 12391 1343
rect 13829 1309 13863 1343
rect 14156 1309 14190 1343
rect 14292 1309 14326 1343
rect 14565 1309 14599 1343
rect 15945 1309 15979 1343
rect 16684 1309 16718 1343
rect 16957 1309 16991 1343
rect 18429 1309 18463 1343
rect 18892 1309 18926 1343
rect 19165 1309 19199 1343
rect 21281 1309 21315 1343
rect 21744 1327 21778 1361
rect 22017 1309 22051 1343
rect 23489 1309 23523 1343
rect 23952 1309 23986 1343
rect 24225 1309 24259 1343
rect 26433 1309 26467 1343
rect 26760 1309 26794 1343
rect 26896 1311 26930 1345
rect 27169 1309 27203 1343
rect 1133 1241 1167 1275
rect 1961 1241 1995 1275
rect 10977 1241 11011 1275
rect 25973 1241 26007 1275
rect 29929 1241 29963 1275
rect 2421 1173 2455 1207
rect 2697 1173 2731 1207
rect 11345 1173 11379 1207
rect 20637 1173 20671 1207
rect 25329 1173 25363 1207
rect 28641 1173 28675 1207
rect 29377 1173 29411 1207
rect 2973 969 3007 1003
rect 7665 969 7699 1003
rect 10241 969 10275 1003
rect 10609 969 10643 1003
rect 10977 969 11011 1003
rect 13277 969 13311 1003
rect 13553 969 13587 1003
rect 16129 969 16163 1003
rect 18705 969 18739 1003
rect 26433 969 26467 1003
rect 28549 969 28583 1003
rect 21281 901 21315 935
rect 949 833 983 867
rect 1445 815 1479 849
rect 1685 833 1719 867
rect 6288 831 6322 865
rect 8401 833 8435 867
rect 8864 833 8898 867
rect 11759 833 11793 867
rect 14335 831 14369 865
rect 16911 833 16945 867
rect 17141 833 17175 867
rect 19487 833 19521 867
rect 21557 833 21591 867
rect 22063 833 22097 867
rect 24320 833 24354 867
rect 24593 833 24627 867
rect 26709 833 26743 867
rect 27215 833 27249 867
rect 27445 833 27479 867
rect 3893 765 3927 799
rect 4997 765 5031 799
rect 5641 765 5675 799
rect 5825 765 5859 799
rect 6561 765 6595 799
rect 9137 765 9171 799
rect 10793 765 10827 799
rect 11161 765 11195 799
rect 11253 765 11287 799
rect 11989 765 12023 799
rect 13729 765 13763 799
rect 13829 765 13863 799
rect 14156 765 14190 799
rect 14565 765 14599 799
rect 16313 765 16347 799
rect 16405 765 16439 799
rect 18889 765 18923 799
rect 18981 765 19015 799
rect 19717 765 19751 799
rect 21465 765 21499 799
rect 21884 765 21918 799
rect 22293 765 22327 799
rect 23673 765 23707 799
rect 23857 765 23891 799
rect 26249 765 26283 799
rect 26617 765 26651 799
rect 27036 765 27070 799
rect 29009 765 29043 799
rect 15945 697 15979 731
rect 1415 629 1449 663
rect 3525 629 3559 663
rect 5365 629 5399 663
rect 5457 629 5491 663
rect 6291 629 6325 663
rect 8867 629 8901 663
rect 11719 629 11753 663
rect 16871 629 16905 663
rect 18245 629 18279 663
rect 19447 629 19481 663
rect 20821 629 20855 663
rect 24323 629 24357 663
rect 25697 629 25731 663
rect 26065 629 26099 663
rect 29193 629 29227 663
<< metal1 >>
rect 1946 22244 1952 22296
rect 2004 22284 2010 22296
rect 8846 22284 8852 22296
rect 2004 22256 8852 22284
rect 2004 22244 2010 22256
rect 8846 22244 8852 22256
rect 8904 22244 8910 22296
rect 9674 22284 9680 22296
rect 9048 22256 9680 22284
rect 4062 22176 4068 22228
rect 4120 22216 4126 22228
rect 9048 22216 9076 22256
rect 9674 22244 9680 22256
rect 9732 22244 9738 22296
rect 18782 22244 18788 22296
rect 18840 22284 18846 22296
rect 23566 22284 23572 22296
rect 18840 22256 23572 22284
rect 18840 22244 18846 22256
rect 23566 22244 23572 22256
rect 23624 22244 23630 22296
rect 25958 22284 25964 22296
rect 23676 22256 25964 22284
rect 4120 22188 9076 22216
rect 4120 22176 4126 22188
rect 9122 22176 9128 22228
rect 9180 22216 9186 22228
rect 9766 22216 9772 22228
rect 9180 22188 9772 22216
rect 9180 22176 9186 22188
rect 9766 22176 9772 22188
rect 9824 22176 9830 22228
rect 10796 22188 12848 22216
rect 3050 22108 3056 22160
rect 3108 22148 3114 22160
rect 10796 22148 10824 22188
rect 12820 22160 12848 22188
rect 12894 22176 12900 22228
rect 12952 22216 12958 22228
rect 12952 22188 18276 22216
rect 12952 22176 12958 22188
rect 3108 22120 10824 22148
rect 3108 22108 3114 22120
rect 12802 22108 12808 22160
rect 12860 22108 12866 22160
rect 5258 22040 5264 22092
rect 5316 22080 5322 22092
rect 5316 22052 6960 22080
rect 5316 22040 5322 22052
rect 6932 22012 6960 22052
rect 9582 22040 9588 22092
rect 9640 22080 9646 22092
rect 12434 22080 12440 22092
rect 9640 22052 12440 22080
rect 9640 22040 9646 22052
rect 12434 22040 12440 22052
rect 12492 22040 12498 22092
rect 18248 22080 18276 22188
rect 18506 22176 18512 22228
rect 18564 22216 18570 22228
rect 22370 22216 22376 22228
rect 18564 22188 22376 22216
rect 18564 22176 18570 22188
rect 22370 22176 22376 22188
rect 22428 22176 22434 22228
rect 22462 22176 22468 22228
rect 22520 22216 22526 22228
rect 23676 22216 23704 22256
rect 25958 22244 25964 22256
rect 26016 22244 26022 22296
rect 22520 22188 23704 22216
rect 22520 22176 22526 22188
rect 23750 22176 23756 22228
rect 23808 22216 23814 22228
rect 28718 22216 28724 22228
rect 23808 22188 28724 22216
rect 23808 22176 23814 22188
rect 28718 22176 28724 22188
rect 28776 22176 28782 22228
rect 18598 22108 18604 22160
rect 18656 22148 18662 22160
rect 28074 22148 28080 22160
rect 18656 22120 28080 22148
rect 18656 22108 18662 22120
rect 28074 22108 28080 22120
rect 28132 22108 28138 22160
rect 28166 22080 28172 22092
rect 18248 22052 28172 22080
rect 28166 22040 28172 22052
rect 28224 22040 28230 22092
rect 12618 22012 12624 22024
rect 6932 21984 12624 22012
rect 12618 21972 12624 21984
rect 12676 21972 12682 22024
rect 28350 22012 28356 22024
rect 18156 21984 19380 22012
rect 2148 21916 6322 21944
rect 2148 21888 2176 21916
rect 2130 21836 2136 21888
rect 2188 21836 2194 21888
rect 2498 21836 2504 21888
rect 2556 21876 2562 21888
rect 3786 21876 3792 21888
rect 2556 21848 3792 21876
rect 2556 21836 2562 21848
rect 3786 21836 3792 21848
rect 3844 21836 3850 21888
rect 6294 21876 6322 21916
rect 7190 21904 7196 21956
rect 7248 21944 7254 21956
rect 16114 21944 16120 21956
rect 7248 21916 16120 21944
rect 7248 21904 7254 21916
rect 16114 21904 16120 21916
rect 16172 21904 16178 21956
rect 18156 21944 18184 21984
rect 16224 21916 18184 21944
rect 8754 21876 8760 21888
rect 6294 21848 8760 21876
rect 8754 21836 8760 21848
rect 8812 21836 8818 21888
rect 8846 21836 8852 21888
rect 8904 21876 8910 21888
rect 12526 21876 12532 21888
rect 8904 21848 12532 21876
rect 8904 21836 8910 21848
rect 12526 21836 12532 21848
rect 12584 21836 12590 21888
rect 13722 21836 13728 21888
rect 13780 21876 13786 21888
rect 16224 21876 16252 21916
rect 18414 21904 18420 21956
rect 18472 21944 18478 21956
rect 19242 21944 19248 21956
rect 18472 21916 19248 21944
rect 18472 21904 18478 21916
rect 19242 21904 19248 21916
rect 19300 21904 19306 21956
rect 19352 21944 19380 21984
rect 23216 21984 28356 22012
rect 23216 21944 23244 21984
rect 28350 21972 28356 21984
rect 28408 21972 28414 22024
rect 19352 21916 23244 21944
rect 23290 21904 23296 21956
rect 23348 21944 23354 21956
rect 23348 21916 30512 21944
rect 23348 21904 23354 21916
rect 30484 21888 30512 21916
rect 13780 21848 16252 21876
rect 13780 21836 13786 21848
rect 16666 21836 16672 21888
rect 16724 21876 16730 21888
rect 21358 21876 21364 21888
rect 16724 21848 21364 21876
rect 16724 21836 16730 21848
rect 21358 21836 21364 21848
rect 21416 21836 21422 21888
rect 22278 21836 22284 21888
rect 22336 21876 22342 21888
rect 26602 21876 26608 21888
rect 22336 21848 26608 21876
rect 22336 21836 22342 21848
rect 26602 21836 26608 21848
rect 26660 21836 26666 21888
rect 30466 21836 30472 21888
rect 30524 21836 30530 21888
rect 552 21786 30912 21808
rect 552 21734 4193 21786
rect 4245 21734 4257 21786
rect 4309 21734 4321 21786
rect 4373 21734 4385 21786
rect 4437 21734 4449 21786
rect 4501 21734 11783 21786
rect 11835 21734 11847 21786
rect 11899 21734 11911 21786
rect 11963 21734 11975 21786
rect 12027 21734 12039 21786
rect 12091 21734 19373 21786
rect 19425 21734 19437 21786
rect 19489 21734 19501 21786
rect 19553 21734 19565 21786
rect 19617 21734 19629 21786
rect 19681 21734 26963 21786
rect 27015 21734 27027 21786
rect 27079 21734 27091 21786
rect 27143 21734 27155 21786
rect 27207 21734 27219 21786
rect 27271 21734 30912 21786
rect 552 21712 30912 21734
rect 2774 21672 2780 21684
rect 952 21644 2780 21672
rect 952 21545 980 21644
rect 2774 21632 2780 21644
rect 2832 21632 2838 21684
rect 8202 21672 8208 21684
rect 3252 21644 5120 21672
rect 937 21539 995 21545
rect 937 21505 949 21539
rect 983 21505 995 21539
rect 937 21499 995 21505
rect 1443 21539 1501 21545
rect 1443 21505 1455 21539
rect 1489 21536 1501 21539
rect 3252 21536 3280 21644
rect 5092 21613 5120 21644
rect 5552 21644 8208 21672
rect 5552 21616 5580 21644
rect 8202 21632 8208 21644
rect 8260 21632 8266 21684
rect 8312 21644 12434 21672
rect 5077 21607 5135 21613
rect 5077 21573 5089 21607
rect 5123 21573 5135 21607
rect 5077 21567 5135 21573
rect 5534 21564 5540 21616
rect 5592 21564 5598 21616
rect 8312 21604 8340 21644
rect 8128 21576 8340 21604
rect 1489 21508 3280 21536
rect 1489 21505 1501 21508
rect 1443 21499 1501 21505
rect 3418 21496 3424 21548
rect 3476 21536 3482 21548
rect 3700 21539 3758 21545
rect 3700 21536 3712 21539
rect 3476 21508 3712 21536
rect 3476 21496 3482 21508
rect 3700 21505 3712 21508
rect 3746 21505 3758 21539
rect 6276 21539 6334 21545
rect 6276 21536 6288 21539
rect 3700 21499 3758 21505
rect 3896 21508 6288 21536
rect 1670 21428 1676 21480
rect 1728 21428 1734 21480
rect 3234 21428 3240 21480
rect 3292 21428 3298 21480
rect 3896 21468 3924 21508
rect 6276 21505 6288 21508
rect 6322 21505 6334 21539
rect 6276 21499 6334 21505
rect 6549 21539 6607 21545
rect 6549 21505 6561 21539
rect 6595 21536 6607 21539
rect 8128 21536 8156 21576
rect 6595 21508 8156 21536
rect 8852 21537 8910 21543
rect 6595 21505 6607 21508
rect 6549 21499 6607 21505
rect 8852 21503 8864 21537
rect 8898 21536 8910 21537
rect 8938 21536 8944 21548
rect 8898 21508 8944 21536
rect 8898 21503 8910 21508
rect 8852 21497 8910 21503
rect 8938 21496 8944 21508
rect 8996 21496 9002 21548
rect 9122 21496 9128 21548
rect 9180 21496 9186 21548
rect 9490 21496 9496 21548
rect 9548 21536 9554 21548
rect 11428 21539 11486 21545
rect 11428 21536 11440 21539
rect 9548 21508 11440 21536
rect 9548 21496 9554 21508
rect 11428 21505 11440 21508
rect 11474 21505 11486 21539
rect 11428 21499 11486 21505
rect 3344 21440 3924 21468
rect 3053 21403 3111 21409
rect 3053 21369 3065 21403
rect 3099 21400 3111 21403
rect 3344 21400 3372 21440
rect 3970 21428 3976 21480
rect 4028 21428 4034 21480
rect 4798 21428 4804 21480
rect 4856 21468 4862 21480
rect 5534 21468 5540 21480
rect 4856 21440 5540 21468
rect 4856 21428 4862 21440
rect 5534 21428 5540 21440
rect 5592 21468 5598 21480
rect 5629 21471 5687 21477
rect 5629 21468 5641 21471
rect 5592 21440 5641 21468
rect 5592 21428 5598 21440
rect 5629 21437 5641 21440
rect 5675 21437 5687 21471
rect 5629 21431 5687 21437
rect 5813 21471 5871 21477
rect 5813 21437 5825 21471
rect 5859 21468 5871 21471
rect 5902 21468 5908 21480
rect 5859 21440 5908 21468
rect 5859 21437 5871 21440
rect 5813 21431 5871 21437
rect 5902 21428 5908 21440
rect 5960 21428 5966 21480
rect 8202 21428 8208 21480
rect 8260 21428 8266 21480
rect 8386 21428 8392 21480
rect 8444 21428 8450 21480
rect 8662 21468 8668 21480
rect 8496 21440 8668 21468
rect 3099 21372 3372 21400
rect 4632 21372 5856 21400
rect 3099 21369 3111 21372
rect 3053 21363 3111 21369
rect 1394 21292 1400 21344
rect 1452 21341 1458 21344
rect 1452 21332 1461 21341
rect 1452 21304 1497 21332
rect 1452 21295 1461 21304
rect 1452 21292 1458 21295
rect 3510 21292 3516 21344
rect 3568 21332 3574 21344
rect 3703 21335 3761 21341
rect 3703 21332 3715 21335
rect 3568 21304 3715 21332
rect 3568 21292 3574 21304
rect 3703 21301 3715 21304
rect 3749 21332 3761 21335
rect 4632 21332 4660 21372
rect 3749 21304 4660 21332
rect 3749 21301 3761 21304
rect 3703 21295 3761 21301
rect 5442 21292 5448 21344
rect 5500 21292 5506 21344
rect 5828 21332 5856 21372
rect 7558 21360 7564 21412
rect 7616 21400 7622 21412
rect 8496 21400 8524 21440
rect 8639 21436 8668 21440
rect 8662 21428 8668 21436
rect 8720 21477 8726 21480
rect 8720 21471 8774 21477
rect 8720 21437 8728 21471
rect 8762 21437 8774 21471
rect 8720 21431 8774 21437
rect 8720 21428 8726 21431
rect 9398 21428 9404 21480
rect 9456 21468 9462 21480
rect 10686 21468 10692 21480
rect 9456 21440 10692 21468
rect 9456 21428 9462 21440
rect 10686 21428 10692 21440
rect 10744 21428 10750 21480
rect 10781 21471 10839 21477
rect 10781 21437 10793 21471
rect 10827 21468 10839 21471
rect 10870 21468 10876 21480
rect 10827 21440 10876 21468
rect 10827 21437 10839 21440
rect 10781 21431 10839 21437
rect 10870 21428 10876 21440
rect 10928 21428 10934 21480
rect 10962 21428 10968 21480
rect 11020 21428 11026 21480
rect 11054 21428 11060 21480
rect 11112 21468 11118 21480
rect 11292 21471 11350 21477
rect 11292 21468 11304 21471
rect 11112 21440 11304 21468
rect 11112 21428 11118 21440
rect 11292 21437 11304 21440
rect 11338 21437 11350 21471
rect 11292 21431 11350 21437
rect 11606 21428 11612 21480
rect 11664 21468 11670 21480
rect 11701 21471 11759 21477
rect 11701 21468 11713 21471
rect 11664 21440 11713 21468
rect 11664 21428 11670 21440
rect 11701 21437 11713 21440
rect 11747 21437 11759 21471
rect 11701 21431 11759 21437
rect 12406 21400 12434 21644
rect 12526 21632 12532 21684
rect 12584 21632 12590 21684
rect 12802 21632 12808 21684
rect 12860 21632 12866 21684
rect 16114 21632 16120 21684
rect 16172 21632 16178 21684
rect 18417 21675 18475 21681
rect 16592 21644 17816 21672
rect 12544 21604 12572 21632
rect 13906 21604 13912 21616
rect 12544 21576 13912 21604
rect 13906 21564 13912 21576
rect 13964 21564 13970 21616
rect 12618 21496 12624 21548
rect 12676 21536 12682 21548
rect 13262 21536 13268 21548
rect 12676 21508 13268 21536
rect 12676 21496 12682 21508
rect 13262 21496 13268 21508
rect 13320 21536 13326 21548
rect 13722 21536 13728 21548
rect 13320 21508 13728 21536
rect 13320 21496 13326 21508
rect 13372 21477 13400 21508
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 16132 21545 16160 21632
rect 14277 21539 14335 21545
rect 14277 21505 14289 21539
rect 14323 21536 14335 21539
rect 16117 21539 16175 21545
rect 14323 21508 14688 21536
rect 14323 21505 14335 21508
rect 14277 21499 14335 21505
rect 14660 21480 14688 21508
rect 16117 21505 16129 21539
rect 16163 21505 16175 21539
rect 16117 21499 16175 21505
rect 13357 21471 13415 21477
rect 13357 21437 13369 21471
rect 13403 21437 13415 21471
rect 14090 21468 14096 21480
rect 13357 21431 13415 21437
rect 13556 21440 14096 21468
rect 13556 21400 13584 21440
rect 14090 21428 14096 21440
rect 14148 21428 14154 21480
rect 14366 21428 14372 21480
rect 14424 21468 14430 21480
rect 14553 21471 14611 21477
rect 14553 21468 14565 21471
rect 14424 21440 14565 21468
rect 14424 21428 14430 21440
rect 14553 21437 14565 21440
rect 14599 21437 14611 21471
rect 14553 21431 14611 21437
rect 14642 21428 14648 21480
rect 14700 21428 14706 21480
rect 7616 21372 8524 21400
rect 9968 21372 11100 21400
rect 12406 21372 13584 21400
rect 13633 21403 13691 21409
rect 7616 21360 7622 21372
rect 6178 21332 6184 21344
rect 5828 21304 6184 21332
rect 6178 21292 6184 21304
rect 6236 21292 6242 21344
rect 6270 21292 6276 21344
rect 6328 21341 6334 21344
rect 6328 21332 6337 21341
rect 6328 21304 6373 21332
rect 6328 21295 6337 21304
rect 6328 21292 6334 21295
rect 6638 21292 6644 21344
rect 6696 21332 6702 21344
rect 7653 21335 7711 21341
rect 7653 21332 7665 21335
rect 6696 21304 7665 21332
rect 6696 21292 6702 21304
rect 7653 21301 7665 21304
rect 7699 21301 7711 21335
rect 7653 21295 7711 21301
rect 7834 21292 7840 21344
rect 7892 21332 7898 21344
rect 8021 21335 8079 21341
rect 8021 21332 8033 21335
rect 7892 21304 8033 21332
rect 7892 21292 7898 21304
rect 8021 21301 8033 21304
rect 8067 21301 8079 21335
rect 8021 21295 8079 21301
rect 8478 21292 8484 21344
rect 8536 21332 8542 21344
rect 9968 21332 9996 21372
rect 8536 21304 9996 21332
rect 8536 21292 8542 21304
rect 10042 21292 10048 21344
rect 10100 21332 10106 21344
rect 10229 21335 10287 21341
rect 10229 21332 10241 21335
rect 10100 21304 10241 21332
rect 10100 21292 10106 21304
rect 10229 21301 10241 21304
rect 10275 21301 10287 21335
rect 10229 21295 10287 21301
rect 10594 21292 10600 21344
rect 10652 21292 10658 21344
rect 11072 21332 11100 21372
rect 13633 21369 13645 21403
rect 13679 21400 13691 21403
rect 13679 21372 14412 21400
rect 13679 21369 13691 21372
rect 13633 21363 13691 21369
rect 11330 21332 11336 21344
rect 11072 21304 11336 21332
rect 11330 21292 11336 21304
rect 11388 21292 11394 21344
rect 13170 21292 13176 21344
rect 13228 21292 13234 21344
rect 13354 21292 13360 21344
rect 13412 21332 13418 21344
rect 13725 21335 13783 21341
rect 13725 21332 13737 21335
rect 13412 21304 13737 21332
rect 13412 21292 13418 21304
rect 13725 21301 13737 21304
rect 13771 21301 13783 21335
rect 14384 21332 14412 21372
rect 15930 21360 15936 21412
rect 15988 21360 15994 21412
rect 16592 21332 16620 21644
rect 16666 21564 16672 21616
rect 16724 21564 16730 21616
rect 17788 21604 17816 21644
rect 18417 21641 18429 21675
rect 18463 21672 18475 21675
rect 18506 21672 18512 21684
rect 18463 21644 18512 21672
rect 18463 21641 18475 21644
rect 18417 21635 18475 21641
rect 18506 21632 18512 21644
rect 18564 21632 18570 21684
rect 19886 21672 19892 21684
rect 18984 21644 19892 21672
rect 18782 21604 18788 21616
rect 17788 21576 18788 21604
rect 18782 21564 18788 21576
rect 18840 21564 18846 21616
rect 18984 21613 19012 21644
rect 19886 21632 19892 21644
rect 19944 21632 19950 21684
rect 21082 21632 21088 21684
rect 21140 21672 21146 21684
rect 23201 21675 23259 21681
rect 21140 21644 22876 21672
rect 21140 21632 21146 21644
rect 18969 21607 19027 21613
rect 18969 21573 18981 21607
rect 19015 21573 19027 21607
rect 21634 21604 21640 21616
rect 18969 21567 19027 21573
rect 21100 21576 21640 21604
rect 16684 21477 16712 21564
rect 16761 21539 16819 21545
rect 16761 21505 16773 21539
rect 16807 21536 16819 21539
rect 21100 21536 21128 21576
rect 21634 21564 21640 21576
rect 21692 21564 21698 21616
rect 21913 21607 21971 21613
rect 21913 21573 21925 21607
rect 21959 21604 21971 21607
rect 22002 21604 22008 21616
rect 21959 21576 22008 21604
rect 21959 21573 21971 21576
rect 21913 21567 21971 21573
rect 22002 21564 22008 21576
rect 22060 21564 22066 21616
rect 16807 21508 18736 21536
rect 16807 21505 16819 21508
rect 16761 21499 16819 21505
rect 16669 21471 16727 21477
rect 16669 21437 16681 21471
rect 16715 21437 16727 21471
rect 16669 21431 16727 21437
rect 16853 21471 16911 21477
rect 16853 21437 16865 21471
rect 16899 21437 16911 21471
rect 16853 21431 16911 21437
rect 17129 21471 17187 21477
rect 17129 21437 17141 21471
rect 17175 21468 17187 21471
rect 18598 21468 18604 21480
rect 17175 21440 18604 21468
rect 17175 21437 17187 21440
rect 17129 21431 17187 21437
rect 14384 21304 16620 21332
rect 16868 21332 16896 21431
rect 18598 21428 18604 21440
rect 18656 21428 18662 21480
rect 18708 21477 18736 21508
rect 19536 21508 21128 21536
rect 18693 21471 18751 21477
rect 18693 21437 18705 21471
rect 18739 21437 18751 21471
rect 18693 21431 18751 21437
rect 19334 21428 19340 21480
rect 19392 21428 19398 21480
rect 19426 21428 19432 21480
rect 19484 21428 19490 21480
rect 19536 21400 19564 21508
rect 21542 21496 21548 21548
rect 21600 21536 21606 21548
rect 22306 21539 22364 21545
rect 22306 21536 22318 21539
rect 21600 21508 22318 21536
rect 21600 21496 21606 21508
rect 22306 21505 22318 21508
rect 22352 21505 22364 21539
rect 22306 21499 22364 21505
rect 22465 21539 22523 21545
rect 22465 21505 22477 21539
rect 22511 21536 22523 21539
rect 22848 21536 22876 21644
rect 23201 21641 23213 21675
rect 23247 21672 23259 21675
rect 23247 21644 28120 21672
rect 23247 21641 23259 21644
rect 23201 21635 23259 21641
rect 23216 21576 24624 21604
rect 23216 21536 23244 21576
rect 24596 21548 24624 21576
rect 25958 21564 25964 21616
rect 26016 21604 26022 21616
rect 26053 21607 26111 21613
rect 26053 21604 26065 21607
rect 26016 21576 26065 21604
rect 26016 21564 26022 21576
rect 26053 21573 26065 21576
rect 26099 21573 26111 21607
rect 26053 21567 26111 21573
rect 23750 21536 23756 21548
rect 22511 21508 23244 21536
rect 23308 21508 23756 21536
rect 22511 21505 22523 21508
rect 22465 21499 22523 21505
rect 19705 21471 19763 21477
rect 19705 21437 19717 21471
rect 19751 21468 19763 21471
rect 19794 21468 19800 21480
rect 19751 21440 19800 21468
rect 19751 21437 19763 21440
rect 19705 21431 19763 21437
rect 19794 21428 19800 21440
rect 19852 21428 19858 21480
rect 21266 21428 21272 21480
rect 21324 21428 21330 21480
rect 21450 21428 21456 21480
rect 21508 21428 21514 21480
rect 22186 21428 22192 21480
rect 22244 21428 22250 21480
rect 23109 21471 23167 21477
rect 23109 21437 23121 21471
rect 23155 21468 23167 21471
rect 23308 21468 23336 21508
rect 23750 21496 23756 21508
rect 23808 21496 23814 21548
rect 23845 21539 23903 21545
rect 23845 21505 23857 21539
rect 23891 21536 23903 21539
rect 23934 21536 23940 21548
rect 23891 21508 23940 21536
rect 23891 21505 23903 21508
rect 23845 21499 23903 21505
rect 23934 21496 23940 21508
rect 23992 21496 23998 21548
rect 24026 21496 24032 21548
rect 24084 21496 24090 21548
rect 24486 21496 24492 21548
rect 24544 21496 24550 21548
rect 24578 21496 24584 21548
rect 24636 21496 24642 21548
rect 24765 21539 24823 21545
rect 24765 21505 24777 21539
rect 24811 21536 24823 21539
rect 25406 21536 25412 21548
rect 24811 21508 25412 21536
rect 24811 21505 24823 21508
rect 24765 21499 24823 21505
rect 25406 21496 25412 21508
rect 25464 21496 25470 21548
rect 26697 21539 26755 21545
rect 26697 21536 26709 21539
rect 26252 21508 26709 21536
rect 26252 21480 26280 21508
rect 26697 21505 26709 21508
rect 26743 21505 26755 21539
rect 26697 21499 26755 21505
rect 27203 21539 27261 21545
rect 27203 21505 27215 21539
rect 27249 21536 27261 21539
rect 27522 21536 27528 21548
rect 27249 21508 27528 21536
rect 27249 21505 27261 21508
rect 27203 21499 27261 21505
rect 27522 21496 27528 21508
rect 27580 21496 27586 21548
rect 23155 21440 23336 21468
rect 23385 21471 23443 21477
rect 23155 21437 23167 21440
rect 23109 21431 23167 21437
rect 23385 21437 23397 21471
rect 23431 21437 23443 21471
rect 23385 21431 23443 21437
rect 18708 21372 19564 21400
rect 18708 21332 18736 21372
rect 23290 21360 23296 21412
rect 23348 21360 23354 21412
rect 23400 21400 23428 21431
rect 23566 21428 23572 21480
rect 23624 21428 23630 21480
rect 23658 21428 23664 21480
rect 23716 21428 23722 21480
rect 24854 21428 24860 21480
rect 24912 21477 24918 21480
rect 24912 21471 24961 21477
rect 24912 21437 24915 21471
rect 24949 21437 24961 21471
rect 24912 21431 24961 21437
rect 24912 21428 24918 21431
rect 25038 21428 25044 21480
rect 25096 21428 25102 21480
rect 25869 21471 25927 21477
rect 25869 21437 25881 21471
rect 25915 21437 25927 21471
rect 25869 21431 25927 21437
rect 23842 21400 23848 21412
rect 23400 21372 23848 21400
rect 23842 21360 23848 21372
rect 23900 21360 23906 21412
rect 16868 21304 18736 21332
rect 13725 21295 13783 21301
rect 19150 21292 19156 21344
rect 19208 21292 19214 21344
rect 20990 21292 20996 21344
rect 21048 21292 21054 21344
rect 22002 21292 22008 21344
rect 22060 21332 22066 21344
rect 23308 21332 23336 21360
rect 25884 21344 25912 21431
rect 26234 21428 26240 21480
rect 26292 21428 26298 21480
rect 26602 21428 26608 21480
rect 26660 21428 26666 21480
rect 26786 21428 26792 21480
rect 26844 21468 26850 21480
rect 27024 21471 27082 21477
rect 27024 21468 27036 21471
rect 26844 21440 27036 21468
rect 26844 21428 26850 21440
rect 27024 21437 27036 21440
rect 27070 21437 27082 21471
rect 27024 21431 27082 21437
rect 27433 21471 27491 21477
rect 27433 21437 27445 21471
rect 27479 21468 27491 21471
rect 27890 21468 27896 21480
rect 27479 21440 27896 21468
rect 27479 21437 27491 21440
rect 27433 21431 27491 21437
rect 27890 21428 27896 21440
rect 27948 21428 27954 21480
rect 28092 21468 28120 21644
rect 29089 21471 29147 21477
rect 29089 21468 29101 21471
rect 28092 21440 29101 21468
rect 29089 21437 29101 21440
rect 29135 21437 29147 21471
rect 30101 21471 30159 21477
rect 30101 21468 30113 21471
rect 29089 21431 29147 21437
rect 29196 21440 30113 21468
rect 26142 21360 26148 21412
rect 26200 21400 26206 21412
rect 29196 21400 29224 21440
rect 30101 21437 30113 21440
rect 30147 21437 30159 21471
rect 30101 21431 30159 21437
rect 26200 21372 26556 21400
rect 26200 21360 26206 21372
rect 22060 21304 23336 21332
rect 22060 21292 22066 21304
rect 24026 21292 24032 21344
rect 24084 21332 24090 21344
rect 25314 21332 25320 21344
rect 24084 21304 25320 21332
rect 24084 21292 24090 21304
rect 25314 21292 25320 21304
rect 25372 21292 25378 21344
rect 25682 21292 25688 21344
rect 25740 21292 25746 21344
rect 25866 21292 25872 21344
rect 25924 21292 25930 21344
rect 26418 21292 26424 21344
rect 26476 21292 26482 21344
rect 26528 21332 26556 21372
rect 28092 21372 29224 21400
rect 29457 21403 29515 21409
rect 28092 21332 28120 21372
rect 29457 21369 29469 21403
rect 29503 21400 29515 21403
rect 29641 21403 29699 21409
rect 29641 21400 29653 21403
rect 29503 21372 29653 21400
rect 29503 21369 29515 21372
rect 29457 21363 29515 21369
rect 29641 21369 29653 21372
rect 29687 21400 29699 21403
rect 29687 21372 31340 21400
rect 29687 21369 29699 21372
rect 29641 21363 29699 21369
rect 31312 21344 31340 21372
rect 26528 21304 28120 21332
rect 28534 21292 28540 21344
rect 28592 21292 28598 21344
rect 29917 21335 29975 21341
rect 29917 21301 29929 21335
rect 29963 21332 29975 21335
rect 30006 21332 30012 21344
rect 29963 21304 30012 21332
rect 29963 21301 29975 21304
rect 29917 21295 29975 21301
rect 30006 21292 30012 21304
rect 30064 21292 30070 21344
rect 30282 21292 30288 21344
rect 30340 21292 30346 21344
rect 31294 21292 31300 21344
rect 31352 21292 31358 21344
rect 552 21242 31072 21264
rect 552 21190 7988 21242
rect 8040 21190 8052 21242
rect 8104 21190 8116 21242
rect 8168 21190 8180 21242
rect 8232 21190 8244 21242
rect 8296 21190 15578 21242
rect 15630 21190 15642 21242
rect 15694 21190 15706 21242
rect 15758 21190 15770 21242
rect 15822 21190 15834 21242
rect 15886 21190 23168 21242
rect 23220 21190 23232 21242
rect 23284 21190 23296 21242
rect 23348 21190 23360 21242
rect 23412 21190 23424 21242
rect 23476 21190 30758 21242
rect 30810 21190 30822 21242
rect 30874 21190 30886 21242
rect 30938 21190 30950 21242
rect 31002 21190 31014 21242
rect 31066 21190 31072 21242
rect 552 21168 31072 21190
rect 7926 21128 7932 21140
rect 1596 21100 7932 21128
rect 1596 21069 1624 21100
rect 7926 21088 7932 21100
rect 7984 21088 7990 21140
rect 8570 21128 8576 21140
rect 8128 21100 8576 21128
rect 1581 21063 1639 21069
rect 1581 21029 1593 21063
rect 1627 21029 1639 21063
rect 1581 21023 1639 21029
rect 1946 21020 1952 21072
rect 2004 21020 2010 21072
rect 2130 21020 2136 21072
rect 2188 21020 2194 21072
rect 5258 21020 5264 21072
rect 5316 21020 5322 21072
rect 5810 21020 5816 21072
rect 5868 21060 5874 21072
rect 5868 21032 6224 21060
rect 5868 21020 5874 21032
rect 937 20995 995 21001
rect 937 20961 949 20995
rect 983 20992 995 20995
rect 1118 20992 1124 21004
rect 983 20964 1124 20992
rect 983 20961 995 20964
rect 937 20955 995 20961
rect 1118 20952 1124 20964
rect 1176 20952 1182 21004
rect 1213 20995 1271 21001
rect 1213 20961 1225 20995
rect 1259 20992 1271 20995
rect 1394 20992 1400 21004
rect 1259 20964 1400 20992
rect 1259 20961 1271 20964
rect 1213 20955 1271 20961
rect 1394 20952 1400 20964
rect 1452 20992 1458 21004
rect 2958 21001 2964 21004
rect 2920 20995 2964 21001
rect 2920 20992 2932 20995
rect 1452 20964 2932 20992
rect 1452 20952 1458 20964
rect 2920 20961 2932 20964
rect 2920 20955 2964 20961
rect 2958 20952 2964 20955
rect 3016 20952 3022 21004
rect 3786 20952 3792 21004
rect 3844 20952 3850 21004
rect 4801 20995 4859 21001
rect 4801 20961 4813 20995
rect 4847 20992 4859 20995
rect 4982 20992 4988 21004
rect 4847 20964 4988 20992
rect 4847 20961 4859 20964
rect 4801 20955 4859 20961
rect 4982 20952 4988 20964
rect 5040 20952 5046 21004
rect 5994 20952 6000 21004
rect 6052 20952 6058 21004
rect 6086 20952 6092 21004
rect 6144 20952 6150 21004
rect 6196 21001 6224 21032
rect 7190 21020 7196 21072
rect 7248 21060 7254 21072
rect 8128 21060 8156 21100
rect 8570 21088 8576 21100
rect 8628 21088 8634 21140
rect 8754 21088 8760 21140
rect 8812 21128 8818 21140
rect 10137 21131 10195 21137
rect 10137 21128 10149 21131
rect 8812 21100 10149 21128
rect 8812 21088 8818 21100
rect 10137 21097 10149 21100
rect 10183 21097 10195 21131
rect 10137 21091 10195 21097
rect 10594 21088 10600 21140
rect 10652 21128 10658 21140
rect 11514 21128 11520 21140
rect 10652 21100 11520 21128
rect 10652 21088 10658 21100
rect 11514 21088 11520 21100
rect 11572 21088 11578 21140
rect 11707 21131 11765 21137
rect 11707 21097 11719 21131
rect 11753 21128 11765 21131
rect 12342 21128 12348 21140
rect 11753 21100 12348 21128
rect 11753 21097 11765 21100
rect 11707 21091 11765 21097
rect 12342 21088 12348 21100
rect 12400 21088 12406 21140
rect 12434 21088 12440 21140
rect 12492 21128 12498 21140
rect 13633 21131 13691 21137
rect 13633 21128 13645 21131
rect 12492 21100 13645 21128
rect 12492 21088 12498 21100
rect 13633 21097 13645 21100
rect 13679 21097 13691 21131
rect 13633 21091 13691 21097
rect 15194 21088 15200 21140
rect 15252 21128 15258 21140
rect 15933 21131 15991 21137
rect 15933 21128 15945 21131
rect 15252 21100 15945 21128
rect 15252 21088 15258 21100
rect 15933 21097 15945 21100
rect 15979 21097 15991 21131
rect 15933 21091 15991 21097
rect 17954 21088 17960 21140
rect 18012 21128 18018 21140
rect 18785 21131 18843 21137
rect 18785 21128 18797 21131
rect 18012 21100 18797 21128
rect 18012 21088 18018 21100
rect 18785 21097 18797 21100
rect 18831 21097 18843 21131
rect 18785 21091 18843 21097
rect 19426 21088 19432 21140
rect 19484 21128 19490 21140
rect 19978 21128 19984 21140
rect 19484 21100 19984 21128
rect 19484 21088 19490 21100
rect 19978 21088 19984 21100
rect 20036 21088 20042 21140
rect 20809 21131 20867 21137
rect 20809 21097 20821 21131
rect 20855 21128 20867 21131
rect 21266 21128 21272 21140
rect 20855 21100 21272 21128
rect 20855 21097 20867 21100
rect 20809 21091 20867 21097
rect 21266 21088 21272 21100
rect 21324 21088 21330 21140
rect 22186 21088 22192 21140
rect 22244 21128 22250 21140
rect 23109 21131 23167 21137
rect 23109 21128 23121 21131
rect 22244 21100 23121 21128
rect 22244 21088 22250 21100
rect 23109 21097 23121 21100
rect 23155 21097 23167 21131
rect 23109 21091 23167 21097
rect 23216 21100 25084 21128
rect 10962 21060 10968 21072
rect 7248 21032 8156 21060
rect 7248 21020 7254 21032
rect 6181 20995 6239 21001
rect 6181 20961 6193 20995
rect 6227 20961 6239 20995
rect 6181 20955 6239 20961
rect 6462 20996 6520 21001
rect 6462 20995 6592 20996
rect 6462 20961 6474 20995
rect 6508 20992 6592 20995
rect 8018 20992 8024 21004
rect 6508 20968 8024 20992
rect 6508 20961 6520 20968
rect 6564 20964 8024 20968
rect 6462 20955 6520 20961
rect 8018 20952 8024 20964
rect 8076 20952 8082 21004
rect 8128 21001 8156 21032
rect 9692 21032 10968 21060
rect 9692 21004 9720 21032
rect 10962 21020 10968 21032
rect 11020 21020 11026 21072
rect 11054 21020 11060 21072
rect 11112 21060 11118 21072
rect 11112 21032 11284 21060
rect 11112 21020 11118 21032
rect 8113 20995 8171 21001
rect 8113 20961 8125 20995
rect 8159 20961 8171 20995
rect 8113 20955 8171 20961
rect 8220 20964 8803 20992
rect 3089 20945 3147 20951
rect 3089 20936 3101 20945
rect 2593 20927 2651 20933
rect 2593 20893 2605 20927
rect 2639 20924 2651 20927
rect 2774 20924 2780 20936
rect 2639 20896 2780 20924
rect 2639 20893 2651 20896
rect 2593 20887 2651 20893
rect 2774 20884 2780 20896
rect 2832 20884 2838 20936
rect 3050 20884 3056 20936
rect 3135 20911 3147 20945
rect 3108 20905 3147 20911
rect 3329 20927 3387 20933
rect 3108 20896 3132 20905
rect 3108 20884 3114 20896
rect 3329 20893 3341 20927
rect 3375 20924 3387 20927
rect 3694 20924 3700 20936
rect 3375 20896 3700 20924
rect 3375 20893 3387 20896
rect 3329 20887 3387 20893
rect 3694 20884 3700 20896
rect 3752 20884 3758 20936
rect 3804 20924 3832 20952
rect 5537 20927 5595 20933
rect 3804 20896 4022 20924
rect 3994 20856 4022 20896
rect 5537 20893 5549 20927
rect 5583 20924 5595 20927
rect 6104 20924 6132 20952
rect 5583 20896 6132 20924
rect 5583 20893 5595 20896
rect 5537 20887 5595 20893
rect 7650 20884 7656 20936
rect 7708 20924 7714 20936
rect 8220 20924 8248 20964
rect 7708 20896 8248 20924
rect 7708 20884 7714 20896
rect 8294 20884 8300 20936
rect 8352 20884 8358 20936
rect 8662 20933 8668 20936
rect 8624 20927 8668 20933
rect 8624 20893 8636 20927
rect 8624 20887 8668 20893
rect 8662 20884 8668 20887
rect 8720 20884 8726 20936
rect 8775 20933 8803 20964
rect 9674 20952 9680 21004
rect 9732 20952 9738 21004
rect 10689 20995 10747 21001
rect 10689 20992 10701 20995
rect 10428 20964 10701 20992
rect 8760 20927 8818 20933
rect 8760 20893 8772 20927
rect 8806 20893 8818 20927
rect 8760 20887 8818 20893
rect 8846 20884 8852 20936
rect 8904 20924 8910 20936
rect 9033 20927 9091 20933
rect 9033 20924 9045 20927
rect 8904 20896 9045 20924
rect 8904 20884 8910 20896
rect 9033 20893 9045 20896
rect 9079 20893 9091 20927
rect 9033 20887 9091 20893
rect 10428 20856 10456 20964
rect 10689 20961 10701 20964
rect 10735 20961 10747 20995
rect 10689 20955 10747 20961
rect 10778 20952 10784 21004
rect 10836 20992 10842 21004
rect 11256 21001 11284 21032
rect 14642 21020 14648 21072
rect 14700 21060 14706 21072
rect 19242 21060 19248 21072
rect 14700 21032 16160 21060
rect 14700 21020 14706 21032
rect 11149 20995 11207 21001
rect 11149 20992 11161 20995
rect 10836 20964 11161 20992
rect 10836 20952 10842 20964
rect 11149 20961 11161 20964
rect 11195 20961 11207 20995
rect 11149 20955 11207 20961
rect 11241 20995 11299 21001
rect 11241 20961 11253 20995
rect 11287 20961 11299 20995
rect 11241 20955 11299 20961
rect 11514 20952 11520 21004
rect 11572 20992 11578 21004
rect 11977 20995 12035 21001
rect 11977 20992 11989 20995
rect 11572 20964 11989 20992
rect 11572 20952 11578 20964
rect 11977 20961 11989 20964
rect 12023 20961 12035 20995
rect 11977 20955 12035 20961
rect 12084 20964 13492 20992
rect 10502 20884 10508 20936
rect 10560 20924 10566 20936
rect 11704 20927 11762 20933
rect 11704 20924 11716 20927
rect 10560 20896 11716 20924
rect 10560 20884 10566 20896
rect 11704 20893 11716 20896
rect 11750 20893 11762 20927
rect 11704 20887 11762 20893
rect 11790 20884 11796 20936
rect 11848 20924 11854 20936
rect 12084 20924 12112 20964
rect 11848 20896 12112 20924
rect 11848 20884 11854 20896
rect 11238 20856 11244 20868
rect 3994 20828 6224 20856
rect 2409 20791 2467 20797
rect 2409 20757 2421 20791
rect 2455 20788 2467 20791
rect 4062 20788 4068 20800
rect 2455 20760 4068 20788
rect 2455 20757 2467 20760
rect 2409 20751 2467 20757
rect 4062 20748 4068 20760
rect 4120 20748 4126 20800
rect 4433 20791 4491 20797
rect 4433 20757 4445 20791
rect 4479 20788 4491 20791
rect 4522 20788 4528 20800
rect 4479 20760 4528 20788
rect 4479 20757 4491 20760
rect 4433 20751 4491 20757
rect 4522 20748 4528 20760
rect 4580 20748 4586 20800
rect 4985 20791 5043 20797
rect 4985 20757 4997 20791
rect 5031 20788 5043 20791
rect 5258 20788 5264 20800
rect 5031 20760 5264 20788
rect 5031 20757 5043 20760
rect 4985 20751 5043 20757
rect 5258 20748 5264 20760
rect 5316 20748 5322 20800
rect 5810 20748 5816 20800
rect 5868 20748 5874 20800
rect 6196 20788 6224 20828
rect 7116 20828 8064 20856
rect 10428 20828 11244 20856
rect 7116 20788 7144 20828
rect 6196 20760 7144 20788
rect 7466 20748 7472 20800
rect 7524 20788 7530 20800
rect 7561 20791 7619 20797
rect 7561 20788 7573 20791
rect 7524 20760 7573 20788
rect 7524 20748 7530 20760
rect 7561 20757 7573 20760
rect 7607 20757 7619 20791
rect 7561 20751 7619 20757
rect 7742 20748 7748 20800
rect 7800 20788 7806 20800
rect 7929 20791 7987 20797
rect 7929 20788 7941 20791
rect 7800 20760 7941 20788
rect 7800 20748 7806 20760
rect 7929 20757 7941 20760
rect 7975 20757 7987 20791
rect 8036 20788 8064 20828
rect 11238 20816 11244 20828
rect 11296 20816 11302 20868
rect 10505 20791 10563 20797
rect 10505 20788 10517 20791
rect 8036 20760 10517 20788
rect 7929 20751 7987 20757
rect 10505 20757 10517 20760
rect 10551 20757 10563 20791
rect 10505 20751 10563 20757
rect 10962 20748 10968 20800
rect 11020 20748 11026 20800
rect 11146 20748 11152 20800
rect 11204 20788 11210 20800
rect 13081 20791 13139 20797
rect 13081 20788 13093 20791
rect 11204 20760 13093 20788
rect 11204 20748 11210 20760
rect 13081 20757 13093 20760
rect 13127 20757 13139 20791
rect 13464 20788 13492 20964
rect 13538 20952 13544 21004
rect 13596 20952 13602 21004
rect 14093 20995 14151 21001
rect 14093 20961 14105 20995
rect 14139 20992 14151 20995
rect 14274 20992 14280 21004
rect 14139 20964 14280 20992
rect 14139 20961 14151 20964
rect 14093 20955 14151 20961
rect 14274 20952 14280 20964
rect 14332 20952 14338 21004
rect 14369 20995 14427 21001
rect 14369 20961 14381 20995
rect 14415 20992 14427 20995
rect 14826 20992 14832 21004
rect 14415 20964 14832 20992
rect 14415 20961 14427 20964
rect 14369 20955 14427 20961
rect 14826 20952 14832 20964
rect 14884 20952 14890 21004
rect 16132 21001 16160 21032
rect 18708 21032 19248 21060
rect 16117 20995 16175 21001
rect 16117 20961 16129 20995
rect 16163 20961 16175 20995
rect 17957 20995 18015 21001
rect 17957 20992 17969 20995
rect 16117 20955 16175 20961
rect 16316 20964 17969 20992
rect 16316 20924 16344 20964
rect 17957 20961 17969 20964
rect 18003 20961 18015 20995
rect 17957 20955 18015 20961
rect 18138 20952 18144 21004
rect 18196 20992 18202 21004
rect 18414 20992 18420 21004
rect 18196 20964 18420 20992
rect 18196 20952 18202 20964
rect 18414 20952 18420 20964
rect 18472 20952 18478 21004
rect 18708 21001 18736 21032
rect 19242 21020 19248 21032
rect 19300 21020 19306 21072
rect 22830 21020 22836 21072
rect 22888 21060 22894 21072
rect 23216 21060 23244 21100
rect 22888 21032 23244 21060
rect 25056 21060 25084 21100
rect 25314 21088 25320 21140
rect 25372 21088 25378 21140
rect 30282 21128 30288 21140
rect 25700 21100 30288 21128
rect 25700 21060 25728 21100
rect 30282 21088 30288 21100
rect 30340 21088 30346 21140
rect 30466 21088 30472 21140
rect 30524 21088 30530 21140
rect 25056 21032 25728 21060
rect 22888 21020 22894 21032
rect 18693 20995 18751 21001
rect 18693 20961 18705 20995
rect 18739 20961 18751 20995
rect 20714 20992 20720 21004
rect 20378 20964 20720 20992
rect 18693 20955 18751 20961
rect 16132 20896 16344 20924
rect 15657 20859 15715 20865
rect 15657 20825 15669 20859
rect 15703 20856 15715 20859
rect 16132 20856 16160 20896
rect 16390 20884 16396 20936
rect 16448 20924 16454 20936
rect 18708 20924 18736 20955
rect 20714 20952 20720 20964
rect 20772 20952 20778 21004
rect 20993 20995 21051 21001
rect 20993 20961 21005 20995
rect 21039 20961 21051 20995
rect 23106 20992 23112 21004
rect 22678 20964 23112 20992
rect 20993 20955 21051 20961
rect 16448 20896 18736 20924
rect 18969 20927 19027 20933
rect 16448 20884 16454 20896
rect 18969 20893 18981 20927
rect 19015 20893 19027 20927
rect 18969 20887 19027 20893
rect 19245 20927 19303 20933
rect 19245 20893 19257 20927
rect 19291 20924 19303 20927
rect 19702 20924 19708 20936
rect 19291 20896 19708 20924
rect 19291 20893 19303 20896
rect 19245 20887 19303 20893
rect 15703 20828 16160 20856
rect 15703 20825 15715 20828
rect 15657 20819 15715 20825
rect 15102 20788 15108 20800
rect 13464 20760 15108 20788
rect 13081 20751 13139 20757
rect 15102 20748 15108 20760
rect 15160 20748 15166 20800
rect 15286 20748 15292 20800
rect 15344 20788 15350 20800
rect 15672 20788 15700 20819
rect 15344 20760 15700 20788
rect 15344 20748 15350 20760
rect 16482 20748 16488 20800
rect 16540 20788 16546 20800
rect 17497 20791 17555 20797
rect 17497 20788 17509 20791
rect 16540 20760 17509 20788
rect 16540 20748 16546 20760
rect 17497 20757 17509 20760
rect 17543 20757 17555 20791
rect 18984 20788 19012 20887
rect 19702 20884 19708 20896
rect 19760 20924 19766 20936
rect 21008 20924 21036 20955
rect 23106 20952 23112 20964
rect 23164 20952 23170 21004
rect 23293 20995 23351 21001
rect 23293 20961 23305 20995
rect 23339 20961 23351 20995
rect 25130 20992 25136 21004
rect 24886 20964 25136 20992
rect 23293 20955 23351 20961
rect 19760 20896 21036 20924
rect 19760 20884 19766 20896
rect 21266 20884 21272 20936
rect 21324 20884 21330 20936
rect 21545 20927 21603 20933
rect 21545 20893 21557 20927
rect 21591 20924 21603 20927
rect 23308 20924 23336 20955
rect 25130 20952 25136 20964
rect 25188 20952 25194 21004
rect 25700 21001 25728 21032
rect 28074 21020 28080 21072
rect 28132 21020 28138 21072
rect 28534 21060 28540 21072
rect 28184 21032 28540 21060
rect 25501 20995 25559 21001
rect 25501 20961 25513 20995
rect 25547 20961 25559 20995
rect 25501 20955 25559 20961
rect 25685 20995 25743 21001
rect 25685 20961 25697 20995
rect 25731 20961 25743 20995
rect 28184 20992 28212 21032
rect 28534 21020 28540 21032
rect 28592 21020 28598 21072
rect 25685 20955 25743 20961
rect 25792 20964 28212 20992
rect 23477 20927 23535 20933
rect 23477 20924 23489 20927
rect 21591 20896 23489 20924
rect 21591 20893 21603 20896
rect 21545 20887 21603 20893
rect 23477 20893 23489 20896
rect 23523 20893 23535 20927
rect 23753 20927 23811 20933
rect 23753 20924 23765 20927
rect 23477 20887 23535 20893
rect 23584 20896 23765 20924
rect 20530 20788 20536 20800
rect 18984 20760 20536 20788
rect 17497 20751 17555 20757
rect 20530 20748 20536 20760
rect 20588 20748 20594 20800
rect 20990 20748 20996 20800
rect 21048 20788 21054 20800
rect 21910 20788 21916 20800
rect 21048 20760 21916 20788
rect 21048 20748 21054 20760
rect 21910 20748 21916 20760
rect 21968 20748 21974 20800
rect 22186 20748 22192 20800
rect 22244 20788 22250 20800
rect 23584 20788 23612 20896
rect 23753 20893 23765 20896
rect 23799 20924 23811 20927
rect 25516 20924 25544 20955
rect 25792 20924 25820 20964
rect 28350 20952 28356 21004
rect 28408 20952 28414 21004
rect 23799 20896 25544 20924
rect 25608 20896 25820 20924
rect 25961 20927 26019 20933
rect 23799 20893 23811 20896
rect 23753 20887 23811 20893
rect 24762 20816 24768 20868
rect 24820 20856 24826 20868
rect 25608 20856 25636 20896
rect 25961 20893 25973 20927
rect 26007 20924 26019 20927
rect 26050 20924 26056 20936
rect 26007 20896 26056 20924
rect 26007 20893 26019 20896
rect 25961 20887 26019 20893
rect 26050 20884 26056 20896
rect 26108 20884 26114 20936
rect 26326 20884 26332 20936
rect 26384 20924 26390 20936
rect 26421 20927 26479 20933
rect 26421 20924 26433 20927
rect 26384 20896 26433 20924
rect 26384 20884 26390 20896
rect 26421 20893 26433 20896
rect 26467 20893 26479 20927
rect 26421 20887 26479 20893
rect 26697 20927 26755 20933
rect 26697 20893 26709 20927
rect 26743 20924 26755 20927
rect 28258 20924 28264 20936
rect 26743 20896 28264 20924
rect 26743 20893 26755 20896
rect 26697 20887 26755 20893
rect 28258 20884 28264 20896
rect 28316 20884 28322 20936
rect 28442 20884 28448 20936
rect 28500 20884 28506 20936
rect 28810 20933 28816 20936
rect 28772 20927 28816 20933
rect 28772 20893 28784 20927
rect 28772 20887 28816 20893
rect 28810 20884 28816 20887
rect 28868 20884 28874 20936
rect 28994 20933 29000 20936
rect 28951 20927 29000 20933
rect 28951 20893 28963 20927
rect 28997 20893 29000 20927
rect 28951 20887 29000 20893
rect 28994 20884 29000 20887
rect 29052 20884 29058 20936
rect 29181 20927 29239 20933
rect 29181 20893 29193 20927
rect 29227 20924 29239 20927
rect 29546 20924 29552 20936
rect 29227 20896 29552 20924
rect 29227 20893 29239 20896
rect 29181 20887 29239 20893
rect 29546 20884 29552 20896
rect 29604 20884 29610 20936
rect 24820 20828 25636 20856
rect 24820 20816 24826 20828
rect 25682 20816 25688 20868
rect 25740 20816 25746 20868
rect 28166 20816 28172 20868
rect 28224 20816 28230 20868
rect 22244 20760 23612 20788
rect 22244 20748 22250 20760
rect 24302 20748 24308 20800
rect 24360 20788 24366 20800
rect 25700 20788 25728 20816
rect 24360 20760 25728 20788
rect 24360 20748 24366 20760
rect 25866 20748 25872 20800
rect 25924 20788 25930 20800
rect 29638 20788 29644 20800
rect 25924 20760 29644 20788
rect 25924 20748 25930 20760
rect 29638 20748 29644 20760
rect 29696 20748 29702 20800
rect 552 20698 30912 20720
rect 552 20646 4193 20698
rect 4245 20646 4257 20698
rect 4309 20646 4321 20698
rect 4373 20646 4385 20698
rect 4437 20646 4449 20698
rect 4501 20646 11783 20698
rect 11835 20646 11847 20698
rect 11899 20646 11911 20698
rect 11963 20646 11975 20698
rect 12027 20646 12039 20698
rect 12091 20646 19373 20698
rect 19425 20646 19437 20698
rect 19489 20646 19501 20698
rect 19553 20646 19565 20698
rect 19617 20646 19629 20698
rect 19681 20646 26963 20698
rect 27015 20646 27027 20698
rect 27079 20646 27091 20698
rect 27143 20646 27155 20698
rect 27207 20646 27219 20698
rect 27271 20646 30912 20698
rect 552 20624 30912 20646
rect 3697 20587 3755 20593
rect 3697 20553 3709 20587
rect 3743 20584 3755 20587
rect 5905 20587 5963 20593
rect 3743 20556 5764 20584
rect 3743 20553 3755 20556
rect 3697 20547 3755 20553
rect 1351 20451 1409 20457
rect 1351 20417 1363 20451
rect 1397 20448 1409 20451
rect 2774 20448 2780 20460
rect 1397 20420 2780 20448
rect 1397 20417 1409 20420
rect 1351 20411 1409 20417
rect 2774 20408 2780 20420
rect 2832 20408 2838 20460
rect 4387 20451 4445 20457
rect 4387 20417 4399 20451
rect 4433 20448 4445 20451
rect 4522 20448 4528 20460
rect 4433 20420 4528 20448
rect 4433 20417 4445 20420
rect 4387 20411 4445 20417
rect 4522 20408 4528 20420
rect 4580 20408 4586 20460
rect 4614 20408 4620 20460
rect 4672 20408 4678 20460
rect 5736 20448 5764 20556
rect 5905 20553 5917 20587
rect 5951 20584 5963 20587
rect 7282 20584 7288 20596
rect 5951 20556 7288 20584
rect 5951 20553 5963 20556
rect 5905 20547 5963 20553
rect 7282 20544 7288 20556
rect 7340 20544 7346 20596
rect 7926 20544 7932 20596
rect 7984 20544 7990 20596
rect 10318 20584 10324 20596
rect 8036 20556 10324 20584
rect 6638 20455 6644 20460
rect 6595 20449 6644 20455
rect 5736 20420 6500 20448
rect 845 20383 903 20389
rect 845 20349 857 20383
rect 891 20380 903 20383
rect 1210 20380 1216 20392
rect 891 20352 1216 20380
rect 891 20349 903 20352
rect 845 20343 903 20349
rect 1210 20340 1216 20352
rect 1268 20340 1274 20392
rect 1578 20340 1584 20392
rect 1636 20340 1642 20392
rect 3881 20383 3939 20389
rect 3881 20349 3893 20383
rect 3927 20380 3939 20383
rect 4706 20380 4712 20392
rect 3927 20352 4712 20380
rect 3927 20349 3939 20352
rect 3881 20343 3939 20349
rect 4706 20340 4712 20352
rect 4764 20340 4770 20392
rect 6089 20383 6147 20389
rect 6089 20349 6101 20383
rect 6135 20380 6147 20383
rect 6178 20380 6184 20392
rect 6135 20352 6184 20380
rect 6135 20349 6147 20352
rect 6089 20343 6147 20349
rect 6178 20340 6184 20352
rect 6236 20340 6242 20392
rect 6472 20380 6500 20420
rect 6595 20415 6607 20449
rect 6641 20415 6644 20449
rect 6595 20409 6644 20415
rect 6638 20408 6644 20409
rect 6696 20408 6702 20460
rect 6822 20408 6828 20460
rect 6880 20408 6886 20460
rect 8036 20380 8064 20556
rect 10318 20544 10324 20556
rect 10376 20544 10382 20596
rect 10502 20544 10508 20596
rect 10560 20544 10566 20596
rect 10612 20556 12480 20584
rect 8846 20448 8852 20460
rect 8496 20420 8852 20448
rect 8496 20389 8524 20420
rect 8846 20408 8852 20420
rect 8904 20408 8910 20460
rect 8987 20451 9045 20457
rect 8987 20417 8999 20451
rect 9033 20448 9045 20451
rect 10226 20448 10232 20460
rect 9033 20420 10232 20448
rect 9033 20417 9045 20420
rect 8987 20411 9045 20417
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 6472 20352 8064 20380
rect 8481 20383 8539 20389
rect 8481 20349 8493 20383
rect 8527 20349 8539 20383
rect 9122 20380 9128 20392
rect 8481 20343 8539 20349
rect 8588 20352 9128 20380
rect 3421 20315 3479 20321
rect 3421 20281 3433 20315
rect 3467 20312 3479 20315
rect 3467 20284 4022 20312
rect 3467 20281 3479 20284
rect 3421 20275 3479 20281
rect 1302 20204 1308 20256
rect 1360 20253 1366 20256
rect 1360 20207 1369 20253
rect 2869 20247 2927 20253
rect 2869 20213 2881 20247
rect 2915 20244 2927 20247
rect 3602 20244 3608 20256
rect 2915 20216 3608 20244
rect 2915 20213 2927 20216
rect 2869 20207 2927 20213
rect 1360 20204 1366 20207
rect 3602 20204 3608 20216
rect 3660 20204 3666 20256
rect 3994 20244 4022 20284
rect 8386 20272 8392 20324
rect 8444 20312 8450 20324
rect 8588 20312 8616 20352
rect 9122 20340 9128 20352
rect 9180 20340 9186 20392
rect 9217 20383 9275 20389
rect 9217 20349 9229 20383
rect 9263 20380 9275 20383
rect 10612 20380 10640 20556
rect 12452 20516 12480 20556
rect 12526 20544 12532 20596
rect 12584 20584 12590 20596
rect 13081 20587 13139 20593
rect 13081 20584 13093 20587
rect 12584 20556 13093 20584
rect 12584 20544 12590 20556
rect 13081 20553 13093 20556
rect 13127 20553 13139 20587
rect 13081 20547 13139 20553
rect 13170 20544 13176 20596
rect 13228 20544 13234 20596
rect 16025 20587 16083 20593
rect 16025 20584 16037 20587
rect 13832 20556 16037 20584
rect 13188 20516 13216 20544
rect 13832 20528 13860 20556
rect 16025 20553 16037 20556
rect 16071 20553 16083 20587
rect 19061 20587 19119 20593
rect 16025 20547 16083 20553
rect 16132 20556 17080 20584
rect 12452 20488 13216 20516
rect 13814 20476 13820 20528
rect 13872 20476 13878 20528
rect 14274 20516 14280 20528
rect 13924 20488 14280 20516
rect 10962 20408 10968 20460
rect 11020 20408 11026 20460
rect 11054 20408 11060 20460
rect 11112 20448 11118 20460
rect 11152 20451 11210 20457
rect 11152 20448 11164 20451
rect 11112 20420 11164 20448
rect 11112 20408 11118 20420
rect 11152 20417 11164 20420
rect 11198 20417 11210 20451
rect 13924 20448 13952 20488
rect 14274 20476 14280 20488
rect 14332 20476 14338 20528
rect 16132 20516 16160 20556
rect 15580 20488 16160 20516
rect 17052 20516 17080 20556
rect 19061 20553 19073 20587
rect 19107 20584 19119 20587
rect 19242 20584 19248 20596
rect 19107 20556 19248 20584
rect 19107 20553 19119 20556
rect 19061 20547 19119 20553
rect 19242 20544 19248 20556
rect 19300 20544 19306 20596
rect 19444 20556 22876 20584
rect 19444 20516 19472 20556
rect 17052 20488 19472 20516
rect 22848 20516 22876 20556
rect 23014 20544 23020 20596
rect 23072 20584 23078 20596
rect 28537 20587 28595 20593
rect 28537 20584 28549 20587
rect 23072 20556 28549 20584
rect 23072 20544 23078 20556
rect 28537 20553 28549 20556
rect 28583 20553 28595 20587
rect 28537 20547 28595 20553
rect 23566 20516 23572 20528
rect 22848 20488 23572 20516
rect 11152 20411 11210 20417
rect 11716 20420 13952 20448
rect 14093 20451 14151 20457
rect 9263 20352 10640 20380
rect 10689 20383 10747 20389
rect 9263 20349 9275 20352
rect 9217 20343 9275 20349
rect 10689 20349 10701 20383
rect 10735 20349 10747 20383
rect 10980 20380 11008 20408
rect 11716 20392 11744 20420
rect 14093 20417 14105 20451
rect 14139 20448 14151 20451
rect 14642 20448 14648 20460
rect 14139 20420 14648 20448
rect 14139 20417 14151 20420
rect 14093 20411 14151 20417
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 15194 20408 15200 20460
rect 15252 20448 15258 20460
rect 15580 20448 15608 20488
rect 23566 20476 23572 20488
rect 23624 20476 23630 20528
rect 25314 20476 25320 20528
rect 25372 20516 25378 20528
rect 26326 20516 26332 20528
rect 25372 20488 26332 20516
rect 25372 20476 25378 20488
rect 26326 20476 26332 20488
rect 26384 20476 26390 20528
rect 15252 20420 15608 20448
rect 15252 20408 15258 20420
rect 15930 20408 15936 20460
rect 15988 20448 15994 20460
rect 16393 20451 16451 20457
rect 16393 20448 16405 20451
rect 15988 20420 16405 20448
rect 15988 20408 15994 20420
rect 16393 20417 16405 20420
rect 16439 20417 16451 20451
rect 16393 20411 16451 20417
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20448 18751 20451
rect 18782 20448 18788 20460
rect 18739 20420 18788 20448
rect 18739 20417 18751 20420
rect 18693 20411 18751 20417
rect 18782 20408 18788 20420
rect 18840 20408 18846 20460
rect 19337 20451 19395 20457
rect 19337 20417 19349 20451
rect 19383 20448 19395 20451
rect 19702 20448 19708 20460
rect 19383 20420 19708 20448
rect 19383 20417 19395 20420
rect 19337 20411 19395 20417
rect 19702 20408 19708 20420
rect 19760 20408 19766 20460
rect 21821 20451 21879 20457
rect 21821 20417 21833 20451
rect 21867 20448 21879 20451
rect 24121 20451 24179 20457
rect 21867 20420 23612 20448
rect 21867 20417 21879 20420
rect 21821 20411 21879 20417
rect 11425 20383 11483 20389
rect 11425 20380 11437 20383
rect 10980 20352 11437 20380
rect 10689 20343 10747 20349
rect 11425 20349 11437 20352
rect 11471 20349 11483 20383
rect 11425 20343 11483 20349
rect 10704 20312 10732 20343
rect 11698 20340 11704 20392
rect 11756 20340 11762 20392
rect 12084 20352 14228 20380
rect 8444 20284 8616 20312
rect 10612 20284 10732 20312
rect 8444 20272 8450 20284
rect 10612 20256 10640 20284
rect 4246 20244 4252 20256
rect 3994 20216 4252 20244
rect 4246 20204 4252 20216
rect 4304 20204 4310 20256
rect 4347 20247 4405 20253
rect 4347 20213 4359 20247
rect 4393 20244 4405 20247
rect 6178 20244 6184 20256
rect 4393 20216 6184 20244
rect 4393 20213 4405 20216
rect 4347 20207 4405 20213
rect 6178 20204 6184 20216
rect 6236 20204 6242 20256
rect 6555 20247 6613 20253
rect 6555 20213 6567 20247
rect 6601 20244 6613 20247
rect 7558 20244 7564 20256
rect 6601 20216 7564 20244
rect 6601 20213 6613 20216
rect 6555 20207 6613 20213
rect 7558 20204 7564 20216
rect 7616 20204 7622 20256
rect 8947 20247 9005 20253
rect 8947 20213 8959 20247
rect 8993 20244 9005 20247
rect 9306 20244 9312 20256
rect 8993 20216 9312 20244
rect 8993 20213 9005 20216
rect 8947 20207 9005 20213
rect 9306 20204 9312 20216
rect 9364 20204 9370 20256
rect 10594 20204 10600 20256
rect 10652 20204 10658 20256
rect 11155 20247 11213 20253
rect 11155 20213 11167 20247
rect 11201 20244 11213 20247
rect 11422 20244 11428 20256
rect 11201 20216 11428 20244
rect 11201 20213 11213 20216
rect 11155 20207 11213 20213
rect 11422 20204 11428 20216
rect 11480 20204 11486 20256
rect 11790 20204 11796 20256
rect 11848 20244 11854 20256
rect 12084 20244 12112 20352
rect 12986 20272 12992 20324
rect 13044 20272 13050 20324
rect 13817 20315 13875 20321
rect 13817 20281 13829 20315
rect 13863 20281 13875 20315
rect 14200 20312 14228 20352
rect 14274 20340 14280 20392
rect 14332 20340 14338 20392
rect 16117 20383 16175 20389
rect 16117 20349 16129 20383
rect 16163 20349 16175 20383
rect 16117 20343 16175 20349
rect 18877 20383 18935 20389
rect 18877 20349 18889 20383
rect 18923 20349 18935 20383
rect 18877 20343 18935 20349
rect 14553 20315 14611 20321
rect 14553 20312 14565 20315
rect 14200 20284 14565 20312
rect 13817 20275 13875 20281
rect 14553 20281 14565 20284
rect 14599 20312 14611 20315
rect 14826 20312 14832 20324
rect 14599 20284 14832 20312
rect 14599 20281 14611 20284
rect 14553 20275 14611 20281
rect 11848 20216 12112 20244
rect 11848 20204 11854 20216
rect 12158 20204 12164 20256
rect 12216 20244 12222 20256
rect 12529 20247 12587 20253
rect 12529 20244 12541 20247
rect 12216 20216 12541 20244
rect 12216 20204 12222 20216
rect 12529 20213 12541 20216
rect 12575 20213 12587 20247
rect 13832 20244 13860 20275
rect 14826 20272 14832 20284
rect 14884 20272 14890 20324
rect 15286 20272 15292 20324
rect 15344 20272 15350 20324
rect 15930 20244 15936 20256
rect 13832 20216 15936 20244
rect 12529 20207 12587 20213
rect 15930 20204 15936 20216
rect 15988 20244 15994 20256
rect 16132 20244 16160 20343
rect 17420 20284 17632 20312
rect 15988 20216 16160 20244
rect 15988 20204 15994 20216
rect 16850 20204 16856 20256
rect 16908 20244 16914 20256
rect 17420 20244 17448 20284
rect 16908 20216 17448 20244
rect 16908 20204 16914 20216
rect 17494 20204 17500 20256
rect 17552 20204 17558 20256
rect 17604 20244 17632 20284
rect 17954 20272 17960 20324
rect 18012 20272 18018 20324
rect 18892 20312 18920 20343
rect 20714 20340 20720 20392
rect 20772 20340 20778 20392
rect 21266 20380 21272 20392
rect 20916 20352 21272 20380
rect 19518 20312 19524 20324
rect 18892 20284 19524 20312
rect 19518 20272 19524 20284
rect 19576 20272 19582 20324
rect 19613 20315 19671 20321
rect 19613 20281 19625 20315
rect 19659 20281 19671 20315
rect 19613 20275 19671 20281
rect 18049 20247 18107 20253
rect 18049 20244 18061 20247
rect 17604 20216 18061 20244
rect 18049 20213 18061 20216
rect 18095 20213 18107 20247
rect 19628 20244 19656 20275
rect 20916 20244 20944 20352
rect 21266 20340 21272 20352
rect 21324 20380 21330 20392
rect 23584 20389 23612 20420
rect 24121 20417 24133 20451
rect 24167 20448 24179 20451
rect 27203 20451 27261 20457
rect 24167 20420 25912 20448
rect 24167 20417 24179 20420
rect 24121 20411 24179 20417
rect 21361 20383 21419 20389
rect 21361 20380 21373 20383
rect 21324 20352 21373 20380
rect 21324 20340 21330 20352
rect 21361 20349 21373 20352
rect 21407 20349 21419 20383
rect 21361 20343 21419 20349
rect 21545 20383 21603 20389
rect 21545 20349 21557 20383
rect 21591 20349 21603 20383
rect 21545 20343 21603 20349
rect 23569 20383 23627 20389
rect 23569 20349 23581 20383
rect 23615 20380 23627 20383
rect 23845 20383 23903 20389
rect 23845 20380 23857 20383
rect 23615 20352 23857 20380
rect 23615 20349 23627 20352
rect 23569 20343 23627 20349
rect 23845 20349 23857 20352
rect 23891 20349 23903 20383
rect 23845 20343 23903 20349
rect 21560 20312 21588 20343
rect 25130 20340 25136 20392
rect 25188 20380 25194 20392
rect 25188 20352 25254 20380
rect 25188 20340 25194 20352
rect 25406 20340 25412 20392
rect 25464 20340 25470 20392
rect 25884 20389 25912 20420
rect 27203 20417 27215 20451
rect 27249 20448 27261 20451
rect 28534 20448 28540 20460
rect 27249 20420 28540 20448
rect 27249 20417 27261 20420
rect 27203 20411 27261 20417
rect 28534 20408 28540 20420
rect 28592 20408 28598 20460
rect 29178 20408 29184 20460
rect 29236 20448 29242 20460
rect 29236 20420 29592 20448
rect 29236 20408 29242 20420
rect 25869 20383 25927 20389
rect 25869 20349 25881 20383
rect 25915 20349 25927 20383
rect 25869 20343 25927 20349
rect 25958 20340 25964 20392
rect 26016 20380 26022 20392
rect 26145 20383 26203 20389
rect 26145 20380 26157 20383
rect 26016 20352 26157 20380
rect 26016 20340 26022 20352
rect 26145 20349 26157 20352
rect 26191 20349 26203 20383
rect 26145 20343 26203 20349
rect 26697 20383 26755 20389
rect 26697 20349 26709 20383
rect 26743 20380 26755 20383
rect 27338 20380 27344 20392
rect 26743 20352 27344 20380
rect 26743 20349 26755 20352
rect 26697 20343 26755 20349
rect 27338 20340 27344 20352
rect 27396 20340 27402 20392
rect 27433 20383 27491 20389
rect 27433 20349 27445 20383
rect 27479 20380 27491 20383
rect 29270 20380 29276 20392
rect 27479 20352 29276 20380
rect 27479 20349 27491 20352
rect 27433 20343 27491 20349
rect 29270 20340 29276 20352
rect 29328 20340 29334 20392
rect 29454 20340 29460 20392
rect 29512 20340 29518 20392
rect 29564 20380 29592 20420
rect 29730 20408 29736 20460
rect 29788 20448 29794 20460
rect 30377 20451 30435 20457
rect 30377 20448 30389 20451
rect 29788 20420 30389 20448
rect 29788 20408 29794 20420
rect 30377 20417 30389 20420
rect 30423 20417 30435 20451
rect 30377 20411 30435 20417
rect 29825 20383 29883 20389
rect 29825 20380 29837 20383
rect 29564 20352 29837 20380
rect 29825 20349 29837 20352
rect 29871 20349 29883 20383
rect 29825 20343 29883 20349
rect 23106 20312 23112 20324
rect 21560 20284 22094 20312
rect 23046 20284 23112 20312
rect 19628 20216 20944 20244
rect 21177 20247 21235 20253
rect 18049 20207 18107 20213
rect 21177 20213 21189 20247
rect 21223 20244 21235 20247
rect 21542 20244 21548 20256
rect 21223 20216 21548 20244
rect 21223 20213 21235 20216
rect 21177 20207 21235 20213
rect 21542 20204 21548 20216
rect 21600 20204 21606 20256
rect 22066 20244 22094 20284
rect 23106 20272 23112 20284
rect 23164 20312 23170 20324
rect 24118 20312 24124 20324
rect 23164 20284 24124 20312
rect 23164 20272 23170 20284
rect 24118 20272 24124 20284
rect 24176 20272 24182 20324
rect 22462 20244 22468 20256
rect 22066 20216 22468 20244
rect 22462 20204 22468 20216
rect 22520 20204 22526 20256
rect 23385 20247 23443 20253
rect 23385 20213 23397 20247
rect 23431 20244 23443 20247
rect 24854 20244 24860 20256
rect 23431 20216 24860 20244
rect 23431 20213 23443 20216
rect 23385 20207 23443 20213
rect 24854 20204 24860 20216
rect 24912 20204 24918 20256
rect 25424 20244 25452 20340
rect 29089 20315 29147 20321
rect 29089 20281 29101 20315
rect 29135 20281 29147 20315
rect 29089 20275 29147 20281
rect 25685 20247 25743 20253
rect 25685 20244 25697 20247
rect 25424 20216 25697 20244
rect 25685 20213 25697 20216
rect 25731 20213 25743 20247
rect 25685 20207 25743 20213
rect 27163 20247 27221 20253
rect 27163 20213 27175 20247
rect 27209 20244 27221 20247
rect 28166 20244 28172 20256
rect 27209 20216 28172 20244
rect 27209 20213 27221 20216
rect 27163 20207 27221 20213
rect 28166 20204 28172 20216
rect 28224 20244 28230 20256
rect 28810 20244 28816 20256
rect 28224 20216 28816 20244
rect 28224 20204 28230 20216
rect 28810 20204 28816 20216
rect 28868 20204 28874 20256
rect 29104 20244 29132 20275
rect 30006 20272 30012 20324
rect 30064 20312 30070 20324
rect 30101 20315 30159 20321
rect 30101 20312 30113 20315
rect 30064 20284 30113 20312
rect 30064 20272 30070 20284
rect 30101 20281 30113 20284
rect 30147 20312 30159 20315
rect 31386 20312 31392 20324
rect 30147 20284 31392 20312
rect 30147 20281 30159 20284
rect 30101 20275 30159 20281
rect 31386 20272 31392 20284
rect 31444 20272 31450 20324
rect 29638 20244 29644 20256
rect 29104 20216 29644 20244
rect 29638 20204 29644 20216
rect 29696 20204 29702 20256
rect 29822 20204 29828 20256
rect 29880 20244 29886 20256
rect 29917 20247 29975 20253
rect 29917 20244 29929 20247
rect 29880 20216 29929 20244
rect 29880 20204 29886 20216
rect 29917 20213 29929 20216
rect 29963 20213 29975 20247
rect 29917 20207 29975 20213
rect 552 20154 31072 20176
rect 552 20102 7988 20154
rect 8040 20102 8052 20154
rect 8104 20102 8116 20154
rect 8168 20102 8180 20154
rect 8232 20102 8244 20154
rect 8296 20102 15578 20154
rect 15630 20102 15642 20154
rect 15694 20102 15706 20154
rect 15758 20102 15770 20154
rect 15822 20102 15834 20154
rect 15886 20102 23168 20154
rect 23220 20102 23232 20154
rect 23284 20102 23296 20154
rect 23348 20102 23360 20154
rect 23412 20102 23424 20154
rect 23476 20102 30758 20154
rect 30810 20102 30822 20154
rect 30874 20102 30886 20154
rect 30938 20102 30950 20154
rect 31002 20102 31014 20154
rect 31066 20102 31072 20154
rect 552 20080 31072 20102
rect 1394 20040 1400 20052
rect 952 20012 1400 20040
rect 952 19904 980 20012
rect 1394 20000 1400 20012
rect 1452 20000 1458 20052
rect 3418 20040 3424 20052
rect 2976 20012 3424 20040
rect 2976 19981 3004 20012
rect 3418 20000 3424 20012
rect 3476 20000 3482 20052
rect 4246 20000 4252 20052
rect 4304 20040 4310 20052
rect 4304 20012 7328 20040
rect 4304 20000 4310 20012
rect 2961 19975 3019 19981
rect 2961 19941 2973 19975
rect 3007 19941 3019 19975
rect 5994 19972 6000 19984
rect 2961 19935 3019 19941
rect 5552 19944 6000 19972
rect 1172 19907 1230 19913
rect 1172 19904 1184 19907
rect 952 19876 1184 19904
rect 1172 19873 1184 19876
rect 1218 19873 1230 19907
rect 5552 19904 5580 19944
rect 5994 19932 6000 19944
rect 6052 19932 6058 19984
rect 1172 19867 1230 19873
rect 1504 19876 2774 19904
rect 842 19796 848 19848
rect 900 19796 906 19848
rect 1351 19839 1409 19845
rect 1351 19805 1363 19839
rect 1397 19836 1409 19839
rect 1504 19836 1532 19876
rect 1397 19808 1532 19836
rect 1397 19805 1409 19808
rect 1351 19799 1409 19805
rect 1578 19796 1584 19848
rect 1636 19796 1642 19848
rect 2746 19700 2774 19876
rect 3712 19876 5580 19904
rect 3712 19848 3740 19876
rect 5626 19864 5632 19916
rect 5684 19864 5690 19916
rect 6294 19904 6411 19908
rect 5736 19880 6411 19904
rect 5736 19876 6322 19880
rect 2958 19796 2964 19848
rect 3016 19836 3022 19848
rect 3053 19839 3111 19845
rect 3053 19836 3065 19839
rect 3016 19808 3065 19836
rect 3016 19796 3022 19808
rect 3053 19805 3065 19808
rect 3099 19805 3111 19839
rect 3053 19799 3111 19805
rect 3234 19796 3240 19848
rect 3292 19836 3298 19848
rect 3602 19847 3608 19848
rect 3380 19839 3438 19845
rect 3380 19836 3392 19839
rect 3292 19808 3392 19836
rect 3292 19796 3298 19808
rect 3380 19805 3392 19808
rect 3426 19805 3438 19839
rect 3380 19799 3438 19805
rect 3559 19841 3608 19847
rect 3559 19807 3571 19841
rect 3605 19807 3608 19841
rect 3559 19801 3608 19807
rect 3602 19796 3608 19801
rect 3660 19796 3666 19848
rect 3694 19796 3700 19848
rect 3752 19796 3758 19848
rect 3789 19839 3847 19845
rect 3789 19805 3801 19839
rect 3835 19836 3847 19839
rect 5258 19836 5264 19848
rect 3835 19808 5264 19836
rect 3835 19805 3847 19808
rect 3789 19799 3847 19805
rect 5258 19796 5264 19808
rect 5316 19796 5322 19848
rect 5350 19796 5356 19848
rect 5408 19836 5414 19848
rect 5736 19836 5764 19876
rect 5408 19808 5764 19836
rect 5408 19796 5414 19808
rect 5902 19796 5908 19848
rect 5960 19836 5966 19848
rect 6086 19836 6092 19848
rect 5960 19808 6092 19836
rect 5960 19796 5966 19808
rect 6086 19796 6092 19808
rect 6144 19796 6150 19848
rect 6270 19845 6276 19848
rect 6232 19839 6276 19845
rect 6232 19805 6244 19839
rect 6232 19799 6276 19805
rect 6270 19796 6276 19799
rect 6328 19796 6334 19848
rect 6383 19845 6411 19880
rect 6368 19839 6426 19845
rect 6368 19805 6380 19839
rect 6414 19805 6426 19839
rect 6368 19799 6426 19805
rect 6638 19796 6644 19848
rect 6696 19796 6702 19848
rect 7300 19836 7328 20012
rect 8938 20000 8944 20052
rect 8996 20049 9002 20052
rect 8996 20040 9005 20049
rect 8996 20012 9041 20040
rect 8996 20003 9005 20012
rect 8996 20000 9002 20003
rect 9214 20000 9220 20052
rect 9272 20040 9278 20052
rect 11146 20040 11152 20052
rect 9272 20012 11152 20040
rect 9272 20000 9278 20012
rect 11146 20000 11152 20012
rect 11204 20000 11210 20052
rect 11885 20043 11943 20049
rect 11885 20009 11897 20043
rect 11931 20040 11943 20043
rect 12250 20040 12256 20052
rect 11931 20012 12256 20040
rect 11931 20009 11943 20012
rect 11885 20003 11943 20009
rect 12250 20000 12256 20012
rect 12308 20000 12314 20052
rect 12434 20000 12440 20052
rect 12492 20040 12498 20052
rect 12627 20043 12685 20049
rect 12627 20040 12639 20043
rect 12492 20012 12639 20040
rect 12492 20000 12498 20012
rect 12627 20009 12639 20012
rect 12673 20009 12685 20043
rect 12627 20003 12685 20009
rect 13538 20000 13544 20052
rect 13596 20040 13602 20052
rect 14001 20043 14059 20049
rect 14001 20040 14013 20043
rect 13596 20012 14013 20040
rect 13596 20000 13602 20012
rect 14001 20009 14013 20012
rect 14047 20009 14059 20043
rect 14001 20003 14059 20009
rect 15194 20000 15200 20052
rect 15252 20000 15258 20052
rect 15286 20000 15292 20052
rect 15344 20040 15350 20052
rect 15473 20043 15531 20049
rect 15473 20040 15485 20043
rect 15344 20012 15485 20040
rect 15344 20000 15350 20012
rect 15473 20009 15485 20012
rect 15519 20009 15531 20043
rect 15473 20003 15531 20009
rect 8021 19975 8079 19981
rect 8021 19941 8033 19975
rect 8067 19972 8079 19975
rect 11698 19972 11704 19984
rect 8067 19944 8616 19972
rect 8067 19941 8079 19944
rect 8021 19935 8079 19941
rect 8113 19907 8171 19913
rect 8113 19873 8125 19907
rect 8159 19904 8171 19907
rect 8294 19904 8300 19916
rect 8159 19876 8300 19904
rect 8159 19873 8171 19876
rect 8113 19867 8171 19873
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 8386 19864 8392 19916
rect 8444 19904 8450 19916
rect 8481 19907 8539 19913
rect 8481 19904 8493 19907
rect 8444 19876 8493 19904
rect 8444 19864 8450 19876
rect 8481 19873 8493 19876
rect 8527 19873 8539 19907
rect 8481 19867 8539 19873
rect 8588 19836 8616 19944
rect 10980 19944 11704 19972
rect 10980 19913 11008 19944
rect 11698 19932 11704 19944
rect 11756 19932 11762 19984
rect 13722 19932 13728 19984
rect 13780 19972 13786 19984
rect 15212 19972 15240 20000
rect 13780 19944 15240 19972
rect 15488 19972 15516 20003
rect 16114 20000 16120 20052
rect 16172 20040 16178 20052
rect 16761 20043 16819 20049
rect 16761 20040 16773 20043
rect 16172 20012 16773 20040
rect 16172 20000 16178 20012
rect 16761 20009 16773 20012
rect 16807 20009 16819 20043
rect 16761 20003 16819 20009
rect 19794 20000 19800 20052
rect 19852 20040 19858 20052
rect 20073 20043 20131 20049
rect 20073 20040 20085 20043
rect 19852 20012 20085 20040
rect 19852 20000 19858 20012
rect 20073 20009 20085 20012
rect 20119 20009 20131 20043
rect 20073 20003 20131 20009
rect 20530 20000 20536 20052
rect 20588 20000 20594 20052
rect 21082 20000 21088 20052
rect 21140 20000 21146 20052
rect 21450 20040 21456 20052
rect 21192 20012 21456 20040
rect 15488 19944 16160 19972
rect 13780 19932 13786 19944
rect 10965 19907 11023 19913
rect 10965 19873 10977 19907
rect 11011 19873 11023 19907
rect 10965 19867 11023 19873
rect 11241 19907 11299 19913
rect 11241 19873 11253 19907
rect 11287 19904 11299 19907
rect 11790 19904 11796 19916
rect 11287 19876 11796 19904
rect 11287 19873 11299 19876
rect 11241 19867 11299 19873
rect 11790 19864 11796 19876
rect 11848 19864 11854 19916
rect 12897 19907 12955 19913
rect 12897 19904 12909 19907
rect 11900 19876 12909 19904
rect 8960 19857 9018 19863
rect 8960 19836 8972 19857
rect 7300 19808 8432 19836
rect 8588 19823 8972 19836
rect 9006 19823 9018 19857
rect 8588 19817 9018 19823
rect 8588 19808 8990 19817
rect 2866 19700 2872 19712
rect 2746 19672 2872 19700
rect 2866 19660 2872 19672
rect 2924 19660 2930 19712
rect 5074 19660 5080 19712
rect 5132 19660 5138 19712
rect 5445 19703 5503 19709
rect 5445 19669 5457 19703
rect 5491 19700 5503 19703
rect 6822 19700 6828 19712
rect 5491 19672 6828 19700
rect 5491 19669 5503 19672
rect 5445 19663 5503 19669
rect 6822 19660 6828 19672
rect 6880 19660 6886 19712
rect 8294 19660 8300 19712
rect 8352 19660 8358 19712
rect 8404 19700 8432 19808
rect 9214 19796 9220 19848
rect 9272 19796 9278 19848
rect 10321 19703 10379 19709
rect 10321 19700 10333 19703
rect 8404 19672 10333 19700
rect 10321 19669 10333 19672
rect 10367 19669 10379 19703
rect 10321 19663 10379 19669
rect 10778 19660 10784 19712
rect 10836 19700 10842 19712
rect 11900 19700 11928 19876
rect 12897 19873 12909 19876
rect 12943 19873 12955 19907
rect 14550 19904 14556 19916
rect 12897 19867 12955 19873
rect 14292 19876 14556 19904
rect 11974 19796 11980 19848
rect 12032 19836 12038 19848
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 12032 19808 12173 19836
rect 12032 19796 12038 19808
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 12618 19796 12624 19848
rect 12676 19836 12682 19848
rect 12676 19808 12721 19836
rect 12676 19796 12682 19808
rect 12802 19796 12808 19848
rect 12860 19836 12866 19848
rect 14292 19836 14320 19876
rect 14550 19864 14556 19876
rect 14608 19864 14614 19916
rect 14645 19907 14703 19913
rect 14645 19873 14657 19907
rect 14691 19904 14703 19907
rect 14826 19904 14832 19916
rect 14691 19876 14832 19904
rect 14691 19873 14703 19876
rect 14645 19867 14703 19873
rect 14826 19864 14832 19876
rect 14884 19904 14890 19916
rect 14884 19876 15516 19904
rect 14884 19864 14890 19876
rect 12860 19808 14320 19836
rect 12860 19796 12866 19808
rect 14366 19796 14372 19848
rect 14424 19796 14430 19848
rect 15488 19836 15516 19876
rect 15562 19864 15568 19916
rect 15620 19904 15626 19916
rect 15933 19907 15991 19913
rect 15933 19904 15945 19907
rect 15620 19876 15945 19904
rect 15620 19864 15626 19876
rect 15933 19873 15945 19876
rect 15979 19873 15991 19907
rect 15933 19867 15991 19873
rect 16132 19848 16160 19944
rect 16206 19932 16212 19984
rect 16264 19932 16270 19984
rect 16390 19932 16396 19984
rect 16448 19972 16454 19984
rect 21192 19972 21220 20012
rect 21450 20000 21456 20012
rect 21508 20000 21514 20052
rect 21542 20000 21548 20052
rect 21600 20040 21606 20052
rect 21600 20012 23796 20040
rect 21600 20000 21606 20012
rect 23768 19972 23796 20012
rect 23934 20000 23940 20052
rect 23992 20040 23998 20052
rect 24029 20043 24087 20049
rect 24029 20040 24041 20043
rect 23992 20012 24041 20040
rect 23992 20000 23998 20012
rect 24029 20009 24041 20012
rect 24075 20009 24087 20043
rect 24029 20003 24087 20009
rect 24118 20000 24124 20052
rect 24176 20040 24182 20052
rect 25130 20040 25136 20052
rect 24176 20012 25136 20040
rect 24176 20000 24182 20012
rect 25130 20000 25136 20012
rect 25188 20000 25194 20052
rect 28810 20000 28816 20052
rect 28868 20049 28874 20052
rect 28868 20040 28877 20049
rect 28868 20012 28913 20040
rect 28868 20003 28877 20012
rect 28868 20000 28874 20003
rect 24136 19972 24164 20000
rect 16448 19944 16528 19972
rect 16448 19932 16454 19944
rect 16224 19904 16252 19932
rect 16500 19913 16528 19944
rect 20640 19944 21220 19972
rect 23690 19944 24164 19972
rect 20640 19916 20668 19944
rect 16301 19907 16359 19913
rect 16301 19904 16313 19907
rect 16224 19876 16313 19904
rect 16301 19873 16313 19876
rect 16347 19873 16359 19907
rect 16301 19867 16359 19873
rect 16485 19907 16543 19913
rect 16485 19873 16497 19907
rect 16531 19873 16543 19907
rect 16485 19867 16543 19873
rect 17954 19864 17960 19916
rect 18012 19864 18018 19916
rect 18601 19907 18659 19913
rect 18601 19873 18613 19907
rect 18647 19904 18659 19907
rect 18969 19907 19027 19913
rect 18969 19904 18981 19907
rect 18647 19876 18981 19904
rect 18647 19873 18659 19876
rect 18601 19867 18659 19873
rect 18969 19873 18981 19876
rect 19015 19873 19027 19907
rect 18969 19867 19027 19873
rect 20622 19864 20628 19916
rect 20680 19864 20686 19916
rect 20898 19864 20904 19916
rect 20956 19864 20962 19916
rect 21542 19864 21548 19916
rect 21600 19864 21606 19916
rect 21821 19907 21879 19913
rect 21821 19873 21833 19907
rect 21867 19873 21879 19907
rect 21821 19867 21879 19873
rect 15488 19808 15884 19836
rect 15856 19768 15884 19808
rect 16114 19796 16120 19848
rect 16172 19836 16178 19848
rect 16209 19839 16267 19845
rect 16209 19836 16221 19839
rect 16172 19808 16221 19836
rect 16172 19796 16178 19808
rect 16209 19805 16221 19808
rect 16255 19805 16267 19839
rect 16209 19799 16267 19805
rect 16850 19796 16856 19848
rect 16908 19836 16914 19848
rect 16945 19839 17003 19845
rect 16945 19836 16957 19839
rect 16908 19808 16957 19836
rect 16908 19796 16914 19808
rect 16945 19805 16957 19808
rect 16991 19805 17003 19839
rect 16945 19799 17003 19805
rect 17218 19796 17224 19848
rect 17276 19796 17282 19848
rect 17972 19836 18000 19864
rect 18690 19836 18696 19848
rect 17972 19808 18696 19836
rect 18690 19796 18696 19808
rect 18748 19796 18754 19848
rect 20714 19796 20720 19848
rect 20772 19836 20778 19848
rect 21560 19836 21588 19864
rect 20772 19808 21588 19836
rect 20772 19796 20778 19808
rect 16298 19768 16304 19780
rect 14936 19740 15792 19768
rect 15856 19740 16304 19768
rect 10836 19672 11928 19700
rect 12069 19703 12127 19709
rect 10836 19660 10842 19672
rect 12069 19669 12081 19703
rect 12115 19700 12127 19703
rect 12802 19700 12808 19712
rect 12115 19672 12808 19700
rect 12115 19669 12127 19672
rect 12069 19663 12127 19669
rect 12802 19660 12808 19672
rect 12860 19660 12866 19712
rect 13078 19660 13084 19712
rect 13136 19700 13142 19712
rect 14936 19700 14964 19740
rect 13136 19672 14964 19700
rect 13136 19660 13142 19672
rect 15286 19660 15292 19712
rect 15344 19700 15350 19712
rect 15764 19709 15792 19740
rect 16298 19728 16304 19740
rect 16356 19728 16362 19780
rect 19886 19728 19892 19780
rect 19944 19768 19950 19780
rect 21836 19768 21864 19867
rect 22186 19864 22192 19916
rect 22244 19864 22250 19916
rect 24213 19907 24271 19913
rect 24213 19873 24225 19907
rect 24259 19873 24271 19907
rect 24213 19867 24271 19873
rect 26053 19907 26111 19913
rect 26053 19873 26065 19907
rect 26099 19904 26111 19907
rect 26697 19907 26755 19913
rect 26697 19904 26709 19907
rect 26099 19876 26709 19904
rect 26099 19873 26111 19876
rect 26053 19867 26111 19873
rect 26697 19873 26709 19876
rect 26743 19873 26755 19907
rect 26697 19867 26755 19873
rect 22462 19796 22468 19848
rect 22520 19836 22526 19848
rect 24228 19836 24256 19867
rect 27338 19864 27344 19916
rect 27396 19904 27402 19916
rect 28353 19907 28411 19913
rect 28353 19904 28365 19907
rect 27396 19876 28365 19904
rect 27396 19864 27402 19876
rect 28353 19873 28365 19876
rect 28399 19904 28411 19907
rect 28442 19904 28448 19916
rect 28399 19876 28448 19904
rect 28399 19873 28411 19876
rect 28353 19867 28411 19873
rect 28442 19864 28448 19876
rect 28500 19864 28506 19916
rect 30469 19907 30527 19913
rect 30469 19904 30481 19907
rect 28552 19876 30481 19904
rect 22520 19808 24256 19836
rect 22520 19796 22526 19808
rect 24394 19796 24400 19848
rect 24452 19796 24458 19848
rect 24670 19796 24676 19848
rect 24728 19796 24734 19848
rect 26421 19839 26479 19845
rect 26421 19805 26433 19839
rect 26467 19836 26479 19839
rect 26878 19836 26884 19848
rect 26467 19808 26884 19836
rect 26467 19805 26479 19808
rect 26421 19799 26479 19805
rect 26878 19796 26884 19808
rect 26936 19796 26942 19848
rect 27522 19796 27528 19848
rect 27580 19836 27586 19848
rect 28552 19836 28580 19876
rect 30469 19873 30481 19876
rect 30515 19873 30527 19907
rect 30469 19867 30527 19873
rect 28902 19845 28908 19848
rect 27580 19808 28580 19836
rect 28859 19839 28908 19845
rect 27580 19796 27586 19808
rect 28859 19805 28871 19839
rect 28905 19805 28908 19839
rect 28859 19799 28908 19805
rect 28902 19796 28908 19799
rect 28960 19796 28966 19848
rect 29086 19796 29092 19848
rect 29144 19796 29150 19848
rect 19944 19740 21864 19768
rect 19944 19728 19950 19740
rect 15657 19703 15715 19709
rect 15657 19700 15669 19703
rect 15344 19672 15669 19700
rect 15344 19660 15350 19672
rect 15657 19669 15669 19672
rect 15703 19669 15715 19703
rect 15657 19663 15715 19669
rect 15749 19703 15807 19709
rect 15749 19669 15761 19703
rect 15795 19669 15807 19703
rect 15749 19663 15807 19669
rect 21358 19660 21364 19712
rect 21416 19660 21422 19712
rect 27982 19660 27988 19712
rect 28040 19660 28046 19712
rect 28074 19660 28080 19712
rect 28132 19700 28138 19712
rect 30466 19700 30472 19712
rect 28132 19672 30472 19700
rect 28132 19660 28138 19672
rect 30466 19660 30472 19672
rect 30524 19660 30530 19712
rect 552 19610 30912 19632
rect 552 19558 4193 19610
rect 4245 19558 4257 19610
rect 4309 19558 4321 19610
rect 4373 19558 4385 19610
rect 4437 19558 4449 19610
rect 4501 19558 11783 19610
rect 11835 19558 11847 19610
rect 11899 19558 11911 19610
rect 11963 19558 11975 19610
rect 12027 19558 12039 19610
rect 12091 19558 19373 19610
rect 19425 19558 19437 19610
rect 19489 19558 19501 19610
rect 19553 19558 19565 19610
rect 19617 19558 19629 19610
rect 19681 19558 26963 19610
rect 27015 19558 27027 19610
rect 27079 19558 27091 19610
rect 27143 19558 27155 19610
rect 27207 19558 27219 19610
rect 27271 19558 30912 19610
rect 552 19536 30912 19558
rect 5074 19456 5080 19508
rect 5132 19456 5138 19508
rect 6086 19456 6092 19508
rect 6144 19496 6150 19508
rect 6144 19468 6868 19496
rect 6144 19456 6150 19468
rect 842 19320 848 19372
rect 900 19360 906 19372
rect 937 19363 995 19369
rect 937 19360 949 19363
rect 900 19332 949 19360
rect 900 19320 906 19332
rect 937 19329 949 19332
rect 983 19329 995 19363
rect 2038 19360 2044 19372
rect 937 19323 995 19329
rect 1412 19345 2044 19360
rect 1412 19314 1445 19345
rect 1433 19311 1445 19314
rect 1479 19332 2044 19345
rect 1479 19311 1491 19332
rect 2038 19320 2044 19332
rect 2096 19320 2102 19372
rect 2958 19320 2964 19372
rect 3016 19360 3022 19372
rect 3234 19360 3240 19372
rect 3016 19332 3240 19360
rect 3016 19320 3022 19332
rect 3234 19320 3240 19332
rect 3292 19320 3298 19372
rect 3743 19363 3801 19369
rect 3743 19329 3755 19363
rect 3789 19360 3801 19363
rect 5092 19360 5120 19456
rect 6840 19428 6868 19468
rect 8294 19456 8300 19508
rect 8352 19496 8358 19508
rect 8352 19468 9812 19496
rect 8352 19456 8358 19468
rect 6840 19400 8340 19428
rect 5908 19363 5966 19369
rect 5908 19360 5920 19363
rect 3789 19332 4292 19360
rect 5092 19332 5920 19360
rect 3789 19329 3801 19332
rect 3743 19323 3801 19329
rect 1433 19305 1491 19311
rect 4264 19304 4292 19332
rect 5908 19329 5920 19332
rect 5954 19329 5966 19363
rect 6086 19360 6092 19372
rect 5908 19323 5966 19329
rect 6012 19332 6092 19360
rect 1673 19295 1731 19301
rect 1673 19261 1685 19295
rect 1719 19292 1731 19295
rect 1946 19292 1952 19304
rect 1719 19264 1952 19292
rect 1719 19261 1731 19264
rect 1673 19255 1731 19261
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 3142 19252 3148 19304
rect 3200 19292 3206 19304
rect 3564 19295 3622 19301
rect 3564 19292 3576 19295
rect 3200 19264 3576 19292
rect 3200 19252 3206 19264
rect 3564 19261 3576 19264
rect 3610 19292 3622 19295
rect 3878 19292 3884 19304
rect 3610 19264 3884 19292
rect 3610 19261 3622 19264
rect 3564 19255 3622 19261
rect 3878 19252 3884 19264
rect 3936 19252 3942 19304
rect 3970 19252 3976 19304
rect 4028 19252 4034 19304
rect 4246 19252 4252 19304
rect 4304 19252 4310 19304
rect 5350 19252 5356 19304
rect 5408 19252 5414 19304
rect 5445 19295 5503 19301
rect 5445 19261 5457 19295
rect 5491 19292 5503 19295
rect 6012 19292 6040 19332
rect 6086 19320 6092 19332
rect 6144 19320 6150 19372
rect 7650 19320 7656 19372
rect 7708 19320 7714 19372
rect 8312 19360 8340 19400
rect 8312 19332 8524 19360
rect 5491 19264 6040 19292
rect 6181 19295 6239 19301
rect 5491 19261 5503 19264
rect 5445 19255 5503 19261
rect 6181 19261 6193 19295
rect 6227 19292 6239 19295
rect 6638 19292 6644 19304
rect 6227 19264 6644 19292
rect 6227 19261 6239 19264
rect 6181 19255 6239 19261
rect 4706 19184 4712 19236
rect 4764 19224 4770 19236
rect 5460 19224 5488 19255
rect 6638 19252 6644 19264
rect 6696 19252 6702 19304
rect 7374 19252 7380 19304
rect 7432 19252 7438 19304
rect 7561 19295 7619 19301
rect 7561 19261 7573 19295
rect 7607 19292 7619 19295
rect 7668 19292 7696 19320
rect 7607 19264 7696 19292
rect 7745 19295 7803 19301
rect 7607 19261 7619 19264
rect 7561 19255 7619 19261
rect 7745 19261 7757 19295
rect 7791 19261 7803 19295
rect 7745 19255 7803 19261
rect 4764 19196 5488 19224
rect 7392 19224 7420 19252
rect 7760 19224 7788 19255
rect 8386 19252 8392 19304
rect 8444 19252 8450 19304
rect 8496 19236 8524 19332
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 8852 19363 8910 19369
rect 8852 19360 8864 19363
rect 8628 19332 8864 19360
rect 8628 19320 8634 19332
rect 8852 19329 8864 19332
rect 8898 19329 8910 19363
rect 8852 19323 8910 19329
rect 8938 19320 8944 19372
rect 8996 19360 9002 19372
rect 9490 19360 9496 19372
rect 8996 19332 9496 19360
rect 8996 19320 9002 19332
rect 9490 19320 9496 19332
rect 9548 19320 9554 19372
rect 9125 19295 9183 19301
rect 9125 19261 9137 19295
rect 9171 19292 9183 19295
rect 9582 19292 9588 19304
rect 9171 19264 9588 19292
rect 9171 19261 9183 19264
rect 9125 19255 9183 19261
rect 9582 19252 9588 19264
rect 9640 19252 9646 19304
rect 9784 19292 9812 19468
rect 10226 19456 10232 19508
rect 10284 19456 10290 19508
rect 11057 19499 11115 19505
rect 11057 19465 11069 19499
rect 11103 19496 11115 19499
rect 11238 19496 11244 19508
rect 11103 19468 11244 19496
rect 11103 19465 11115 19468
rect 11057 19459 11115 19465
rect 11238 19456 11244 19468
rect 11296 19496 11302 19508
rect 11974 19496 11980 19508
rect 11296 19468 11980 19496
rect 11296 19456 11302 19468
rect 11974 19456 11980 19468
rect 12032 19456 12038 19508
rect 12342 19456 12348 19508
rect 12400 19496 12406 19508
rect 12400 19468 12940 19496
rect 12400 19456 12406 19468
rect 12912 19428 12940 19468
rect 12986 19456 12992 19508
rect 13044 19496 13050 19508
rect 13081 19499 13139 19505
rect 13081 19496 13093 19499
rect 13044 19468 13093 19496
rect 13044 19456 13050 19468
rect 13081 19465 13093 19468
rect 13127 19465 13139 19499
rect 14458 19496 14464 19508
rect 13081 19459 13139 19465
rect 13188 19468 14464 19496
rect 13188 19428 13216 19468
rect 14458 19456 14464 19468
rect 14516 19456 14522 19508
rect 18046 19456 18052 19508
rect 18104 19456 18110 19508
rect 22462 19456 22468 19508
rect 22520 19496 22526 19508
rect 23014 19496 23020 19508
rect 22520 19468 23020 19496
rect 22520 19456 22526 19468
rect 23014 19456 23020 19468
rect 23072 19456 23078 19508
rect 26418 19496 26424 19508
rect 24504 19468 26424 19496
rect 12912 19400 13216 19428
rect 11747 19363 11805 19369
rect 11747 19329 11759 19363
rect 11793 19360 11805 19363
rect 12158 19360 12164 19372
rect 11793 19332 12164 19360
rect 11793 19329 11805 19332
rect 11747 19323 11805 19329
rect 12158 19320 12164 19332
rect 12216 19320 12222 19372
rect 14004 19363 14062 19369
rect 14004 19360 14016 19363
rect 13188 19332 14016 19360
rect 13188 19304 13216 19332
rect 14004 19329 14016 19332
rect 14050 19329 14062 19363
rect 14004 19323 14062 19329
rect 14366 19320 14372 19372
rect 14424 19360 14430 19372
rect 14424 19332 15232 19360
rect 14424 19320 14430 19332
rect 11054 19292 11060 19304
rect 9784 19264 11060 19292
rect 11054 19252 11060 19264
rect 11112 19252 11118 19304
rect 11241 19295 11299 19301
rect 11241 19261 11253 19295
rect 11287 19292 11299 19295
rect 11882 19292 11888 19304
rect 11287 19264 11888 19292
rect 11287 19261 11299 19264
rect 11241 19255 11299 19261
rect 7392 19196 7788 19224
rect 8021 19227 8079 19233
rect 4764 19184 4770 19196
rect 8021 19193 8033 19227
rect 8067 19193 8079 19227
rect 8021 19187 8079 19193
rect 1394 19116 1400 19168
rect 1452 19165 1458 19168
rect 1452 19156 1461 19165
rect 2961 19159 3019 19165
rect 1452 19128 1497 19156
rect 1452 19119 1461 19128
rect 2961 19125 2973 19159
rect 3007 19156 3019 19159
rect 5166 19156 5172 19168
rect 3007 19128 5172 19156
rect 3007 19125 3019 19128
rect 2961 19119 3019 19125
rect 1452 19116 1458 19119
rect 5166 19116 5172 19128
rect 5224 19116 5230 19168
rect 5911 19159 5969 19165
rect 5911 19125 5923 19159
rect 5957 19156 5969 19159
rect 6270 19156 6276 19168
rect 5957 19128 6276 19156
rect 5957 19125 5969 19128
rect 5911 19119 5969 19125
rect 6270 19116 6276 19128
rect 6328 19116 6334 19168
rect 8036 19156 8064 19187
rect 8478 19184 8484 19236
rect 8536 19184 8542 19236
rect 10226 19184 10232 19236
rect 10284 19224 10290 19236
rect 10781 19227 10839 19233
rect 10781 19224 10793 19227
rect 10284 19196 10793 19224
rect 10284 19184 10290 19196
rect 10781 19193 10793 19196
rect 10827 19193 10839 19227
rect 10781 19187 10839 19193
rect 10870 19184 10876 19236
rect 10928 19224 10934 19236
rect 11256 19224 11284 19255
rect 11882 19252 11888 19264
rect 11940 19252 11946 19304
rect 11977 19295 12035 19301
rect 11977 19261 11989 19295
rect 12023 19292 12035 19295
rect 13078 19292 13084 19304
rect 12023 19264 13084 19292
rect 12023 19261 12035 19264
rect 11977 19255 12035 19261
rect 13078 19252 13084 19264
rect 13136 19252 13142 19304
rect 13170 19252 13176 19304
rect 13228 19252 13234 19304
rect 13538 19252 13544 19304
rect 13596 19252 13602 19304
rect 14274 19252 14280 19304
rect 14332 19252 14338 19304
rect 15204 19292 15232 19332
rect 15930 19320 15936 19372
rect 15988 19320 15994 19372
rect 18693 19363 18751 19369
rect 18693 19360 18705 19363
rect 16868 19332 18705 19360
rect 16868 19304 16896 19332
rect 18693 19329 18705 19332
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 22002 19320 22008 19372
rect 22060 19369 22066 19372
rect 24504 19369 24532 19468
rect 26418 19456 26424 19468
rect 26476 19456 26482 19508
rect 22060 19363 22109 19369
rect 22060 19329 22063 19363
rect 22097 19360 22109 19363
rect 24489 19363 24547 19369
rect 22097 19332 22153 19360
rect 23768 19332 23980 19360
rect 22097 19329 22109 19332
rect 22060 19323 22109 19329
rect 22060 19320 22066 19323
rect 23768 19304 23796 19332
rect 16022 19292 16028 19304
rect 15204 19264 16028 19292
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 16206 19252 16212 19304
rect 16264 19252 16270 19304
rect 16850 19252 16856 19304
rect 16908 19252 16914 19304
rect 17589 19295 17647 19301
rect 17589 19261 17601 19295
rect 17635 19292 17647 19295
rect 17635 19264 18184 19292
rect 17635 19261 17647 19264
rect 17589 19255 17647 19261
rect 10928 19196 11284 19224
rect 10928 19184 10934 19196
rect 15102 19184 15108 19236
rect 15160 19224 15166 19236
rect 15160 19196 15884 19224
rect 15160 19184 15166 19196
rect 8754 19156 8760 19168
rect 8036 19128 8760 19156
rect 8754 19116 8760 19128
rect 8812 19116 8818 19168
rect 8846 19116 8852 19168
rect 8904 19165 8910 19168
rect 8904 19156 8913 19165
rect 8904 19128 8949 19156
rect 8904 19119 8913 19128
rect 8904 19116 8910 19119
rect 9030 19116 9036 19168
rect 9088 19156 9094 19168
rect 11707 19159 11765 19165
rect 11707 19156 11719 19159
rect 9088 19128 11719 19156
rect 9088 19116 9094 19128
rect 11707 19125 11719 19128
rect 11753 19156 11765 19159
rect 12342 19156 12348 19168
rect 11753 19128 12348 19156
rect 11753 19125 11765 19128
rect 11707 19119 11765 19125
rect 12342 19116 12348 19128
rect 12400 19116 12406 19168
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 14007 19159 14065 19165
rect 14007 19156 14019 19159
rect 12492 19128 14019 19156
rect 12492 19116 12498 19128
rect 14007 19125 14019 19128
rect 14053 19125 14065 19159
rect 14007 19119 14065 19125
rect 14182 19116 14188 19168
rect 14240 19156 14246 19168
rect 15381 19159 15439 19165
rect 15381 19156 15393 19159
rect 14240 19128 15393 19156
rect 14240 19116 14246 19128
rect 15381 19125 15393 19128
rect 15427 19125 15439 19159
rect 15856 19156 15884 19196
rect 17770 19184 17776 19236
rect 17828 19184 17834 19236
rect 18156 19224 18184 19264
rect 18230 19252 18236 19304
rect 18288 19252 18294 19304
rect 18322 19252 18328 19304
rect 18380 19292 18386 19304
rect 18509 19295 18567 19301
rect 18509 19292 18521 19295
rect 18380 19264 18521 19292
rect 18380 19252 18386 19264
rect 18509 19261 18521 19264
rect 18555 19261 18567 19295
rect 18969 19295 19027 19301
rect 18969 19292 18981 19295
rect 18509 19255 18567 19261
rect 18800 19264 18981 19292
rect 18800 19224 18828 19264
rect 18969 19261 18981 19264
rect 19015 19261 19027 19295
rect 18969 19255 19027 19261
rect 20533 19295 20591 19301
rect 20533 19261 20545 19295
rect 20579 19292 20591 19295
rect 21174 19292 21180 19304
rect 20579 19264 21180 19292
rect 20579 19261 20591 19264
rect 20533 19255 20591 19261
rect 21174 19252 21180 19264
rect 21232 19252 21238 19304
rect 21545 19295 21603 19301
rect 21545 19261 21557 19295
rect 21591 19292 21603 19295
rect 21818 19292 21824 19304
rect 21591 19264 21824 19292
rect 21591 19261 21603 19264
rect 21545 19255 21603 19261
rect 21818 19252 21824 19264
rect 21876 19252 21882 19304
rect 22281 19295 22339 19301
rect 22281 19261 22293 19295
rect 22327 19292 22339 19295
rect 22327 19264 23704 19292
rect 22327 19261 22339 19264
rect 22281 19255 22339 19261
rect 18156 19196 18828 19224
rect 20717 19227 20775 19233
rect 20717 19193 20729 19227
rect 20763 19224 20775 19227
rect 21358 19224 21364 19236
rect 20763 19196 21364 19224
rect 20763 19193 20775 19196
rect 20717 19187 20775 19193
rect 21358 19184 21364 19196
rect 21416 19184 21422 19236
rect 17865 19159 17923 19165
rect 17865 19156 17877 19159
rect 15856 19128 17877 19156
rect 15381 19119 15439 19125
rect 17865 19125 17877 19128
rect 17911 19125 17923 19159
rect 17865 19119 17923 19125
rect 18322 19116 18328 19168
rect 18380 19116 18386 19168
rect 20070 19116 20076 19168
rect 20128 19116 20134 19168
rect 20806 19116 20812 19168
rect 20864 19116 20870 19168
rect 21082 19116 21088 19168
rect 21140 19116 21146 19168
rect 22011 19159 22069 19165
rect 22011 19125 22023 19159
rect 22057 19156 22069 19159
rect 22186 19156 22192 19168
rect 22057 19128 22192 19156
rect 22057 19125 22069 19128
rect 22011 19119 22069 19125
rect 22186 19116 22192 19128
rect 22244 19116 22250 19168
rect 23566 19116 23572 19168
rect 23624 19116 23630 19168
rect 23676 19156 23704 19264
rect 23750 19252 23756 19304
rect 23808 19252 23814 19304
rect 23842 19252 23848 19304
rect 23900 19252 23906 19304
rect 23952 19292 23980 19332
rect 24489 19329 24501 19363
rect 24535 19329 24547 19363
rect 24489 19323 24547 19329
rect 25179 19363 25237 19369
rect 25179 19329 25191 19363
rect 25225 19360 25237 19363
rect 25225 19332 25728 19360
rect 25225 19329 25237 19332
rect 25179 19323 25237 19329
rect 25700 19304 25728 19332
rect 26804 19332 27292 19360
rect 24213 19295 24271 19301
rect 24213 19292 24225 19295
rect 23952 19264 24225 19292
rect 24213 19261 24225 19264
rect 24259 19261 24271 19295
rect 24213 19255 24271 19261
rect 24302 19252 24308 19304
rect 24360 19252 24366 19304
rect 24578 19252 24584 19304
rect 24636 19292 24642 19304
rect 24673 19295 24731 19301
rect 24673 19292 24685 19295
rect 24636 19264 24685 19292
rect 24636 19252 24642 19264
rect 24673 19261 24685 19264
rect 24719 19261 24731 19295
rect 25409 19295 25467 19301
rect 25409 19292 25421 19295
rect 24673 19255 24731 19261
rect 24780 19264 25421 19292
rect 23750 19156 23756 19168
rect 23676 19128 23756 19156
rect 23750 19116 23756 19128
rect 23808 19116 23814 19168
rect 23860 19165 23888 19252
rect 24118 19184 24124 19236
rect 24176 19224 24182 19236
rect 24780 19224 24808 19264
rect 25409 19261 25421 19264
rect 25455 19261 25467 19295
rect 25409 19255 25467 19261
rect 25682 19252 25688 19304
rect 25740 19252 25746 19304
rect 26050 19252 26056 19304
rect 26108 19292 26114 19304
rect 26804 19292 26832 19332
rect 26108 19264 26832 19292
rect 26108 19252 26114 19264
rect 26878 19252 26884 19304
rect 26936 19252 26942 19304
rect 27157 19295 27215 19301
rect 27157 19292 27169 19295
rect 26988 19264 27169 19292
rect 24176 19196 24808 19224
rect 24176 19184 24182 19196
rect 26234 19184 26240 19236
rect 26292 19224 26298 19236
rect 26988 19224 27016 19264
rect 27157 19261 27169 19264
rect 27203 19261 27215 19295
rect 27264 19292 27292 19332
rect 28629 19295 28687 19301
rect 28629 19292 28641 19295
rect 27264 19264 28641 19292
rect 27157 19255 27215 19261
rect 28629 19261 28641 19264
rect 28675 19261 28687 19295
rect 28629 19255 28687 19261
rect 28718 19252 28724 19304
rect 28776 19252 28782 19304
rect 28997 19295 29055 19301
rect 28997 19261 29009 19295
rect 29043 19261 29055 19295
rect 28997 19255 29055 19261
rect 29012 19224 29040 19255
rect 29178 19252 29184 19304
rect 29236 19292 29242 19304
rect 29273 19295 29331 19301
rect 29273 19292 29285 19295
rect 29236 19264 29285 19292
rect 29236 19252 29242 19264
rect 29273 19261 29285 19264
rect 29319 19261 29331 19295
rect 29273 19255 29331 19261
rect 30558 19252 30564 19304
rect 30616 19252 30622 19304
rect 29454 19224 29460 19236
rect 26292 19196 27016 19224
rect 28644 19196 29460 19224
rect 26292 19184 26298 19196
rect 28644 19168 28672 19196
rect 29454 19184 29460 19196
rect 29512 19184 29518 19236
rect 29638 19184 29644 19236
rect 29696 19224 29702 19236
rect 29917 19227 29975 19233
rect 29917 19224 29929 19227
rect 29696 19196 29929 19224
rect 29696 19184 29702 19196
rect 29917 19193 29929 19196
rect 29963 19224 29975 19227
rect 29963 19196 30236 19224
rect 29963 19193 29975 19196
rect 29917 19187 29975 19193
rect 30208 19168 30236 19196
rect 23845 19159 23903 19165
rect 23845 19125 23857 19159
rect 23891 19125 23903 19159
rect 23845 19119 23903 19125
rect 25130 19116 25136 19168
rect 25188 19165 25194 19168
rect 25188 19119 25197 19165
rect 25188 19116 25194 19119
rect 26510 19116 26516 19168
rect 26568 19116 26574 19168
rect 26694 19116 26700 19168
rect 26752 19156 26758 19168
rect 28261 19159 28319 19165
rect 28261 19156 28273 19159
rect 26752 19128 28273 19156
rect 26752 19116 26758 19128
rect 28261 19125 28273 19128
rect 28307 19125 28319 19159
rect 28261 19119 28319 19125
rect 28626 19116 28632 19168
rect 28684 19116 28690 19168
rect 30098 19116 30104 19168
rect 30156 19116 30162 19168
rect 30190 19116 30196 19168
rect 30248 19116 30254 19168
rect 30374 19116 30380 19168
rect 30432 19116 30438 19168
rect 552 19066 31072 19088
rect 552 19014 7988 19066
rect 8040 19014 8052 19066
rect 8104 19014 8116 19066
rect 8168 19014 8180 19066
rect 8232 19014 8244 19066
rect 8296 19014 15578 19066
rect 15630 19014 15642 19066
rect 15694 19014 15706 19066
rect 15758 19014 15770 19066
rect 15822 19014 15834 19066
rect 15886 19014 23168 19066
rect 23220 19014 23232 19066
rect 23284 19014 23296 19066
rect 23348 19014 23360 19066
rect 23412 19014 23424 19066
rect 23476 19014 30758 19066
rect 30810 19014 30822 19066
rect 30874 19014 30886 19066
rect 30938 19014 30950 19066
rect 31002 19014 31014 19066
rect 31066 19014 31072 19066
rect 552 18992 31072 19014
rect 845 18955 903 18961
rect 845 18921 857 18955
rect 891 18952 903 18955
rect 891 18924 4200 18952
rect 891 18921 903 18924
rect 845 18915 903 18921
rect 1210 18844 1216 18896
rect 1268 18844 1274 18896
rect 1302 18844 1308 18896
rect 1360 18884 1366 18896
rect 1397 18887 1455 18893
rect 1397 18884 1409 18887
rect 1360 18856 1409 18884
rect 1360 18844 1366 18856
rect 1397 18853 1409 18856
rect 1443 18884 1455 18887
rect 4172 18884 4200 18924
rect 4246 18912 4252 18964
rect 4304 18912 4310 18964
rect 6270 18952 6276 18964
rect 5460 18924 6276 18952
rect 4614 18884 4620 18896
rect 1443 18856 1900 18884
rect 4172 18856 4620 18884
rect 1443 18853 1455 18856
rect 1397 18847 1455 18853
rect 1026 18776 1032 18828
rect 1084 18776 1090 18828
rect 1118 18776 1124 18828
rect 1176 18776 1182 18828
rect 1228 18816 1256 18844
rect 1765 18819 1823 18825
rect 1765 18816 1777 18819
rect 1228 18788 1777 18816
rect 1765 18785 1777 18788
rect 1811 18785 1823 18819
rect 1872 18816 1900 18856
rect 4614 18844 4620 18856
rect 4672 18844 4678 18896
rect 4706 18844 4712 18896
rect 4764 18844 4770 18896
rect 5460 18893 5488 18924
rect 6270 18912 6276 18924
rect 6328 18952 6334 18964
rect 9131 18955 9189 18961
rect 9131 18952 9143 18955
rect 6328 18924 9143 18952
rect 6328 18912 6334 18924
rect 9131 18921 9143 18924
rect 9177 18952 9189 18955
rect 9306 18952 9312 18964
rect 9177 18924 9312 18952
rect 9177 18921 9189 18924
rect 9131 18915 9189 18921
rect 9306 18912 9312 18924
rect 9364 18952 9370 18964
rect 10689 18955 10747 18961
rect 9364 18924 10088 18952
rect 9364 18912 9370 18924
rect 5445 18887 5503 18893
rect 5445 18853 5457 18887
rect 5491 18853 5503 18887
rect 5445 18847 5503 18853
rect 7650 18844 7656 18896
rect 7708 18884 7714 18896
rect 8021 18887 8079 18893
rect 7708 18856 7880 18884
rect 7708 18844 7714 18856
rect 2736 18819 2794 18825
rect 2736 18816 2748 18819
rect 1872 18788 2748 18816
rect 1765 18779 1823 18785
rect 2736 18785 2748 18788
rect 2782 18816 2794 18819
rect 3510 18816 3516 18828
rect 2782 18788 3516 18816
rect 2782 18785 2794 18788
rect 2736 18779 2794 18785
rect 1136 18748 1164 18776
rect 1578 18748 1584 18760
rect 1136 18720 1584 18748
rect 1578 18708 1584 18720
rect 1636 18708 1642 18760
rect 1780 18748 1808 18779
rect 3510 18776 3516 18788
rect 3568 18776 3574 18828
rect 3786 18776 3792 18828
rect 3844 18816 3850 18828
rect 5169 18819 5227 18825
rect 5169 18816 5181 18819
rect 3844 18788 5181 18816
rect 3844 18776 3850 18788
rect 5169 18785 5181 18788
rect 5215 18816 5227 18819
rect 5350 18816 5356 18828
rect 5215 18788 5356 18816
rect 5215 18785 5227 18788
rect 5169 18779 5227 18785
rect 5350 18776 5356 18788
rect 5408 18776 5414 18828
rect 6641 18819 6699 18825
rect 5828 18788 6598 18816
rect 2406 18748 2412 18760
rect 1780 18720 2412 18748
rect 2406 18708 2412 18720
rect 2464 18708 2470 18760
rect 2872 18753 2930 18759
rect 2872 18719 2884 18753
rect 2918 18748 2930 18753
rect 2958 18748 2964 18760
rect 2918 18720 2964 18748
rect 2918 18719 2930 18720
rect 2872 18713 2930 18719
rect 2958 18708 2964 18720
rect 3016 18708 3022 18760
rect 3145 18751 3203 18757
rect 3145 18717 3157 18751
rect 3191 18748 3203 18751
rect 5534 18748 5540 18760
rect 3191 18720 5540 18748
rect 3191 18717 3203 18720
rect 3145 18711 3203 18717
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 842 18640 848 18692
rect 900 18680 906 18692
rect 1949 18683 2007 18689
rect 1949 18680 1961 18683
rect 900 18652 1961 18680
rect 900 18640 906 18652
rect 1949 18649 1961 18652
rect 1995 18649 2007 18683
rect 5828 18680 5856 18788
rect 6270 18757 6276 18760
rect 5905 18751 5963 18757
rect 5905 18717 5917 18751
rect 5951 18717 5963 18751
rect 5905 18711 5963 18717
rect 6232 18751 6276 18757
rect 6232 18717 6244 18751
rect 6232 18711 6276 18717
rect 1949 18643 2007 18649
rect 4816 18652 5856 18680
rect 1964 18612 1992 18643
rect 3878 18612 3884 18624
rect 1964 18584 3884 18612
rect 3878 18572 3884 18584
rect 3936 18572 3942 18624
rect 4062 18572 4068 18624
rect 4120 18612 4126 18624
rect 4816 18621 4844 18652
rect 4801 18615 4859 18621
rect 4801 18612 4813 18615
rect 4120 18584 4813 18612
rect 4120 18572 4126 18584
rect 4801 18581 4813 18584
rect 4847 18581 4859 18615
rect 5920 18612 5948 18711
rect 6270 18708 6276 18711
rect 6328 18708 6334 18760
rect 6362 18708 6368 18760
rect 6420 18708 6426 18760
rect 6570 18748 6598 18788
rect 6641 18785 6653 18819
rect 6687 18816 6699 18819
rect 7742 18816 7748 18828
rect 6687 18788 7748 18816
rect 6687 18785 6699 18788
rect 6641 18779 6699 18785
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 7852 18816 7880 18856
rect 8021 18853 8033 18887
rect 8067 18884 8079 18887
rect 8754 18884 8760 18896
rect 8067 18856 8760 18884
rect 8067 18853 8079 18856
rect 8021 18847 8079 18853
rect 8754 18844 8760 18856
rect 8812 18844 8818 18896
rect 10060 18884 10088 18924
rect 10689 18921 10701 18955
rect 10735 18952 10747 18955
rect 13170 18952 13176 18964
rect 10735 18924 13176 18952
rect 10735 18921 10747 18924
rect 10689 18915 10747 18921
rect 13170 18912 13176 18924
rect 13228 18912 13234 18964
rect 13446 18912 13452 18964
rect 13504 18952 13510 18964
rect 14182 18952 14188 18964
rect 13504 18924 14188 18952
rect 13504 18912 13510 18924
rect 14182 18912 14188 18924
rect 14240 18912 14246 18964
rect 15286 18952 15292 18964
rect 14384 18924 15292 18952
rect 14384 18884 14412 18924
rect 15286 18912 15292 18924
rect 15344 18912 15350 18964
rect 15841 18955 15899 18961
rect 15841 18921 15853 18955
rect 15887 18952 15899 18955
rect 16206 18952 16212 18964
rect 15887 18924 16212 18952
rect 15887 18921 15899 18924
rect 15841 18915 15899 18921
rect 16206 18912 16212 18924
rect 16264 18912 16270 18964
rect 18046 18952 18052 18964
rect 16500 18924 18052 18952
rect 16500 18884 16528 18924
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 21453 18955 21511 18961
rect 21453 18952 21465 18955
rect 20548 18924 21465 18952
rect 10060 18856 11008 18884
rect 8205 18819 8263 18825
rect 8205 18816 8217 18819
rect 7852 18788 8217 18816
rect 8205 18785 8217 18788
rect 8251 18785 8263 18819
rect 8205 18779 8263 18785
rect 8294 18776 8300 18828
rect 8352 18816 8358 18828
rect 8573 18819 8631 18825
rect 8573 18816 8585 18819
rect 8352 18788 8585 18816
rect 8352 18776 8358 18788
rect 8573 18785 8585 18788
rect 8619 18816 8631 18819
rect 8938 18816 8944 18828
rect 8619 18788 8944 18816
rect 8619 18785 8631 18788
rect 8573 18779 8631 18785
rect 8938 18776 8944 18788
rect 8996 18776 9002 18828
rect 10502 18816 10508 18828
rect 9324 18788 10508 18816
rect 8386 18748 8392 18760
rect 6570 18720 8392 18748
rect 8386 18708 8392 18720
rect 8444 18708 8450 18760
rect 8478 18708 8484 18760
rect 8536 18748 8542 18760
rect 8665 18751 8723 18757
rect 8665 18748 8677 18751
rect 8536 18720 8677 18748
rect 8536 18708 8542 18720
rect 8665 18717 8677 18720
rect 8711 18748 8723 18751
rect 9030 18748 9036 18760
rect 8711 18720 9036 18748
rect 8711 18717 8723 18720
rect 8665 18711 8723 18717
rect 9030 18708 9036 18720
rect 9088 18708 9094 18760
rect 9171 18751 9229 18757
rect 9171 18717 9183 18751
rect 9217 18748 9229 18751
rect 9324 18748 9352 18788
rect 10502 18776 10508 18788
rect 10560 18776 10566 18828
rect 9217 18720 9352 18748
rect 9401 18751 9459 18757
rect 9217 18717 9229 18720
rect 9171 18711 9229 18717
rect 9401 18717 9413 18751
rect 9447 18748 9459 18751
rect 10870 18748 10876 18760
rect 9447 18720 10876 18748
rect 9447 18717 9459 18720
rect 9401 18711 9459 18717
rect 10870 18708 10876 18720
rect 10928 18708 10934 18760
rect 10980 18748 11008 18856
rect 14052 18856 14412 18884
rect 16408 18856 16528 18884
rect 11146 18776 11152 18828
rect 11204 18776 11210 18828
rect 11238 18776 11244 18828
rect 11296 18816 11302 18828
rect 11333 18819 11391 18825
rect 11333 18816 11345 18819
rect 11296 18788 11345 18816
rect 11296 18776 11302 18788
rect 11333 18785 11345 18788
rect 11379 18785 11391 18819
rect 14052 18816 14080 18856
rect 11333 18779 11391 18785
rect 12452 18788 14080 18816
rect 11422 18748 11428 18760
rect 10980 18720 11428 18748
rect 11422 18708 11428 18720
rect 11480 18708 11486 18760
rect 11698 18708 11704 18760
rect 11756 18748 11762 18760
rect 12158 18757 12164 18760
rect 11793 18751 11851 18757
rect 11793 18748 11805 18751
rect 11756 18720 11805 18748
rect 11756 18708 11762 18720
rect 11793 18717 11805 18720
rect 11839 18717 11851 18751
rect 11793 18711 11851 18717
rect 12120 18751 12164 18757
rect 12120 18717 12132 18751
rect 12120 18711 12164 18717
rect 12158 18708 12164 18711
rect 12216 18708 12222 18760
rect 12299 18751 12357 18757
rect 12299 18717 12311 18751
rect 12345 18748 12357 18751
rect 12452 18748 12480 18788
rect 14182 18776 14188 18828
rect 14240 18776 14246 18828
rect 14277 18819 14335 18825
rect 14277 18785 14289 18819
rect 14323 18816 14335 18819
rect 14642 18816 14648 18828
rect 14323 18788 14648 18816
rect 14323 18785 14335 18788
rect 14277 18779 14335 18785
rect 14642 18776 14648 18788
rect 14700 18776 14706 18828
rect 16022 18776 16028 18828
rect 16080 18816 16086 18828
rect 16408 18825 16436 18856
rect 19978 18844 19984 18896
rect 20036 18884 20042 18896
rect 20548 18893 20576 18924
rect 21453 18921 21465 18924
rect 21499 18921 21511 18955
rect 21453 18915 21511 18921
rect 22186 18912 22192 18964
rect 22244 18952 22250 18964
rect 22379 18955 22437 18961
rect 22379 18952 22391 18955
rect 22244 18924 22391 18952
rect 22244 18912 22250 18924
rect 22379 18921 22391 18924
rect 22425 18952 22437 18955
rect 22425 18924 23428 18952
rect 22425 18921 22437 18924
rect 22379 18915 22437 18921
rect 20533 18887 20591 18893
rect 20533 18884 20545 18887
rect 20036 18856 20545 18884
rect 20036 18844 20042 18856
rect 20533 18853 20545 18856
rect 20579 18853 20591 18887
rect 23400 18884 23428 18924
rect 23474 18912 23480 18964
rect 23532 18952 23538 18964
rect 23842 18952 23848 18964
rect 23532 18924 23848 18952
rect 23532 18912 23538 18924
rect 23842 18912 23848 18924
rect 23900 18952 23906 18964
rect 24394 18952 24400 18964
rect 23900 18924 24400 18952
rect 23900 18912 23906 18924
rect 24394 18912 24400 18924
rect 24452 18912 24458 18964
rect 24486 18912 24492 18964
rect 24544 18952 24550 18964
rect 24587 18955 24645 18961
rect 24587 18952 24599 18955
rect 24544 18924 24599 18952
rect 24544 18912 24550 18924
rect 24587 18921 24599 18924
rect 24633 18952 24645 18955
rect 24633 18924 25544 18952
rect 24633 18921 24645 18924
rect 24587 18915 24645 18921
rect 25516 18884 25544 18924
rect 25682 18912 25688 18964
rect 25740 18952 25746 18964
rect 25961 18955 26019 18961
rect 25961 18952 25973 18955
rect 25740 18924 25973 18952
rect 25740 18912 25746 18924
rect 25961 18921 25973 18924
rect 26007 18921 26019 18955
rect 26786 18952 26792 18964
rect 25961 18915 26019 18921
rect 26068 18924 26792 18952
rect 26068 18884 26096 18924
rect 26786 18912 26792 18924
rect 26844 18952 26850 18964
rect 26887 18955 26945 18961
rect 26887 18952 26899 18955
rect 26844 18924 26899 18952
rect 26844 18912 26850 18924
rect 26887 18921 26899 18924
rect 26933 18921 26945 18955
rect 26887 18915 26945 18921
rect 30374 18912 30380 18964
rect 30432 18912 30438 18964
rect 30466 18912 30472 18964
rect 30524 18912 30530 18964
rect 30392 18884 30420 18912
rect 23400 18856 24256 18884
rect 25516 18856 26096 18884
rect 27816 18856 30420 18884
rect 20533 18847 20591 18853
rect 16393 18819 16451 18825
rect 16393 18816 16405 18819
rect 16080 18788 16405 18816
rect 16080 18776 16086 18788
rect 16393 18785 16405 18788
rect 16439 18785 16451 18819
rect 16393 18779 16451 18785
rect 16485 18819 16543 18825
rect 16485 18785 16497 18819
rect 16531 18816 16543 18819
rect 17221 18819 17279 18825
rect 16531 18788 17172 18816
rect 16531 18785 16543 18788
rect 16485 18779 16543 18785
rect 12345 18720 12480 18748
rect 12345 18717 12357 18720
rect 12299 18711 12357 18717
rect 12526 18708 12532 18760
rect 12584 18708 12590 18760
rect 14458 18708 14464 18760
rect 14516 18748 14522 18760
rect 14553 18751 14611 18757
rect 14553 18748 14565 18751
rect 14516 18720 14565 18748
rect 14516 18708 14522 18720
rect 14553 18717 14565 18720
rect 14599 18748 14611 18751
rect 16206 18748 16212 18760
rect 14599 18720 16212 18748
rect 14599 18717 14611 18720
rect 14553 18711 14611 18717
rect 16206 18708 16212 18720
rect 16264 18708 16270 18760
rect 16298 18708 16304 18760
rect 16356 18748 16362 18760
rect 16500 18748 16528 18779
rect 16356 18720 16528 18748
rect 16356 18708 16362 18720
rect 16850 18708 16856 18760
rect 16908 18748 16914 18760
rect 16945 18751 17003 18757
rect 16945 18748 16957 18751
rect 16908 18720 16957 18748
rect 16908 18708 16914 18720
rect 16945 18717 16957 18720
rect 16991 18717 17003 18751
rect 17144 18748 17172 18788
rect 17221 18785 17233 18819
rect 17267 18816 17279 18819
rect 17494 18816 17500 18828
rect 17267 18788 17500 18816
rect 17267 18785 17279 18788
rect 17221 18779 17279 18785
rect 17494 18776 17500 18788
rect 17552 18776 17558 18828
rect 18601 18819 18659 18825
rect 18601 18785 18613 18819
rect 18647 18816 18659 18819
rect 18969 18819 19027 18825
rect 18969 18816 18981 18819
rect 18647 18788 18981 18816
rect 18647 18785 18659 18788
rect 18601 18779 18659 18785
rect 18969 18785 18981 18788
rect 19015 18785 19027 18819
rect 18969 18779 19027 18785
rect 21361 18819 21419 18825
rect 21361 18785 21373 18819
rect 21407 18785 21419 18819
rect 21361 18779 21419 18785
rect 18138 18748 18144 18760
rect 17144 18720 18144 18748
rect 16945 18711 17003 18717
rect 18138 18708 18144 18720
rect 18196 18708 18202 18760
rect 18690 18708 18696 18760
rect 18748 18748 18754 18760
rect 20809 18751 20867 18757
rect 20809 18748 20821 18751
rect 18748 18720 20821 18748
rect 18748 18708 18754 18720
rect 20809 18717 20821 18720
rect 20855 18717 20867 18751
rect 20809 18711 20867 18717
rect 7558 18640 7564 18692
rect 7616 18680 7622 18692
rect 7616 18652 8432 18680
rect 7616 18640 7622 18652
rect 6086 18612 6092 18624
rect 5920 18584 6092 18612
rect 4801 18575 4859 18581
rect 6086 18572 6092 18584
rect 6144 18612 6150 18624
rect 8202 18612 8208 18624
rect 6144 18584 8208 18612
rect 6144 18572 6150 18584
rect 8202 18572 8208 18584
rect 8260 18572 8266 18624
rect 8404 18612 8432 18652
rect 10778 18640 10784 18692
rect 10836 18640 10842 18692
rect 15378 18640 15384 18692
rect 15436 18680 15442 18692
rect 16761 18683 16819 18689
rect 16761 18680 16773 18683
rect 15436 18652 16773 18680
rect 15436 18640 15442 18652
rect 16761 18649 16773 18652
rect 16807 18649 16819 18683
rect 21376 18680 21404 18779
rect 21818 18776 21824 18828
rect 21876 18816 21882 18828
rect 21913 18819 21971 18825
rect 21913 18816 21925 18819
rect 21876 18788 21925 18816
rect 21876 18776 21882 18788
rect 21913 18785 21925 18788
rect 21959 18816 21971 18819
rect 24228 18816 24256 18856
rect 24394 18816 24400 18828
rect 21959 18788 24164 18816
rect 24228 18788 24400 18816
rect 21959 18785 21971 18788
rect 21913 18779 21971 18785
rect 22376 18753 22434 18759
rect 22376 18719 22388 18753
rect 22422 18748 22434 18753
rect 22462 18748 22468 18760
rect 22422 18720 22468 18748
rect 22422 18719 22434 18720
rect 22376 18713 22434 18719
rect 22462 18708 22468 18720
rect 22520 18708 22526 18760
rect 22646 18708 22652 18760
rect 22704 18708 22710 18760
rect 24136 18757 24164 18788
rect 24394 18776 24400 18788
rect 24452 18776 24458 18828
rect 24857 18819 24915 18825
rect 24504 18788 24808 18816
rect 24121 18751 24179 18757
rect 24121 18717 24133 18751
rect 24167 18748 24179 18751
rect 24504 18748 24532 18788
rect 24670 18757 24676 18760
rect 24167 18720 24532 18748
rect 24627 18751 24676 18757
rect 24167 18717 24179 18720
rect 24121 18711 24179 18717
rect 24627 18717 24639 18751
rect 24673 18717 24676 18751
rect 24627 18711 24676 18717
rect 24670 18708 24676 18711
rect 24728 18708 24734 18760
rect 24780 18748 24808 18788
rect 24857 18785 24869 18819
rect 24903 18816 24915 18819
rect 27816 18816 27844 18856
rect 24903 18788 27844 18816
rect 28629 18819 28687 18825
rect 24903 18785 24915 18788
rect 24857 18779 24915 18785
rect 28629 18785 28641 18819
rect 28675 18785 28687 18819
rect 28629 18779 28687 18785
rect 26326 18748 26332 18760
rect 24780 18720 26332 18748
rect 26326 18708 26332 18720
rect 26384 18748 26390 18760
rect 26421 18751 26479 18757
rect 26421 18748 26433 18751
rect 26384 18720 26433 18748
rect 26384 18708 26390 18720
rect 26421 18717 26433 18720
rect 26467 18717 26479 18751
rect 26421 18711 26479 18717
rect 26927 18751 26985 18757
rect 26927 18717 26939 18751
rect 26973 18748 26985 18751
rect 27062 18748 27068 18760
rect 26973 18720 27068 18748
rect 26973 18717 26985 18720
rect 26927 18711 26985 18717
rect 27062 18708 27068 18720
rect 27120 18708 27126 18760
rect 27157 18751 27215 18757
rect 27157 18717 27169 18751
rect 27203 18748 27215 18751
rect 27203 18720 28580 18748
rect 27203 18717 27215 18720
rect 27157 18711 27215 18717
rect 21376 18652 21864 18680
rect 16761 18643 16819 18649
rect 9766 18612 9772 18624
rect 8404 18584 9772 18612
rect 9766 18572 9772 18584
rect 9824 18572 9830 18624
rect 10796 18612 10824 18640
rect 10965 18615 11023 18621
rect 10965 18612 10977 18615
rect 10796 18584 10977 18612
rect 10965 18581 10977 18584
rect 11011 18581 11023 18615
rect 10965 18575 11023 18581
rect 11054 18572 11060 18624
rect 11112 18612 11118 18624
rect 11425 18615 11483 18621
rect 11425 18612 11437 18615
rect 11112 18584 11437 18612
rect 11112 18572 11118 18584
rect 11425 18581 11437 18584
rect 11471 18581 11483 18615
rect 11425 18575 11483 18581
rect 12986 18572 12992 18624
rect 13044 18612 13050 18624
rect 13633 18615 13691 18621
rect 13633 18612 13645 18615
rect 13044 18584 13645 18612
rect 13044 18572 13050 18584
rect 13633 18581 13645 18584
rect 13679 18581 13691 18615
rect 13633 18575 13691 18581
rect 14001 18615 14059 18621
rect 14001 18581 14013 18615
rect 14047 18612 14059 18615
rect 14550 18612 14556 18624
rect 14047 18584 14556 18612
rect 14047 18581 14059 18584
rect 14001 18575 14059 18581
rect 14550 18572 14556 18584
rect 14608 18572 14614 18624
rect 19794 18572 19800 18624
rect 19852 18612 19858 18624
rect 20073 18615 20131 18621
rect 20073 18612 20085 18615
rect 19852 18584 20085 18612
rect 19852 18572 19858 18584
rect 20073 18581 20085 18584
rect 20119 18581 20131 18615
rect 20073 18575 20131 18581
rect 20254 18572 20260 18624
rect 20312 18612 20318 18624
rect 21726 18612 21732 18624
rect 20312 18584 21732 18612
rect 20312 18572 20318 18584
rect 21726 18572 21732 18584
rect 21784 18572 21790 18624
rect 21836 18612 21864 18652
rect 26142 18640 26148 18692
rect 26200 18640 26206 18692
rect 22278 18612 22284 18624
rect 21836 18584 22284 18612
rect 22278 18572 22284 18584
rect 22336 18612 22342 18624
rect 23474 18612 23480 18624
rect 22336 18584 23480 18612
rect 22336 18572 22342 18584
rect 23474 18572 23480 18584
rect 23532 18572 23538 18624
rect 23937 18615 23995 18621
rect 23937 18581 23949 18615
rect 23983 18612 23995 18615
rect 24394 18612 24400 18624
rect 23983 18584 24400 18612
rect 23983 18581 23995 18584
rect 23937 18575 23995 18581
rect 24394 18572 24400 18584
rect 24452 18572 24458 18624
rect 24486 18572 24492 18624
rect 24544 18612 24550 18624
rect 26160 18612 26188 18640
rect 24544 18584 26188 18612
rect 24544 18572 24550 18584
rect 27062 18572 27068 18624
rect 27120 18612 27126 18624
rect 27614 18612 27620 18624
rect 27120 18584 27620 18612
rect 27120 18572 27126 18584
rect 27614 18572 27620 18584
rect 27672 18572 27678 18624
rect 27798 18572 27804 18624
rect 27856 18612 27862 18624
rect 28261 18615 28319 18621
rect 28261 18612 28273 18615
rect 27856 18584 28273 18612
rect 27856 18572 27862 18584
rect 28261 18581 28273 18584
rect 28307 18581 28319 18615
rect 28552 18612 28580 18720
rect 28644 18692 28672 18779
rect 28810 18776 28816 18828
rect 28868 18816 28874 18828
rect 28905 18819 28963 18825
rect 28905 18816 28917 18819
rect 28868 18788 28917 18816
rect 28868 18776 28874 18788
rect 28905 18785 28917 18788
rect 28951 18816 28963 18819
rect 29178 18816 29184 18828
rect 28951 18788 29184 18816
rect 28951 18785 28963 18788
rect 28905 18779 28963 18785
rect 29178 18776 29184 18788
rect 29236 18776 29242 18828
rect 28626 18640 28632 18692
rect 28684 18640 28690 18692
rect 30190 18640 30196 18692
rect 30248 18640 30254 18692
rect 30374 18612 30380 18624
rect 28552 18584 30380 18612
rect 28261 18575 28319 18581
rect 30374 18572 30380 18584
rect 30432 18572 30438 18624
rect 552 18522 30912 18544
rect 552 18470 4193 18522
rect 4245 18470 4257 18522
rect 4309 18470 4321 18522
rect 4373 18470 4385 18522
rect 4437 18470 4449 18522
rect 4501 18470 11783 18522
rect 11835 18470 11847 18522
rect 11899 18470 11911 18522
rect 11963 18470 11975 18522
rect 12027 18470 12039 18522
rect 12091 18470 19373 18522
rect 19425 18470 19437 18522
rect 19489 18470 19501 18522
rect 19553 18470 19565 18522
rect 19617 18470 19629 18522
rect 19681 18470 26963 18522
rect 27015 18470 27027 18522
rect 27079 18470 27091 18522
rect 27143 18470 27155 18522
rect 27207 18470 27219 18522
rect 27271 18470 30912 18522
rect 552 18448 30912 18470
rect 2406 18368 2412 18420
rect 2464 18408 2470 18420
rect 2464 18380 2774 18408
rect 2464 18368 2470 18380
rect 2746 18340 2774 18380
rect 2958 18368 2964 18420
rect 3016 18368 3022 18420
rect 3326 18368 3332 18420
rect 3384 18368 3390 18420
rect 3510 18368 3516 18420
rect 3568 18408 3574 18420
rect 5718 18408 5724 18420
rect 3568 18380 5724 18408
rect 3568 18368 3574 18380
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 5905 18411 5963 18417
rect 5905 18377 5917 18411
rect 5951 18408 5963 18411
rect 6362 18408 6368 18420
rect 5951 18380 6368 18408
rect 5951 18377 5963 18380
rect 5905 18371 5963 18377
rect 6362 18368 6368 18380
rect 6420 18368 6426 18420
rect 6454 18368 6460 18420
rect 6512 18408 6518 18420
rect 10686 18408 10692 18420
rect 6512 18380 10692 18408
rect 6512 18368 6518 18380
rect 10686 18368 10692 18380
rect 10744 18368 10750 18420
rect 12618 18368 12624 18420
rect 12676 18368 12682 18420
rect 12728 18380 16804 18408
rect 3344 18340 3372 18368
rect 2746 18312 3372 18340
rect 12250 18300 12256 18352
rect 12308 18340 12314 18352
rect 12728 18340 12756 18380
rect 12308 18312 12756 18340
rect 16776 18340 16804 18380
rect 17218 18368 17224 18420
rect 17276 18368 17282 18420
rect 17494 18368 17500 18420
rect 17552 18408 17558 18420
rect 22189 18411 22247 18417
rect 22189 18408 22201 18411
rect 17552 18380 22201 18408
rect 17552 18368 17558 18380
rect 22189 18377 22201 18380
rect 22235 18377 22247 18411
rect 22189 18371 22247 18377
rect 22738 18368 22744 18420
rect 22796 18368 22802 18420
rect 22925 18411 22983 18417
rect 22925 18377 22937 18411
rect 22971 18408 22983 18411
rect 23474 18408 23480 18420
rect 22971 18380 23480 18408
rect 22971 18377 22983 18380
rect 22925 18371 22983 18377
rect 23474 18368 23480 18380
rect 23532 18368 23538 18420
rect 23750 18368 23756 18420
rect 23808 18408 23814 18420
rect 23808 18380 27844 18408
rect 23808 18368 23814 18380
rect 18230 18340 18236 18352
rect 16776 18312 18236 18340
rect 12308 18300 12314 18312
rect 18230 18300 18236 18312
rect 18288 18300 18294 18352
rect 19886 18340 19892 18352
rect 19812 18312 19892 18340
rect 842 18232 848 18284
rect 900 18272 906 18284
rect 937 18275 995 18281
rect 937 18272 949 18275
rect 900 18244 949 18272
rect 900 18232 906 18244
rect 937 18241 949 18244
rect 983 18241 995 18275
rect 937 18235 995 18241
rect 1443 18275 1501 18281
rect 1443 18241 1455 18275
rect 1489 18272 1501 18275
rect 3142 18272 3148 18284
rect 1489 18244 3148 18272
rect 1489 18241 1501 18244
rect 1443 18235 1501 18241
rect 3142 18232 3148 18244
rect 3200 18232 3206 18284
rect 4062 18272 4068 18284
rect 3344 18244 4068 18272
rect 1673 18207 1731 18213
rect 1673 18173 1685 18207
rect 1719 18204 1731 18207
rect 2406 18204 2412 18216
rect 1719 18176 2412 18204
rect 1719 18173 1731 18176
rect 1673 18167 1731 18173
rect 2406 18164 2412 18176
rect 2464 18164 2470 18216
rect 3234 18164 3240 18216
rect 3292 18204 3298 18216
rect 3344 18213 3372 18244
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 4246 18281 4252 18284
rect 4208 18275 4252 18281
rect 4208 18241 4220 18275
rect 4208 18235 4252 18241
rect 4246 18232 4252 18235
rect 4304 18232 4310 18284
rect 4338 18232 4344 18284
rect 4396 18272 4402 18284
rect 4617 18275 4675 18281
rect 4396 18244 4441 18272
rect 4396 18232 4402 18244
rect 4617 18241 4629 18275
rect 4663 18272 4675 18275
rect 5350 18272 5356 18284
rect 4663 18244 5356 18272
rect 4663 18241 4675 18244
rect 4617 18235 4675 18241
rect 5350 18232 5356 18244
rect 5408 18232 5414 18284
rect 5626 18232 5632 18284
rect 5684 18272 5690 18284
rect 6552 18275 6610 18281
rect 6552 18272 6564 18275
rect 5684 18244 6564 18272
rect 5684 18232 5690 18244
rect 6552 18241 6564 18244
rect 6598 18241 6610 18275
rect 6552 18235 6610 18241
rect 8386 18232 8392 18284
rect 8444 18272 8450 18284
rect 8570 18272 8576 18284
rect 8444 18244 8576 18272
rect 8444 18232 8450 18244
rect 8570 18232 8576 18244
rect 8628 18232 8634 18284
rect 8754 18232 8760 18284
rect 8812 18272 8818 18284
rect 9036 18275 9094 18281
rect 9036 18272 9048 18275
rect 8812 18244 9048 18272
rect 8812 18232 8818 18244
rect 9036 18241 9048 18244
rect 9082 18241 9094 18275
rect 9036 18235 9094 18241
rect 9122 18232 9128 18284
rect 9180 18272 9186 18284
rect 10689 18275 10747 18281
rect 9180 18244 9444 18272
rect 9180 18232 9186 18244
rect 3329 18207 3387 18213
rect 3329 18204 3341 18207
rect 3292 18176 3341 18204
rect 3292 18164 3298 18176
rect 3329 18173 3341 18176
rect 3375 18173 3387 18207
rect 3329 18167 3387 18173
rect 3878 18164 3884 18216
rect 3936 18164 3942 18216
rect 6086 18164 6092 18216
rect 6144 18164 6150 18216
rect 6730 18164 6736 18216
rect 6788 18204 6794 18216
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6788 18176 6837 18204
rect 6788 18164 6794 18176
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 9309 18207 9367 18213
rect 9309 18204 9321 18207
rect 6825 18167 6883 18173
rect 8680 18176 9321 18204
rect 8205 18139 8263 18145
rect 8205 18105 8217 18139
rect 8251 18136 8263 18139
rect 8478 18136 8484 18148
rect 8251 18108 8484 18136
rect 8251 18105 8263 18108
rect 8205 18099 8263 18105
rect 8478 18096 8484 18108
rect 8536 18096 8542 18148
rect 1394 18028 1400 18080
rect 1452 18077 1458 18080
rect 1452 18068 1461 18077
rect 1452 18040 1497 18068
rect 1452 18031 1461 18040
rect 1452 18028 1458 18031
rect 3326 18028 3332 18080
rect 3384 18068 3390 18080
rect 3605 18071 3663 18077
rect 3605 18068 3617 18071
rect 3384 18040 3617 18068
rect 3384 18028 3390 18040
rect 3605 18037 3617 18040
rect 3651 18068 3663 18071
rect 6178 18068 6184 18080
rect 3651 18040 6184 18068
rect 3651 18037 3663 18040
rect 3605 18031 3663 18037
rect 6178 18028 6184 18040
rect 6236 18028 6242 18080
rect 6454 18028 6460 18080
rect 6512 18068 6518 18080
rect 6555 18071 6613 18077
rect 6555 18068 6567 18071
rect 6512 18040 6567 18068
rect 6512 18028 6518 18040
rect 6555 18037 6567 18040
rect 6601 18068 6613 18071
rect 6822 18068 6828 18080
rect 6601 18040 6828 18068
rect 6601 18037 6613 18040
rect 6555 18031 6613 18037
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 8386 18028 8392 18080
rect 8444 18068 8450 18080
rect 8680 18068 8708 18176
rect 9309 18173 9321 18176
rect 9355 18173 9367 18207
rect 9416 18204 9444 18244
rect 10689 18241 10701 18275
rect 10735 18272 10747 18275
rect 11244 18275 11302 18281
rect 11244 18272 11256 18275
rect 10735 18244 11256 18272
rect 10735 18241 10747 18244
rect 10689 18235 10747 18241
rect 11244 18241 11256 18244
rect 11290 18241 11302 18275
rect 11244 18235 11302 18241
rect 11330 18232 11336 18284
rect 11388 18272 11394 18284
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 11388 18244 11529 18272
rect 11388 18232 11394 18244
rect 11517 18241 11529 18244
rect 11563 18241 11575 18275
rect 13722 18272 13728 18284
rect 11517 18235 11575 18241
rect 13372 18244 13728 18272
rect 10778 18204 10784 18216
rect 9416 18176 10784 18204
rect 9309 18167 9367 18173
rect 10778 18164 10784 18176
rect 10836 18164 10842 18216
rect 13372 18213 13400 18244
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 13998 18232 14004 18284
rect 14056 18263 14062 18284
rect 14056 18257 14095 18263
rect 14016 18226 14049 18232
rect 14037 18223 14049 18226
rect 14083 18223 14095 18257
rect 15838 18232 15844 18284
rect 15896 18272 15902 18284
rect 16022 18272 16028 18284
rect 15896 18244 16028 18272
rect 15896 18232 15902 18244
rect 16022 18232 16028 18244
rect 16080 18232 16086 18284
rect 16117 18275 16175 18281
rect 16117 18241 16129 18275
rect 16163 18272 16175 18275
rect 16482 18272 16488 18284
rect 16163 18244 16488 18272
rect 16163 18241 16175 18244
rect 16117 18235 16175 18241
rect 16482 18232 16488 18244
rect 16540 18232 16546 18284
rect 18509 18275 18567 18281
rect 18509 18272 18521 18275
rect 17512 18244 18521 18272
rect 14037 18217 14095 18223
rect 13357 18207 13415 18213
rect 13357 18204 13369 18207
rect 10888 18176 13369 18204
rect 10226 18096 10232 18148
rect 10284 18136 10290 18148
rect 10888 18136 10916 18176
rect 13357 18173 13369 18176
rect 13403 18173 13415 18207
rect 13357 18167 13415 18173
rect 13538 18164 13544 18216
rect 13596 18164 13602 18216
rect 14277 18207 14335 18213
rect 14277 18173 14289 18207
rect 14323 18204 14335 18207
rect 14642 18204 14648 18216
rect 14323 18176 14648 18204
rect 14323 18173 14335 18176
rect 14277 18167 14335 18173
rect 14642 18164 14648 18176
rect 14700 18164 14706 18216
rect 16390 18164 16396 18216
rect 16448 18204 16454 18216
rect 17512 18204 17540 18244
rect 18509 18241 18521 18244
rect 18555 18241 18567 18275
rect 18509 18235 18567 18241
rect 16448 18176 17540 18204
rect 16448 18164 16454 18176
rect 18046 18164 18052 18216
rect 18104 18164 18110 18216
rect 18138 18164 18144 18216
rect 18196 18204 18202 18216
rect 18417 18207 18475 18213
rect 18417 18204 18429 18207
rect 18196 18176 18429 18204
rect 18196 18164 18202 18176
rect 18417 18173 18429 18176
rect 18463 18173 18475 18207
rect 19812 18190 19840 18312
rect 19886 18300 19892 18312
rect 19944 18300 19950 18352
rect 22756 18340 22784 18368
rect 23293 18343 23351 18349
rect 23293 18340 23305 18343
rect 22756 18312 23305 18340
rect 23293 18309 23305 18312
rect 23339 18309 23351 18343
rect 23293 18303 23351 18309
rect 24228 18312 24491 18340
rect 24228 18284 24256 18312
rect 20165 18275 20223 18281
rect 20165 18241 20177 18275
rect 20211 18272 20223 18275
rect 20622 18272 20628 18284
rect 20211 18244 20628 18272
rect 20211 18241 20223 18244
rect 20165 18235 20223 18241
rect 20622 18232 20628 18244
rect 20680 18232 20686 18284
rect 20855 18275 20913 18281
rect 20855 18241 20867 18275
rect 20901 18272 20913 18275
rect 22830 18272 22836 18284
rect 20901 18244 22836 18272
rect 20901 18241 20913 18244
rect 20855 18235 20913 18241
rect 22830 18232 22836 18244
rect 22888 18232 22894 18284
rect 24210 18232 24216 18284
rect 24268 18232 24274 18284
rect 18417 18167 18475 18173
rect 20254 18164 20260 18216
rect 20312 18164 20318 18216
rect 20349 18207 20407 18213
rect 20349 18173 20361 18207
rect 20395 18173 20407 18207
rect 20349 18167 20407 18173
rect 10284 18108 10916 18136
rect 17681 18139 17739 18145
rect 10284 18096 10290 18108
rect 17681 18105 17693 18139
rect 17727 18105 17739 18139
rect 17681 18099 17739 18105
rect 19061 18139 19119 18145
rect 19061 18105 19073 18139
rect 19107 18136 19119 18139
rect 19150 18136 19156 18148
rect 19107 18108 19156 18136
rect 19107 18105 19119 18108
rect 19061 18099 19119 18105
rect 8444 18040 8708 18068
rect 8444 18028 8450 18040
rect 8846 18028 8852 18080
rect 8904 18068 8910 18080
rect 9039 18071 9097 18077
rect 9039 18068 9051 18071
rect 8904 18040 9051 18068
rect 8904 18028 8910 18040
rect 9039 18037 9051 18040
rect 9085 18037 9097 18071
rect 9039 18031 9097 18037
rect 11247 18071 11305 18077
rect 11247 18037 11259 18071
rect 11293 18068 11305 18071
rect 11422 18068 11428 18080
rect 11293 18040 11428 18068
rect 11293 18037 11305 18040
rect 11247 18031 11305 18037
rect 11422 18028 11428 18040
rect 11480 18028 11486 18080
rect 13173 18071 13231 18077
rect 13173 18037 13185 18071
rect 13219 18068 13231 18071
rect 13814 18068 13820 18080
rect 13219 18040 13820 18068
rect 13219 18037 13231 18040
rect 13173 18031 13231 18037
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 14007 18071 14065 18077
rect 14007 18037 14019 18071
rect 14053 18068 14065 18071
rect 15102 18068 15108 18080
rect 14053 18040 15108 18068
rect 14053 18037 14065 18040
rect 14007 18031 14065 18037
rect 15102 18028 15108 18040
rect 15160 18028 15166 18080
rect 15562 18028 15568 18080
rect 15620 18028 15626 18080
rect 16206 18028 16212 18080
rect 16264 18068 16270 18080
rect 17696 18068 17724 18099
rect 19150 18096 19156 18108
rect 19208 18096 19214 18148
rect 19886 18096 19892 18148
rect 19944 18136 19950 18148
rect 20070 18136 20076 18148
rect 19944 18108 20076 18136
rect 19944 18096 19950 18108
rect 20070 18096 20076 18108
rect 20128 18096 20134 18148
rect 20272 18068 20300 18164
rect 20364 18080 20392 18167
rect 20990 18164 20996 18216
rect 21048 18204 21054 18216
rect 21085 18207 21143 18213
rect 21085 18204 21097 18207
rect 21048 18176 21097 18204
rect 21048 18164 21054 18176
rect 21085 18173 21097 18176
rect 21131 18173 21143 18207
rect 21085 18167 21143 18173
rect 22922 18164 22928 18216
rect 22980 18204 22986 18216
rect 23109 18207 23167 18213
rect 23109 18204 23121 18207
rect 22980 18176 23121 18204
rect 22980 18164 22986 18176
rect 23109 18173 23121 18176
rect 23155 18173 23167 18207
rect 23109 18167 23167 18173
rect 23658 18164 23664 18216
rect 23716 18164 23722 18216
rect 24305 18207 24363 18213
rect 24305 18204 24317 18207
rect 23868 18176 24317 18204
rect 22649 18139 22707 18145
rect 22649 18105 22661 18139
rect 22695 18136 22707 18139
rect 23868 18136 23896 18176
rect 24305 18173 24317 18176
rect 24351 18173 24363 18207
rect 24463 18204 24491 18312
rect 24578 18300 24584 18352
rect 24636 18340 24642 18352
rect 27816 18340 27844 18380
rect 28258 18368 28264 18420
rect 28316 18368 28322 18420
rect 30377 18411 30435 18417
rect 30377 18408 30389 18411
rect 28920 18380 30389 18408
rect 28629 18343 28687 18349
rect 28629 18340 28641 18343
rect 24636 18312 24716 18340
rect 27816 18312 28641 18340
rect 24636 18300 24642 18312
rect 24688 18281 24716 18312
rect 28629 18309 28641 18312
rect 28675 18309 28687 18343
rect 28629 18303 28687 18309
rect 24673 18275 24731 18281
rect 24673 18241 24685 18275
rect 24719 18241 24731 18275
rect 24673 18235 24731 18241
rect 24854 18232 24860 18284
rect 24912 18272 24918 18284
rect 25136 18275 25194 18281
rect 25136 18272 25148 18275
rect 24912 18244 25148 18272
rect 24912 18232 24918 18244
rect 25136 18241 25148 18244
rect 25182 18241 25194 18275
rect 26878 18272 26884 18284
rect 25136 18235 25194 18241
rect 25332 18244 26884 18272
rect 24581 18207 24639 18213
rect 24581 18204 24593 18207
rect 24463 18176 24593 18204
rect 24305 18167 24363 18173
rect 24581 18173 24593 18176
rect 24627 18173 24639 18207
rect 25332 18204 25360 18244
rect 26878 18232 26884 18244
rect 26936 18232 26942 18284
rect 27890 18232 27896 18284
rect 27948 18272 27954 18284
rect 28920 18272 28948 18380
rect 30377 18377 30389 18380
rect 30423 18377 30435 18411
rect 30377 18371 30435 18377
rect 27948 18244 28948 18272
rect 27948 18232 27954 18244
rect 24581 18167 24639 18173
rect 24780 18176 25360 18204
rect 22695 18108 23896 18136
rect 22695 18105 22707 18108
rect 22649 18099 22707 18105
rect 23934 18096 23940 18148
rect 23992 18096 23998 18148
rect 24320 18136 24348 18167
rect 24780 18136 24808 18176
rect 25406 18164 25412 18216
rect 25464 18164 25470 18216
rect 26602 18164 26608 18216
rect 26660 18204 26666 18216
rect 27157 18207 27215 18213
rect 27157 18204 27169 18207
rect 26660 18176 27169 18204
rect 26660 18164 26666 18176
rect 27157 18173 27169 18176
rect 27203 18173 27215 18207
rect 27157 18167 27215 18173
rect 28718 18164 28724 18216
rect 28776 18204 28782 18216
rect 28813 18207 28871 18213
rect 28813 18204 28825 18207
rect 28776 18176 28825 18204
rect 28776 18164 28782 18176
rect 28813 18173 28825 18176
rect 28859 18173 28871 18207
rect 28813 18167 28871 18173
rect 28997 18207 29055 18213
rect 28997 18173 29009 18207
rect 29043 18173 29055 18207
rect 28997 18167 29055 18173
rect 24320 18108 24808 18136
rect 28626 18096 28632 18148
rect 28684 18136 28690 18148
rect 29012 18136 29040 18167
rect 29178 18164 29184 18216
rect 29236 18204 29242 18216
rect 29273 18207 29331 18213
rect 29273 18204 29285 18207
rect 29236 18176 29285 18204
rect 29236 18164 29242 18176
rect 29273 18173 29285 18176
rect 29319 18173 29331 18207
rect 29273 18167 29331 18173
rect 29362 18164 29368 18216
rect 29420 18204 29426 18216
rect 30101 18207 30159 18213
rect 30101 18204 30113 18207
rect 29420 18176 30113 18204
rect 29420 18164 29426 18176
rect 30101 18173 30113 18176
rect 30147 18204 30159 18207
rect 30190 18204 30196 18216
rect 30147 18176 30196 18204
rect 30147 18173 30159 18176
rect 30101 18167 30159 18173
rect 30190 18164 30196 18176
rect 30248 18164 30254 18216
rect 30561 18207 30619 18213
rect 30561 18173 30573 18207
rect 30607 18173 30619 18207
rect 30561 18167 30619 18173
rect 30576 18136 30604 18167
rect 28684 18108 29684 18136
rect 28684 18096 28690 18108
rect 29656 18080 29684 18108
rect 29932 18108 30604 18136
rect 29932 18080 29960 18108
rect 16264 18040 20300 18068
rect 16264 18028 16270 18040
rect 20346 18028 20352 18080
rect 20404 18028 20410 18080
rect 20815 18071 20873 18077
rect 20815 18037 20827 18071
rect 20861 18068 20873 18071
rect 21542 18068 21548 18080
rect 20861 18040 21548 18068
rect 20861 18037 20873 18040
rect 20815 18031 20873 18037
rect 21542 18028 21548 18040
rect 21600 18028 21606 18080
rect 21726 18028 21732 18080
rect 21784 18068 21790 18080
rect 23382 18068 23388 18080
rect 21784 18040 23388 18068
rect 21784 18028 21790 18040
rect 23382 18028 23388 18040
rect 23440 18028 23446 18080
rect 23477 18071 23535 18077
rect 23477 18037 23489 18071
rect 23523 18068 23535 18071
rect 24302 18068 24308 18080
rect 23523 18040 24308 18068
rect 23523 18037 23535 18040
rect 23477 18031 23535 18037
rect 24302 18028 24308 18040
rect 24360 18028 24366 18080
rect 24397 18071 24455 18077
rect 24397 18037 24409 18071
rect 24443 18068 24455 18071
rect 24946 18068 24952 18080
rect 24443 18040 24952 18068
rect 24443 18037 24455 18040
rect 24397 18031 24455 18037
rect 24946 18028 24952 18040
rect 25004 18028 25010 18080
rect 25130 18028 25136 18080
rect 25188 18077 25194 18080
rect 25188 18068 25197 18077
rect 25188 18040 25233 18068
rect 25188 18031 25197 18040
rect 25188 18028 25194 18031
rect 26418 18028 26424 18080
rect 26476 18068 26482 18080
rect 26513 18071 26571 18077
rect 26513 18068 26525 18071
rect 26476 18040 26525 18068
rect 26476 18028 26482 18040
rect 26513 18037 26525 18040
rect 26559 18037 26571 18071
rect 26513 18031 26571 18037
rect 29638 18028 29644 18080
rect 29696 18028 29702 18080
rect 29914 18028 29920 18080
rect 29972 18028 29978 18080
rect 30282 18028 30288 18080
rect 30340 18028 30346 18080
rect 552 17978 31072 18000
rect 552 17926 7988 17978
rect 8040 17926 8052 17978
rect 8104 17926 8116 17978
rect 8168 17926 8180 17978
rect 8232 17926 8244 17978
rect 8296 17926 15578 17978
rect 15630 17926 15642 17978
rect 15694 17926 15706 17978
rect 15758 17926 15770 17978
rect 15822 17926 15834 17978
rect 15886 17926 23168 17978
rect 23220 17926 23232 17978
rect 23284 17926 23296 17978
rect 23348 17926 23360 17978
rect 23412 17926 23424 17978
rect 23476 17926 30758 17978
rect 30810 17926 30822 17978
rect 30874 17926 30886 17978
rect 30938 17926 30950 17978
rect 31002 17926 31014 17978
rect 31066 17926 31072 17978
rect 552 17904 31072 17926
rect 1394 17824 1400 17876
rect 1452 17873 1458 17876
rect 1452 17864 1461 17873
rect 1452 17836 2360 17864
rect 1452 17827 1461 17836
rect 1452 17824 1458 17827
rect 2332 17796 2360 17836
rect 2774 17824 2780 17876
rect 2832 17824 2838 17876
rect 3145 17867 3203 17873
rect 3145 17833 3157 17867
rect 3191 17864 3203 17867
rect 3510 17864 3516 17876
rect 3191 17836 3516 17864
rect 3191 17833 3203 17836
rect 3145 17827 3203 17833
rect 3510 17824 3516 17836
rect 3568 17824 3574 17876
rect 3979 17867 4037 17873
rect 3979 17864 3991 17867
rect 3620 17836 3991 17864
rect 3620 17796 3648 17836
rect 3979 17833 3991 17836
rect 4025 17864 4037 17867
rect 4246 17864 4252 17876
rect 4025 17836 4252 17864
rect 4025 17833 4037 17836
rect 3979 17827 4037 17833
rect 4246 17824 4252 17836
rect 4304 17864 4310 17876
rect 4522 17864 4528 17876
rect 4304 17836 4528 17864
rect 4304 17824 4310 17836
rect 4522 17824 4528 17836
rect 4580 17824 4586 17876
rect 6181 17867 6239 17873
rect 6181 17833 6193 17867
rect 6227 17864 6239 17867
rect 8386 17864 8392 17876
rect 6227 17836 8392 17864
rect 6227 17833 6239 17836
rect 6181 17827 6239 17833
rect 8386 17824 8392 17836
rect 8444 17824 8450 17876
rect 10965 17867 11023 17873
rect 8496 17836 10180 17864
rect 2332 17768 3648 17796
rect 5626 17756 5632 17808
rect 5684 17756 5690 17808
rect 8496 17796 8524 17836
rect 5736 17768 6500 17796
rect 842 17688 848 17740
rect 900 17728 906 17740
rect 937 17731 995 17737
rect 937 17728 949 17731
rect 900 17700 949 17728
rect 900 17688 906 17700
rect 937 17697 949 17700
rect 983 17697 995 17731
rect 2958 17728 2964 17740
rect 937 17691 995 17697
rect 1596 17700 2964 17728
rect 1433 17681 1491 17687
rect 1433 17678 1445 17681
rect 1412 17647 1445 17678
rect 1479 17660 1491 17681
rect 1596 17660 1624 17700
rect 2958 17688 2964 17700
rect 3016 17688 3022 17740
rect 3329 17731 3387 17737
rect 3329 17697 3341 17731
rect 3375 17728 3387 17731
rect 3602 17728 3608 17740
rect 3375 17700 3608 17728
rect 3375 17697 3387 17700
rect 3329 17691 3387 17697
rect 3602 17688 3608 17700
rect 3660 17688 3666 17740
rect 4338 17688 4344 17740
rect 4396 17728 4402 17740
rect 4890 17728 4896 17740
rect 4396 17700 4896 17728
rect 4396 17688 4402 17700
rect 4890 17688 4896 17700
rect 4948 17688 4954 17740
rect 3976 17681 4034 17687
rect 1479 17647 1624 17660
rect 1412 17632 1624 17647
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 3418 17660 3424 17672
rect 1719 17632 3424 17660
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 3418 17620 3424 17632
rect 3476 17620 3482 17672
rect 3513 17663 3571 17669
rect 3513 17629 3525 17663
rect 3559 17660 3571 17663
rect 3878 17660 3884 17672
rect 3559 17632 3884 17660
rect 3559 17629 3571 17632
rect 3513 17623 3571 17629
rect 3878 17620 3884 17632
rect 3936 17620 3942 17672
rect 3976 17647 3988 17681
rect 4022 17660 4034 17681
rect 4062 17660 4068 17672
rect 4022 17647 4068 17660
rect 3976 17641 4068 17647
rect 3991 17632 4068 17641
rect 4062 17620 4068 17632
rect 4120 17620 4126 17672
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 5166 17660 5172 17672
rect 4295 17632 5172 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 3786 17484 3792 17536
rect 3844 17524 3850 17536
rect 5736 17524 5764 17768
rect 6089 17731 6147 17737
rect 6089 17697 6101 17731
rect 6135 17728 6147 17731
rect 6270 17728 6276 17740
rect 6135 17700 6276 17728
rect 6135 17697 6147 17700
rect 6089 17691 6147 17697
rect 6270 17688 6276 17700
rect 6328 17688 6334 17740
rect 6362 17688 6368 17740
rect 6420 17688 6426 17740
rect 6472 17728 6500 17768
rect 7852 17768 8524 17796
rect 8573 17799 8631 17805
rect 7852 17728 7880 17768
rect 8573 17765 8585 17799
rect 8619 17796 8631 17799
rect 8754 17796 8760 17808
rect 8619 17768 8760 17796
rect 8619 17765 8631 17768
rect 8573 17759 8631 17765
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 10152 17740 10180 17836
rect 10965 17833 10977 17867
rect 11011 17833 11023 17867
rect 10965 17827 11023 17833
rect 11609 17867 11667 17873
rect 11609 17833 11621 17867
rect 11655 17864 11667 17867
rect 12342 17864 12348 17876
rect 11655 17836 12348 17864
rect 11655 17833 11667 17836
rect 11609 17827 11667 17833
rect 10980 17796 11008 17827
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 16022 17824 16028 17876
rect 16080 17864 16086 17876
rect 16577 17867 16635 17873
rect 16577 17864 16589 17867
rect 16080 17836 16589 17864
rect 16080 17824 16086 17836
rect 16577 17833 16589 17836
rect 16623 17833 16635 17867
rect 16577 17827 16635 17833
rect 16758 17824 16764 17876
rect 16816 17864 16822 17876
rect 18322 17864 18328 17876
rect 16816 17836 18328 17864
rect 16816 17824 16822 17836
rect 18322 17824 18328 17836
rect 18380 17824 18386 17876
rect 23569 17867 23627 17873
rect 18616 17836 21128 17864
rect 16301 17799 16359 17805
rect 10980 17768 11744 17796
rect 6472 17700 7880 17728
rect 8478 17688 8484 17740
rect 8536 17728 8542 17740
rect 8536 17700 9171 17728
rect 8536 17688 8542 17700
rect 6178 17620 6184 17672
rect 6236 17660 6242 17672
rect 6822 17669 6828 17672
rect 6457 17663 6515 17669
rect 6457 17660 6469 17663
rect 6236 17632 6469 17660
rect 6236 17620 6242 17632
rect 6457 17629 6469 17632
rect 6503 17629 6515 17663
rect 6457 17623 6515 17629
rect 6784 17663 6828 17669
rect 6784 17629 6796 17663
rect 6784 17623 6828 17629
rect 6822 17620 6828 17623
rect 6880 17620 6886 17672
rect 6920 17665 6978 17671
rect 6920 17631 6932 17665
rect 6966 17660 6978 17665
rect 7006 17660 7012 17672
rect 6966 17632 7012 17660
rect 6966 17631 6978 17632
rect 6920 17625 6978 17631
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 7190 17620 7196 17672
rect 7248 17620 7254 17672
rect 8570 17620 8576 17672
rect 8628 17660 8634 17672
rect 8665 17663 8723 17669
rect 8665 17660 8677 17663
rect 8628 17632 8677 17660
rect 8628 17620 8634 17632
rect 8665 17629 8677 17632
rect 8711 17629 8723 17663
rect 8665 17623 8723 17629
rect 8846 17620 8852 17672
rect 8904 17660 8910 17672
rect 9030 17669 9036 17672
rect 8992 17663 9036 17669
rect 8992 17660 9004 17663
rect 8904 17632 9004 17660
rect 8904 17620 8910 17632
rect 8992 17629 9004 17632
rect 8992 17623 9036 17629
rect 9030 17620 9036 17623
rect 9088 17620 9094 17672
rect 9143 17671 9171 17700
rect 10134 17688 10140 17740
rect 10192 17688 10198 17740
rect 10781 17731 10839 17737
rect 10781 17697 10793 17731
rect 10827 17728 10839 17731
rect 10962 17728 10968 17740
rect 10827 17700 10968 17728
rect 10827 17697 10839 17700
rect 10781 17691 10839 17697
rect 10962 17688 10968 17700
rect 11020 17688 11026 17740
rect 11146 17688 11152 17740
rect 11204 17688 11210 17740
rect 11333 17731 11391 17737
rect 11333 17697 11345 17731
rect 11379 17697 11391 17731
rect 11716 17728 11744 17768
rect 16301 17765 16313 17799
rect 16347 17796 16359 17799
rect 16850 17796 16856 17808
rect 16347 17768 16856 17796
rect 16347 17765 16359 17768
rect 16301 17759 16359 17765
rect 16850 17756 16856 17768
rect 16908 17756 16914 17808
rect 12529 17731 12587 17737
rect 12529 17728 12541 17731
rect 11716 17700 12541 17728
rect 11333 17691 11391 17697
rect 12529 17697 12541 17700
rect 12575 17697 12587 17731
rect 12529 17691 12587 17697
rect 9128 17665 9186 17671
rect 9128 17631 9140 17665
rect 9174 17631 9186 17665
rect 9128 17625 9186 17631
rect 9214 17620 9220 17672
rect 9272 17660 9278 17672
rect 9401 17663 9459 17669
rect 9401 17660 9413 17663
rect 9272 17632 9413 17660
rect 9272 17620 9278 17632
rect 9401 17629 9413 17632
rect 9447 17629 9459 17663
rect 9401 17623 9459 17629
rect 5905 17595 5963 17601
rect 5905 17561 5917 17595
rect 5951 17592 5963 17595
rect 11348 17592 11376 17691
rect 13906 17688 13912 17740
rect 13964 17728 13970 17740
rect 14185 17731 14243 17737
rect 13964 17700 14136 17728
rect 13964 17688 13970 17700
rect 11514 17620 11520 17672
rect 11572 17660 11578 17672
rect 11698 17660 11704 17672
rect 11572 17632 11704 17660
rect 11572 17620 11578 17632
rect 11698 17620 11704 17632
rect 11756 17660 11762 17672
rect 12158 17669 12164 17672
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11756 17632 11805 17660
rect 11756 17620 11762 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 12120 17663 12164 17669
rect 12120 17629 12132 17663
rect 12120 17623 12164 17629
rect 12158 17620 12164 17623
rect 12216 17620 12222 17672
rect 12299 17663 12357 17669
rect 12299 17629 12311 17663
rect 12345 17660 12357 17663
rect 14108 17660 14136 17700
rect 14185 17697 14197 17731
rect 14231 17728 14243 17731
rect 14826 17728 14832 17740
rect 14231 17700 14832 17728
rect 14231 17697 14243 17700
rect 14185 17691 14243 17697
rect 14826 17688 14832 17700
rect 14884 17688 14890 17740
rect 16390 17688 16396 17740
rect 16448 17728 16454 17740
rect 17681 17731 17739 17737
rect 17681 17728 17693 17731
rect 16448 17700 17693 17728
rect 16448 17688 16454 17700
rect 17681 17697 17693 17700
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 14274 17660 14280 17672
rect 12345 17632 13952 17660
rect 14108 17632 14280 17660
rect 12345 17629 12357 17632
rect 12299 17623 12357 17629
rect 5951 17564 6500 17592
rect 11348 17564 11836 17592
rect 5951 17561 5963 17564
rect 5905 17555 5963 17561
rect 3844 17496 5764 17524
rect 6472 17524 6500 17564
rect 9214 17524 9220 17536
rect 6472 17496 9220 17524
rect 3844 17484 3850 17496
rect 9214 17484 9220 17496
rect 9272 17484 9278 17536
rect 11808 17524 11836 17564
rect 13924 17536 13952 17632
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 14553 17663 14611 17669
rect 14553 17629 14565 17663
rect 14599 17660 14611 17663
rect 14918 17660 14924 17672
rect 14599 17632 14924 17660
rect 14599 17629 14611 17632
rect 14553 17623 14611 17629
rect 14918 17620 14924 17632
rect 14976 17620 14982 17672
rect 16482 17620 16488 17672
rect 16540 17660 16546 17672
rect 17310 17669 17316 17672
rect 16945 17663 17003 17669
rect 16945 17660 16957 17663
rect 16540 17632 16957 17660
rect 16540 17620 16546 17632
rect 16945 17629 16957 17632
rect 16991 17629 17003 17663
rect 16945 17623 17003 17629
rect 17272 17663 17316 17669
rect 17272 17629 17284 17663
rect 17272 17623 17316 17629
rect 17310 17620 17316 17623
rect 17368 17620 17374 17672
rect 17494 17671 17500 17672
rect 17451 17665 17500 17671
rect 17451 17631 17463 17665
rect 17497 17631 17500 17665
rect 17451 17625 17500 17631
rect 17494 17620 17500 17625
rect 17552 17620 17558 17672
rect 15841 17595 15899 17601
rect 15841 17561 15853 17595
rect 15887 17592 15899 17595
rect 16758 17592 16764 17604
rect 15887 17564 16764 17592
rect 15887 17561 15899 17564
rect 15841 17555 15899 17561
rect 16758 17552 16764 17564
rect 16816 17552 16822 17604
rect 13446 17524 13452 17536
rect 11808 17496 13452 17524
rect 13446 17484 13452 17496
rect 13504 17484 13510 17536
rect 13630 17484 13636 17536
rect 13688 17484 13694 17536
rect 13906 17484 13912 17536
rect 13964 17484 13970 17536
rect 14001 17527 14059 17533
rect 14001 17493 14013 17527
rect 14047 17524 14059 17527
rect 14458 17524 14464 17536
rect 14047 17496 14464 17524
rect 14047 17493 14059 17496
rect 14001 17487 14059 17493
rect 14458 17484 14464 17496
rect 14516 17484 14522 17536
rect 16298 17484 16304 17536
rect 16356 17524 16362 17536
rect 18616 17524 18644 17836
rect 21100 17740 21128 17836
rect 23569 17833 23581 17867
rect 23615 17833 23627 17867
rect 23569 17827 23627 17833
rect 23845 17867 23903 17873
rect 23845 17833 23857 17867
rect 23891 17864 23903 17867
rect 23891 17836 24256 17864
rect 23891 17833 23903 17836
rect 23845 17827 23903 17833
rect 23584 17796 23612 17827
rect 24118 17796 24124 17808
rect 23584 17768 24124 17796
rect 24118 17756 24124 17768
rect 24176 17756 24182 17808
rect 18690 17688 18696 17740
rect 18748 17728 18754 17740
rect 19153 17731 19211 17737
rect 19153 17728 19165 17731
rect 18748 17700 19165 17728
rect 18748 17688 18754 17700
rect 19153 17697 19165 17700
rect 19199 17697 19211 17731
rect 19153 17691 19211 17697
rect 19429 17731 19487 17737
rect 19429 17697 19441 17731
rect 19475 17728 19487 17731
rect 19886 17728 19892 17740
rect 19475 17700 19892 17728
rect 19475 17697 19487 17700
rect 19429 17691 19487 17697
rect 19886 17688 19892 17700
rect 19944 17688 19950 17740
rect 20346 17688 20352 17740
rect 20404 17728 20410 17740
rect 20404 17700 20944 17728
rect 20404 17688 20410 17700
rect 20916 17660 20944 17700
rect 21082 17688 21088 17740
rect 21140 17688 21146 17740
rect 21634 17737 21640 17740
rect 21269 17731 21327 17737
rect 21269 17728 21281 17731
rect 21192 17700 21281 17728
rect 21192 17660 21220 17700
rect 21269 17697 21281 17700
rect 21315 17697 21327 17731
rect 21269 17691 21327 17697
rect 21596 17731 21640 17737
rect 21596 17697 21608 17731
rect 21596 17691 21640 17697
rect 21634 17688 21640 17691
rect 21692 17688 21698 17740
rect 22005 17731 22063 17737
rect 22005 17697 22017 17731
rect 22051 17728 22063 17731
rect 22094 17728 22100 17740
rect 22051 17700 22100 17728
rect 22051 17697 22063 17700
rect 22005 17691 22063 17697
rect 22094 17688 22100 17700
rect 22152 17688 22158 17740
rect 23750 17688 23756 17740
rect 23808 17688 23814 17740
rect 24026 17688 24032 17740
rect 24084 17688 24090 17740
rect 24228 17728 24256 17836
rect 24394 17824 24400 17876
rect 24452 17864 24458 17876
rect 24587 17867 24645 17873
rect 24587 17864 24599 17867
rect 24452 17836 24599 17864
rect 24452 17824 24458 17836
rect 24587 17833 24599 17836
rect 24633 17864 24645 17867
rect 25130 17864 25136 17876
rect 24633 17836 25136 17864
rect 24633 17833 24645 17836
rect 24587 17827 24645 17833
rect 25130 17824 25136 17836
rect 25188 17824 25194 17876
rect 26510 17824 26516 17876
rect 26568 17864 26574 17876
rect 27154 17864 27160 17876
rect 26568 17836 27160 17864
rect 26568 17824 26574 17836
rect 27154 17824 27160 17836
rect 27212 17824 27218 17876
rect 28718 17824 28724 17876
rect 28776 17864 28782 17876
rect 30650 17864 30656 17876
rect 28776 17836 30656 17864
rect 28776 17824 28782 17836
rect 30650 17824 30656 17836
rect 30708 17824 30714 17876
rect 28626 17756 28632 17808
rect 28684 17796 28690 17808
rect 28810 17796 28816 17808
rect 28684 17768 28816 17796
rect 28684 17756 28690 17768
rect 28810 17756 28816 17768
rect 28868 17796 28874 17808
rect 28905 17799 28963 17805
rect 28905 17796 28917 17799
rect 28868 17768 28917 17796
rect 28868 17756 28874 17768
rect 28905 17765 28917 17768
rect 28951 17765 28963 17799
rect 28905 17759 28963 17765
rect 29362 17756 29368 17808
rect 29420 17756 29426 17808
rect 26786 17737 26792 17740
rect 24857 17731 24915 17737
rect 24857 17728 24869 17731
rect 24228 17700 24869 17728
rect 24857 17697 24869 17700
rect 24903 17697 24915 17731
rect 24857 17691 24915 17697
rect 26421 17731 26479 17737
rect 26421 17697 26433 17731
rect 26467 17697 26479 17731
rect 26421 17691 26479 17697
rect 26748 17731 26792 17737
rect 26748 17697 26760 17731
rect 26748 17691 26792 17697
rect 21726 17660 21732 17672
rect 20916 17632 21220 17660
rect 21690 17632 21732 17660
rect 21726 17620 21732 17632
rect 21784 17620 21790 17672
rect 24044 17660 24072 17688
rect 22664 17632 24072 17660
rect 24121 17663 24179 17669
rect 16356 17496 18644 17524
rect 16356 17484 16362 17496
rect 18782 17484 18788 17536
rect 18840 17484 18846 17536
rect 18966 17484 18972 17536
rect 19024 17524 19030 17536
rect 20622 17524 20628 17536
rect 19024 17496 20628 17524
rect 19024 17484 19030 17496
rect 20622 17484 20628 17496
rect 20680 17484 20686 17536
rect 20714 17484 20720 17536
rect 20772 17484 20778 17536
rect 20901 17527 20959 17533
rect 20901 17493 20913 17527
rect 20947 17524 20959 17527
rect 20990 17524 20996 17536
rect 20947 17496 20996 17524
rect 20947 17493 20959 17496
rect 20901 17487 20959 17493
rect 20990 17484 20996 17496
rect 21048 17484 21054 17536
rect 21082 17484 21088 17536
rect 21140 17524 21146 17536
rect 22664 17524 22692 17632
rect 24121 17629 24133 17663
rect 24167 17660 24179 17663
rect 24486 17660 24492 17672
rect 24167 17632 24492 17660
rect 24167 17629 24179 17632
rect 24121 17623 24179 17629
rect 23014 17552 23020 17604
rect 23072 17592 23078 17604
rect 23072 17564 23704 17592
rect 23072 17552 23078 17564
rect 21140 17496 22692 17524
rect 21140 17484 21146 17496
rect 23106 17484 23112 17536
rect 23164 17484 23170 17536
rect 23676 17524 23704 17564
rect 24026 17552 24032 17604
rect 24084 17592 24090 17604
rect 24136 17592 24164 17623
rect 24486 17620 24492 17632
rect 24544 17620 24550 17672
rect 24627 17665 24685 17671
rect 24627 17631 24639 17665
rect 24673 17660 24685 17665
rect 24762 17660 24768 17672
rect 24673 17632 24768 17660
rect 24673 17631 24685 17632
rect 24627 17625 24685 17631
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25958 17620 25964 17672
rect 26016 17660 26022 17672
rect 26326 17660 26332 17672
rect 26016 17632 26332 17660
rect 26016 17620 26022 17632
rect 26326 17620 26332 17632
rect 26384 17660 26390 17672
rect 26436 17660 26464 17691
rect 26786 17688 26792 17691
rect 26844 17688 26850 17740
rect 27154 17688 27160 17740
rect 27212 17688 27218 17740
rect 26384 17632 26464 17660
rect 26384 17620 26390 17632
rect 26878 17620 26884 17672
rect 26936 17620 26942 17672
rect 28629 17663 28687 17669
rect 28629 17629 28641 17663
rect 28675 17660 28687 17663
rect 29638 17660 29644 17672
rect 28675 17632 29644 17660
rect 28675 17629 28687 17632
rect 28629 17623 28687 17629
rect 29638 17620 29644 17632
rect 29696 17620 29702 17672
rect 24084 17564 24164 17592
rect 24084 17552 24090 17564
rect 25961 17527 26019 17533
rect 25961 17524 25973 17527
rect 23676 17496 25973 17524
rect 25961 17493 25973 17496
rect 26007 17493 26019 17527
rect 25961 17487 26019 17493
rect 26326 17484 26332 17536
rect 26384 17524 26390 17536
rect 28261 17527 28319 17533
rect 28261 17524 28273 17527
rect 26384 17496 28273 17524
rect 26384 17484 26390 17496
rect 28261 17493 28273 17496
rect 28307 17493 28319 17527
rect 28261 17487 28319 17493
rect 28350 17484 28356 17536
rect 28408 17524 28414 17536
rect 29914 17524 29920 17536
rect 28408 17496 29920 17524
rect 28408 17484 28414 17496
rect 29914 17484 29920 17496
rect 29972 17484 29978 17536
rect 30006 17484 30012 17536
rect 30064 17524 30070 17536
rect 30377 17527 30435 17533
rect 30377 17524 30389 17527
rect 30064 17496 30389 17524
rect 30064 17484 30070 17496
rect 30377 17493 30389 17496
rect 30423 17493 30435 17527
rect 30377 17487 30435 17493
rect 552 17434 30912 17456
rect 552 17382 4193 17434
rect 4245 17382 4257 17434
rect 4309 17382 4321 17434
rect 4373 17382 4385 17434
rect 4437 17382 4449 17434
rect 4501 17382 11783 17434
rect 11835 17382 11847 17434
rect 11899 17382 11911 17434
rect 11963 17382 11975 17434
rect 12027 17382 12039 17434
rect 12091 17382 19373 17434
rect 19425 17382 19437 17434
rect 19489 17382 19501 17434
rect 19553 17382 19565 17434
rect 19617 17382 19629 17434
rect 19681 17382 26963 17434
rect 27015 17382 27027 17434
rect 27079 17382 27091 17434
rect 27143 17382 27155 17434
rect 27207 17382 27219 17434
rect 27271 17382 30912 17434
rect 552 17360 30912 17382
rect 2777 17323 2835 17329
rect 2777 17289 2789 17323
rect 2823 17320 2835 17323
rect 2866 17320 2872 17332
rect 2823 17292 2872 17320
rect 2823 17289 2835 17292
rect 2777 17283 2835 17289
rect 2866 17280 2872 17292
rect 2924 17280 2930 17332
rect 3786 17280 3792 17332
rect 3844 17280 3850 17332
rect 3878 17280 3884 17332
rect 3936 17320 3942 17332
rect 3936 17292 5856 17320
rect 3936 17280 3942 17292
rect 3804 17252 3832 17280
rect 2746 17224 3832 17252
rect 1443 17187 1501 17193
rect 1443 17153 1455 17187
rect 1489 17184 1501 17187
rect 2746 17184 2774 17224
rect 1489 17156 2774 17184
rect 1489 17153 1501 17156
rect 1443 17147 1501 17153
rect 3326 17144 3332 17196
rect 3384 17184 3390 17196
rect 3896 17193 3924 17280
rect 5276 17224 5672 17252
rect 3881 17187 3939 17193
rect 3881 17184 3893 17187
rect 3384 17156 3893 17184
rect 3384 17144 3390 17156
rect 3881 17153 3893 17156
rect 3927 17153 3939 17187
rect 3881 17147 3939 17153
rect 4387 17187 4445 17193
rect 4387 17153 4399 17187
rect 4433 17184 4445 17187
rect 5276 17184 5304 17224
rect 4433 17156 5304 17184
rect 4433 17153 4445 17156
rect 4387 17147 4445 17153
rect 5442 17144 5448 17196
rect 5500 17144 5506 17196
rect 937 17119 995 17125
rect 937 17085 949 17119
rect 983 17116 995 17119
rect 1302 17116 1308 17128
rect 983 17088 1308 17116
rect 983 17085 995 17088
rect 937 17079 995 17085
rect 1302 17076 1308 17088
rect 1360 17076 1366 17128
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17116 1731 17119
rect 2130 17116 2136 17128
rect 1719 17088 2136 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 2130 17076 2136 17088
rect 2188 17076 2194 17128
rect 3237 17119 3295 17125
rect 3237 17085 3249 17119
rect 3283 17116 3295 17119
rect 3694 17116 3700 17128
rect 3283 17088 3700 17116
rect 3283 17085 3295 17088
rect 3237 17079 3295 17085
rect 3694 17076 3700 17088
rect 3752 17076 3758 17128
rect 4617 17119 4675 17125
rect 4617 17085 4629 17119
rect 4663 17116 4675 17119
rect 5460 17116 5488 17144
rect 4663 17088 5488 17116
rect 4663 17085 4675 17088
rect 4617 17079 4675 17085
rect 5644 17060 5672 17224
rect 5828 17060 5856 17292
rect 7190 17280 7196 17332
rect 7248 17320 7254 17332
rect 7248 17292 10456 17320
rect 7248 17280 7254 17292
rect 8386 17212 8392 17264
rect 8444 17212 8450 17264
rect 8570 17212 8576 17264
rect 8628 17212 8634 17264
rect 10428 17252 10456 17292
rect 10502 17280 10508 17332
rect 10560 17280 10566 17332
rect 10870 17280 10876 17332
rect 10928 17280 10934 17332
rect 10980 17292 13860 17320
rect 10980 17252 11008 17292
rect 10428 17224 11008 17252
rect 5997 17187 6055 17193
rect 5997 17153 6009 17187
rect 6043 17184 6055 17187
rect 6552 17187 6610 17193
rect 6552 17184 6564 17187
rect 6043 17156 6564 17184
rect 6043 17153 6055 17156
rect 5997 17147 6055 17153
rect 6552 17153 6564 17156
rect 6598 17153 6610 17187
rect 8588 17184 8616 17212
rect 8665 17187 8723 17193
rect 8665 17184 8677 17187
rect 8588 17156 8677 17184
rect 6552 17147 6610 17153
rect 8665 17153 8677 17156
rect 8711 17153 8723 17187
rect 9128 17185 9186 17191
rect 9128 17184 9140 17185
rect 8665 17147 8723 17153
rect 8772 17156 9140 17184
rect 6089 17119 6147 17125
rect 6089 17085 6101 17119
rect 6135 17116 6147 17119
rect 6178 17116 6184 17128
rect 6135 17088 6184 17116
rect 6135 17085 6147 17088
rect 6089 17079 6147 17085
rect 6178 17076 6184 17088
rect 6236 17076 6242 17128
rect 6454 17125 6460 17128
rect 6416 17119 6460 17125
rect 6416 17085 6428 17119
rect 6416 17079 6460 17085
rect 6454 17076 6460 17079
rect 6512 17076 6518 17128
rect 6822 17076 6828 17128
rect 6880 17076 6886 17128
rect 8478 17076 8484 17128
rect 8536 17116 8542 17128
rect 8573 17119 8631 17125
rect 8573 17116 8585 17119
rect 8536 17088 8585 17116
rect 8536 17076 8542 17088
rect 8573 17085 8585 17088
rect 8619 17085 8631 17119
rect 8573 17079 8631 17085
rect 3513 17051 3571 17057
rect 3513 17017 3525 17051
rect 3559 17017 3571 17051
rect 3513 17011 3571 17017
rect 1394 16940 1400 16992
rect 1452 16989 1458 16992
rect 1452 16943 1461 16989
rect 3528 16980 3556 17011
rect 5626 17008 5632 17060
rect 5684 17008 5690 17060
rect 5810 17008 5816 17060
rect 5868 17008 5874 17060
rect 8205 17051 8263 17057
rect 8205 17017 8217 17051
rect 8251 17048 8263 17051
rect 8772 17048 8800 17156
rect 9128 17151 9140 17156
rect 9174 17151 9186 17185
rect 9128 17145 9186 17151
rect 9398 17144 9404 17196
rect 9456 17144 9462 17196
rect 11241 17187 11299 17193
rect 11241 17153 11253 17187
rect 11287 17184 11299 17187
rect 11514 17184 11520 17196
rect 11287 17156 11520 17184
rect 11287 17153 11299 17156
rect 11241 17147 11299 17153
rect 11514 17144 11520 17156
rect 11572 17144 11578 17196
rect 11747 17187 11805 17193
rect 11747 17153 11759 17187
rect 11793 17184 11805 17187
rect 13446 17184 13452 17196
rect 11793 17156 13452 17184
rect 11793 17153 11805 17156
rect 11747 17147 11805 17153
rect 13446 17144 13452 17156
rect 13504 17144 13510 17196
rect 13832 17184 13860 17292
rect 13906 17280 13912 17332
rect 13964 17320 13970 17332
rect 16025 17323 16083 17329
rect 16025 17320 16037 17323
rect 13964 17292 16037 17320
rect 13964 17280 13970 17292
rect 16025 17289 16037 17292
rect 16071 17289 16083 17323
rect 16025 17283 16083 17289
rect 16408 17292 18828 17320
rect 14001 17255 14059 17261
rect 14001 17221 14013 17255
rect 14047 17252 14059 17255
rect 14182 17252 14188 17264
rect 14047 17224 14188 17252
rect 14047 17221 14059 17224
rect 14001 17215 14059 17221
rect 14182 17212 14188 17224
rect 14240 17212 14246 17264
rect 14691 17187 14749 17193
rect 13832 17156 14596 17184
rect 9674 17076 9680 17128
rect 9732 17116 9738 17128
rect 10594 17116 10600 17128
rect 9732 17088 10600 17116
rect 9732 17076 9738 17088
rect 10594 17076 10600 17088
rect 10652 17116 10658 17128
rect 11057 17119 11115 17125
rect 11057 17116 11069 17119
rect 10652 17088 11069 17116
rect 10652 17076 10658 17088
rect 11057 17085 11069 17088
rect 11103 17085 11115 17119
rect 11977 17119 12035 17125
rect 11977 17116 11989 17119
rect 11057 17079 11115 17085
rect 11348 17088 11989 17116
rect 8251 17020 8800 17048
rect 8251 17017 8263 17020
rect 8205 17011 8263 17017
rect 10870 17008 10876 17060
rect 10928 17048 10934 17060
rect 11348 17048 11376 17088
rect 11977 17085 11989 17088
rect 12023 17085 12035 17119
rect 11977 17079 12035 17085
rect 13998 17076 14004 17128
rect 14056 17116 14062 17128
rect 14185 17119 14243 17125
rect 14185 17116 14197 17119
rect 14056 17088 14197 17116
rect 14056 17076 14062 17088
rect 14185 17085 14197 17088
rect 14231 17085 14243 17119
rect 14568 17116 14596 17156
rect 14691 17153 14703 17187
rect 14737 17184 14749 17187
rect 16408 17184 16436 17292
rect 18800 17252 18828 17292
rect 18966 17280 18972 17332
rect 19024 17280 19030 17332
rect 19245 17323 19303 17329
rect 19245 17289 19257 17323
rect 19291 17320 19303 17323
rect 21910 17320 21916 17332
rect 19291 17292 21916 17320
rect 19291 17289 19303 17292
rect 19245 17283 19303 17289
rect 21910 17280 21916 17292
rect 21968 17280 21974 17332
rect 22002 17280 22008 17332
rect 22060 17320 22066 17332
rect 22060 17292 23152 17320
rect 22060 17280 22066 17292
rect 19058 17252 19064 17264
rect 18800 17224 19064 17252
rect 19058 17212 19064 17224
rect 19116 17212 19122 17264
rect 19518 17212 19524 17264
rect 19576 17212 19582 17264
rect 19702 17212 19708 17264
rect 19760 17252 19766 17264
rect 23014 17252 23020 17264
rect 19760 17224 20116 17252
rect 19760 17212 19766 17224
rect 14737 17156 16436 17184
rect 16899 17187 16957 17193
rect 14737 17153 14749 17156
rect 14691 17147 14749 17153
rect 16899 17153 16911 17187
rect 16945 17184 16957 17187
rect 17862 17184 17868 17196
rect 16945 17156 17868 17184
rect 16945 17153 16957 17156
rect 16899 17147 16957 17153
rect 17862 17144 17868 17156
rect 17920 17144 17926 17196
rect 18690 17144 18696 17196
rect 18748 17144 18754 17196
rect 18984 17156 19472 17184
rect 14826 17116 14832 17128
rect 14568 17088 14832 17116
rect 14185 17079 14243 17085
rect 14826 17076 14832 17088
rect 14884 17076 14890 17128
rect 14921 17119 14979 17125
rect 14921 17085 14933 17119
rect 14967 17116 14979 17119
rect 15930 17116 15936 17128
rect 14967 17088 15936 17116
rect 14967 17085 14979 17088
rect 14921 17079 14979 17085
rect 15930 17076 15936 17088
rect 15988 17076 15994 17128
rect 16393 17119 16451 17125
rect 16393 17085 16405 17119
rect 16439 17116 16451 17119
rect 16482 17116 16488 17128
rect 16439 17088 16488 17116
rect 16439 17085 16451 17088
rect 16393 17079 16451 17085
rect 16482 17076 16488 17088
rect 16540 17076 16546 17128
rect 16758 17125 16764 17128
rect 16720 17119 16764 17125
rect 16720 17085 16732 17119
rect 16816 17116 16822 17128
rect 17034 17116 17040 17128
rect 16816 17088 17040 17116
rect 16720 17079 16764 17085
rect 16758 17076 16764 17079
rect 16816 17076 16822 17088
rect 17034 17076 17040 17088
rect 17092 17076 17098 17128
rect 17129 17119 17187 17125
rect 17129 17085 17141 17119
rect 17175 17116 17187 17119
rect 18138 17116 18144 17128
rect 17175 17088 18144 17116
rect 17175 17085 17187 17088
rect 17129 17079 17187 17085
rect 18138 17076 18144 17088
rect 18196 17076 18202 17128
rect 10928 17020 11376 17048
rect 10928 17008 10934 17020
rect 13170 17008 13176 17060
rect 13228 17048 13234 17060
rect 13725 17051 13783 17057
rect 13725 17048 13737 17051
rect 13228 17020 13737 17048
rect 13228 17008 13234 17020
rect 13725 17017 13737 17020
rect 13771 17048 13783 17051
rect 13906 17048 13912 17060
rect 13771 17020 13912 17048
rect 13771 17017 13783 17020
rect 13725 17011 13783 17017
rect 13906 17008 13912 17020
rect 13964 17008 13970 17060
rect 18984 17048 19012 17156
rect 19153 17119 19211 17125
rect 19153 17085 19165 17119
rect 19199 17116 19211 17119
rect 19334 17116 19340 17128
rect 19199 17088 19340 17116
rect 19199 17085 19211 17088
rect 19153 17079 19211 17085
rect 19334 17076 19340 17088
rect 19392 17076 19398 17128
rect 19444 17125 19472 17156
rect 19429 17119 19487 17125
rect 19429 17085 19441 17119
rect 19475 17085 19487 17119
rect 19429 17079 19487 17085
rect 19705 17119 19763 17125
rect 19705 17085 19717 17119
rect 19751 17085 19763 17119
rect 19705 17079 19763 17085
rect 19797 17119 19855 17125
rect 19797 17085 19809 17119
rect 19843 17116 19855 17119
rect 20088 17116 20116 17224
rect 22066 17224 23020 17252
rect 20855 17187 20913 17193
rect 20855 17153 20867 17187
rect 20901 17184 20913 17187
rect 22066 17184 22094 17224
rect 23014 17212 23020 17224
rect 23072 17212 23078 17264
rect 23124 17252 23152 17292
rect 23198 17280 23204 17332
rect 23256 17320 23262 17332
rect 23256 17292 25268 17320
rect 23256 17280 23262 17292
rect 23124 17224 23704 17252
rect 20901 17156 22094 17184
rect 23477 17187 23535 17193
rect 20901 17153 20913 17156
rect 20855 17147 20913 17153
rect 23477 17153 23489 17187
rect 23523 17184 23535 17187
rect 23566 17184 23572 17196
rect 23523 17156 23572 17184
rect 23523 17153 23535 17156
rect 23477 17147 23535 17153
rect 23566 17144 23572 17156
rect 23624 17144 23630 17196
rect 23676 17184 23704 17224
rect 24121 17187 24179 17193
rect 24121 17184 24133 17187
rect 23676 17156 24133 17184
rect 24121 17153 24133 17156
rect 24167 17153 24179 17187
rect 24121 17147 24179 17153
rect 20254 17116 20260 17128
rect 19843 17088 20260 17116
rect 19843 17085 19855 17088
rect 19797 17079 19855 17085
rect 18156 17020 19012 17048
rect 4347 16983 4405 16989
rect 4347 16980 4359 16983
rect 3528 16952 4359 16980
rect 4347 16949 4359 16952
rect 4393 16980 4405 16983
rect 4522 16980 4528 16992
rect 4393 16952 4528 16980
rect 4393 16949 4405 16952
rect 4347 16943 4405 16949
rect 1452 16940 1458 16943
rect 4522 16940 4528 16952
rect 4580 16980 4586 16992
rect 6178 16980 6184 16992
rect 4580 16952 6184 16980
rect 4580 16940 4586 16952
rect 6178 16940 6184 16952
rect 6236 16940 6242 16992
rect 9030 16940 9036 16992
rect 9088 16980 9094 16992
rect 9131 16983 9189 16989
rect 9131 16980 9143 16983
rect 9088 16952 9143 16980
rect 9088 16940 9094 16952
rect 9131 16949 9143 16952
rect 9177 16949 9189 16983
rect 9131 16943 9189 16949
rect 11707 16983 11765 16989
rect 11707 16949 11719 16983
rect 11753 16980 11765 16983
rect 12066 16980 12072 16992
rect 11753 16952 12072 16980
rect 11753 16949 11765 16952
rect 11707 16943 11765 16949
rect 12066 16940 12072 16952
rect 12124 16940 12130 16992
rect 13078 16940 13084 16992
rect 13136 16940 13142 16992
rect 14182 16940 14188 16992
rect 14240 16980 14246 16992
rect 14651 16983 14709 16989
rect 14651 16980 14663 16983
rect 14240 16952 14663 16980
rect 14240 16940 14246 16952
rect 14651 16949 14663 16952
rect 14697 16949 14709 16983
rect 14651 16943 14709 16949
rect 14826 16940 14832 16992
rect 14884 16980 14890 16992
rect 16666 16980 16672 16992
rect 14884 16952 16672 16980
rect 14884 16940 14890 16952
rect 16666 16940 16672 16952
rect 16724 16940 16730 16992
rect 17034 16940 17040 16992
rect 17092 16980 17098 16992
rect 18156 16980 18184 17020
rect 17092 16952 18184 16980
rect 17092 16940 17098 16952
rect 18230 16940 18236 16992
rect 18288 16940 18294 16992
rect 19444 16980 19472 17079
rect 19720 17048 19748 17079
rect 20254 17076 20260 17088
rect 20312 17076 20318 17128
rect 20346 17076 20352 17128
rect 20404 17076 20410 17128
rect 20622 17116 20628 17128
rect 20456 17088 20628 17116
rect 19886 17048 19892 17060
rect 19720 17020 19892 17048
rect 19886 17008 19892 17020
rect 19944 17008 19950 17060
rect 19978 17008 19984 17060
rect 20036 17048 20042 17060
rect 20073 17051 20131 17057
rect 20073 17048 20085 17051
rect 20036 17020 20085 17048
rect 20036 17008 20042 17020
rect 20073 17017 20085 17020
rect 20119 17048 20131 17051
rect 20456 17048 20484 17088
rect 20622 17076 20628 17088
rect 20680 17125 20686 17128
rect 20680 17119 20734 17125
rect 20680 17085 20688 17119
rect 20722 17116 20734 17119
rect 20722 17088 20773 17116
rect 20722 17085 20734 17088
rect 20680 17079 20734 17085
rect 20680 17076 20686 17079
rect 20990 17076 20996 17128
rect 21048 17116 21054 17128
rect 21085 17119 21143 17125
rect 21085 17116 21097 17119
rect 21048 17088 21097 17116
rect 21048 17076 21054 17088
rect 21085 17085 21097 17088
rect 21131 17085 21143 17119
rect 23106 17116 23112 17128
rect 21085 17079 21143 17085
rect 21928 17088 23112 17116
rect 20119 17020 20484 17048
rect 20119 17017 20131 17020
rect 20073 17011 20131 17017
rect 21928 16980 21956 17088
rect 23106 17076 23112 17088
rect 23164 17076 23170 17128
rect 23201 17119 23259 17125
rect 23201 17085 23213 17119
rect 23247 17085 23259 17119
rect 23201 17079 23259 17085
rect 22646 17008 22652 17060
rect 22704 17008 22710 17060
rect 23014 17008 23020 17060
rect 23072 17048 23078 17060
rect 23216 17048 23244 17079
rect 23842 17076 23848 17128
rect 23900 17076 23906 17128
rect 24210 17076 24216 17128
rect 24268 17116 24274 17128
rect 25240 17116 25268 17292
rect 25406 17280 25412 17332
rect 25464 17320 25470 17332
rect 25593 17323 25651 17329
rect 25593 17320 25605 17323
rect 25464 17292 25605 17320
rect 25464 17280 25470 17292
rect 25593 17289 25605 17292
rect 25639 17289 25651 17323
rect 26234 17320 26240 17332
rect 25593 17283 25651 17289
rect 25884 17292 26240 17320
rect 25501 17187 25559 17193
rect 25501 17153 25513 17187
rect 25547 17184 25559 17187
rect 25884 17184 25912 17292
rect 26234 17280 26240 17292
rect 26292 17280 26298 17332
rect 27246 17280 27252 17332
rect 27304 17280 27310 17332
rect 28718 17320 28724 17332
rect 28184 17292 28724 17320
rect 27264 17252 27292 17280
rect 28184 17252 28212 17292
rect 28718 17280 28724 17292
rect 28776 17320 28782 17332
rect 29362 17320 29368 17332
rect 28776 17292 29368 17320
rect 28776 17280 28782 17292
rect 29362 17280 29368 17292
rect 29420 17280 29426 17332
rect 30377 17323 30435 17329
rect 30377 17289 30389 17323
rect 30423 17320 30435 17323
rect 30558 17320 30564 17332
rect 30423 17292 30564 17320
rect 30423 17289 30435 17292
rect 30377 17283 30435 17289
rect 30558 17280 30564 17292
rect 30616 17280 30622 17332
rect 27264 17224 28212 17252
rect 25547 17156 25912 17184
rect 26375 17187 26433 17193
rect 25547 17153 25559 17156
rect 25501 17147 25559 17153
rect 26375 17153 26387 17187
rect 26421 17184 26433 17187
rect 27522 17184 27528 17196
rect 26421 17156 27528 17184
rect 26421 17153 26433 17156
rect 26375 17147 26433 17153
rect 27522 17144 27528 17156
rect 27580 17144 27586 17196
rect 28184 17193 28212 17224
rect 28626 17212 28632 17264
rect 28684 17252 28690 17264
rect 28684 17224 29868 17252
rect 28684 17212 28690 17224
rect 29840 17193 29868 17224
rect 28169 17187 28227 17193
rect 28169 17153 28181 17187
rect 28215 17153 28227 17187
rect 29825 17187 29883 17193
rect 28169 17147 28227 17153
rect 28368 17156 29684 17184
rect 25774 17116 25780 17128
rect 24268 17088 25176 17116
rect 25240 17088 25780 17116
rect 24268 17076 24274 17088
rect 25148 17060 25176 17088
rect 25774 17076 25780 17088
rect 25832 17076 25838 17128
rect 25869 17119 25927 17125
rect 25869 17085 25881 17119
rect 25915 17116 25927 17119
rect 25958 17116 25964 17128
rect 25915 17088 25964 17116
rect 25915 17085 25927 17088
rect 25869 17079 25927 17085
rect 25958 17076 25964 17088
rect 26016 17076 26022 17128
rect 26605 17119 26663 17125
rect 26605 17085 26617 17119
rect 26651 17116 26663 17119
rect 27338 17116 27344 17128
rect 26651 17088 27344 17116
rect 26651 17085 26663 17088
rect 26605 17079 26663 17085
rect 27338 17076 27344 17088
rect 27396 17076 27402 17128
rect 28368 17125 28396 17156
rect 29656 17128 29684 17156
rect 29825 17153 29837 17187
rect 29871 17184 29883 17187
rect 30282 17184 30288 17196
rect 29871 17156 30288 17184
rect 29871 17153 29883 17156
rect 29825 17147 29883 17153
rect 30282 17144 30288 17156
rect 30340 17144 30346 17196
rect 28353 17119 28411 17125
rect 28353 17085 28365 17119
rect 28399 17085 28411 17119
rect 28353 17079 28411 17085
rect 28445 17119 28503 17125
rect 28445 17085 28457 17119
rect 28491 17116 28503 17119
rect 28491 17088 28672 17116
rect 28491 17085 28503 17088
rect 28445 17079 28503 17085
rect 28644 17060 28672 17088
rect 28718 17076 28724 17128
rect 28776 17116 28782 17128
rect 29089 17119 29147 17125
rect 29089 17116 29101 17119
rect 28776 17088 29101 17116
rect 28776 17076 28782 17088
rect 29089 17085 29101 17088
rect 29135 17085 29147 17119
rect 29089 17079 29147 17085
rect 29638 17076 29644 17128
rect 29696 17076 29702 17128
rect 23072 17020 23983 17048
rect 23072 17008 23078 17020
rect 19444 16952 21956 16980
rect 22186 16940 22192 16992
rect 22244 16940 22250 16992
rect 22925 16983 22983 16989
rect 22925 16949 22937 16983
rect 22971 16980 22983 16983
rect 23842 16980 23848 16992
rect 22971 16952 23848 16980
rect 22971 16949 22983 16952
rect 22925 16943 22983 16949
rect 23842 16940 23848 16952
rect 23900 16940 23906 16992
rect 23955 16980 23983 17020
rect 25130 17008 25136 17060
rect 25188 17008 25194 17060
rect 28258 17048 28264 17060
rect 27264 17020 28264 17048
rect 27264 16992 27292 17020
rect 28258 17008 28264 17020
rect 28316 17008 28322 17060
rect 28626 17008 28632 17060
rect 28684 17008 28690 17060
rect 30098 17048 30104 17060
rect 29840 17020 30104 17048
rect 26142 16980 26148 16992
rect 23955 16952 26148 16980
rect 26142 16940 26148 16952
rect 26200 16940 26206 16992
rect 26335 16983 26393 16989
rect 26335 16949 26347 16983
rect 26381 16980 26393 16983
rect 26694 16980 26700 16992
rect 26381 16952 26700 16980
rect 26381 16949 26393 16952
rect 26335 16943 26393 16949
rect 26694 16940 26700 16952
rect 26752 16940 26758 16992
rect 27246 16940 27252 16992
rect 27304 16940 27310 16992
rect 27706 16940 27712 16992
rect 27764 16940 27770 16992
rect 28718 16940 28724 16992
rect 28776 16940 28782 16992
rect 29362 16940 29368 16992
rect 29420 16980 29426 16992
rect 29840 16980 29868 17020
rect 30098 17008 30104 17020
rect 30156 17008 30162 17060
rect 29420 16952 29868 16980
rect 29420 16940 29426 16952
rect 29914 16940 29920 16992
rect 29972 16940 29978 16992
rect 552 16890 31072 16912
rect 552 16838 7988 16890
rect 8040 16838 8052 16890
rect 8104 16838 8116 16890
rect 8168 16838 8180 16890
rect 8232 16838 8244 16890
rect 8296 16838 15578 16890
rect 15630 16838 15642 16890
rect 15694 16838 15706 16890
rect 15758 16838 15770 16890
rect 15822 16838 15834 16890
rect 15886 16838 23168 16890
rect 23220 16838 23232 16890
rect 23284 16838 23296 16890
rect 23348 16838 23360 16890
rect 23412 16838 23424 16890
rect 23476 16838 30758 16890
rect 30810 16838 30822 16890
rect 30874 16838 30886 16890
rect 30938 16838 30950 16890
rect 31002 16838 31014 16890
rect 31066 16838 31072 16890
rect 552 16816 31072 16838
rect 1403 16779 1461 16785
rect 1403 16745 1415 16779
rect 1449 16776 1461 16779
rect 2866 16776 2872 16788
rect 1449 16748 2872 16776
rect 1449 16745 1461 16748
rect 1403 16739 1461 16745
rect 2866 16736 2872 16748
rect 2924 16736 2930 16788
rect 3145 16779 3203 16785
rect 3145 16745 3157 16779
rect 3191 16776 3203 16779
rect 3191 16748 3648 16776
rect 3191 16745 3203 16748
rect 3145 16739 3203 16745
rect 934 16600 940 16652
rect 992 16600 998 16652
rect 3329 16643 3387 16649
rect 3329 16640 3341 16643
rect 1596 16612 2820 16640
rect 1433 16593 1491 16599
rect 1433 16559 1445 16593
rect 1479 16572 1491 16593
rect 1596 16572 1624 16612
rect 2792 16584 2820 16612
rect 3252 16612 3341 16640
rect 3252 16584 3280 16612
rect 3329 16609 3341 16612
rect 3375 16609 3387 16643
rect 3620 16640 3648 16748
rect 4154 16736 4160 16788
rect 4212 16776 4218 16788
rect 4706 16776 4712 16788
rect 4212 16748 4712 16776
rect 4212 16736 4218 16748
rect 4706 16736 4712 16748
rect 4764 16736 4770 16788
rect 4890 16736 4896 16788
rect 4948 16776 4954 16788
rect 5353 16779 5411 16785
rect 5353 16776 5365 16779
rect 4948 16748 5365 16776
rect 4948 16736 4954 16748
rect 5353 16745 5365 16748
rect 5399 16745 5411 16779
rect 6914 16776 6920 16788
rect 5353 16739 5411 16745
rect 5460 16748 6920 16776
rect 4249 16643 4307 16649
rect 4249 16640 4261 16643
rect 3620 16612 4261 16640
rect 3329 16603 3387 16609
rect 4249 16609 4261 16612
rect 4295 16609 4307 16643
rect 5460 16640 5488 16748
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 7006 16736 7012 16788
rect 7064 16776 7070 16788
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 7064 16748 7665 16776
rect 7064 16736 7070 16748
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 7653 16739 7711 16745
rect 8389 16779 8447 16785
rect 8389 16745 8401 16779
rect 8435 16776 8447 16779
rect 8570 16776 8576 16788
rect 8435 16748 8576 16776
rect 8435 16745 8447 16748
rect 8389 16739 8447 16745
rect 8570 16736 8576 16748
rect 8628 16736 8634 16788
rect 8680 16748 10088 16776
rect 8113 16711 8171 16717
rect 8113 16677 8125 16711
rect 8159 16708 8171 16711
rect 8680 16708 8708 16748
rect 10060 16720 10088 16748
rect 10962 16736 10968 16788
rect 11020 16776 11026 16788
rect 12342 16776 12348 16788
rect 11020 16748 12348 16776
rect 11020 16736 11026 16748
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 12802 16736 12808 16788
rect 12860 16776 12866 16788
rect 13449 16779 13507 16785
rect 13449 16776 13461 16779
rect 12860 16748 13461 16776
rect 12860 16736 12866 16748
rect 13449 16745 13461 16748
rect 13495 16745 13507 16779
rect 15657 16779 15715 16785
rect 15657 16776 15669 16779
rect 13449 16739 13507 16745
rect 13556 16748 15669 16776
rect 8159 16680 8708 16708
rect 8159 16677 8171 16680
rect 8113 16671 8171 16677
rect 10042 16668 10048 16720
rect 10100 16668 10106 16720
rect 11422 16708 11428 16720
rect 10980 16680 11428 16708
rect 4249 16603 4307 16609
rect 4356 16612 5488 16640
rect 1479 16559 1624 16572
rect 1433 16553 1624 16559
rect 1448 16544 1624 16553
rect 1670 16532 1676 16584
rect 1728 16532 1734 16584
rect 2774 16532 2780 16584
rect 2832 16532 2838 16584
rect 3234 16532 3240 16584
rect 3292 16532 3298 16584
rect 3510 16532 3516 16584
rect 3568 16532 3574 16584
rect 3878 16581 3884 16584
rect 3840 16575 3884 16581
rect 3840 16541 3852 16575
rect 3840 16535 3884 16541
rect 3878 16532 3884 16535
rect 3936 16532 3942 16584
rect 3976 16577 4034 16583
rect 3976 16543 3988 16577
rect 4022 16572 4034 16577
rect 4356 16572 4384 16612
rect 5718 16600 5724 16652
rect 5776 16640 5782 16652
rect 6549 16643 6607 16649
rect 6549 16640 6561 16643
rect 5776 16612 6561 16640
rect 5776 16600 5782 16612
rect 6549 16609 6561 16612
rect 6595 16609 6607 16643
rect 6549 16603 6607 16609
rect 8573 16643 8631 16649
rect 8573 16609 8585 16643
rect 8619 16640 8631 16643
rect 8662 16640 8668 16652
rect 8619 16612 8668 16640
rect 8619 16609 8631 16612
rect 8573 16603 8631 16609
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 9306 16600 9312 16652
rect 9364 16600 9370 16652
rect 10980 16640 11008 16680
rect 11422 16668 11428 16680
rect 11480 16668 11486 16720
rect 9646 16612 11008 16640
rect 11057 16643 11115 16649
rect 9069 16593 9127 16599
rect 4022 16544 4384 16572
rect 4022 16543 4034 16544
rect 3976 16537 4034 16543
rect 5810 16532 5816 16584
rect 5868 16532 5874 16584
rect 6178 16581 6184 16584
rect 6140 16575 6184 16581
rect 6140 16541 6152 16575
rect 6140 16535 6184 16541
rect 6178 16532 6184 16535
rect 6236 16532 6242 16584
rect 6270 16532 6276 16584
rect 6328 16532 6334 16584
rect 6638 16532 6644 16584
rect 6696 16572 6702 16584
rect 8938 16581 8944 16584
rect 8900 16575 8944 16581
rect 6696 16544 8616 16572
rect 6696 16532 6702 16544
rect 2406 16464 2412 16516
rect 2464 16504 2470 16516
rect 2464 16476 3556 16504
rect 2464 16464 2470 16476
rect 2314 16396 2320 16448
rect 2372 16436 2378 16448
rect 2777 16439 2835 16445
rect 2777 16436 2789 16439
rect 2372 16408 2789 16436
rect 2372 16396 2378 16408
rect 2777 16405 2789 16408
rect 2823 16405 2835 16439
rect 3528 16436 3556 16476
rect 7282 16436 7288 16448
rect 3528 16408 7288 16436
rect 2777 16399 2835 16405
rect 7282 16396 7288 16408
rect 7340 16396 7346 16448
rect 8588 16436 8616 16544
rect 8900 16541 8912 16575
rect 8900 16535 8944 16541
rect 8938 16532 8944 16535
rect 8996 16532 9002 16584
rect 9069 16559 9081 16593
rect 9115 16590 9127 16593
rect 9115 16572 9214 16590
rect 9646 16572 9674 16612
rect 11057 16609 11069 16643
rect 11103 16640 11115 16643
rect 11103 16612 11468 16640
rect 11103 16609 11115 16612
rect 11057 16603 11115 16609
rect 9115 16562 9674 16572
rect 9115 16559 9127 16562
rect 9069 16553 9127 16559
rect 9186 16544 9674 16562
rect 9766 16532 9772 16584
rect 9824 16572 9830 16584
rect 11146 16572 11152 16584
rect 9824 16544 11152 16572
rect 9824 16532 9830 16544
rect 11146 16532 11152 16544
rect 11204 16572 11210 16584
rect 11333 16575 11391 16581
rect 11333 16572 11345 16575
rect 11204 16544 11345 16572
rect 11204 16532 11210 16544
rect 11333 16541 11345 16544
rect 11379 16541 11391 16575
rect 11333 16535 11391 16541
rect 11440 16516 11468 16612
rect 11514 16600 11520 16652
rect 11572 16640 11578 16652
rect 11609 16643 11667 16649
rect 11609 16640 11621 16643
rect 11572 16612 11621 16640
rect 11572 16600 11578 16612
rect 11609 16609 11621 16612
rect 11655 16609 11667 16643
rect 13556 16640 13584 16748
rect 15657 16745 15669 16748
rect 15703 16745 15715 16779
rect 15657 16739 15715 16745
rect 16390 16736 16396 16788
rect 16448 16736 16454 16788
rect 16574 16736 16580 16788
rect 16632 16736 16638 16788
rect 16669 16779 16727 16785
rect 16669 16745 16681 16779
rect 16715 16745 16727 16779
rect 16669 16739 16727 16745
rect 11609 16603 11667 16609
rect 12268 16612 13584 16640
rect 11974 16581 11980 16584
rect 11936 16575 11980 16581
rect 11936 16541 11948 16575
rect 11936 16535 11980 16541
rect 11974 16532 11980 16535
rect 12032 16532 12038 16584
rect 12115 16575 12173 16581
rect 12115 16541 12127 16575
rect 12161 16572 12173 16575
rect 12268 16572 12296 16612
rect 14458 16600 14464 16652
rect 14516 16640 14522 16652
rect 14553 16643 14611 16649
rect 14553 16640 14565 16643
rect 14516 16612 14565 16640
rect 14516 16600 14522 16612
rect 14553 16609 14565 16612
rect 14599 16609 14611 16643
rect 14553 16603 14611 16609
rect 14660 16612 16252 16640
rect 12161 16544 12296 16572
rect 12161 16541 12173 16544
rect 12115 16535 12173 16541
rect 12342 16532 12348 16584
rect 12400 16532 12406 16584
rect 13817 16575 13875 16581
rect 13817 16541 13829 16575
rect 13863 16572 13875 16575
rect 13998 16572 14004 16584
rect 13863 16544 14004 16572
rect 13863 16541 13875 16544
rect 13817 16535 13875 16541
rect 13998 16532 14004 16544
rect 14056 16532 14062 16584
rect 14182 16581 14188 16584
rect 14144 16575 14188 16581
rect 14144 16541 14156 16575
rect 14144 16535 14188 16541
rect 14182 16532 14188 16535
rect 14240 16532 14246 16584
rect 14280 16577 14338 16583
rect 14280 16543 14292 16577
rect 14326 16572 14338 16577
rect 14660 16572 14688 16612
rect 14326 16544 14688 16572
rect 16224 16572 16252 16612
rect 16298 16600 16304 16652
rect 16356 16600 16362 16652
rect 16592 16649 16620 16736
rect 16684 16708 16712 16739
rect 17310 16736 17316 16788
rect 17368 16776 17374 16788
rect 17411 16779 17469 16785
rect 17411 16776 17423 16779
rect 17368 16748 17423 16776
rect 17368 16736 17374 16748
rect 17411 16745 17423 16748
rect 17457 16745 17469 16779
rect 17411 16739 17469 16745
rect 18138 16736 18144 16788
rect 18196 16776 18202 16788
rect 19153 16779 19211 16785
rect 19153 16776 19165 16779
rect 18196 16748 19165 16776
rect 18196 16736 18202 16748
rect 19153 16745 19165 16748
rect 19199 16745 19211 16779
rect 23109 16779 23167 16785
rect 23109 16776 23121 16779
rect 19153 16739 19211 16745
rect 19306 16748 23121 16776
rect 16684 16680 17080 16708
rect 16577 16643 16635 16649
rect 16577 16609 16589 16643
rect 16623 16609 16635 16643
rect 16577 16603 16635 16609
rect 16850 16600 16856 16652
rect 16908 16600 16914 16652
rect 17052 16640 17080 16680
rect 19058 16668 19064 16720
rect 19116 16668 19122 16720
rect 19306 16708 19334 16748
rect 23109 16745 23121 16748
rect 23155 16745 23167 16779
rect 23109 16739 23167 16745
rect 23753 16779 23811 16785
rect 23753 16745 23765 16779
rect 23799 16776 23811 16779
rect 24118 16776 24124 16788
rect 23799 16748 24124 16776
rect 23799 16745 23811 16748
rect 23753 16739 23811 16745
rect 24118 16736 24124 16748
rect 24176 16736 24182 16788
rect 26418 16776 26424 16788
rect 24228 16748 26424 16776
rect 19168 16680 19334 16708
rect 17681 16643 17739 16649
rect 17681 16640 17693 16643
rect 17052 16612 17693 16640
rect 17681 16609 17693 16612
rect 17727 16609 17739 16643
rect 17681 16603 17739 16609
rect 16945 16575 17003 16581
rect 16224 16544 16620 16572
rect 14326 16543 14338 16544
rect 14280 16537 14338 16543
rect 10042 16464 10048 16516
rect 10100 16504 10106 16516
rect 11422 16504 11428 16516
rect 10100 16476 11428 16504
rect 10100 16464 10106 16476
rect 11422 16464 11428 16476
rect 11480 16464 11486 16516
rect 9030 16436 9036 16448
rect 8588 16408 9036 16436
rect 9030 16396 9036 16408
rect 9088 16396 9094 16448
rect 9490 16396 9496 16448
rect 9548 16436 9554 16448
rect 10413 16439 10471 16445
rect 10413 16436 10425 16439
rect 9548 16408 10425 16436
rect 9548 16396 9554 16408
rect 10413 16405 10425 16408
rect 10459 16405 10471 16439
rect 10413 16399 10471 16405
rect 13814 16396 13820 16448
rect 13872 16436 13878 16448
rect 14458 16436 14464 16448
rect 13872 16408 14464 16436
rect 13872 16396 13878 16408
rect 14458 16396 14464 16408
rect 14516 16396 14522 16448
rect 16114 16396 16120 16448
rect 16172 16396 16178 16448
rect 16592 16436 16620 16544
rect 16945 16541 16957 16575
rect 16991 16572 17003 16575
rect 17218 16572 17224 16584
rect 16991 16544 17224 16572
rect 16991 16541 17003 16544
rect 16945 16535 17003 16541
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 17451 16577 17509 16583
rect 17451 16543 17463 16577
rect 17497 16572 17509 16577
rect 19168 16572 19196 16680
rect 20622 16668 20628 16720
rect 20680 16708 20686 16720
rect 24228 16708 24256 16748
rect 26418 16736 26424 16748
rect 26476 16736 26482 16788
rect 26988 16748 29132 16776
rect 26513 16711 26571 16717
rect 26513 16708 26525 16711
rect 20680 16680 21220 16708
rect 20680 16668 20686 16680
rect 19334 16600 19340 16652
rect 19392 16640 19398 16652
rect 19705 16643 19763 16649
rect 19392 16612 19656 16640
rect 19392 16600 19398 16612
rect 17497 16544 19196 16572
rect 19429 16575 19487 16581
rect 17497 16543 17509 16544
rect 17451 16537 17509 16543
rect 19429 16541 19441 16575
rect 19475 16541 19487 16575
rect 19628 16572 19656 16612
rect 19705 16609 19717 16643
rect 19751 16640 19763 16643
rect 19794 16640 19800 16652
rect 19751 16612 19800 16640
rect 19751 16609 19763 16612
rect 19705 16603 19763 16609
rect 19794 16600 19800 16612
rect 19852 16600 19858 16652
rect 21082 16640 21088 16652
rect 19904 16612 21088 16640
rect 19904 16572 19932 16612
rect 21082 16600 21088 16612
rect 21140 16600 21146 16652
rect 21192 16640 21220 16680
rect 23584 16680 24256 16708
rect 25516 16680 26525 16708
rect 23584 16640 23612 16680
rect 21192 16612 21639 16640
rect 21611 16584 21639 16612
rect 21790 16612 23612 16640
rect 23661 16643 23719 16649
rect 19628 16544 19932 16572
rect 19429 16535 19487 16541
rect 17126 16436 17132 16448
rect 16592 16408 17132 16436
rect 17126 16396 17132 16408
rect 17184 16396 17190 16448
rect 19444 16436 19472 16535
rect 20346 16532 20352 16584
rect 20404 16572 20410 16584
rect 21611 16581 21640 16584
rect 21269 16575 21327 16581
rect 21269 16572 21281 16575
rect 20404 16544 21281 16572
rect 20404 16532 20410 16544
rect 21269 16541 21281 16544
rect 21315 16541 21327 16575
rect 21269 16535 21327 16541
rect 21596 16575 21640 16581
rect 21596 16541 21608 16575
rect 21596 16535 21640 16541
rect 21284 16448 21312 16535
rect 21634 16532 21640 16535
rect 21692 16532 21698 16584
rect 21790 16583 21818 16612
rect 23661 16609 23673 16643
rect 23707 16609 23719 16643
rect 23661 16603 23719 16609
rect 21775 16577 21833 16583
rect 21775 16543 21787 16577
rect 21821 16543 21833 16577
rect 21775 16537 21833 16543
rect 21910 16532 21916 16584
rect 21968 16574 21974 16584
rect 22005 16575 22063 16581
rect 22005 16574 22017 16575
rect 21968 16546 22017 16574
rect 21968 16532 21974 16546
rect 22005 16541 22017 16546
rect 22051 16541 22063 16575
rect 22005 16535 22063 16541
rect 22646 16532 22652 16584
rect 22704 16532 22710 16584
rect 23676 16572 23704 16603
rect 23934 16600 23940 16652
rect 23992 16600 23998 16652
rect 24026 16600 24032 16652
rect 24084 16640 24090 16652
rect 24121 16643 24179 16649
rect 24121 16640 24133 16643
rect 24084 16612 24133 16640
rect 24084 16600 24090 16612
rect 24121 16609 24133 16612
rect 24167 16640 24179 16643
rect 24857 16643 24915 16649
rect 24167 16612 24808 16640
rect 24167 16609 24179 16612
rect 24121 16603 24179 16609
rect 22756 16544 23704 16572
rect 19702 16436 19708 16448
rect 19444 16408 19708 16436
rect 19702 16396 19708 16408
rect 19760 16436 19766 16448
rect 20070 16436 20076 16448
rect 19760 16408 20076 16436
rect 19760 16396 19766 16408
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 20990 16396 20996 16448
rect 21048 16396 21054 16448
rect 21266 16396 21272 16448
rect 21324 16436 21330 16448
rect 22664 16436 22692 16532
rect 22756 16448 22784 16544
rect 24302 16532 24308 16584
rect 24360 16572 24366 16584
rect 24448 16575 24506 16581
rect 24448 16572 24460 16575
rect 24360 16544 24460 16572
rect 24360 16532 24366 16544
rect 24448 16541 24460 16544
rect 24494 16541 24506 16575
rect 24448 16535 24506 16541
rect 24578 16532 24584 16584
rect 24636 16574 24642 16584
rect 24636 16546 24679 16574
rect 24780 16572 24808 16612
rect 24857 16609 24869 16643
rect 24903 16640 24915 16643
rect 24946 16640 24952 16652
rect 24903 16612 24952 16640
rect 24903 16609 24915 16612
rect 24857 16603 24915 16609
rect 24946 16600 24952 16612
rect 25004 16600 25010 16652
rect 25516 16640 25544 16680
rect 26513 16677 26525 16680
rect 26559 16677 26571 16711
rect 26513 16671 26571 16677
rect 25056 16612 25544 16640
rect 25056 16572 25084 16612
rect 25866 16600 25872 16652
rect 25924 16640 25930 16652
rect 26988 16649 27016 16748
rect 28810 16668 28816 16720
rect 28868 16668 28874 16720
rect 29104 16708 29132 16748
rect 29178 16736 29184 16788
rect 29236 16736 29242 16788
rect 29914 16776 29920 16788
rect 29564 16748 29920 16776
rect 29564 16708 29592 16748
rect 29914 16736 29920 16748
rect 29972 16736 29978 16788
rect 30374 16736 30380 16788
rect 30432 16736 30438 16788
rect 29104 16680 29592 16708
rect 29638 16668 29644 16720
rect 29696 16708 29702 16720
rect 29696 16680 31156 16708
rect 29696 16668 29702 16680
rect 26973 16643 27031 16649
rect 26973 16640 26985 16643
rect 25924 16612 26985 16640
rect 25924 16600 25930 16612
rect 26973 16609 26985 16612
rect 27019 16609 27031 16643
rect 26973 16603 27031 16609
rect 27341 16643 27399 16649
rect 27341 16609 27353 16643
rect 27387 16640 27399 16643
rect 27430 16640 27436 16652
rect 27387 16612 27436 16640
rect 27387 16609 27399 16612
rect 27341 16603 27399 16609
rect 27430 16600 27436 16612
rect 27488 16600 27494 16652
rect 27668 16643 27726 16649
rect 27668 16609 27680 16643
rect 27714 16640 27726 16643
rect 27714 16612 28028 16640
rect 27714 16609 27726 16612
rect 27668 16603 27726 16609
rect 27890 16583 27896 16584
rect 24636 16532 24642 16546
rect 24780 16544 25084 16572
rect 27847 16577 27896 16583
rect 27847 16543 27859 16577
rect 27893 16543 27896 16577
rect 27847 16537 27896 16543
rect 27890 16532 27896 16537
rect 27948 16532 27954 16584
rect 28000 16572 28028 16612
rect 28074 16600 28080 16652
rect 28132 16600 28138 16652
rect 28166 16600 28172 16652
rect 28224 16600 28230 16652
rect 28828 16640 28856 16668
rect 29840 16649 29868 16680
rect 31128 16652 31156 16680
rect 29825 16643 29883 16649
rect 28828 16612 29684 16640
rect 28184 16572 28212 16600
rect 29656 16581 29684 16612
rect 29825 16609 29837 16643
rect 29871 16609 29883 16643
rect 29825 16603 29883 16609
rect 29917 16643 29975 16649
rect 29917 16609 29929 16643
rect 29963 16640 29975 16643
rect 30282 16640 30288 16652
rect 29963 16612 30288 16640
rect 29963 16609 29975 16612
rect 29917 16603 29975 16609
rect 30282 16600 30288 16612
rect 30340 16600 30346 16652
rect 30374 16600 30380 16652
rect 30432 16640 30438 16652
rect 30561 16643 30619 16649
rect 30561 16640 30573 16643
rect 30432 16612 30573 16640
rect 30432 16600 30438 16612
rect 30561 16609 30573 16612
rect 30607 16609 30619 16643
rect 30561 16603 30619 16609
rect 31110 16600 31116 16652
rect 31168 16600 31174 16652
rect 28000 16544 28212 16572
rect 29641 16575 29699 16581
rect 29641 16541 29653 16575
rect 29687 16541 29699 16575
rect 29641 16535 29699 16541
rect 22830 16464 22836 16516
rect 22888 16504 22894 16516
rect 22888 16476 23704 16504
rect 22888 16464 22894 16476
rect 21324 16408 22692 16436
rect 21324 16396 21330 16408
rect 22738 16396 22744 16448
rect 22796 16396 22802 16448
rect 23477 16439 23535 16445
rect 23477 16405 23489 16439
rect 23523 16436 23535 16439
rect 23566 16436 23572 16448
rect 23523 16408 23572 16436
rect 23523 16405 23535 16408
rect 23477 16399 23535 16405
rect 23566 16396 23572 16408
rect 23624 16396 23630 16448
rect 23676 16436 23704 16476
rect 23750 16464 23756 16516
rect 23808 16504 23814 16516
rect 23934 16504 23940 16516
rect 23808 16476 23940 16504
rect 23808 16464 23814 16476
rect 23934 16464 23940 16476
rect 23992 16464 23998 16516
rect 25961 16507 26019 16513
rect 25961 16473 25973 16507
rect 26007 16473 26019 16507
rect 25961 16467 26019 16473
rect 26068 16476 27292 16504
rect 25976 16436 26004 16467
rect 26068 16448 26096 16476
rect 23676 16408 26004 16436
rect 26050 16396 26056 16448
rect 26108 16396 26114 16448
rect 26326 16396 26332 16448
rect 26384 16436 26390 16448
rect 26786 16436 26792 16448
rect 26384 16408 26792 16436
rect 26384 16396 26390 16408
rect 26786 16396 26792 16408
rect 26844 16396 26850 16448
rect 27154 16396 27160 16448
rect 27212 16396 27218 16448
rect 27264 16436 27292 16476
rect 30193 16439 30251 16445
rect 30193 16436 30205 16439
rect 27264 16408 30205 16436
rect 30193 16405 30205 16408
rect 30239 16405 30251 16439
rect 30193 16399 30251 16405
rect 552 16346 30912 16368
rect 552 16294 4193 16346
rect 4245 16294 4257 16346
rect 4309 16294 4321 16346
rect 4373 16294 4385 16346
rect 4437 16294 4449 16346
rect 4501 16294 11783 16346
rect 11835 16294 11847 16346
rect 11899 16294 11911 16346
rect 11963 16294 11975 16346
rect 12027 16294 12039 16346
rect 12091 16294 19373 16346
rect 19425 16294 19437 16346
rect 19489 16294 19501 16346
rect 19553 16294 19565 16346
rect 19617 16294 19629 16346
rect 19681 16294 26963 16346
rect 27015 16294 27027 16346
rect 27079 16294 27091 16346
rect 27143 16294 27155 16346
rect 27207 16294 27219 16346
rect 27271 16294 30912 16346
rect 552 16272 30912 16294
rect 2038 16192 2044 16244
rect 2096 16232 2102 16244
rect 2777 16235 2835 16241
rect 2777 16232 2789 16235
rect 2096 16204 2789 16232
rect 2096 16192 2102 16204
rect 2777 16201 2789 16204
rect 2823 16201 2835 16235
rect 2777 16195 2835 16201
rect 4246 16192 4252 16244
rect 4304 16232 4310 16244
rect 4614 16232 4620 16244
rect 4304 16204 4620 16232
rect 4304 16192 4310 16204
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 4706 16192 4712 16244
rect 4764 16232 4770 16244
rect 5629 16235 5687 16241
rect 5629 16232 5641 16235
rect 4764 16204 5641 16232
rect 4764 16192 4770 16204
rect 5629 16201 5641 16204
rect 5675 16201 5687 16235
rect 7929 16235 7987 16241
rect 7929 16232 7941 16235
rect 5629 16195 5687 16201
rect 6104 16204 7941 16232
rect 4295 16099 4353 16105
rect 1412 16081 4200 16096
rect 1412 16050 1445 16081
rect 1433 16047 1445 16050
rect 1479 16068 4200 16081
rect 1479 16047 1491 16068
rect 1433 16041 1491 16047
rect 937 16031 995 16037
rect 937 15997 949 16031
rect 983 16028 995 16031
rect 1302 16028 1308 16040
rect 983 16000 1308 16028
rect 983 15997 995 16000
rect 937 15991 995 15997
rect 1302 15988 1308 16000
rect 1360 15988 1366 16040
rect 1673 16031 1731 16037
rect 1673 15997 1685 16031
rect 1719 16028 1731 16031
rect 2498 16028 2504 16040
rect 1719 16000 2504 16028
rect 1719 15997 1731 16000
rect 1673 15991 1731 15997
rect 2498 15988 2504 16000
rect 2556 15988 2562 16040
rect 3326 15988 3332 16040
rect 3384 15988 3390 16040
rect 3789 16031 3847 16037
rect 3789 16028 3801 16031
rect 3620 16000 3801 16028
rect 3620 15904 3648 16000
rect 3789 15997 3801 16000
rect 3835 15997 3847 16031
rect 4172 16028 4200 16068
rect 4295 16065 4307 16099
rect 4341 16096 4353 16099
rect 6104 16096 6132 16204
rect 7929 16201 7941 16204
rect 7975 16201 7987 16235
rect 9766 16232 9772 16244
rect 7929 16195 7987 16201
rect 8588 16204 9772 16232
rect 4341 16068 6132 16096
rect 4341 16065 4353 16068
rect 4295 16059 4353 16065
rect 6454 16056 6460 16108
rect 6512 16096 6518 16108
rect 6595 16097 6653 16103
rect 6595 16096 6607 16097
rect 6512 16068 6607 16096
rect 6512 16056 6518 16068
rect 6595 16063 6607 16068
rect 6641 16063 6653 16097
rect 6595 16057 6653 16063
rect 4430 16028 4436 16040
rect 4172 16000 4436 16028
rect 3789 15991 3847 15997
rect 4430 15988 4436 16000
rect 4488 15988 4494 16040
rect 4522 15988 4528 16040
rect 4580 15988 4586 16040
rect 6086 15988 6092 16040
rect 6144 15988 6150 16040
rect 8588 16037 8616 16204
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 13078 16232 13084 16244
rect 10796 16204 13084 16232
rect 9171 16099 9229 16105
rect 9171 16065 9183 16099
rect 9217 16096 9229 16099
rect 10796 16096 10824 16204
rect 13078 16192 13084 16204
rect 13136 16192 13142 16244
rect 14366 16192 14372 16244
rect 14424 16232 14430 16244
rect 14826 16232 14832 16244
rect 14424 16204 14832 16232
rect 14424 16192 14430 16204
rect 14826 16192 14832 16204
rect 14884 16192 14890 16244
rect 18230 16232 18236 16244
rect 16040 16204 18236 16232
rect 10962 16124 10968 16176
rect 11020 16124 11026 16176
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 11112 16136 11192 16164
rect 11112 16124 11118 16136
rect 9217 16068 10824 16096
rect 9217 16065 9229 16068
rect 9171 16059 9229 16065
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6196 16000 6837 16028
rect 5258 15920 5264 15972
rect 5316 15960 5322 15972
rect 6196 15960 6224 16000
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 6825 15991 6883 15997
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 15997 8631 16031
rect 8573 15991 8631 15997
rect 8662 15988 8668 16040
rect 8720 15988 8726 16040
rect 8938 15988 8944 16040
rect 8996 16028 9002 16040
rect 9401 16031 9459 16037
rect 9401 16028 9413 16031
rect 8996 16000 9413 16028
rect 8996 15988 9002 16000
rect 9401 15997 9413 16000
rect 9447 15997 9459 16031
rect 9401 15991 9459 15997
rect 9858 15988 9864 16040
rect 9916 16028 9922 16040
rect 11164 16037 11192 16136
rect 11241 16099 11299 16105
rect 11241 16065 11253 16099
rect 11287 16096 11299 16099
rect 11514 16096 11520 16108
rect 11287 16068 11520 16096
rect 11287 16065 11299 16068
rect 11241 16059 11299 16065
rect 11514 16056 11520 16068
rect 11572 16056 11578 16108
rect 11698 16056 11704 16108
rect 11756 16094 11762 16108
rect 11756 16066 11799 16094
rect 11900 16068 13676 16096
rect 11756 16056 11762 16066
rect 11149 16031 11207 16037
rect 9916 16000 11100 16028
rect 9916 15988 9922 16000
rect 5316 15932 6224 15960
rect 8312 15932 8800 15960
rect 5316 15920 5322 15932
rect 1394 15852 1400 15904
rect 1452 15901 1458 15904
rect 1452 15892 1461 15901
rect 1452 15864 1497 15892
rect 1452 15855 1461 15864
rect 1452 15852 1458 15855
rect 3602 15852 3608 15904
rect 3660 15852 3666 15904
rect 3878 15852 3884 15904
rect 3936 15892 3942 15904
rect 4255 15895 4313 15901
rect 4255 15892 4267 15895
rect 3936 15864 4267 15892
rect 3936 15852 3942 15864
rect 4255 15861 4267 15864
rect 4301 15861 4313 15895
rect 4255 15855 4313 15861
rect 6454 15852 6460 15904
rect 6512 15892 6518 15904
rect 6555 15895 6613 15901
rect 6555 15892 6567 15895
rect 6512 15864 6567 15892
rect 6512 15852 6518 15864
rect 6555 15861 6567 15864
rect 6601 15892 6613 15895
rect 8312 15892 8340 15932
rect 6601 15864 8340 15892
rect 6601 15861 6613 15864
rect 6555 15855 6613 15861
rect 8386 15852 8392 15904
rect 8444 15852 8450 15904
rect 8772 15892 8800 15932
rect 9030 15892 9036 15904
rect 8772 15864 9036 15892
rect 9030 15852 9036 15864
rect 9088 15892 9094 15904
rect 9131 15895 9189 15901
rect 9131 15892 9143 15895
rect 9088 15864 9143 15892
rect 9088 15852 9094 15864
rect 9131 15861 9143 15864
rect 9177 15861 9189 15895
rect 9131 15855 9189 15861
rect 10502 15852 10508 15904
rect 10560 15852 10566 15904
rect 11072 15892 11100 16000
rect 11149 15997 11161 16031
rect 11195 15997 11207 16031
rect 11532 16028 11560 16056
rect 11900 16028 11928 16068
rect 11532 16000 11928 16028
rect 11977 16031 12035 16037
rect 11149 15991 11207 15997
rect 11977 15997 11989 16031
rect 12023 16028 12035 16031
rect 12710 16028 12716 16040
rect 12023 16000 12716 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 12710 15988 12716 16000
rect 12768 15988 12774 16040
rect 13648 16037 13676 16068
rect 14550 16056 14556 16108
rect 14608 16056 14614 16108
rect 14691 16099 14749 16105
rect 14691 16065 14703 16099
rect 14737 16096 14749 16099
rect 16040 16096 16068 16204
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 19794 16232 19800 16244
rect 19628 16204 19800 16232
rect 14737 16068 16068 16096
rect 14737 16065 14749 16068
rect 14691 16059 14749 16065
rect 16114 16056 16120 16108
rect 16172 16096 16178 16108
rect 16899 16099 16957 16105
rect 16172 16068 16712 16096
rect 16172 16056 16178 16068
rect 13633 16031 13691 16037
rect 13633 15997 13645 16031
rect 13679 15997 13691 16031
rect 14185 16031 14243 16037
rect 14185 16028 14197 16031
rect 13633 15991 13691 15997
rect 14016 16000 14197 16028
rect 14016 15904 14044 16000
rect 14185 15997 14197 16000
rect 14231 15997 14243 16031
rect 14568 16028 14596 16056
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 14568 16000 14933 16028
rect 14185 15991 14243 15997
rect 14921 15997 14933 16000
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 16393 16031 16451 16037
rect 16393 15997 16405 16031
rect 16439 16028 16451 16031
rect 16482 16028 16488 16040
rect 16439 16000 16488 16028
rect 16439 15997 16451 16000
rect 16393 15991 16451 15997
rect 16482 15988 16488 16000
rect 16540 15988 16546 16040
rect 16684 16028 16712 16068
rect 16899 16065 16911 16099
rect 16945 16096 16957 16099
rect 17862 16096 17868 16108
rect 16945 16068 17868 16096
rect 16945 16065 16957 16068
rect 16899 16059 16957 16065
rect 17862 16056 17868 16068
rect 17920 16056 17926 16108
rect 19628 16105 19656 16204
rect 19794 16192 19800 16204
rect 19852 16232 19858 16244
rect 20346 16232 20352 16244
rect 19852 16204 20352 16232
rect 19852 16192 19858 16204
rect 20346 16192 20352 16204
rect 20404 16192 20410 16244
rect 23385 16235 23443 16241
rect 23385 16201 23397 16235
rect 23431 16232 23443 16235
rect 26602 16232 26608 16244
rect 23431 16204 26608 16232
rect 23431 16201 23443 16204
rect 23385 16195 23443 16201
rect 26602 16192 26608 16204
rect 26660 16192 26666 16244
rect 26786 16192 26792 16244
rect 26844 16232 26850 16244
rect 27706 16232 27712 16244
rect 26844 16204 27712 16232
rect 26844 16192 26850 16204
rect 27706 16192 27712 16204
rect 27764 16192 27770 16244
rect 30374 16232 30380 16244
rect 28966 16204 30380 16232
rect 25685 16167 25743 16173
rect 25685 16133 25697 16167
rect 25731 16133 25743 16167
rect 25685 16127 25743 16133
rect 19978 16105 19984 16108
rect 19613 16099 19671 16105
rect 19613 16096 19625 16099
rect 19168 16068 19625 16096
rect 17129 16031 17187 16037
rect 17129 16028 17141 16031
rect 16684 16000 17141 16028
rect 17129 15997 17141 16000
rect 17175 15997 17187 16031
rect 17129 15991 17187 15997
rect 17218 15988 17224 16040
rect 17276 16028 17282 16040
rect 19168 16037 19196 16068
rect 19613 16065 19625 16068
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 19940 16099 19984 16105
rect 19940 16065 19952 16099
rect 19940 16059 19984 16065
rect 19978 16056 19984 16059
rect 20036 16056 20042 16108
rect 20088 16081 20944 16096
rect 20088 16050 20121 16081
rect 20109 16047 20121 16050
rect 20155 16068 20944 16081
rect 20155 16047 20167 16068
rect 20109 16041 20167 16047
rect 18785 16031 18843 16037
rect 18785 16028 18797 16031
rect 17276 16000 18797 16028
rect 17276 15988 17282 16000
rect 18785 15997 18797 16000
rect 18831 15997 18843 16031
rect 18785 15991 18843 15997
rect 19153 16031 19211 16037
rect 19153 15997 19165 16031
rect 19199 15997 19211 16031
rect 19153 15991 19211 15997
rect 19426 15988 19432 16040
rect 19484 15988 19490 16040
rect 20254 15988 20260 16040
rect 20312 16028 20318 16040
rect 20349 16031 20407 16037
rect 20349 16028 20361 16031
rect 20312 16000 20361 16028
rect 20312 15988 20318 16000
rect 20349 15997 20361 16000
rect 20395 15997 20407 16031
rect 20916 16028 20944 16068
rect 20990 16056 20996 16108
rect 21048 16096 21054 16108
rect 22097 16099 22155 16105
rect 22097 16096 22109 16099
rect 21048 16068 22109 16096
rect 21048 16056 21054 16068
rect 22097 16065 22109 16068
rect 22143 16065 22155 16099
rect 22097 16059 22155 16065
rect 22278 16056 22284 16108
rect 22336 16056 22342 16108
rect 23750 16056 23756 16108
rect 23808 16096 23814 16108
rect 24210 16096 24216 16108
rect 23808 16068 24216 16096
rect 23808 16056 23814 16068
rect 24210 16056 24216 16068
rect 24268 16056 24274 16108
rect 24308 16097 24366 16103
rect 24308 16063 24320 16097
rect 24354 16096 24366 16097
rect 24394 16096 24400 16108
rect 24354 16068 24400 16096
rect 24354 16063 24366 16068
rect 24308 16057 24366 16063
rect 24394 16056 24400 16068
rect 24452 16056 24458 16108
rect 25700 16096 25728 16127
rect 24504 16068 25728 16096
rect 26559 16099 26617 16105
rect 21821 16031 21879 16037
rect 20916 16000 21588 16028
rect 20349 15991 20407 15997
rect 11146 15892 11152 15904
rect 11072 15864 11152 15892
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 11707 15895 11765 15901
rect 11707 15861 11719 15895
rect 11753 15892 11765 15895
rect 11882 15892 11888 15904
rect 11753 15864 11888 15892
rect 11753 15861 11765 15864
rect 11707 15855 11765 15861
rect 11882 15852 11888 15864
rect 11940 15892 11946 15904
rect 12066 15892 12072 15904
rect 11940 15864 12072 15892
rect 11940 15852 11946 15864
rect 12066 15852 12072 15864
rect 12124 15852 12130 15904
rect 13078 15852 13084 15904
rect 13136 15852 13142 15904
rect 13909 15895 13967 15901
rect 13909 15861 13921 15895
rect 13955 15892 13967 15895
rect 13998 15892 14004 15904
rect 13955 15864 14004 15892
rect 13955 15861 13967 15864
rect 13909 15855 13967 15861
rect 13998 15852 14004 15864
rect 14056 15852 14062 15904
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 14458 15892 14464 15904
rect 14240 15864 14464 15892
rect 14240 15852 14246 15864
rect 14458 15852 14464 15864
rect 14516 15892 14522 15904
rect 14651 15895 14709 15901
rect 14651 15892 14663 15895
rect 14516 15864 14663 15892
rect 14516 15852 14522 15864
rect 14651 15861 14663 15864
rect 14697 15892 14709 15895
rect 14918 15892 14924 15904
rect 14697 15864 14924 15892
rect 14697 15861 14709 15864
rect 14651 15855 14709 15861
rect 14918 15852 14924 15864
rect 14976 15852 14982 15904
rect 15286 15852 15292 15904
rect 15344 15892 15350 15904
rect 16025 15895 16083 15901
rect 16025 15892 16037 15895
rect 15344 15864 16037 15892
rect 15344 15852 15350 15864
rect 16025 15861 16037 15864
rect 16071 15861 16083 15895
rect 16025 15855 16083 15861
rect 16758 15852 16764 15904
rect 16816 15892 16822 15904
rect 16859 15895 16917 15901
rect 16859 15892 16871 15895
rect 16816 15864 16871 15892
rect 16816 15852 16822 15864
rect 16859 15861 16871 15864
rect 16905 15892 16917 15895
rect 17034 15892 17040 15904
rect 16905 15864 17040 15892
rect 16905 15861 16917 15864
rect 16859 15855 16917 15861
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 17126 15852 17132 15904
rect 17184 15892 17190 15904
rect 18233 15895 18291 15901
rect 18233 15892 18245 15895
rect 17184 15864 18245 15892
rect 17184 15852 17190 15864
rect 18233 15861 18245 15864
rect 18279 15861 18291 15895
rect 18233 15855 18291 15861
rect 19242 15852 19248 15904
rect 19300 15852 19306 15904
rect 20346 15852 20352 15904
rect 20404 15892 20410 15904
rect 21453 15895 21511 15901
rect 21453 15892 21465 15895
rect 20404 15864 21465 15892
rect 20404 15852 20410 15864
rect 21453 15861 21465 15864
rect 21499 15861 21511 15895
rect 21560 15892 21588 16000
rect 21821 15997 21833 16031
rect 21867 16028 21879 16031
rect 22296 16028 22324 16056
rect 21867 16000 22324 16028
rect 21867 15997 21879 16000
rect 21821 15991 21879 15997
rect 22738 15988 22744 16040
rect 22796 16028 22802 16040
rect 23474 16028 23480 16040
rect 22796 16000 23480 16028
rect 22796 15988 22802 16000
rect 23474 15988 23480 16000
rect 23532 15988 23538 16040
rect 23658 15988 23664 16040
rect 23716 16028 23722 16040
rect 23842 16028 23848 16040
rect 23716 16000 23848 16028
rect 23716 15988 23722 16000
rect 23842 15988 23848 16000
rect 23900 15988 23906 16040
rect 24504 16028 24532 16068
rect 26559 16065 26571 16099
rect 26605 16096 26617 16099
rect 28258 16096 28264 16108
rect 26605 16068 28264 16096
rect 26605 16065 26617 16068
rect 26559 16059 26617 16065
rect 28258 16056 28264 16068
rect 28316 16056 28322 16108
rect 23952 16000 24532 16028
rect 23952 15960 23980 16000
rect 24578 15988 24584 16040
rect 24636 15988 24642 16040
rect 25958 15988 25964 16040
rect 26016 16028 26022 16040
rect 26053 16031 26111 16037
rect 26053 16028 26065 16031
rect 26016 16000 26065 16028
rect 26016 15988 26022 16000
rect 26053 15997 26065 16000
rect 26099 15997 26111 16031
rect 26053 15991 26111 15997
rect 26380 16031 26438 16037
rect 26380 15997 26392 16031
rect 26426 16028 26438 16031
rect 26694 16028 26700 16040
rect 26426 16000 26700 16028
rect 26426 15997 26438 16000
rect 26380 15991 26438 15997
rect 23124 15932 23980 15960
rect 23124 15892 23152 15932
rect 21560 15864 23152 15892
rect 21453 15855 21511 15861
rect 23842 15852 23848 15904
rect 23900 15892 23906 15904
rect 24302 15892 24308 15904
rect 24360 15901 24366 15904
rect 23900 15864 24308 15892
rect 23900 15852 23906 15864
rect 24302 15852 24308 15864
rect 24360 15892 24369 15901
rect 26068 15892 26096 15991
rect 26694 15988 26700 16000
rect 26752 15988 26758 16040
rect 26786 15988 26792 16040
rect 26844 15988 26850 16040
rect 27246 15988 27252 16040
rect 27304 16028 27310 16040
rect 27430 16028 27436 16040
rect 27304 16000 27436 16028
rect 27304 15988 27310 16000
rect 27430 15988 27436 16000
rect 27488 15988 27494 16040
rect 28353 16031 28411 16037
rect 28353 16028 28365 16031
rect 27816 16000 28365 16028
rect 27816 15972 27844 16000
rect 28353 15997 28365 16000
rect 28399 15997 28411 16031
rect 28353 15991 28411 15997
rect 27798 15920 27804 15972
rect 27856 15920 27862 15972
rect 26326 15892 26332 15904
rect 24360 15864 24405 15892
rect 26068 15864 26332 15892
rect 24360 15855 24369 15864
rect 24360 15852 24366 15855
rect 26326 15852 26332 15864
rect 26384 15852 26390 15904
rect 26694 15852 26700 15904
rect 26752 15892 26758 15904
rect 27893 15895 27951 15901
rect 27893 15892 27905 15895
rect 26752 15864 27905 15892
rect 26752 15852 26758 15864
rect 27893 15861 27905 15864
rect 27939 15861 27951 15895
rect 27893 15855 27951 15861
rect 28629 15895 28687 15901
rect 28629 15861 28641 15895
rect 28675 15892 28687 15895
rect 28810 15892 28816 15904
rect 28675 15864 28816 15892
rect 28675 15861 28687 15864
rect 28629 15855 28687 15861
rect 28810 15852 28816 15864
rect 28868 15892 28874 15904
rect 28966 15892 28994 16204
rect 30374 16192 30380 16204
rect 30432 16192 30438 16244
rect 30466 16192 30472 16244
rect 30524 16192 30530 16244
rect 30484 16164 30512 16192
rect 29104 16136 30512 16164
rect 29104 15960 29132 16136
rect 30098 16056 30104 16108
rect 30156 16056 30162 16108
rect 29178 15988 29184 16040
rect 29236 16028 29242 16040
rect 29730 16028 29736 16040
rect 29236 16000 29736 16028
rect 29236 15988 29242 16000
rect 29730 15988 29736 16000
rect 29788 15988 29794 16040
rect 29825 16031 29883 16037
rect 29825 15997 29837 16031
rect 29871 16028 29883 16031
rect 30190 16028 30196 16040
rect 29871 16000 30196 16028
rect 29871 15997 29883 16000
rect 29825 15991 29883 15997
rect 30190 15988 30196 16000
rect 30248 15988 30254 16040
rect 30285 16031 30343 16037
rect 30285 15997 30297 16031
rect 30331 15997 30343 16031
rect 30285 15991 30343 15997
rect 29273 15963 29331 15969
rect 29273 15960 29285 15963
rect 29104 15932 29285 15960
rect 29273 15929 29285 15932
rect 29319 15929 29331 15963
rect 29748 15960 29776 15988
rect 30300 15960 30328 15991
rect 29748 15932 30328 15960
rect 29273 15923 29331 15929
rect 28868 15864 28994 15892
rect 29549 15895 29607 15901
rect 28868 15852 28874 15864
rect 29549 15861 29561 15895
rect 29595 15892 29607 15895
rect 30190 15892 30196 15904
rect 29595 15864 30196 15892
rect 29595 15861 29607 15864
rect 29549 15855 29607 15861
rect 30190 15852 30196 15864
rect 30248 15852 30254 15904
rect 30466 15852 30472 15904
rect 30524 15852 30530 15904
rect 552 15802 31072 15824
rect 552 15750 7988 15802
rect 8040 15750 8052 15802
rect 8104 15750 8116 15802
rect 8168 15750 8180 15802
rect 8232 15750 8244 15802
rect 8296 15750 15578 15802
rect 15630 15750 15642 15802
rect 15694 15750 15706 15802
rect 15758 15750 15770 15802
rect 15822 15750 15834 15802
rect 15886 15750 23168 15802
rect 23220 15750 23232 15802
rect 23284 15750 23296 15802
rect 23348 15750 23360 15802
rect 23412 15750 23424 15802
rect 23476 15750 30758 15802
rect 30810 15750 30822 15802
rect 30874 15750 30886 15802
rect 30938 15750 30950 15802
rect 31002 15750 31014 15802
rect 31066 15750 31072 15802
rect 552 15728 31072 15750
rect 1394 15648 1400 15700
rect 1452 15688 1458 15700
rect 1771 15691 1829 15697
rect 1771 15688 1783 15691
rect 1452 15660 1783 15688
rect 1452 15648 1458 15660
rect 1771 15657 1783 15660
rect 1817 15657 1829 15691
rect 1771 15651 1829 15657
rect 3142 15648 3148 15700
rect 3200 15648 3206 15700
rect 13078 15688 13084 15700
rect 3436 15660 4936 15688
rect 1121 15555 1179 15561
rect 1121 15521 1133 15555
rect 1167 15552 1179 15555
rect 3436 15552 3464 15660
rect 4908 15620 4936 15660
rect 5460 15660 7972 15688
rect 5460 15620 5488 15660
rect 7944 15632 7972 15660
rect 8312 15660 13084 15688
rect 4908 15592 5488 15620
rect 5626 15580 5632 15632
rect 5684 15580 5690 15632
rect 6454 15580 6460 15632
rect 6512 15580 6518 15632
rect 7926 15580 7932 15632
rect 7984 15580 7990 15632
rect 1167 15524 1716 15552
rect 1167 15521 1179 15524
rect 1121 15515 1179 15521
rect 1688 15496 1716 15524
rect 1964 15524 3464 15552
rect 3513 15555 3571 15561
rect 1801 15505 1859 15511
rect 1305 15487 1363 15493
rect 1305 15453 1317 15487
rect 1351 15453 1363 15487
rect 1305 15447 1363 15453
rect 1320 15360 1348 15447
rect 1670 15444 1676 15496
rect 1728 15444 1734 15496
rect 1801 15471 1813 15505
rect 1847 15484 1859 15505
rect 1964 15484 1992 15524
rect 3513 15521 3525 15555
rect 3559 15552 3571 15555
rect 3602 15552 3608 15564
rect 3559 15524 3608 15552
rect 3559 15521 3571 15524
rect 3513 15515 3571 15521
rect 1847 15471 1992 15484
rect 1801 15465 1992 15471
rect 1826 15456 1992 15465
rect 2041 15487 2099 15493
rect 2041 15453 2053 15487
rect 2087 15484 2099 15487
rect 2406 15484 2412 15496
rect 2087 15456 2412 15484
rect 2087 15453 2099 15456
rect 2041 15447 2099 15453
rect 2406 15444 2412 15456
rect 2464 15444 2470 15496
rect 934 15308 940 15360
rect 992 15308 998 15360
rect 1302 15308 1308 15360
rect 1360 15348 1366 15360
rect 3528 15348 3556 15515
rect 3602 15512 3608 15524
rect 3660 15512 3666 15564
rect 4246 15512 4252 15564
rect 4304 15512 4310 15564
rect 4338 15512 4344 15564
rect 4396 15552 4402 15564
rect 5905 15555 5963 15561
rect 5905 15552 5917 15555
rect 4396 15524 5917 15552
rect 4396 15512 4402 15524
rect 5905 15521 5917 15524
rect 5951 15521 5963 15555
rect 6472 15552 6500 15580
rect 6784 15555 6842 15561
rect 6784 15552 6796 15555
rect 6472 15524 6796 15552
rect 5905 15515 5963 15521
rect 6784 15521 6796 15524
rect 6830 15521 6842 15555
rect 8312 15552 8340 15660
rect 13078 15648 13084 15660
rect 13136 15648 13142 15700
rect 13446 15648 13452 15700
rect 13504 15688 13510 15700
rect 15657 15691 15715 15697
rect 15657 15688 15669 15691
rect 13504 15660 15669 15688
rect 13504 15648 13510 15660
rect 15657 15657 15669 15660
rect 15703 15657 15715 15691
rect 15657 15651 15715 15657
rect 15930 15648 15936 15700
rect 15988 15648 15994 15700
rect 16390 15648 16396 15700
rect 16448 15688 16454 15700
rect 18782 15688 18788 15700
rect 16448 15660 18788 15688
rect 16448 15648 16454 15660
rect 18782 15648 18788 15660
rect 18840 15648 18846 15700
rect 20346 15648 20352 15700
rect 20404 15648 20410 15700
rect 23109 15691 23167 15697
rect 23109 15688 23121 15691
rect 20824 15660 23121 15688
rect 11330 15580 11336 15632
rect 11388 15620 11394 15632
rect 11425 15623 11483 15629
rect 11425 15620 11437 15623
rect 11388 15592 11437 15620
rect 11388 15580 11394 15592
rect 11425 15589 11437 15592
rect 11471 15620 11483 15623
rect 11514 15620 11520 15632
rect 11471 15592 11520 15620
rect 11471 15589 11483 15592
rect 11425 15583 11483 15589
rect 6784 15515 6842 15521
rect 7116 15524 8340 15552
rect 6953 15505 7011 15511
rect 3878 15493 3884 15496
rect 3840 15487 3884 15493
rect 3840 15453 3852 15487
rect 3840 15447 3884 15453
rect 3878 15444 3884 15447
rect 3936 15444 3942 15496
rect 4019 15487 4077 15493
rect 4019 15453 4031 15487
rect 4065 15484 4077 15487
rect 5994 15484 6000 15496
rect 4065 15456 6000 15484
rect 4065 15453 4077 15456
rect 4019 15447 4077 15453
rect 5994 15444 6000 15456
rect 6052 15444 6058 15496
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15453 6515 15487
rect 6953 15471 6965 15505
rect 6999 15484 7011 15505
rect 7116 15484 7144 15524
rect 8386 15512 8392 15564
rect 8444 15552 8450 15564
rect 9401 15555 9459 15561
rect 9401 15552 9413 15555
rect 8444 15524 9413 15552
rect 8444 15512 8450 15524
rect 9401 15521 9413 15524
rect 9447 15521 9459 15555
rect 9401 15515 9459 15521
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15521 11115 15555
rect 11057 15515 11115 15521
rect 6999 15471 7144 15484
rect 6953 15465 7144 15471
rect 6968 15456 7144 15465
rect 6457 15447 6515 15453
rect 6086 15376 6092 15428
rect 6144 15416 6150 15428
rect 6181 15419 6239 15425
rect 6181 15416 6193 15419
rect 6144 15388 6193 15416
rect 6144 15376 6150 15388
rect 6181 15385 6193 15388
rect 6227 15416 6239 15419
rect 6472 15416 6500 15447
rect 7190 15444 7196 15496
rect 7248 15444 7254 15496
rect 9030 15493 9036 15496
rect 8665 15487 8723 15493
rect 8665 15453 8677 15487
rect 8711 15453 8723 15487
rect 8665 15447 8723 15453
rect 8992 15487 9036 15493
rect 8992 15453 9004 15487
rect 8992 15447 9036 15453
rect 8680 15416 8708 15447
rect 9030 15444 9036 15447
rect 9088 15444 9094 15496
rect 9214 15495 9220 15496
rect 9171 15489 9220 15495
rect 9171 15455 9183 15489
rect 9217 15455 9220 15489
rect 9171 15449 9220 15455
rect 9214 15444 9220 15449
rect 9272 15444 9278 15496
rect 9490 15444 9496 15496
rect 9548 15484 9554 15496
rect 10962 15484 10968 15496
rect 9548 15456 10968 15484
rect 9548 15444 9554 15456
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 11072 15416 11100 15515
rect 11443 15484 11471 15583
rect 11514 15580 11520 15592
rect 11572 15580 11578 15632
rect 15948 15620 15976 15648
rect 15948 15592 16712 15620
rect 11882 15561 11888 15564
rect 11844 15555 11888 15561
rect 11844 15521 11856 15555
rect 11844 15515 11888 15521
rect 11882 15512 11888 15515
rect 11940 15512 11946 15564
rect 14458 15552 14464 15564
rect 12176 15524 12434 15552
rect 11517 15487 11575 15493
rect 11517 15484 11529 15487
rect 11443 15456 11529 15484
rect 11517 15453 11529 15456
rect 11563 15453 11575 15487
rect 11517 15447 11575 15453
rect 12023 15487 12081 15493
rect 12023 15453 12035 15487
rect 12069 15484 12081 15487
rect 12176 15484 12204 15524
rect 12069 15456 12204 15484
rect 12069 15453 12081 15456
rect 12023 15447 12081 15453
rect 12250 15444 12256 15496
rect 12308 15444 12314 15496
rect 12406 15484 12434 15524
rect 14159 15524 14464 15552
rect 13817 15487 13875 15493
rect 12406 15456 13676 15484
rect 6227 15388 6500 15416
rect 6227 15385 6239 15388
rect 6181 15379 6239 15385
rect 3786 15348 3792 15360
rect 1360 15320 3792 15348
rect 1360 15308 1366 15320
rect 3786 15308 3792 15320
rect 3844 15348 3850 15360
rect 4338 15348 4344 15360
rect 3844 15320 4344 15348
rect 3844 15308 3850 15320
rect 4338 15308 4344 15320
rect 4396 15308 4402 15360
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 4890 15348 4896 15360
rect 4764 15320 4896 15348
rect 4764 15308 4770 15320
rect 4890 15308 4896 15320
rect 4948 15308 4954 15360
rect 6472 15348 6500 15388
rect 7852 15388 8708 15416
rect 7852 15348 7880 15388
rect 8680 15360 8708 15388
rect 10060 15388 11100 15416
rect 6472 15320 7880 15348
rect 8294 15308 8300 15360
rect 8352 15308 8358 15360
rect 8662 15308 8668 15360
rect 8720 15348 8726 15360
rect 10060 15348 10088 15388
rect 13648 15360 13676 15456
rect 13817 15453 13829 15487
rect 13863 15484 13875 15487
rect 13998 15484 14004 15496
rect 13863 15456 14004 15484
rect 13863 15453 13875 15456
rect 13817 15447 13875 15453
rect 13998 15444 14004 15456
rect 14056 15444 14062 15496
rect 14159 15493 14187 15524
rect 14458 15512 14464 15524
rect 14516 15512 14522 15564
rect 14550 15512 14556 15564
rect 14608 15512 14614 15564
rect 14826 15512 14832 15564
rect 14884 15552 14890 15564
rect 16301 15555 16359 15561
rect 16301 15552 16313 15555
rect 14884 15524 16313 15552
rect 14884 15512 14890 15524
rect 16301 15521 16313 15524
rect 16347 15521 16359 15555
rect 16301 15515 16359 15521
rect 16574 15512 16580 15564
rect 16632 15512 16638 15564
rect 14144 15487 14202 15493
rect 14144 15453 14156 15487
rect 14190 15453 14202 15487
rect 14144 15447 14202 15453
rect 14323 15487 14381 15493
rect 14323 15453 14335 15487
rect 14369 15484 14381 15487
rect 16390 15484 16396 15496
rect 14369 15456 16396 15484
rect 14369 15453 14381 15456
rect 14323 15447 14381 15453
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 13722 15376 13728 15428
rect 13780 15376 13786 15428
rect 15204 15388 15792 15416
rect 8720 15320 10088 15348
rect 8720 15308 8726 15320
rect 10134 15308 10140 15360
rect 10192 15348 10198 15360
rect 10505 15351 10563 15357
rect 10505 15348 10517 15351
rect 10192 15320 10517 15348
rect 10192 15308 10198 15320
rect 10505 15317 10517 15320
rect 10551 15317 10563 15351
rect 10505 15311 10563 15317
rect 11054 15308 11060 15360
rect 11112 15348 11118 15360
rect 12158 15348 12164 15360
rect 11112 15320 12164 15348
rect 11112 15308 11118 15320
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 13354 15308 13360 15360
rect 13412 15308 13418 15360
rect 13630 15308 13636 15360
rect 13688 15308 13694 15360
rect 13740 15348 13768 15376
rect 15204 15348 15232 15388
rect 13740 15320 15232 15348
rect 15764 15348 15792 15388
rect 16114 15376 16120 15428
rect 16172 15376 16178 15428
rect 16684 15357 16712 15592
rect 17034 15580 17040 15632
rect 17092 15580 17098 15632
rect 16853 15555 16911 15561
rect 16853 15521 16865 15555
rect 16899 15521 16911 15555
rect 17052 15552 17080 15580
rect 17364 15555 17422 15561
rect 17364 15552 17376 15555
rect 17052 15524 17376 15552
rect 16853 15515 16911 15521
rect 17364 15521 17376 15524
rect 17410 15521 17422 15555
rect 20364 15552 20392 15648
rect 17364 15515 17422 15521
rect 17696 15524 20392 15552
rect 16868 15428 16896 15515
rect 17037 15487 17095 15493
rect 17037 15453 17049 15487
rect 17083 15484 17095 15487
rect 17218 15484 17224 15496
rect 17083 15456 17224 15484
rect 17083 15453 17095 15456
rect 17037 15447 17095 15453
rect 17218 15444 17224 15456
rect 17276 15444 17282 15496
rect 17543 15487 17601 15493
rect 17543 15453 17555 15487
rect 17589 15484 17601 15487
rect 17696 15484 17724 15524
rect 20714 15512 20720 15564
rect 20772 15512 20778 15564
rect 17589 15456 17724 15484
rect 17773 15487 17831 15493
rect 17589 15453 17601 15456
rect 17543 15447 17601 15453
rect 17773 15453 17785 15487
rect 17819 15484 17831 15487
rect 18966 15484 18972 15496
rect 17819 15456 18972 15484
rect 17819 15453 17831 15456
rect 17773 15447 17831 15453
rect 18966 15444 18972 15456
rect 19024 15444 19030 15496
rect 19429 15487 19487 15493
rect 19429 15453 19441 15487
rect 19475 15484 19487 15487
rect 19610 15484 19616 15496
rect 19475 15456 19616 15484
rect 19475 15453 19487 15456
rect 19429 15447 19487 15453
rect 19610 15444 19616 15456
rect 19668 15444 19674 15496
rect 19705 15487 19763 15493
rect 19705 15453 19717 15487
rect 19751 15484 19763 15487
rect 20732 15484 20760 15512
rect 19751 15456 20760 15484
rect 19751 15453 19763 15456
rect 19705 15447 19763 15453
rect 16850 15376 16856 15428
rect 16908 15376 16914 15428
rect 18432 15388 19472 15416
rect 16393 15351 16451 15357
rect 16393 15348 16405 15351
rect 15764 15320 16405 15348
rect 16393 15317 16405 15320
rect 16439 15317 16451 15351
rect 16393 15311 16451 15317
rect 16669 15351 16727 15357
rect 16669 15317 16681 15351
rect 16715 15317 16727 15351
rect 16669 15311 16727 15317
rect 17402 15308 17408 15360
rect 17460 15348 17466 15360
rect 18432 15348 18460 15388
rect 17460 15320 18460 15348
rect 17460 15308 17466 15320
rect 18874 15308 18880 15360
rect 18932 15308 18938 15360
rect 19444 15348 19472 15388
rect 20824 15348 20852 15660
rect 23109 15657 23121 15660
rect 23155 15657 23167 15691
rect 24578 15688 24584 15700
rect 23109 15651 23167 15657
rect 23216 15660 24584 15688
rect 23014 15580 23020 15632
rect 23072 15620 23078 15632
rect 23216 15620 23244 15660
rect 24578 15648 24584 15660
rect 24636 15648 24642 15700
rect 25685 15691 25743 15697
rect 25685 15657 25697 15691
rect 25731 15688 25743 15691
rect 26786 15688 26792 15700
rect 25731 15660 26792 15688
rect 25731 15657 25743 15660
rect 25685 15651 25743 15657
rect 26786 15648 26792 15660
rect 26844 15648 26850 15700
rect 27338 15648 27344 15700
rect 27396 15688 27402 15700
rect 27709 15691 27767 15697
rect 27709 15688 27721 15691
rect 27396 15660 27721 15688
rect 27396 15648 27402 15660
rect 27709 15657 27721 15660
rect 27755 15657 27767 15691
rect 27709 15651 27767 15657
rect 27798 15648 27804 15700
rect 27856 15688 27862 15700
rect 30377 15691 30435 15697
rect 30377 15688 30389 15691
rect 27856 15660 30389 15688
rect 27856 15648 27862 15660
rect 30377 15657 30389 15660
rect 30423 15657 30435 15691
rect 30377 15651 30435 15657
rect 23072 15592 23244 15620
rect 23072 15580 23078 15592
rect 23474 15580 23480 15632
rect 23532 15580 23538 15632
rect 26234 15620 26240 15632
rect 25976 15592 26240 15620
rect 21085 15555 21143 15561
rect 21085 15521 21097 15555
rect 21131 15552 21143 15555
rect 23492 15552 23520 15580
rect 21131 15524 21496 15552
rect 21131 15521 21143 15524
rect 21085 15515 21143 15521
rect 21468 15496 21496 15524
rect 21928 15524 23520 15552
rect 21765 15505 21823 15511
rect 21266 15444 21272 15496
rect 21324 15444 21330 15496
rect 21450 15444 21456 15496
rect 21508 15444 21514 15496
rect 21634 15493 21640 15496
rect 21596 15487 21640 15493
rect 21596 15453 21608 15487
rect 21596 15447 21640 15453
rect 21634 15444 21640 15447
rect 21692 15444 21698 15496
rect 21765 15471 21777 15505
rect 21811 15484 21823 15505
rect 21928 15484 21956 15524
rect 23566 15512 23572 15564
rect 23624 15552 23630 15564
rect 24213 15555 24271 15561
rect 24213 15552 24225 15555
rect 23624 15524 24225 15552
rect 23624 15512 23630 15524
rect 24213 15521 24225 15524
rect 24259 15521 24271 15555
rect 24213 15515 24271 15521
rect 24302 15512 24308 15564
rect 24360 15552 24366 15564
rect 25976 15561 26004 15592
rect 26234 15580 26240 15592
rect 26292 15580 26298 15632
rect 26602 15580 26608 15632
rect 26660 15620 26666 15632
rect 26660 15592 27384 15620
rect 26660 15580 26666 15592
rect 25869 15555 25927 15561
rect 25869 15552 25881 15555
rect 24360 15524 25881 15552
rect 24360 15512 24366 15524
rect 25869 15521 25881 15524
rect 25915 15521 25927 15555
rect 25869 15515 25927 15521
rect 25961 15555 26019 15561
rect 25961 15521 25973 15555
rect 26007 15521 26019 15555
rect 25961 15515 26019 15521
rect 21811 15471 21956 15484
rect 21765 15465 21956 15471
rect 21790 15456 21956 15465
rect 22002 15444 22008 15496
rect 22060 15444 22066 15496
rect 23477 15487 23535 15493
rect 23477 15453 23489 15487
rect 23523 15484 23535 15487
rect 23658 15484 23664 15496
rect 23523 15456 23664 15484
rect 23523 15453 23535 15456
rect 23477 15447 23535 15453
rect 23658 15444 23664 15456
rect 23716 15444 23722 15496
rect 23842 15493 23848 15496
rect 23804 15487 23848 15493
rect 23804 15453 23816 15487
rect 23804 15447 23848 15453
rect 23842 15444 23848 15447
rect 23900 15444 23906 15496
rect 23983 15487 24041 15493
rect 23983 15453 23995 15487
rect 24029 15484 24041 15487
rect 24670 15484 24676 15496
rect 24029 15456 24676 15484
rect 24029 15453 24041 15456
rect 23983 15447 24041 15453
rect 24670 15444 24676 15456
rect 24728 15444 24734 15496
rect 25884 15416 25912 15515
rect 26050 15512 26056 15564
rect 26108 15552 26114 15564
rect 26697 15555 26755 15561
rect 26697 15552 26709 15555
rect 26108 15524 26709 15552
rect 26108 15512 26114 15524
rect 26697 15521 26709 15524
rect 26743 15521 26755 15555
rect 26697 15515 26755 15521
rect 27157 15555 27215 15561
rect 27157 15521 27169 15555
rect 27203 15521 27215 15555
rect 27157 15515 27215 15521
rect 26234 15444 26240 15496
rect 26292 15484 26298 15496
rect 27172 15484 27200 15515
rect 27356 15493 27384 15592
rect 27586 15592 28028 15620
rect 26292 15456 27200 15484
rect 27341 15487 27399 15493
rect 26292 15444 26298 15456
rect 27341 15453 27353 15487
rect 27387 15453 27399 15487
rect 27341 15447 27399 15453
rect 26145 15419 26203 15425
rect 26145 15416 26157 15419
rect 22848 15388 23244 15416
rect 25884 15388 26157 15416
rect 19444 15320 20852 15348
rect 21910 15308 21916 15360
rect 21968 15348 21974 15360
rect 22848 15348 22876 15388
rect 21968 15320 22876 15348
rect 23216 15348 23244 15388
rect 26145 15385 26157 15388
rect 26191 15385 26203 15419
rect 26145 15379 26203 15385
rect 25317 15351 25375 15357
rect 25317 15348 25329 15351
rect 23216 15320 25329 15348
rect 21968 15308 21974 15320
rect 25317 15317 25329 15320
rect 25363 15317 25375 15351
rect 25317 15311 25375 15317
rect 25958 15308 25964 15360
rect 26016 15348 26022 15360
rect 26252 15348 26280 15444
rect 26786 15376 26792 15428
rect 26844 15416 26850 15428
rect 27586 15416 27614 15592
rect 28000 15561 28028 15592
rect 28350 15561 28356 15564
rect 27869 15555 27927 15561
rect 27869 15552 27881 15555
rect 26844 15388 27614 15416
rect 27862 15521 27881 15552
rect 27915 15521 27927 15555
rect 27862 15515 27927 15521
rect 27985 15555 28043 15561
rect 27985 15521 27997 15555
rect 28031 15521 28043 15555
rect 27985 15515 28043 15521
rect 28312 15555 28356 15561
rect 28312 15521 28324 15555
rect 28312 15515 28356 15521
rect 26844 15376 26850 15388
rect 26016 15320 26280 15348
rect 26973 15351 27031 15357
rect 26016 15308 26022 15320
rect 26973 15317 26985 15351
rect 27019 15348 27031 15351
rect 27862 15348 27890 15515
rect 28350 15512 28356 15515
rect 28408 15512 28414 15564
rect 29362 15512 29368 15564
rect 29420 15552 29426 15564
rect 30285 15555 30343 15561
rect 30285 15552 30297 15555
rect 29420 15524 30297 15552
rect 29420 15512 29426 15524
rect 30285 15521 30297 15524
rect 30331 15521 30343 15555
rect 30285 15515 30343 15521
rect 28491 15487 28549 15493
rect 28491 15453 28503 15487
rect 28537 15484 28549 15487
rect 28626 15484 28632 15496
rect 28537 15456 28632 15484
rect 28537 15453 28549 15456
rect 28491 15447 28549 15453
rect 28626 15444 28632 15456
rect 28684 15444 28690 15496
rect 28721 15487 28779 15493
rect 28721 15453 28733 15487
rect 28767 15484 28779 15487
rect 29822 15484 29828 15496
rect 28767 15456 29828 15484
rect 28767 15453 28779 15456
rect 28721 15447 28779 15453
rect 29822 15444 29828 15456
rect 29880 15444 29886 15496
rect 29546 15376 29552 15428
rect 29604 15416 29610 15428
rect 29730 15416 29736 15428
rect 29604 15388 29736 15416
rect 29604 15376 29610 15388
rect 29730 15376 29736 15388
rect 29788 15376 29794 15428
rect 28350 15348 28356 15360
rect 27019 15320 28356 15348
rect 27019 15317 27031 15320
rect 26973 15311 27031 15317
rect 28350 15308 28356 15320
rect 28408 15308 28414 15360
rect 28534 15308 28540 15360
rect 28592 15348 28598 15360
rect 29825 15351 29883 15357
rect 29825 15348 29837 15351
rect 28592 15320 29837 15348
rect 28592 15308 28598 15320
rect 29825 15317 29837 15320
rect 29871 15317 29883 15351
rect 29825 15311 29883 15317
rect 552 15258 30912 15280
rect 552 15206 4193 15258
rect 4245 15206 4257 15258
rect 4309 15206 4321 15258
rect 4373 15206 4385 15258
rect 4437 15206 4449 15258
rect 4501 15206 11783 15258
rect 11835 15206 11847 15258
rect 11899 15206 11911 15258
rect 11963 15206 11975 15258
rect 12027 15206 12039 15258
rect 12091 15206 19373 15258
rect 19425 15206 19437 15258
rect 19489 15206 19501 15258
rect 19553 15206 19565 15258
rect 19617 15206 19629 15258
rect 19681 15206 26963 15258
rect 27015 15206 27027 15258
rect 27079 15206 27091 15258
rect 27143 15206 27155 15258
rect 27207 15206 27219 15258
rect 27271 15206 30912 15258
rect 552 15184 30912 15206
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 1728 15116 2360 15144
rect 1728 15104 1734 15116
rect 2332 15076 2360 15116
rect 2958 15104 2964 15156
rect 3016 15104 3022 15156
rect 4246 15144 4252 15156
rect 3068 15116 4252 15144
rect 3068 15076 3096 15116
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 8294 15144 8300 15156
rect 6104 15116 8300 15144
rect 2332 15048 3096 15076
rect 937 15011 995 15017
rect 937 14977 949 15011
rect 983 15008 995 15011
rect 1302 15008 1308 15020
rect 983 14980 1308 15008
rect 983 14977 995 14980
rect 937 14971 995 14977
rect 1302 14968 1308 14980
rect 1360 14968 1366 15020
rect 1443 15011 1501 15017
rect 1443 14977 1455 15011
rect 1489 15008 1501 15011
rect 3510 15008 3516 15020
rect 1489 14980 3516 15008
rect 1489 14977 1501 14980
rect 1443 14971 1501 14977
rect 3510 14968 3516 14980
rect 3568 14968 3574 15020
rect 3786 14968 3792 15020
rect 3844 15008 3850 15020
rect 3881 15011 3939 15017
rect 3881 15008 3893 15011
rect 3844 14980 3893 15008
rect 3844 14968 3850 14980
rect 3881 14977 3893 14980
rect 3927 14977 3939 15011
rect 3881 14971 3939 14977
rect 4387 15011 4445 15017
rect 4387 14977 4399 15011
rect 4433 15008 4445 15011
rect 6104 15008 6132 15116
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 10505 15147 10563 15153
rect 10505 15144 10517 15147
rect 8404 15116 10517 15144
rect 7926 15036 7932 15088
rect 7984 15076 7990 15088
rect 8404 15076 8432 15116
rect 10505 15113 10517 15116
rect 10551 15113 10563 15147
rect 10505 15107 10563 15113
rect 10870 15104 10876 15156
rect 10928 15144 10934 15156
rect 10965 15147 11023 15153
rect 10965 15144 10977 15147
rect 10928 15116 10977 15144
rect 10928 15104 10934 15116
rect 10965 15113 10977 15116
rect 11011 15113 11023 15147
rect 10965 15107 11023 15113
rect 11790 15104 11796 15156
rect 11848 15144 11854 15156
rect 15378 15144 15384 15156
rect 11848 15116 15384 15144
rect 11848 15104 11854 15116
rect 15378 15104 15384 15116
rect 15436 15104 15442 15156
rect 16206 15104 16212 15156
rect 16264 15144 16270 15156
rect 17126 15144 17132 15156
rect 16264 15116 17132 15144
rect 16264 15104 16270 15116
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 19337 15147 19395 15153
rect 19337 15113 19349 15147
rect 19383 15144 19395 15147
rect 20254 15144 20260 15156
rect 19383 15116 20260 15144
rect 19383 15113 19395 15116
rect 19337 15107 19395 15113
rect 20254 15104 20260 15116
rect 20312 15104 20318 15156
rect 20346 15104 20352 15156
rect 20404 15144 20410 15156
rect 23382 15144 23388 15156
rect 20404 15116 23388 15144
rect 20404 15104 20410 15116
rect 23382 15104 23388 15116
rect 23440 15104 23446 15156
rect 23474 15104 23480 15156
rect 23532 15144 23538 15156
rect 25685 15147 25743 15153
rect 25685 15144 25697 15147
rect 23532 15116 25697 15144
rect 23532 15104 23538 15116
rect 25685 15113 25697 15116
rect 25731 15113 25743 15147
rect 25685 15107 25743 15113
rect 26053 15147 26111 15153
rect 26053 15113 26065 15147
rect 26099 15144 26111 15147
rect 26510 15144 26516 15156
rect 26099 15116 26516 15144
rect 26099 15113 26111 15116
rect 26053 15107 26111 15113
rect 26510 15104 26516 15116
rect 26568 15104 26574 15156
rect 27338 15144 27344 15156
rect 26620 15116 27344 15144
rect 7984 15048 8432 15076
rect 13081 15079 13139 15085
rect 7984 15036 7990 15048
rect 13081 15045 13093 15079
rect 13127 15045 13139 15079
rect 13081 15039 13139 15045
rect 4433 14980 6132 15008
rect 4433 14977 4445 14980
rect 4387 14971 4445 14977
rect 6270 14968 6276 15020
rect 6328 14968 6334 15020
rect 9030 15017 9036 15020
rect 6595 15011 6653 15017
rect 6595 14977 6607 15011
rect 6641 15008 6653 15011
rect 8992 15011 9036 15017
rect 6641 14980 8892 15008
rect 6641 14977 6653 14980
rect 6595 14971 6653 14977
rect 1673 14943 1731 14949
rect 1673 14909 1685 14943
rect 1719 14940 1731 14943
rect 2682 14940 2688 14952
rect 1719 14912 2688 14940
rect 1719 14909 1731 14912
rect 1673 14903 1731 14909
rect 2682 14900 2688 14912
rect 2740 14900 2746 14952
rect 3237 14943 3295 14949
rect 3237 14909 3249 14943
rect 3283 14940 3295 14943
rect 3694 14940 3700 14952
rect 3283 14912 3700 14940
rect 3283 14909 3295 14912
rect 3237 14903 3295 14909
rect 3694 14900 3700 14912
rect 3752 14900 3758 14952
rect 4154 14900 4160 14952
rect 4212 14940 4218 14952
rect 4617 14943 4675 14949
rect 4617 14940 4629 14943
rect 4212 14912 4629 14940
rect 4212 14900 4218 14912
rect 4617 14909 4629 14912
rect 4663 14909 4675 14943
rect 4617 14903 4675 14909
rect 6086 14900 6092 14952
rect 6144 14900 6150 14952
rect 6288 14940 6316 14968
rect 6196 14912 6316 14940
rect 3513 14875 3571 14881
rect 3513 14841 3525 14875
rect 3559 14841 3571 14875
rect 3513 14835 3571 14841
rect 5997 14875 6055 14881
rect 5997 14841 6009 14875
rect 6043 14872 6055 14875
rect 6196 14872 6224 14912
rect 6822 14900 6828 14952
rect 6880 14900 6886 14952
rect 7282 14900 7288 14952
rect 7340 14940 7346 14952
rect 7340 14912 7512 14940
rect 7340 14900 7346 14912
rect 6043 14844 6224 14872
rect 7484 14872 7512 14912
rect 8478 14900 8484 14952
rect 8536 14940 8542 14952
rect 8573 14943 8631 14949
rect 8573 14940 8585 14943
rect 8536 14912 8585 14940
rect 8536 14900 8542 14912
rect 8573 14909 8585 14912
rect 8619 14909 8631 14943
rect 8573 14903 8631 14909
rect 7484 14844 8432 14872
rect 6043 14841 6055 14844
rect 5997 14835 6055 14841
rect 1394 14764 1400 14816
rect 1452 14813 1458 14816
rect 1452 14804 1461 14813
rect 3528 14804 3556 14835
rect 3878 14804 3884 14816
rect 1452 14776 3884 14804
rect 1452 14767 1461 14776
rect 1452 14764 1458 14767
rect 3878 14764 3884 14776
rect 3936 14804 3942 14816
rect 4347 14807 4405 14813
rect 4347 14804 4359 14807
rect 3936 14776 4359 14804
rect 3936 14764 3942 14776
rect 4347 14773 4359 14776
rect 4393 14773 4405 14807
rect 4347 14767 4405 14773
rect 6454 14764 6460 14816
rect 6512 14804 6518 14816
rect 6555 14807 6613 14813
rect 6555 14804 6567 14807
rect 6512 14776 6567 14804
rect 6512 14764 6518 14776
rect 6555 14773 6567 14776
rect 6601 14773 6613 14807
rect 6555 14767 6613 14773
rect 6914 14764 6920 14816
rect 6972 14804 6978 14816
rect 8404 14813 8432 14844
rect 7929 14807 7987 14813
rect 7929 14804 7941 14807
rect 6972 14776 7941 14804
rect 6972 14764 6978 14776
rect 7929 14773 7941 14776
rect 7975 14773 7987 14807
rect 7929 14767 7987 14773
rect 8389 14807 8447 14813
rect 8389 14773 8401 14807
rect 8435 14773 8447 14807
rect 8588 14804 8616 14903
rect 8662 14900 8668 14952
rect 8720 14900 8726 14952
rect 8864 14940 8892 14980
rect 8992 14977 9004 15011
rect 8992 14971 9036 14977
rect 9030 14968 9036 14971
rect 9088 14968 9094 15020
rect 9214 15017 9220 15020
rect 9171 15011 9220 15017
rect 9171 14977 9183 15011
rect 9217 14977 9220 15011
rect 9171 14971 9220 14977
rect 9214 14968 9220 14971
rect 9272 14968 9278 15020
rect 11790 15017 11796 15020
rect 11747 15011 11796 15017
rect 9324 14980 11468 15008
rect 9324 14940 9352 14980
rect 8864 14912 9352 14940
rect 9398 14900 9404 14952
rect 9456 14900 9462 14952
rect 10318 14900 10324 14952
rect 10376 14940 10382 14952
rect 10870 14940 10876 14952
rect 10376 14912 10876 14940
rect 10376 14900 10382 14912
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 11054 14900 11060 14952
rect 11112 14940 11118 14952
rect 11149 14943 11207 14949
rect 11149 14940 11161 14943
rect 11112 14912 11161 14940
rect 11112 14900 11118 14912
rect 11149 14909 11161 14912
rect 11195 14909 11207 14943
rect 11149 14903 11207 14909
rect 11241 14943 11299 14949
rect 11241 14909 11253 14943
rect 11287 14940 11299 14943
rect 11330 14940 11336 14952
rect 11287 14912 11336 14940
rect 11287 14909 11299 14912
rect 11241 14903 11299 14909
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 11440 14940 11468 14980
rect 11747 14977 11759 15011
rect 11793 14977 11796 15011
rect 11747 14971 11796 14977
rect 11790 14968 11796 14971
rect 11848 14968 11854 15020
rect 13096 15008 13124 15039
rect 13906 15036 13912 15088
rect 13964 15036 13970 15088
rect 14090 15036 14096 15088
rect 14148 15076 14154 15088
rect 14185 15079 14243 15085
rect 14185 15076 14197 15079
rect 14148 15048 14197 15076
rect 14148 15036 14154 15048
rect 14185 15045 14197 15048
rect 14231 15045 14243 15079
rect 19426 15076 19432 15088
rect 14185 15039 14243 15045
rect 18432 15048 19432 15076
rect 11900 14980 13124 15008
rect 11900 14940 11928 14980
rect 13630 14968 13636 15020
rect 13688 15008 13694 15020
rect 15059 15011 15117 15017
rect 13688 14980 14688 15008
rect 13688 14968 13694 14980
rect 11440 14912 11928 14940
rect 11977 14943 12035 14949
rect 11977 14909 11989 14943
rect 12023 14940 12035 14943
rect 12434 14940 12440 14952
rect 12023 14912 12440 14940
rect 12023 14909 12035 14912
rect 11977 14903 12035 14909
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 12618 14900 12624 14952
rect 12676 14940 12682 14952
rect 14093 14943 14151 14949
rect 14093 14940 14105 14943
rect 12676 14912 14105 14940
rect 12676 14900 12682 14912
rect 13446 14832 13452 14884
rect 13504 14872 13510 14884
rect 13633 14875 13691 14881
rect 13633 14872 13645 14875
rect 13504 14844 13645 14872
rect 13504 14832 13510 14844
rect 13633 14841 13645 14844
rect 13679 14841 13691 14875
rect 13633 14835 13691 14841
rect 13722 14832 13728 14884
rect 13780 14872 13786 14884
rect 13817 14875 13875 14881
rect 13817 14872 13829 14875
rect 13780 14844 13829 14872
rect 13780 14832 13786 14844
rect 13817 14841 13829 14844
rect 13863 14841 13875 14875
rect 13817 14835 13875 14841
rect 11330 14804 11336 14816
rect 8588 14776 11336 14804
rect 8389 14767 8447 14773
rect 11330 14764 11336 14776
rect 11388 14764 11394 14816
rect 11698 14764 11704 14816
rect 11756 14813 11762 14816
rect 11756 14804 11765 14813
rect 13924 14804 13952 14912
rect 14093 14909 14105 14912
rect 14139 14909 14151 14943
rect 14093 14903 14151 14909
rect 14274 14900 14280 14952
rect 14332 14900 14338 14952
rect 14369 14943 14427 14949
rect 14369 14909 14381 14943
rect 14415 14940 14427 14943
rect 14458 14940 14464 14952
rect 14415 14912 14464 14940
rect 14415 14909 14427 14912
rect 14369 14903 14427 14909
rect 14458 14900 14464 14912
rect 14516 14900 14522 14952
rect 14553 14943 14611 14949
rect 14553 14909 14565 14943
rect 14599 14909 14611 14943
rect 14660 14940 14688 14980
rect 15059 14977 15071 15011
rect 15105 15008 15117 15011
rect 15105 14980 16804 15008
rect 15105 14977 15117 14980
rect 15059 14971 15117 14977
rect 15194 14940 15200 14952
rect 14660 14912 15200 14940
rect 14553 14903 14611 14909
rect 13998 14832 14004 14884
rect 14056 14872 14062 14884
rect 14292 14872 14320 14900
rect 14568 14872 14596 14903
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 15286 14900 15292 14952
rect 15344 14900 15350 14952
rect 14056 14844 14596 14872
rect 14056 14832 14062 14844
rect 14090 14804 14096 14816
rect 11756 14776 11801 14804
rect 13924 14776 14096 14804
rect 11756 14767 11765 14776
rect 11756 14764 11762 14767
rect 14090 14764 14096 14776
rect 14148 14804 14154 14816
rect 14366 14804 14372 14816
rect 14148 14776 14372 14804
rect 14148 14764 14154 14776
rect 14366 14764 14372 14776
rect 14424 14764 14430 14816
rect 14918 14764 14924 14816
rect 14976 14804 14982 14816
rect 15019 14807 15077 14813
rect 15019 14804 15031 14807
rect 14976 14776 15031 14804
rect 14976 14764 14982 14776
rect 15019 14773 15031 14776
rect 15065 14773 15077 14807
rect 15019 14767 15077 14773
rect 16390 14764 16396 14816
rect 16448 14764 16454 14816
rect 16776 14804 16804 14980
rect 17126 14968 17132 15020
rect 17184 14968 17190 15020
rect 18432 15008 18460 15048
rect 19426 15036 19432 15048
rect 19484 15036 19490 15088
rect 23842 15036 23848 15088
rect 23900 15036 23906 15088
rect 26418 15036 26424 15088
rect 26476 15076 26482 15088
rect 26620 15076 26648 15116
rect 27338 15104 27344 15116
rect 27396 15144 27402 15156
rect 27396 15116 28120 15144
rect 27396 15104 27402 15116
rect 26476 15048 26648 15076
rect 28092 15076 28120 15116
rect 28350 15104 28356 15156
rect 28408 15144 28414 15156
rect 28534 15144 28540 15156
rect 28408 15116 28540 15144
rect 28408 15104 28414 15116
rect 28534 15104 28540 15116
rect 28592 15104 28598 15156
rect 28721 15147 28779 15153
rect 28721 15113 28733 15147
rect 28767 15144 28779 15147
rect 28994 15144 29000 15156
rect 28767 15116 29000 15144
rect 28767 15113 28779 15116
rect 28721 15107 28779 15113
rect 28994 15104 29000 15116
rect 29052 15104 29058 15156
rect 29454 15104 29460 15156
rect 29512 15144 29518 15156
rect 30193 15147 30251 15153
rect 30193 15144 30205 15147
rect 29512 15116 30205 15144
rect 29512 15104 29518 15116
rect 30193 15113 30205 15116
rect 30239 15113 30251 15147
rect 30193 15107 30251 15113
rect 30650 15104 30656 15156
rect 30708 15104 30714 15156
rect 29273 15079 29331 15085
rect 29273 15076 29285 15079
rect 28092 15048 29285 15076
rect 26476 15036 26482 15048
rect 29273 15045 29285 15048
rect 29319 15076 29331 15079
rect 29362 15076 29368 15088
rect 29319 15048 29368 15076
rect 29319 15045 29331 15048
rect 29273 15039 29331 15045
rect 29362 15036 29368 15048
rect 29420 15036 29426 15088
rect 29914 15036 29920 15088
rect 29972 15076 29978 15088
rect 30668 15076 30696 15104
rect 29972 15048 30696 15076
rect 29972 15036 29978 15048
rect 17236 14980 18460 15008
rect 18509 15011 18567 15017
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14940 16911 14943
rect 17236 14940 17264 14980
rect 18509 14977 18521 15011
rect 18555 15008 18567 15011
rect 19978 15008 19984 15020
rect 18555 14980 19984 15008
rect 18555 14977 18567 14980
rect 18509 14971 18567 14977
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 22281 15011 22339 15017
rect 20088 14993 21128 15008
rect 20088 14962 20121 14993
rect 20109 14959 20121 14962
rect 20155 14980 21128 14993
rect 20155 14959 20167 14980
rect 20109 14953 20167 14959
rect 16899 14912 17264 14940
rect 16899 14909 16911 14912
rect 16853 14903 16911 14909
rect 17586 14900 17592 14952
rect 17644 14940 17650 14952
rect 18693 14943 18751 14949
rect 18693 14940 18705 14943
rect 17644 14912 18705 14940
rect 17644 14900 17650 14912
rect 18693 14909 18705 14912
rect 18739 14940 18751 14943
rect 18782 14940 18788 14952
rect 18739 14912 18788 14940
rect 18739 14909 18751 14912
rect 18693 14903 18751 14909
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 19521 14943 19579 14949
rect 19521 14940 19533 14943
rect 19168 14912 19533 14940
rect 17954 14832 17960 14884
rect 18012 14872 18018 14884
rect 18969 14875 19027 14881
rect 18969 14872 18981 14875
rect 18012 14844 18981 14872
rect 18012 14832 18018 14844
rect 18969 14841 18981 14844
rect 19015 14841 19027 14875
rect 18969 14835 19027 14841
rect 19168 14816 19196 14912
rect 19521 14909 19533 14912
rect 19567 14909 19579 14943
rect 19521 14903 19579 14909
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14940 19671 14943
rect 19702 14940 19708 14952
rect 19659 14912 19708 14940
rect 19659 14909 19671 14912
rect 19613 14903 19671 14909
rect 19702 14900 19708 14912
rect 19760 14900 19766 14952
rect 20346 14900 20352 14952
rect 20404 14900 20410 14952
rect 21100 14872 21128 14980
rect 22281 14977 22293 15011
rect 22327 15008 22339 15011
rect 22922 15008 22928 15020
rect 22327 14980 22928 15008
rect 22327 14977 22339 14980
rect 22281 14971 22339 14977
rect 22922 14968 22928 14980
rect 22980 14968 22986 15020
rect 23658 14968 23664 15020
rect 23716 14968 23722 15020
rect 23860 15008 23888 15036
rect 24172 15011 24230 15017
rect 24172 15008 24184 15011
rect 23860 14980 24184 15008
rect 24172 14977 24184 14980
rect 24218 14977 24230 15011
rect 24172 14971 24230 14977
rect 24351 15011 24409 15017
rect 24351 14977 24363 15011
rect 24397 15008 24409 15011
rect 24762 15008 24768 15020
rect 24397 14980 24768 15008
rect 24397 14977 24409 14980
rect 24351 14971 24409 14977
rect 24762 14968 24768 14980
rect 24820 14968 24826 15020
rect 24946 14968 24952 15020
rect 25004 15008 25010 15020
rect 27062 15008 27068 15020
rect 25004 14980 27068 15008
rect 25004 14968 25010 14980
rect 22005 14943 22063 14949
rect 22005 14909 22017 14943
rect 22051 14940 22063 14943
rect 23566 14940 23572 14952
rect 22051 14912 23572 14940
rect 22051 14909 22063 14912
rect 22005 14903 22063 14909
rect 23566 14900 23572 14912
rect 23624 14900 23630 14952
rect 23676 14940 23704 14968
rect 23845 14943 23903 14949
rect 23845 14940 23857 14943
rect 23676 14912 23857 14940
rect 23845 14909 23857 14912
rect 23891 14909 23903 14943
rect 24581 14943 24639 14949
rect 24581 14940 24593 14943
rect 23845 14903 23903 14909
rect 23952 14912 24593 14940
rect 22094 14872 22100 14884
rect 21100 14844 22100 14872
rect 22094 14832 22100 14844
rect 22152 14832 22158 14884
rect 23952 14872 23980 14912
rect 24581 14909 24593 14912
rect 24627 14909 24639 14943
rect 24581 14903 24639 14909
rect 24670 14900 24676 14952
rect 24728 14940 24734 14952
rect 26344 14949 26372 14980
rect 27062 14968 27068 14980
rect 27120 14968 27126 15020
rect 27160 15009 27218 15015
rect 27160 14975 27172 15009
rect 27206 14975 27218 15009
rect 27160 14969 27218 14975
rect 26237 14943 26295 14949
rect 26237 14940 26249 14943
rect 24728 14912 26249 14940
rect 24728 14900 24734 14912
rect 26237 14909 26249 14912
rect 26283 14909 26295 14943
rect 26237 14903 26295 14909
rect 26329 14943 26387 14949
rect 26329 14909 26341 14943
rect 26375 14909 26387 14943
rect 26329 14903 26387 14909
rect 22940 14844 23980 14872
rect 22940 14816 22968 14844
rect 18782 14804 18788 14816
rect 16776 14776 18788 14804
rect 18782 14764 18788 14776
rect 18840 14764 18846 14816
rect 19150 14764 19156 14816
rect 19208 14764 19214 14816
rect 20079 14807 20137 14813
rect 20079 14773 20091 14807
rect 20125 14804 20137 14807
rect 20622 14804 20628 14816
rect 20125 14776 20628 14804
rect 20125 14773 20137 14776
rect 20079 14767 20137 14773
rect 20622 14764 20628 14776
rect 20680 14764 20686 14816
rect 21174 14764 21180 14816
rect 21232 14804 21238 14816
rect 21453 14807 21511 14813
rect 21453 14804 21465 14807
rect 21232 14776 21465 14804
rect 21232 14764 21238 14776
rect 21453 14773 21465 14776
rect 21499 14773 21511 14807
rect 21453 14767 21511 14773
rect 21542 14764 21548 14816
rect 21600 14804 21606 14816
rect 22738 14804 22744 14816
rect 21600 14776 22744 14804
rect 21600 14764 21606 14776
rect 22738 14764 22744 14776
rect 22796 14764 22802 14816
rect 22922 14764 22928 14816
rect 22980 14764 22986 14816
rect 23569 14807 23627 14813
rect 23569 14773 23581 14807
rect 23615 14804 23627 14807
rect 26142 14804 26148 14816
rect 23615 14776 26148 14804
rect 23615 14773 23627 14776
rect 23569 14767 23627 14773
rect 26142 14764 26148 14776
rect 26200 14764 26206 14816
rect 26252 14804 26280 14903
rect 26602 14900 26608 14952
rect 26660 14940 26666 14952
rect 26697 14943 26755 14949
rect 26697 14940 26709 14943
rect 26660 14912 26709 14940
rect 26660 14900 26666 14912
rect 26697 14909 26709 14912
rect 26743 14940 26755 14943
rect 26786 14940 26792 14952
rect 26743 14912 26792 14940
rect 26743 14909 26755 14912
rect 26697 14903 26755 14909
rect 26786 14900 26792 14912
rect 26844 14900 26850 14952
rect 27172 14936 27200 14969
rect 27246 14968 27252 15020
rect 27304 15008 27310 15020
rect 27304 14980 30512 15008
rect 27304 14968 27310 14980
rect 30484 14952 30512 14980
rect 27338 14940 27344 14952
rect 27264 14936 27344 14940
rect 27172 14912 27344 14936
rect 27172 14908 27292 14912
rect 27338 14900 27344 14912
rect 27396 14900 27402 14952
rect 27433 14943 27491 14949
rect 27433 14909 27445 14943
rect 27479 14940 27491 14943
rect 28994 14940 29000 14952
rect 27479 14912 29000 14940
rect 27479 14909 27491 14912
rect 27433 14903 27491 14909
rect 28994 14900 29000 14912
rect 29052 14900 29058 14952
rect 29178 14900 29184 14952
rect 29236 14940 29242 14952
rect 29641 14943 29699 14949
rect 29641 14940 29653 14943
rect 29236 14912 29653 14940
rect 29236 14900 29242 14912
rect 29641 14909 29653 14912
rect 29687 14940 29699 14943
rect 30006 14940 30012 14952
rect 29687 14912 30012 14940
rect 29687 14909 29699 14912
rect 29641 14903 29699 14909
rect 30006 14900 30012 14912
rect 30064 14900 30070 14952
rect 30190 14900 30196 14952
rect 30248 14940 30254 14952
rect 30377 14943 30435 14949
rect 30377 14940 30389 14943
rect 30248 14912 30389 14940
rect 30248 14900 30254 14912
rect 30377 14909 30389 14912
rect 30423 14909 30435 14943
rect 30377 14903 30435 14909
rect 30466 14900 30472 14952
rect 30524 14900 30530 14952
rect 29089 14875 29147 14881
rect 29089 14841 29101 14875
rect 29135 14841 29147 14875
rect 29089 14835 29147 14841
rect 26513 14807 26571 14813
rect 26513 14804 26525 14807
rect 26252 14776 26525 14804
rect 26513 14773 26525 14776
rect 26559 14773 26571 14807
rect 26513 14767 26571 14773
rect 27163 14807 27221 14813
rect 27163 14773 27175 14807
rect 27209 14804 27221 14807
rect 27430 14804 27436 14816
rect 27209 14776 27436 14804
rect 27209 14773 27221 14776
rect 27163 14767 27221 14773
rect 27430 14764 27436 14776
rect 27488 14764 27494 14816
rect 27706 14764 27712 14816
rect 27764 14804 27770 14816
rect 29104 14804 29132 14835
rect 27764 14776 29132 14804
rect 27764 14764 27770 14776
rect 552 14714 31072 14736
rect 552 14662 7988 14714
rect 8040 14662 8052 14714
rect 8104 14662 8116 14714
rect 8168 14662 8180 14714
rect 8232 14662 8244 14714
rect 8296 14662 15578 14714
rect 15630 14662 15642 14714
rect 15694 14662 15706 14714
rect 15758 14662 15770 14714
rect 15822 14662 15834 14714
rect 15886 14662 23168 14714
rect 23220 14662 23232 14714
rect 23284 14662 23296 14714
rect 23348 14662 23360 14714
rect 23412 14662 23424 14714
rect 23476 14662 30758 14714
rect 30810 14662 30822 14714
rect 30874 14662 30886 14714
rect 30938 14662 30950 14714
rect 31002 14662 31014 14714
rect 31066 14662 31072 14714
rect 552 14640 31072 14662
rect 1213 14603 1271 14609
rect 1213 14569 1225 14603
rect 1259 14600 1271 14603
rect 1259 14572 4022 14600
rect 1259 14569 1271 14572
rect 1213 14563 1271 14569
rect 1118 14424 1124 14476
rect 1176 14424 1182 14476
rect 1394 14424 1400 14476
rect 1452 14424 1458 14476
rect 1816 14467 1874 14473
rect 1816 14433 1828 14467
rect 1862 14433 1874 14467
rect 1816 14427 1874 14433
rect 3881 14467 3939 14473
rect 3881 14433 3893 14467
rect 3927 14433 3939 14467
rect 3994 14464 4022 14572
rect 4062 14560 4068 14612
rect 4120 14560 4126 14612
rect 4341 14603 4399 14609
rect 4341 14569 4353 14603
rect 4387 14600 4399 14603
rect 4522 14600 4528 14612
rect 4387 14572 4528 14600
rect 4387 14569 4399 14572
rect 4341 14563 4399 14569
rect 4522 14560 4528 14572
rect 4580 14560 4586 14612
rect 4893 14603 4951 14609
rect 4893 14569 4905 14603
rect 4939 14600 4951 14603
rect 5074 14600 5080 14612
rect 4939 14572 5080 14600
rect 4939 14569 4951 14572
rect 4893 14563 4951 14569
rect 5074 14560 5080 14572
rect 5132 14560 5138 14612
rect 5169 14603 5227 14609
rect 5169 14569 5181 14603
rect 5215 14569 5227 14603
rect 5169 14563 5227 14569
rect 5445 14603 5503 14609
rect 5445 14569 5457 14603
rect 5491 14569 5503 14603
rect 5445 14563 5503 14569
rect 6273 14603 6331 14609
rect 6273 14569 6285 14603
rect 6319 14600 6331 14603
rect 6822 14600 6828 14612
rect 6319 14572 6828 14600
rect 6319 14569 6331 14572
rect 6273 14563 6331 14569
rect 4614 14532 4620 14544
rect 4172 14504 4620 14532
rect 4172 14464 4200 14504
rect 4614 14492 4620 14504
rect 4672 14492 4678 14544
rect 4724 14504 5120 14532
rect 3994 14436 4200 14464
rect 3881 14427 3939 14433
rect 1816 14408 1844 14427
rect 1486 14356 1492 14408
rect 1544 14356 1550 14408
rect 1762 14356 1768 14408
rect 1820 14368 1844 14408
rect 2038 14407 2044 14408
rect 1995 14401 2044 14407
rect 1820 14356 1826 14368
rect 1995 14367 2007 14401
rect 2041 14367 2044 14401
rect 1995 14361 2044 14367
rect 2038 14356 2044 14361
rect 2096 14356 2102 14408
rect 2222 14356 2228 14408
rect 2280 14356 2286 14408
rect 3234 14356 3240 14408
rect 3292 14396 3298 14408
rect 3896 14396 3924 14427
rect 4246 14424 4252 14476
rect 4304 14424 4310 14476
rect 4430 14424 4436 14476
rect 4488 14464 4494 14476
rect 4525 14467 4583 14473
rect 4525 14464 4537 14467
rect 4488 14436 4537 14464
rect 4488 14424 4494 14436
rect 4525 14433 4537 14436
rect 4571 14464 4583 14467
rect 4724 14464 4752 14504
rect 5092 14473 5120 14504
rect 5184 14476 5212 14563
rect 5460 14532 5488 14563
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 9030 14560 9036 14612
rect 9088 14560 9094 14612
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 9953 14603 10011 14609
rect 9953 14600 9965 14603
rect 9916 14572 9965 14600
rect 9916 14560 9922 14572
rect 9953 14569 9965 14572
rect 9999 14569 10011 14603
rect 9953 14563 10011 14569
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14569 10655 14603
rect 10597 14563 10655 14569
rect 5810 14532 5816 14544
rect 5460 14504 5816 14532
rect 5810 14492 5816 14504
rect 5868 14492 5874 14544
rect 9048 14532 9076 14560
rect 9309 14535 9367 14541
rect 9309 14532 9321 14535
rect 9048 14504 9321 14532
rect 9309 14501 9321 14504
rect 9355 14501 9367 14535
rect 10318 14532 10324 14544
rect 9309 14495 9367 14501
rect 9646 14504 10324 14532
rect 4571 14436 4752 14464
rect 4801 14467 4859 14473
rect 4571 14433 4583 14436
rect 4525 14427 4583 14433
rect 4801 14433 4813 14467
rect 4847 14433 4859 14467
rect 4801 14427 4859 14433
rect 5077 14467 5135 14473
rect 5077 14433 5089 14467
rect 5123 14433 5135 14467
rect 5077 14427 5135 14433
rect 3292 14368 3924 14396
rect 4264 14396 4292 14424
rect 4816 14396 4844 14427
rect 5166 14424 5172 14476
rect 5224 14424 5230 14476
rect 5258 14424 5264 14476
rect 5316 14464 5322 14476
rect 5353 14471 5411 14477
rect 5353 14464 5365 14471
rect 5316 14437 5365 14464
rect 5399 14464 5411 14471
rect 5442 14464 5448 14476
rect 5399 14437 5448 14464
rect 5316 14436 5448 14437
rect 5316 14424 5322 14436
rect 5353 14431 5411 14436
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 5629 14467 5687 14473
rect 5629 14433 5641 14467
rect 5675 14464 5687 14467
rect 5997 14467 6055 14473
rect 5997 14464 6009 14467
rect 5675 14436 6009 14464
rect 5675 14433 5687 14436
rect 5629 14427 5687 14433
rect 5997 14433 6009 14436
rect 6043 14433 6055 14467
rect 5997 14427 6055 14433
rect 4264 14368 4844 14396
rect 3292 14356 3298 14368
rect 4816 14328 4844 14368
rect 5644 14328 5672 14427
rect 6012 14396 6040 14427
rect 6178 14424 6184 14476
rect 6236 14464 6242 14476
rect 6457 14467 6515 14473
rect 6457 14464 6469 14467
rect 6236 14436 6469 14464
rect 6236 14424 6242 14436
rect 6457 14433 6469 14436
rect 6503 14433 6515 14467
rect 6457 14427 6515 14433
rect 6270 14396 6276 14408
rect 6012 14368 6276 14396
rect 6270 14356 6276 14368
rect 6328 14356 6334 14408
rect 6472 14396 6500 14427
rect 6638 14424 6644 14476
rect 6696 14464 6702 14476
rect 6733 14467 6791 14473
rect 6733 14464 6745 14467
rect 6696 14436 6745 14464
rect 6696 14424 6702 14436
rect 6733 14433 6745 14436
rect 6779 14464 6791 14467
rect 8478 14464 8484 14476
rect 6779 14436 8484 14464
rect 6779 14433 6791 14436
rect 6733 14427 6791 14433
rect 8478 14424 8484 14436
rect 8536 14424 8542 14476
rect 8754 14424 8760 14476
rect 8812 14464 8818 14476
rect 9033 14467 9091 14473
rect 9033 14464 9045 14467
rect 8812 14436 9045 14464
rect 8812 14424 8818 14436
rect 9033 14433 9045 14436
rect 9079 14464 9091 14467
rect 9646 14464 9674 14504
rect 10318 14492 10324 14504
rect 10376 14492 10382 14544
rect 10612 14532 10640 14563
rect 10778 14560 10784 14612
rect 10836 14600 10842 14612
rect 11149 14603 11207 14609
rect 11149 14600 11161 14603
rect 10836 14572 11161 14600
rect 10836 14560 10842 14572
rect 11149 14569 11161 14572
rect 11195 14569 11207 14603
rect 11149 14563 11207 14569
rect 11262 14572 11468 14600
rect 11262 14532 11290 14572
rect 10612 14504 11290 14532
rect 11440 14532 11468 14572
rect 12158 14560 12164 14612
rect 12216 14600 12222 14612
rect 13354 14600 13360 14612
rect 12216 14572 13360 14600
rect 12216 14560 12222 14572
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 16390 14600 16396 14612
rect 13740 14572 16396 14600
rect 11440 14504 11560 14532
rect 9079 14436 9674 14464
rect 9079 14433 9091 14436
rect 9033 14427 9091 14433
rect 9766 14424 9772 14476
rect 9824 14424 9830 14476
rect 10505 14467 10563 14473
rect 9876 14436 10088 14464
rect 6472 14368 6776 14396
rect 6748 14340 6776 14368
rect 6822 14356 6828 14408
rect 6880 14356 6886 14408
rect 7190 14405 7196 14408
rect 7152 14399 7196 14405
rect 7152 14365 7164 14399
rect 7152 14359 7196 14365
rect 7190 14356 7196 14359
rect 7248 14356 7254 14408
rect 7282 14356 7288 14408
rect 7340 14356 7346 14408
rect 7558 14356 7564 14408
rect 7616 14356 7622 14408
rect 8570 14356 8576 14408
rect 8628 14396 8634 14408
rect 9876 14396 9904 14436
rect 10060 14405 10088 14436
rect 10505 14433 10517 14467
rect 10551 14464 10563 14467
rect 10594 14464 10600 14476
rect 10551 14436 10600 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 10686 14424 10692 14476
rect 10744 14464 10750 14476
rect 10781 14467 10839 14473
rect 10781 14464 10793 14467
rect 10744 14436 10793 14464
rect 10744 14424 10750 14436
rect 10781 14433 10793 14436
rect 10827 14433 10839 14467
rect 10781 14427 10839 14433
rect 10870 14424 10876 14476
rect 10928 14464 10934 14476
rect 11057 14467 11115 14473
rect 11057 14464 11069 14467
rect 10928 14436 11069 14464
rect 10928 14424 10934 14436
rect 11057 14433 11069 14436
rect 11103 14433 11115 14467
rect 11057 14427 11115 14433
rect 11422 14424 11428 14476
rect 11480 14424 11486 14476
rect 11532 14464 11560 14504
rect 12345 14467 12403 14473
rect 12345 14464 12357 14467
rect 11532 14436 12357 14464
rect 12345 14433 12357 14436
rect 12391 14433 12403 14467
rect 12345 14427 12403 14433
rect 12618 14424 12624 14476
rect 12676 14464 12682 14476
rect 13170 14464 13176 14476
rect 12676 14436 13176 14464
rect 12676 14424 12682 14436
rect 13170 14424 13176 14436
rect 13228 14424 13234 14476
rect 8628 14368 9904 14396
rect 10045 14399 10103 14405
rect 8628 14356 8634 14368
rect 10045 14365 10057 14399
rect 10091 14365 10103 14399
rect 10612 14396 10640 14424
rect 11330 14396 11336 14408
rect 10612 14368 11336 14396
rect 10045 14359 10103 14365
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 11440 14396 11468 14424
rect 11609 14399 11667 14405
rect 11609 14396 11621 14399
rect 11440 14368 11621 14396
rect 11609 14365 11621 14368
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 11790 14356 11796 14408
rect 11848 14396 11854 14408
rect 11936 14399 11994 14405
rect 11936 14396 11948 14399
rect 11848 14368 11948 14396
rect 11848 14356 11854 14368
rect 11936 14365 11948 14368
rect 11982 14365 11994 14399
rect 11936 14359 11994 14365
rect 12115 14399 12173 14405
rect 12115 14365 12127 14399
rect 12161 14396 12173 14399
rect 13740 14396 13768 14572
rect 16390 14560 16396 14572
rect 16448 14560 16454 14612
rect 16482 14560 16488 14612
rect 16540 14560 16546 14612
rect 16666 14560 16672 14612
rect 16724 14560 16730 14612
rect 17034 14560 17040 14612
rect 17092 14600 17098 14612
rect 17411 14603 17469 14609
rect 17411 14600 17423 14603
rect 17092 14572 17423 14600
rect 17092 14560 17098 14572
rect 17411 14569 17423 14572
rect 17457 14600 17469 14603
rect 17954 14600 17960 14612
rect 17457 14572 17960 14600
rect 17457 14569 17469 14572
rect 17411 14563 17469 14569
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 18782 14560 18788 14612
rect 18840 14560 18846 14612
rect 20993 14603 21051 14609
rect 20993 14569 21005 14603
rect 21039 14600 21051 14603
rect 21542 14600 21548 14612
rect 21039 14572 21548 14600
rect 21039 14569 21051 14572
rect 20993 14563 21051 14569
rect 21542 14560 21548 14572
rect 21600 14560 21606 14612
rect 21634 14560 21640 14612
rect 21692 14600 21698 14612
rect 21735 14603 21793 14609
rect 21735 14600 21747 14603
rect 21692 14572 21747 14600
rect 21692 14560 21698 14572
rect 21735 14569 21747 14572
rect 21781 14569 21793 14603
rect 21735 14563 21793 14569
rect 22094 14560 22100 14612
rect 22152 14600 22158 14612
rect 25317 14603 25375 14609
rect 25317 14600 25329 14603
rect 22152 14572 25329 14600
rect 22152 14560 22158 14572
rect 25317 14569 25329 14572
rect 25363 14569 25375 14603
rect 25317 14563 25375 14569
rect 25406 14560 25412 14612
rect 25464 14600 25470 14612
rect 26970 14600 26976 14612
rect 25464 14572 26976 14600
rect 25464 14560 25470 14572
rect 26970 14560 26976 14572
rect 27028 14560 27034 14612
rect 27614 14560 27620 14612
rect 27672 14600 27678 14612
rect 28261 14603 28319 14609
rect 28261 14600 28273 14603
rect 27672 14572 28273 14600
rect 27672 14560 27678 14572
rect 28261 14569 28273 14572
rect 28307 14569 28319 14603
rect 28261 14563 28319 14569
rect 28350 14560 28356 14612
rect 28408 14600 28414 14612
rect 29178 14600 29184 14612
rect 28408 14572 29184 14600
rect 28408 14560 28414 14572
rect 29178 14560 29184 14572
rect 29236 14560 29242 14612
rect 29270 14560 29276 14612
rect 29328 14600 29334 14612
rect 30377 14603 30435 14609
rect 30377 14600 30389 14603
rect 29328 14572 30389 14600
rect 29328 14560 29334 14572
rect 30377 14569 30389 14572
rect 30423 14569 30435 14603
rect 30377 14563 30435 14569
rect 15378 14492 15384 14544
rect 15436 14532 15442 14544
rect 15933 14535 15991 14541
rect 15933 14532 15945 14535
rect 15436 14504 15945 14532
rect 15436 14492 15442 14504
rect 15933 14501 15945 14504
rect 15979 14501 15991 14535
rect 28166 14532 28172 14544
rect 15933 14495 15991 14501
rect 18340 14504 19564 14532
rect 18340 14476 18368 14504
rect 13906 14424 13912 14476
rect 13964 14464 13970 14476
rect 14553 14468 14611 14473
rect 14108 14467 14611 14468
rect 14108 14464 14565 14467
rect 13964 14440 14565 14464
rect 13964 14436 14136 14440
rect 13964 14424 13970 14436
rect 14553 14433 14565 14440
rect 14599 14433 14611 14467
rect 14553 14427 14611 14433
rect 15010 14424 15016 14476
rect 15068 14464 15074 14476
rect 16209 14467 16267 14473
rect 16209 14464 16221 14467
rect 15068 14436 16221 14464
rect 15068 14424 15074 14436
rect 16209 14433 16221 14436
rect 16255 14433 16267 14467
rect 16209 14427 16267 14433
rect 16853 14467 16911 14473
rect 16853 14433 16865 14467
rect 16899 14433 16911 14467
rect 16853 14427 16911 14433
rect 12161 14368 13768 14396
rect 13817 14399 13875 14405
rect 12161 14365 12173 14368
rect 12115 14359 12173 14365
rect 13817 14365 13829 14399
rect 13863 14365 13875 14399
rect 13817 14359 13875 14365
rect 952 14300 1532 14328
rect 952 14269 980 14300
rect 937 14263 995 14269
rect 937 14229 949 14263
rect 983 14229 995 14263
rect 1504 14260 1532 14300
rect 3436 14300 4108 14328
rect 4816 14300 5672 14328
rect 3436 14260 3464 14300
rect 4080 14272 4108 14300
rect 6362 14288 6368 14340
rect 6420 14328 6426 14340
rect 6420 14300 6684 14328
rect 6420 14288 6426 14300
rect 1504 14232 3464 14260
rect 937 14223 995 14229
rect 3510 14220 3516 14272
rect 3568 14220 3574 14272
rect 3697 14263 3755 14269
rect 3697 14229 3709 14263
rect 3743 14260 3755 14263
rect 3786 14260 3792 14272
rect 3743 14232 3792 14260
rect 3743 14229 3755 14232
rect 3697 14223 3755 14229
rect 3786 14220 3792 14232
rect 3844 14220 3850 14272
rect 4062 14220 4068 14272
rect 4120 14220 4126 14272
rect 4617 14263 4675 14269
rect 4617 14229 4629 14263
rect 4663 14260 4675 14263
rect 5718 14260 5724 14272
rect 4663 14232 5724 14260
rect 4663 14229 4675 14232
rect 4617 14223 4675 14229
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 5810 14220 5816 14272
rect 5868 14220 5874 14272
rect 5902 14220 5908 14272
rect 5960 14260 5966 14272
rect 6549 14263 6607 14269
rect 6549 14260 6561 14263
rect 5960 14232 6561 14260
rect 5960 14220 5966 14232
rect 6549 14229 6561 14232
rect 6595 14229 6607 14263
rect 6656 14260 6684 14300
rect 6730 14288 6736 14340
rect 6788 14288 6794 14340
rect 8849 14331 8907 14337
rect 8849 14297 8861 14331
rect 8895 14328 8907 14331
rect 9674 14328 9680 14340
rect 8895 14300 9680 14328
rect 8895 14297 8907 14300
rect 8849 14291 8907 14297
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 10321 14331 10379 14337
rect 10321 14297 10333 14331
rect 10367 14328 10379 14331
rect 10367 14300 11100 14328
rect 10367 14297 10379 14300
rect 10321 14291 10379 14297
rect 8754 14260 8760 14272
rect 6656 14232 8760 14260
rect 6549 14223 6607 14229
rect 8754 14220 8760 14232
rect 8812 14260 8818 14272
rect 10686 14260 10692 14272
rect 8812 14232 10692 14260
rect 8812 14220 8818 14232
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 11072 14260 11100 14300
rect 12250 14260 12256 14272
rect 11072 14232 12256 14260
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 12342 14220 12348 14272
rect 12400 14260 12406 14272
rect 13449 14263 13507 14269
rect 13449 14260 13461 14263
rect 12400 14232 13461 14260
rect 12400 14220 12406 14232
rect 13449 14229 13461 14232
rect 13495 14229 13507 14263
rect 13832 14260 13860 14359
rect 13998 14356 14004 14408
rect 14056 14396 14062 14408
rect 14366 14407 14372 14408
rect 14144 14399 14202 14405
rect 14144 14396 14156 14399
rect 14056 14368 14156 14396
rect 14056 14356 14062 14368
rect 14144 14365 14156 14368
rect 14190 14365 14202 14399
rect 14144 14359 14202 14365
rect 14323 14401 14372 14407
rect 14323 14367 14335 14401
rect 14369 14367 14372 14401
rect 14323 14361 14372 14367
rect 14366 14356 14372 14361
rect 14424 14356 14430 14408
rect 14458 14356 14464 14408
rect 14516 14396 14522 14408
rect 16298 14396 16304 14408
rect 14516 14368 16304 14396
rect 14516 14356 14522 14368
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 16868 14328 16896 14427
rect 18322 14424 18328 14476
rect 18380 14424 18386 14476
rect 19337 14467 19395 14473
rect 19337 14433 19349 14467
rect 19383 14433 19395 14467
rect 19337 14427 19395 14433
rect 16945 14399 17003 14405
rect 16945 14365 16957 14399
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 16040 14300 16896 14328
rect 16040 14272 16068 14300
rect 14182 14260 14188 14272
rect 13832 14232 14188 14260
rect 13449 14223 13507 14229
rect 14182 14220 14188 14232
rect 14240 14260 14246 14272
rect 15010 14260 15016 14272
rect 14240 14232 15016 14260
rect 14240 14220 14246 14232
rect 15010 14220 15016 14232
rect 15068 14220 15074 14272
rect 16022 14220 16028 14272
rect 16080 14220 16086 14272
rect 16482 14220 16488 14272
rect 16540 14260 16546 14272
rect 16960 14260 16988 14359
rect 17402 14356 17408 14408
rect 17460 14407 17466 14408
rect 17460 14401 17509 14407
rect 17460 14367 17463 14401
rect 17497 14367 17509 14401
rect 17460 14361 17509 14367
rect 17681 14399 17739 14405
rect 17681 14365 17693 14399
rect 17727 14396 17739 14399
rect 19352 14396 19380 14427
rect 19426 14424 19432 14476
rect 19484 14424 19490 14476
rect 19536 14464 19564 14504
rect 27816 14504 28172 14532
rect 19705 14467 19763 14473
rect 19705 14464 19717 14467
rect 19536 14436 19717 14464
rect 19705 14433 19717 14436
rect 19751 14433 19763 14467
rect 19705 14427 19763 14433
rect 21266 14424 21272 14476
rect 21324 14424 21330 14476
rect 23842 14473 23848 14476
rect 23804 14467 23848 14473
rect 23804 14433 23816 14467
rect 23804 14427 23848 14433
rect 23842 14424 23848 14427
rect 23900 14424 23906 14476
rect 24118 14424 24124 14476
rect 24176 14464 24182 14476
rect 24213 14467 24271 14473
rect 24213 14464 24225 14467
rect 24176 14436 24225 14464
rect 24176 14424 24182 14436
rect 24213 14433 24225 14436
rect 24259 14433 24271 14467
rect 24213 14427 24271 14433
rect 24486 14424 24492 14476
rect 24544 14424 24550 14476
rect 25777 14467 25835 14473
rect 25777 14433 25789 14467
rect 25823 14464 25835 14467
rect 25958 14464 25964 14476
rect 25823 14436 25964 14464
rect 25823 14433 25835 14436
rect 25777 14427 25835 14433
rect 25958 14424 25964 14436
rect 26016 14424 26022 14476
rect 26418 14424 26424 14476
rect 26476 14424 26482 14476
rect 26694 14464 26700 14476
rect 26528 14436 26700 14464
rect 21765 14417 21823 14423
rect 17727 14368 19196 14396
rect 19352 14368 20576 14396
rect 17727 14365 17739 14368
rect 17460 14356 17466 14361
rect 17681 14359 17739 14365
rect 19168 14337 19196 14368
rect 20548 14340 20576 14368
rect 21174 14356 21180 14408
rect 21232 14356 21238 14408
rect 21765 14383 21777 14417
rect 21811 14396 21823 14417
rect 21910 14396 21916 14408
rect 21811 14383 21916 14396
rect 21765 14377 21916 14383
rect 21790 14368 21916 14377
rect 21910 14356 21916 14368
rect 21968 14356 21974 14408
rect 22002 14356 22008 14408
rect 22060 14356 22066 14408
rect 23477 14399 23535 14405
rect 23477 14365 23489 14399
rect 23523 14396 23535 14399
rect 23658 14396 23664 14408
rect 23523 14368 23664 14396
rect 23523 14365 23535 14368
rect 23477 14359 23535 14365
rect 23658 14356 23664 14368
rect 23716 14356 23722 14408
rect 23983 14399 24041 14405
rect 23983 14365 23995 14399
rect 24029 14396 24041 14399
rect 24504 14396 24532 14424
rect 24029 14368 24532 14396
rect 24029 14365 24041 14368
rect 23983 14359 24041 14365
rect 24854 14356 24860 14408
rect 24912 14396 24918 14408
rect 26053 14399 26111 14405
rect 26053 14396 26065 14399
rect 24912 14368 26065 14396
rect 24912 14356 24918 14368
rect 26053 14365 26065 14368
rect 26099 14396 26111 14399
rect 26528 14396 26556 14436
rect 26694 14424 26700 14436
rect 26752 14473 26758 14476
rect 26752 14467 26806 14473
rect 26752 14433 26760 14467
rect 26794 14464 26806 14467
rect 27816 14464 27844 14504
rect 28166 14492 28172 14504
rect 28224 14492 28230 14544
rect 31294 14532 31300 14544
rect 29932 14504 31300 14532
rect 26794 14436 27844 14464
rect 26794 14433 26806 14436
rect 26752 14427 26806 14433
rect 26752 14424 26758 14427
rect 27982 14424 27988 14476
rect 28040 14464 28046 14476
rect 28905 14467 28963 14473
rect 28905 14464 28917 14467
rect 28040 14436 28917 14464
rect 28040 14424 28046 14436
rect 28905 14433 28917 14436
rect 28951 14433 28963 14467
rect 28905 14427 28963 14433
rect 29178 14424 29184 14476
rect 29236 14464 29242 14476
rect 29932 14464 29960 14504
rect 31294 14492 31300 14504
rect 31352 14492 31358 14544
rect 29236 14436 29960 14464
rect 29236 14424 29242 14436
rect 30006 14424 30012 14476
rect 30064 14464 30070 14476
rect 30190 14464 30196 14476
rect 30064 14436 30196 14464
rect 30064 14424 30070 14436
rect 30190 14424 30196 14436
rect 30248 14464 30254 14476
rect 30561 14467 30619 14473
rect 30561 14464 30573 14467
rect 30248 14436 30573 14464
rect 30248 14424 30254 14436
rect 30561 14433 30573 14436
rect 30607 14433 30619 14467
rect 30561 14427 30619 14433
rect 26099 14368 26556 14396
rect 26927 14399 26985 14405
rect 26099 14365 26111 14368
rect 26053 14359 26111 14365
rect 26927 14365 26939 14399
rect 26973 14396 26985 14399
rect 27062 14396 27068 14408
rect 26973 14368 27068 14396
rect 26973 14365 26985 14368
rect 26927 14359 26985 14365
rect 27062 14356 27068 14368
rect 27120 14356 27126 14408
rect 27157 14399 27215 14405
rect 27157 14365 27169 14399
rect 27203 14396 27215 14399
rect 27522 14396 27528 14408
rect 27203 14368 27528 14396
rect 27203 14365 27215 14368
rect 27157 14359 27215 14365
rect 27522 14356 27528 14368
rect 27580 14356 27586 14408
rect 28629 14399 28687 14405
rect 28629 14396 28641 14399
rect 27816 14368 28641 14396
rect 19153 14331 19211 14337
rect 19153 14297 19165 14331
rect 19199 14297 19211 14331
rect 19153 14291 19211 14297
rect 20530 14288 20536 14340
rect 20588 14288 20594 14340
rect 16540 14232 16988 14260
rect 16540 14220 16546 14232
rect 18138 14220 18144 14272
rect 18196 14260 18202 14272
rect 21192 14260 21220 14356
rect 18196 14232 21220 14260
rect 18196 14220 18202 14232
rect 21266 14220 21272 14272
rect 21324 14260 21330 14272
rect 23109 14263 23167 14269
rect 23109 14260 23121 14263
rect 21324 14232 23121 14260
rect 21324 14220 21330 14232
rect 23109 14229 23121 14232
rect 23155 14229 23167 14263
rect 23109 14223 23167 14229
rect 24026 14220 24032 14272
rect 24084 14260 24090 14272
rect 26786 14260 26792 14272
rect 24084 14232 26792 14260
rect 24084 14220 24090 14232
rect 26786 14220 26792 14232
rect 26844 14220 26850 14272
rect 26970 14220 26976 14272
rect 27028 14260 27034 14272
rect 27816 14260 27844 14368
rect 28629 14365 28641 14368
rect 28675 14365 28687 14399
rect 28629 14359 28687 14365
rect 27028 14232 27844 14260
rect 27028 14220 27034 14232
rect 28626 14220 28632 14272
rect 28684 14260 28690 14272
rect 30009 14263 30067 14269
rect 30009 14260 30021 14263
rect 28684 14232 30021 14260
rect 28684 14220 28690 14232
rect 30009 14229 30021 14232
rect 30055 14229 30067 14263
rect 30009 14223 30067 14229
rect 552 14170 30912 14192
rect 552 14118 4193 14170
rect 4245 14118 4257 14170
rect 4309 14118 4321 14170
rect 4373 14118 4385 14170
rect 4437 14118 4449 14170
rect 4501 14118 11783 14170
rect 11835 14118 11847 14170
rect 11899 14118 11911 14170
rect 11963 14118 11975 14170
rect 12027 14118 12039 14170
rect 12091 14118 19373 14170
rect 19425 14118 19437 14170
rect 19489 14118 19501 14170
rect 19553 14118 19565 14170
rect 19617 14118 19629 14170
rect 19681 14118 26963 14170
rect 27015 14118 27027 14170
rect 27079 14118 27091 14170
rect 27143 14118 27155 14170
rect 27207 14118 27219 14170
rect 27271 14118 30912 14170
rect 552 14096 30912 14118
rect 1118 14016 1124 14068
rect 1176 14056 1182 14068
rect 1176 14028 2360 14056
rect 1176 14016 1182 14028
rect 2038 13920 2044 13932
rect 1412 13905 2044 13920
rect 1412 13874 1445 13905
rect 1433 13871 1445 13874
rect 1479 13892 2044 13905
rect 1479 13871 1491 13892
rect 2038 13880 2044 13892
rect 2096 13880 2102 13932
rect 2332 13920 2360 14028
rect 2774 14016 2780 14068
rect 2832 14016 2838 14068
rect 3418 14016 3424 14068
rect 3476 14056 3482 14068
rect 5718 14056 5724 14068
rect 3476 14028 5724 14056
rect 3476 14016 3482 14028
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 5810 14016 5816 14068
rect 5868 14016 5874 14068
rect 6914 14056 6920 14068
rect 5920 14028 6920 14056
rect 3329 13991 3387 13997
rect 3329 13957 3341 13991
rect 3375 13988 3387 13991
rect 3602 13988 3608 14000
rect 3375 13960 3608 13988
rect 3375 13957 3387 13960
rect 3329 13951 3387 13957
rect 3602 13948 3608 13960
rect 3660 13948 3666 14000
rect 4522 13920 4528 13932
rect 2332 13892 3832 13920
rect 1433 13865 1491 13871
rect 937 13855 995 13861
rect 937 13821 949 13855
rect 983 13852 995 13855
rect 1210 13852 1216 13864
rect 983 13824 1216 13852
rect 983 13821 995 13824
rect 937 13815 995 13821
rect 1210 13812 1216 13824
rect 1268 13812 1274 13864
rect 1670 13812 1676 13864
rect 1728 13812 1734 13864
rect 2498 13812 2504 13864
rect 2556 13852 2562 13864
rect 3804 13861 3832 13892
rect 4356 13905 4528 13920
rect 4356 13874 4389 13905
rect 4377 13871 4389 13874
rect 4423 13892 4528 13905
rect 4423 13871 4435 13892
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 4617 13923 4675 13929
rect 4617 13889 4629 13923
rect 4663 13920 4675 13923
rect 5828 13920 5856 14016
rect 5920 13997 5948 14028
rect 6914 14016 6920 14028
rect 6972 14016 6978 14068
rect 7006 14016 7012 14068
rect 7064 14056 7070 14068
rect 7064 14028 7512 14056
rect 7064 14016 7070 14028
rect 5905 13991 5963 13997
rect 5905 13957 5917 13991
rect 5951 13957 5963 13991
rect 7484 13988 7512 14028
rect 7742 14016 7748 14068
rect 7800 14056 7806 14068
rect 7929 14059 7987 14065
rect 7929 14056 7941 14059
rect 7800 14028 7941 14056
rect 7800 14016 7806 14028
rect 7929 14025 7941 14028
rect 7975 14025 7987 14059
rect 7929 14019 7987 14025
rect 8481 14059 8539 14065
rect 8481 14025 8493 14059
rect 8527 14056 8539 14059
rect 8938 14056 8944 14068
rect 8527 14028 8944 14056
rect 8527 14025 8539 14028
rect 8481 14019 8539 14025
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 9214 14016 9220 14068
rect 9272 14016 9278 14068
rect 9306 14016 9312 14068
rect 9364 14056 9370 14068
rect 9401 14059 9459 14065
rect 9401 14056 9413 14059
rect 9364 14028 9413 14056
rect 9364 14016 9370 14028
rect 9401 14025 9413 14028
rect 9447 14025 9459 14059
rect 12342 14056 12348 14068
rect 9401 14019 9459 14025
rect 9692 14028 12348 14056
rect 8757 13991 8815 13997
rect 8757 13988 8769 13991
rect 7484 13960 8769 13988
rect 5905 13951 5963 13957
rect 8757 13957 8769 13960
rect 8803 13957 8815 13991
rect 8757 13951 8815 13957
rect 8846 13948 8852 14000
rect 8904 13988 8910 14000
rect 9692 13988 9720 14028
rect 12342 14016 12348 14028
rect 12400 14016 12406 14068
rect 12434 14016 12440 14068
rect 12492 14016 12498 14068
rect 12526 14016 12532 14068
rect 12584 14056 12590 14068
rect 12989 14059 13047 14065
rect 12989 14056 13001 14059
rect 12584 14028 13001 14056
rect 12584 14016 12590 14028
rect 12989 14025 13001 14028
rect 13035 14025 13047 14059
rect 12989 14019 13047 14025
rect 13464 14028 13768 14056
rect 8904 13960 9720 13988
rect 8904 13948 8910 13960
rect 11698 13948 11704 14000
rect 11756 13988 11762 14000
rect 11756 13960 12204 13988
rect 11756 13948 11762 13960
rect 6454 13929 6460 13932
rect 6416 13923 6460 13929
rect 4663 13892 5856 13920
rect 6012 13892 6224 13920
rect 4663 13889 4675 13892
rect 4617 13883 4675 13889
rect 4377 13865 4435 13871
rect 3513 13855 3571 13861
rect 2556 13824 3464 13852
rect 2556 13812 2562 13824
rect 3436 13784 3464 13824
rect 3513 13821 3525 13855
rect 3559 13852 3571 13855
rect 3789 13855 3847 13861
rect 3559 13824 3746 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 3718 13784 3746 13824
rect 3789 13821 3801 13855
rect 3835 13821 3847 13855
rect 3789 13815 3847 13821
rect 3878 13812 3884 13864
rect 3936 13812 3942 13864
rect 4246 13852 4252 13864
rect 3994 13824 4252 13852
rect 3994 13784 4022 13824
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 5074 13812 5080 13864
rect 5132 13852 5138 13864
rect 6012 13852 6040 13892
rect 5132 13824 6040 13852
rect 5132 13812 5138 13824
rect 6086 13812 6092 13864
rect 6144 13812 6150 13864
rect 6196 13852 6224 13892
rect 6416 13889 6428 13923
rect 6416 13883 6460 13889
rect 6454 13880 6460 13883
rect 6512 13880 6518 13932
rect 6595 13923 6653 13929
rect 6595 13889 6607 13923
rect 6641 13920 6653 13923
rect 6641 13892 10088 13920
rect 6641 13889 6653 13892
rect 6595 13883 6653 13889
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6196 13824 6837 13852
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13852 8723 13855
rect 8711 13824 8892 13852
rect 8711 13821 8723 13824
rect 8665 13815 8723 13821
rect 3436 13756 3648 13784
rect 3718 13756 4022 13784
rect 8864 13784 8892 13824
rect 8938 13812 8944 13864
rect 8996 13812 9002 13864
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13852 9091 13855
rect 9079 13824 9352 13852
rect 9079 13821 9091 13824
rect 9033 13815 9091 13821
rect 9048 13784 9076 13815
rect 8864 13756 9076 13784
rect 9324 13784 9352 13824
rect 9398 13812 9404 13864
rect 9456 13852 9462 13864
rect 9585 13855 9643 13861
rect 9585 13852 9597 13855
rect 9456 13824 9597 13852
rect 9456 13812 9462 13824
rect 9585 13821 9597 13824
rect 9631 13821 9643 13855
rect 9585 13815 9643 13821
rect 9674 13812 9680 13864
rect 9732 13812 9738 13864
rect 9950 13852 9956 13864
rect 9784 13824 9956 13852
rect 9784 13784 9812 13824
rect 9950 13812 9956 13824
rect 10008 13812 10014 13864
rect 10060 13852 10088 13892
rect 10134 13880 10140 13932
rect 10192 13880 10198 13932
rect 12066 13920 12072 13932
rect 10244 13892 12072 13920
rect 10244 13852 10272 13892
rect 12066 13880 12072 13892
rect 12124 13880 12130 13932
rect 10060 13824 10272 13852
rect 10410 13812 10416 13864
rect 10468 13812 10474 13864
rect 11514 13812 11520 13864
rect 11572 13812 11578 13864
rect 11790 13812 11796 13864
rect 11848 13812 11854 13864
rect 12176 13861 12204 13960
rect 12710 13948 12716 14000
rect 12768 13948 12774 14000
rect 11885 13855 11943 13861
rect 11885 13821 11897 13855
rect 11931 13852 11943 13855
rect 12161 13855 12219 13861
rect 11931 13824 12118 13852
rect 11931 13821 11943 13824
rect 11885 13815 11943 13821
rect 9324 13756 9812 13784
rect 11532 13784 11560 13812
rect 12090 13784 12118 13824
rect 12161 13821 12173 13855
rect 12207 13821 12219 13855
rect 12161 13815 12219 13821
rect 12618 13812 12624 13864
rect 12676 13812 12682 13864
rect 12894 13812 12900 13864
rect 12952 13812 12958 13864
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13852 13231 13855
rect 13464 13852 13492 14028
rect 13633 13991 13691 13997
rect 13633 13957 13645 13991
rect 13679 13957 13691 13991
rect 13740 13988 13768 14028
rect 13906 14016 13912 14068
rect 13964 14016 13970 14068
rect 18874 14056 18880 14068
rect 16408 14028 18880 14056
rect 14090 13988 14096 14000
rect 13740 13960 14096 13988
rect 13633 13951 13691 13957
rect 13648 13920 13676 13951
rect 14090 13948 14096 13960
rect 14148 13948 14154 14000
rect 14691 13923 14749 13929
rect 13648 13892 14320 13920
rect 13219 13824 13492 13852
rect 13817 13855 13875 13861
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 13817 13821 13829 13855
rect 13863 13821 13875 13855
rect 13817 13815 13875 13821
rect 11532 13756 12118 13784
rect 1394 13676 1400 13728
rect 1452 13725 1458 13728
rect 3620 13725 3648 13756
rect 1452 13679 1461 13725
rect 3605 13719 3663 13725
rect 3605 13685 3617 13719
rect 3651 13685 3663 13719
rect 3605 13679 3663 13685
rect 1452 13676 1458 13679
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 4347 13719 4405 13725
rect 4347 13716 4359 13719
rect 4028 13688 4359 13716
rect 4028 13676 4034 13688
rect 4347 13685 4359 13688
rect 4393 13685 4405 13719
rect 4347 13679 4405 13685
rect 9582 13676 9588 13728
rect 9640 13716 9646 13728
rect 10143 13719 10201 13725
rect 10143 13716 10155 13719
rect 9640 13688 10155 13716
rect 9640 13676 9646 13688
rect 10143 13685 10155 13688
rect 10189 13685 10201 13719
rect 10143 13679 10201 13685
rect 10686 13676 10692 13728
rect 10744 13716 10750 13728
rect 11514 13716 11520 13728
rect 10744 13688 11520 13716
rect 10744 13676 10750 13688
rect 11514 13676 11520 13688
rect 11572 13676 11578 13728
rect 12090 13716 12118 13756
rect 12710 13744 12716 13796
rect 12768 13784 12774 13796
rect 13722 13784 13728 13796
rect 12768 13756 13728 13784
rect 12768 13744 12774 13756
rect 13722 13744 13728 13756
rect 13780 13784 13786 13796
rect 13832 13784 13860 13815
rect 14090 13812 14096 13864
rect 14148 13812 14154 13864
rect 14182 13812 14188 13864
rect 14240 13812 14246 13864
rect 14292 13852 14320 13892
rect 14691 13889 14703 13923
rect 14737 13920 14749 13923
rect 16408 13920 16436 14028
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 18966 14016 18972 14068
rect 19024 14016 19030 14068
rect 19613 14059 19671 14065
rect 19613 14025 19625 14059
rect 19659 14056 19671 14059
rect 20346 14056 20352 14068
rect 19659 14028 20352 14056
rect 19659 14025 19671 14028
rect 19613 14019 19671 14025
rect 20346 14016 20352 14028
rect 20404 14016 20410 14068
rect 22741 14059 22799 14065
rect 22741 14025 22753 14059
rect 22787 14056 22799 14059
rect 22922 14056 22928 14068
rect 22787 14028 22928 14056
rect 22787 14025 22799 14028
rect 22741 14019 22799 14025
rect 22922 14016 22928 14028
rect 22980 14016 22986 14068
rect 23014 14016 23020 14068
rect 23072 14016 23078 14068
rect 24213 14059 24271 14065
rect 24213 14025 24225 14059
rect 24259 14056 24271 14059
rect 26513 14059 26571 14065
rect 24259 14028 25912 14056
rect 24259 14025 24271 14028
rect 24213 14019 24271 14025
rect 19245 13991 19303 13997
rect 19245 13957 19257 13991
rect 19291 13957 19303 13991
rect 19245 13951 19303 13957
rect 22189 13991 22247 13997
rect 22189 13957 22201 13991
rect 22235 13988 22247 13991
rect 23566 13988 23572 14000
rect 22235 13960 23572 13988
rect 22235 13957 22247 13960
rect 22189 13951 22247 13957
rect 16942 13929 16948 13932
rect 14737 13892 16436 13920
rect 16899 13923 16948 13929
rect 14737 13889 14749 13892
rect 14691 13883 14749 13889
rect 16899 13889 16911 13923
rect 16945 13889 16948 13923
rect 16899 13883 16948 13889
rect 16942 13880 16948 13883
rect 17000 13880 17006 13932
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13920 17187 13923
rect 19260 13920 19288 13951
rect 23566 13948 23572 13960
rect 23624 13948 23630 14000
rect 23937 13991 23995 13997
rect 23937 13957 23949 13991
rect 23983 13957 23995 13991
rect 23937 13951 23995 13957
rect 20352 13923 20410 13929
rect 20352 13920 20364 13923
rect 17175 13892 19288 13920
rect 20180 13892 20364 13920
rect 17175 13889 17187 13892
rect 17129 13883 17187 13889
rect 20180 13864 20208 13892
rect 20352 13889 20364 13892
rect 20398 13889 20410 13923
rect 23750 13920 23756 13932
rect 20352 13883 20410 13889
rect 20548 13892 23756 13920
rect 14921 13855 14979 13861
rect 14921 13852 14933 13855
rect 14292 13824 14933 13852
rect 14921 13821 14933 13824
rect 14967 13821 14979 13855
rect 14921 13815 14979 13821
rect 15194 13812 15200 13864
rect 15252 13852 15258 13864
rect 16301 13855 16359 13861
rect 16301 13852 16313 13855
rect 15252 13824 16313 13852
rect 15252 13812 15258 13824
rect 16301 13821 16313 13824
rect 16347 13821 16359 13855
rect 16301 13815 16359 13821
rect 16393 13855 16451 13861
rect 16393 13821 16405 13855
rect 16439 13852 16451 13855
rect 16482 13852 16488 13864
rect 16439 13824 16488 13852
rect 16439 13821 16451 13824
rect 16393 13815 16451 13821
rect 16482 13812 16488 13824
rect 16540 13852 16546 13864
rect 17034 13852 17040 13864
rect 16540 13824 17040 13852
rect 16540 13812 16546 13824
rect 17034 13812 17040 13824
rect 17092 13812 17098 13864
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 18874 13852 18880 13864
rect 18012 13824 18880 13852
rect 18012 13812 18018 13824
rect 18874 13812 18880 13824
rect 18932 13812 18938 13864
rect 19150 13812 19156 13864
rect 19208 13852 19214 13864
rect 19429 13855 19487 13861
rect 19208 13824 19288 13852
rect 19208 13812 19214 13824
rect 13780 13756 13860 13784
rect 13780 13744 13786 13756
rect 13906 13744 13912 13796
rect 13964 13744 13970 13796
rect 13924 13716 13952 13744
rect 12090 13688 13952 13716
rect 14200 13716 14228 13812
rect 19260 13728 19288 13824
rect 19429 13821 19441 13855
rect 19475 13852 19487 13855
rect 19797 13855 19855 13861
rect 19797 13852 19809 13855
rect 19475 13824 19809 13852
rect 19475 13821 19487 13824
rect 19429 13815 19487 13821
rect 19797 13821 19809 13824
rect 19843 13821 19855 13855
rect 19797 13815 19855 13821
rect 19812 13728 19840 13815
rect 19886 13812 19892 13864
rect 19944 13812 19950 13864
rect 20162 13812 20168 13864
rect 20220 13812 20226 13864
rect 20254 13812 20260 13864
rect 20312 13852 20318 13864
rect 20548 13852 20576 13892
rect 20312 13824 20576 13852
rect 20312 13812 20318 13824
rect 20622 13812 20628 13864
rect 20680 13812 20686 13864
rect 22005 13855 22063 13861
rect 22005 13821 22017 13855
rect 22051 13852 22063 13855
rect 22278 13852 22284 13864
rect 22051 13824 22284 13852
rect 22051 13821 22063 13824
rect 22005 13815 22063 13821
rect 22278 13812 22284 13824
rect 22336 13812 22342 13864
rect 22388 13861 22416 13892
rect 23676 13861 23704 13892
rect 23750 13880 23756 13892
rect 23808 13880 23814 13932
rect 23952 13920 23980 13951
rect 24854 13929 24860 13932
rect 24816 13923 24860 13929
rect 23952 13892 24624 13920
rect 22373 13855 22431 13861
rect 22373 13821 22385 13855
rect 22419 13821 22431 13855
rect 22373 13815 22431 13821
rect 22925 13855 22983 13861
rect 22925 13821 22937 13855
rect 22971 13821 22983 13855
rect 22925 13815 22983 13821
rect 23201 13855 23259 13861
rect 23201 13821 23213 13855
rect 23247 13821 23259 13855
rect 23201 13815 23259 13821
rect 23661 13855 23719 13861
rect 23661 13821 23673 13855
rect 23707 13821 23719 13855
rect 23661 13815 23719 13821
rect 24121 13855 24179 13861
rect 24121 13821 24133 13855
rect 24167 13821 24179 13855
rect 24121 13815 24179 13821
rect 22940 13784 22968 13815
rect 23014 13784 23020 13796
rect 22940 13756 23020 13784
rect 23014 13744 23020 13756
rect 23072 13744 23078 13796
rect 23216 13784 23244 13815
rect 24136 13784 24164 13815
rect 24394 13812 24400 13864
rect 24452 13812 24458 13864
rect 24489 13855 24547 13861
rect 24489 13821 24501 13855
rect 24535 13821 24547 13855
rect 24596 13852 24624 13892
rect 24816 13889 24828 13923
rect 24816 13883 24860 13889
rect 24854 13880 24860 13883
rect 24912 13880 24918 13932
rect 24995 13923 25053 13929
rect 24995 13889 25007 13923
rect 25041 13920 25053 13923
rect 25884 13920 25912 14028
rect 26513 14025 26525 14059
rect 26559 14056 26571 14059
rect 26878 14056 26884 14068
rect 26559 14028 26884 14056
rect 26559 14025 26571 14028
rect 26513 14019 26571 14025
rect 26878 14016 26884 14028
rect 26936 14016 26942 14068
rect 28074 14016 28080 14068
rect 28132 14056 28138 14068
rect 28997 14059 29055 14065
rect 28997 14056 29009 14059
rect 28132 14028 29009 14056
rect 28132 14016 28138 14028
rect 28997 14025 29009 14028
rect 29043 14025 29055 14059
rect 28997 14019 29055 14025
rect 29086 14016 29092 14068
rect 29144 14056 29150 14068
rect 29273 14059 29331 14065
rect 29273 14056 29285 14059
rect 29144 14028 29285 14056
rect 29144 14016 29150 14028
rect 29273 14025 29285 14028
rect 29319 14025 29331 14059
rect 29273 14019 29331 14025
rect 29549 14059 29607 14065
rect 29549 14025 29561 14059
rect 29595 14056 29607 14059
rect 29730 14056 29736 14068
rect 29595 14028 29736 14056
rect 29595 14025 29607 14028
rect 29549 14019 29607 14025
rect 29730 14016 29736 14028
rect 29788 14016 29794 14068
rect 30558 14016 30564 14068
rect 30616 14016 30622 14068
rect 28537 13991 28595 13997
rect 28537 13957 28549 13991
rect 28583 13957 28595 13991
rect 29638 13988 29644 14000
rect 28537 13951 28595 13957
rect 29196 13960 29644 13988
rect 25041 13892 25728 13920
rect 25884 13892 26832 13920
rect 25041 13889 25053 13892
rect 24995 13883 25053 13889
rect 25700 13864 25728 13892
rect 25225 13855 25283 13861
rect 25225 13852 25237 13855
rect 24596 13824 25237 13852
rect 24489 13815 24547 13821
rect 25225 13821 25237 13824
rect 25271 13821 25283 13855
rect 25225 13815 25283 13821
rect 24302 13784 24308 13796
rect 23216 13756 24308 13784
rect 14550 13716 14556 13728
rect 14200 13688 14556 13716
rect 14550 13676 14556 13688
rect 14608 13676 14614 13728
rect 14651 13719 14709 13725
rect 14651 13685 14663 13719
rect 14697 13716 14709 13719
rect 14918 13716 14924 13728
rect 14697 13688 14924 13716
rect 14697 13685 14709 13688
rect 14651 13679 14709 13685
rect 14918 13676 14924 13688
rect 14976 13676 14982 13728
rect 16859 13719 16917 13725
rect 16859 13685 16871 13719
rect 16905 13716 16917 13719
rect 17126 13716 17132 13728
rect 16905 13688 17132 13716
rect 16905 13685 16917 13688
rect 16859 13679 16917 13685
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 18230 13676 18236 13728
rect 18288 13676 18294 13728
rect 18690 13676 18696 13728
rect 18748 13676 18754 13728
rect 19242 13676 19248 13728
rect 19300 13676 19306 13728
rect 19794 13676 19800 13728
rect 19852 13716 19858 13728
rect 20254 13716 20260 13728
rect 19852 13688 20260 13716
rect 19852 13676 19858 13688
rect 20254 13676 20260 13688
rect 20312 13676 20318 13728
rect 20355 13719 20413 13725
rect 20355 13685 20367 13719
rect 20401 13716 20413 13719
rect 20898 13716 20904 13728
rect 20401 13688 20904 13716
rect 20401 13685 20413 13688
rect 20355 13679 20413 13685
rect 20898 13676 20904 13688
rect 20956 13676 20962 13728
rect 22830 13676 22836 13728
rect 22888 13716 22894 13728
rect 23216 13716 23244 13756
rect 24302 13744 24308 13756
rect 24360 13744 24366 13796
rect 24504 13784 24532 13815
rect 25682 13812 25688 13864
rect 25740 13812 25746 13864
rect 26142 13812 26148 13864
rect 26200 13812 26206 13864
rect 26418 13812 26424 13864
rect 26476 13852 26482 13864
rect 26697 13855 26755 13861
rect 26697 13852 26709 13855
rect 26476 13824 26709 13852
rect 26476 13812 26482 13824
rect 26697 13821 26709 13824
rect 26743 13821 26755 13855
rect 26804 13852 26832 13892
rect 26878 13880 26884 13932
rect 26936 13920 26942 13932
rect 27160 13923 27218 13929
rect 27160 13920 27172 13923
rect 26936 13892 27172 13920
rect 26936 13880 26942 13892
rect 27160 13889 27172 13892
rect 27206 13889 27218 13923
rect 27160 13883 27218 13889
rect 27614 13880 27620 13932
rect 27672 13920 27678 13932
rect 28552 13920 28580 13951
rect 27672 13892 28580 13920
rect 27672 13880 27678 13892
rect 27433 13855 27491 13861
rect 27433 13852 27445 13855
rect 26804 13824 27445 13852
rect 26697 13815 26755 13821
rect 27433 13821 27445 13824
rect 27479 13821 27491 13855
rect 28166 13852 28172 13864
rect 27433 13815 27491 13821
rect 28092 13824 28172 13852
rect 24578 13784 24584 13796
rect 24504 13756 24584 13784
rect 24578 13744 24584 13756
rect 24636 13744 24642 13796
rect 22888 13688 23244 13716
rect 23477 13719 23535 13725
rect 22888 13676 22894 13688
rect 23477 13685 23489 13719
rect 23523 13716 23535 13719
rect 25314 13716 25320 13728
rect 23523 13688 25320 13716
rect 23523 13685 23535 13688
rect 23477 13679 23535 13685
rect 25314 13676 25320 13688
rect 25372 13676 25378 13728
rect 25590 13676 25596 13728
rect 25648 13716 25654 13728
rect 26050 13716 26056 13728
rect 25648 13688 26056 13716
rect 25648 13676 25654 13688
rect 26050 13676 26056 13688
rect 26108 13676 26114 13728
rect 26160 13716 26188 13812
rect 27062 13716 27068 13728
rect 26160 13688 27068 13716
rect 27062 13676 27068 13688
rect 27120 13676 27126 13728
rect 27163 13719 27221 13725
rect 27163 13685 27175 13719
rect 27209 13716 27221 13719
rect 28092 13716 28120 13824
rect 28166 13812 28172 13824
rect 28224 13812 28230 13864
rect 29196 13861 29224 13960
rect 29638 13948 29644 13960
rect 29696 13988 29702 14000
rect 30576 13988 30604 14016
rect 29696 13960 30604 13988
rect 29696 13948 29702 13960
rect 29914 13920 29920 13932
rect 29748 13892 29920 13920
rect 29748 13861 29776 13892
rect 29914 13880 29920 13892
rect 29972 13920 29978 13932
rect 30466 13920 30472 13932
rect 29972 13892 30472 13920
rect 29972 13880 29978 13892
rect 30466 13880 30472 13892
rect 30524 13880 30530 13932
rect 29181 13855 29239 13861
rect 29181 13821 29193 13855
rect 29227 13821 29239 13855
rect 29181 13815 29239 13821
rect 29457 13855 29515 13861
rect 29457 13821 29469 13855
rect 29503 13852 29515 13855
rect 29733 13855 29791 13861
rect 29503 13824 29592 13852
rect 29503 13821 29515 13824
rect 29457 13815 29515 13821
rect 29564 13796 29592 13824
rect 29733 13821 29745 13855
rect 29779 13821 29791 13855
rect 29733 13815 29791 13821
rect 29546 13744 29552 13796
rect 29604 13784 29610 13796
rect 30098 13784 30104 13796
rect 29604 13756 30104 13784
rect 29604 13744 29610 13756
rect 30098 13744 30104 13756
rect 30156 13744 30162 13796
rect 27209 13688 28120 13716
rect 27209 13685 27221 13688
rect 27163 13679 27221 13685
rect 28166 13676 28172 13728
rect 28224 13716 28230 13728
rect 28810 13716 28816 13728
rect 28224 13688 28816 13716
rect 28224 13676 28230 13688
rect 28810 13676 28816 13688
rect 28868 13676 28874 13728
rect 552 13626 31072 13648
rect 552 13574 7988 13626
rect 8040 13574 8052 13626
rect 8104 13574 8116 13626
rect 8168 13574 8180 13626
rect 8232 13574 8244 13626
rect 8296 13574 15578 13626
rect 15630 13574 15642 13626
rect 15694 13574 15706 13626
rect 15758 13574 15770 13626
rect 15822 13574 15834 13626
rect 15886 13574 23168 13626
rect 23220 13574 23232 13626
rect 23284 13574 23296 13626
rect 23348 13574 23360 13626
rect 23412 13574 23424 13626
rect 23476 13574 30758 13626
rect 30810 13574 30822 13626
rect 30874 13574 30886 13626
rect 30938 13574 30950 13626
rect 31002 13574 31014 13626
rect 31066 13574 31072 13626
rect 552 13552 31072 13574
rect 1762 13472 1768 13524
rect 1820 13521 1826 13524
rect 1820 13512 1829 13521
rect 1820 13484 1865 13512
rect 1820 13475 1829 13484
rect 1820 13472 1826 13475
rect 3970 13472 3976 13524
rect 4028 13521 4034 13524
rect 4028 13512 4037 13521
rect 4028 13484 4073 13512
rect 4028 13475 4037 13484
rect 4028 13472 4034 13475
rect 6546 13472 6552 13524
rect 6604 13472 6610 13524
rect 8754 13472 8760 13524
rect 8812 13472 8818 13524
rect 9398 13472 9404 13524
rect 9456 13472 9462 13524
rect 9769 13515 9827 13521
rect 9769 13481 9781 13515
rect 9815 13512 9827 13515
rect 9858 13512 9864 13524
rect 9815 13484 9864 13512
rect 9815 13481 9827 13484
rect 9769 13475 9827 13481
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 10870 13512 10876 13524
rect 10244 13484 10876 13512
rect 3436 13416 3648 13444
rect 1213 13379 1271 13385
rect 1213 13376 1225 13379
rect 1136 13348 1225 13376
rect 1136 13320 1164 13348
rect 1213 13345 1225 13348
rect 1259 13345 1271 13379
rect 3142 13376 3148 13388
rect 1213 13339 1271 13345
rect 1826 13348 3148 13376
rect 1118 13268 1124 13320
rect 1176 13268 1182 13320
rect 1302 13268 1308 13320
rect 1360 13308 1366 13320
rect 1486 13308 1492 13320
rect 1360 13280 1492 13308
rect 1360 13268 1366 13280
rect 1486 13268 1492 13280
rect 1544 13268 1550 13320
rect 1826 13319 1854 13348
rect 3142 13336 3148 13348
rect 3200 13336 3206 13388
rect 3436 13385 3464 13416
rect 3421 13379 3479 13385
rect 3421 13345 3433 13379
rect 3467 13345 3479 13379
rect 3421 13339 3479 13345
rect 3513 13379 3571 13385
rect 3513 13345 3525 13379
rect 3559 13345 3571 13379
rect 3513 13339 3571 13345
rect 1811 13313 1869 13319
rect 1811 13279 1823 13313
rect 1857 13279 1869 13313
rect 1811 13273 1869 13279
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13308 2099 13311
rect 3326 13308 3332 13320
rect 2087 13280 3332 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 3528 13240 3556 13339
rect 3620 13308 3648 13416
rect 5626 13404 5632 13456
rect 5684 13404 5690 13456
rect 6270 13404 6276 13456
rect 6328 13444 6334 13456
rect 8772 13444 8800 13472
rect 6328 13416 6960 13444
rect 8772 13416 9260 13444
rect 6328 13404 6334 13416
rect 6472 13385 6500 13416
rect 6181 13379 6239 13385
rect 6181 13345 6193 13379
rect 6227 13345 6239 13379
rect 6181 13339 6239 13345
rect 6457 13379 6515 13385
rect 6457 13345 6469 13379
rect 6503 13345 6515 13379
rect 6457 13339 6515 13345
rect 3976 13311 4034 13317
rect 3976 13308 3988 13311
rect 3620 13280 3988 13308
rect 3976 13277 3988 13280
rect 4022 13277 4034 13311
rect 3976 13271 4034 13277
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13308 4307 13311
rect 5074 13308 5080 13320
rect 4295 13280 5080 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 5074 13268 5080 13280
rect 5132 13268 5138 13320
rect 5350 13268 5356 13320
rect 5408 13308 5414 13320
rect 6196 13308 6224 13339
rect 6822 13336 6828 13388
rect 6880 13336 6886 13388
rect 6932 13376 6960 13416
rect 9232 13385 9260 13416
rect 9306 13404 9312 13456
rect 9364 13404 9370 13456
rect 9416 13444 9444 13472
rect 10244 13444 10272 13484
rect 9416 13416 10272 13444
rect 9217 13379 9275 13385
rect 6932 13348 9168 13376
rect 6638 13308 6644 13320
rect 5408 13280 6040 13308
rect 6196 13280 6644 13308
rect 5408 13268 5414 13280
rect 6012 13249 6040 13280
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 3344 13212 3556 13240
rect 5997 13243 6055 13249
rect 3344 13184 3372 13212
rect 5997 13209 6009 13243
rect 6043 13209 6055 13243
rect 5997 13203 6055 13209
rect 6362 13200 6368 13252
rect 6420 13240 6426 13252
rect 6840 13240 6868 13336
rect 7190 13317 7196 13320
rect 7152 13311 7196 13317
rect 7152 13277 7164 13311
rect 7152 13271 7196 13277
rect 7190 13268 7196 13271
rect 7248 13268 7254 13320
rect 7282 13268 7288 13320
rect 7340 13268 7346 13320
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13308 7619 13311
rect 7607 13280 9076 13308
rect 7607 13277 7619 13280
rect 7561 13271 7619 13277
rect 9048 13249 9076 13280
rect 9033 13243 9091 13249
rect 6420 13212 6868 13240
rect 8772 13212 8984 13240
rect 6420 13200 6426 13212
rect 1026 13132 1032 13184
rect 1084 13132 1090 13184
rect 3326 13132 3332 13184
rect 3384 13172 3390 13184
rect 3878 13172 3884 13184
rect 3384 13144 3884 13172
rect 3384 13132 3390 13144
rect 3878 13132 3884 13144
rect 3936 13132 3942 13184
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 5902 13172 5908 13184
rect 4304 13144 5908 13172
rect 4304 13132 4310 13144
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 6270 13132 6276 13184
rect 6328 13132 6334 13184
rect 7466 13132 7472 13184
rect 7524 13172 7530 13184
rect 8772 13172 8800 13212
rect 7524 13144 8800 13172
rect 7524 13132 7530 13144
rect 8846 13132 8852 13184
rect 8904 13132 8910 13184
rect 8956 13172 8984 13212
rect 9033 13209 9045 13243
rect 9079 13209 9091 13243
rect 9140 13240 9168 13348
rect 9217 13345 9229 13379
rect 9263 13345 9275 13379
rect 9416 13376 9444 13416
rect 9585 13379 9643 13385
rect 9585 13376 9597 13379
rect 9416 13348 9597 13376
rect 9217 13339 9275 13345
rect 9585 13345 9597 13348
rect 9631 13345 9643 13379
rect 9585 13339 9643 13345
rect 9858 13336 9864 13388
rect 9916 13336 9922 13388
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13345 10195 13379
rect 10137 13339 10195 13345
rect 10413 13379 10471 13385
rect 10413 13345 10425 13379
rect 10459 13376 10471 13379
rect 10520 13376 10548 13484
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 10962 13472 10968 13524
rect 11020 13472 11026 13524
rect 11425 13515 11483 13521
rect 11425 13481 11437 13515
rect 11471 13512 11483 13515
rect 11606 13512 11612 13524
rect 11471 13484 11612 13512
rect 11471 13481 11483 13484
rect 11425 13475 11483 13481
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 11698 13472 11704 13524
rect 11756 13512 11762 13524
rect 12710 13512 12716 13524
rect 11756 13484 12716 13512
rect 11756 13472 11762 13484
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 12903 13515 12961 13521
rect 12903 13481 12915 13515
rect 12949 13512 12961 13515
rect 13262 13512 13268 13524
rect 12949 13484 13268 13512
rect 12949 13481 12961 13484
rect 12903 13475 12961 13481
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 14274 13472 14280 13524
rect 14332 13512 14338 13524
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 14332 13484 16313 13512
rect 14332 13472 14338 13484
rect 16301 13481 16313 13484
rect 16347 13512 16359 13515
rect 16390 13512 16396 13524
rect 16347 13484 16396 13512
rect 16347 13481 16359 13484
rect 16301 13475 16359 13481
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 16669 13515 16727 13521
rect 16669 13512 16681 13515
rect 16632 13484 16681 13512
rect 16632 13472 16638 13484
rect 16669 13481 16681 13484
rect 16715 13481 16727 13515
rect 16669 13475 16727 13481
rect 17126 13472 17132 13524
rect 17184 13512 17190 13524
rect 17503 13515 17561 13521
rect 17503 13512 17515 13515
rect 17184 13484 17515 13512
rect 17184 13472 17190 13484
rect 17503 13481 17515 13484
rect 17549 13481 17561 13515
rect 17503 13475 17561 13481
rect 17678 13472 17684 13524
rect 17736 13512 17742 13524
rect 18877 13515 18935 13521
rect 18877 13512 18889 13515
rect 17736 13484 18889 13512
rect 17736 13472 17742 13484
rect 18877 13481 18889 13484
rect 18923 13481 18935 13515
rect 18877 13475 18935 13481
rect 21637 13515 21695 13521
rect 21637 13481 21649 13515
rect 21683 13481 21695 13515
rect 21637 13475 21695 13481
rect 22379 13515 22437 13521
rect 22379 13481 22391 13515
rect 22425 13512 22437 13515
rect 24587 13515 24645 13521
rect 24587 13512 24599 13515
rect 22425 13484 24599 13512
rect 22425 13481 22437 13484
rect 22379 13475 22437 13481
rect 10980 13444 11008 13472
rect 10980 13416 11284 13444
rect 10965 13379 11023 13385
rect 10965 13376 10977 13379
rect 10459 13348 10548 13376
rect 10612 13348 10977 13376
rect 10459 13345 10471 13348
rect 10413 13339 10471 13345
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 10152 13308 10180 13339
rect 10612 13308 10640 13348
rect 10965 13345 10977 13348
rect 11011 13376 11023 13379
rect 11146 13376 11152 13388
rect 11011 13348 11152 13376
rect 11011 13345 11023 13348
rect 10965 13339 11023 13345
rect 11146 13336 11152 13348
rect 11204 13336 11210 13388
rect 11256 13385 11284 13416
rect 11514 13404 11520 13456
rect 11572 13444 11578 13456
rect 11572 13416 11652 13444
rect 11572 13404 11578 13416
rect 11624 13400 11652 13416
rect 11882 13404 11888 13456
rect 11940 13444 11946 13456
rect 12526 13444 12532 13456
rect 11940 13416 12532 13444
rect 11940 13404 11946 13416
rect 11624 13385 11750 13400
rect 11241 13379 11299 13385
rect 11241 13345 11253 13379
rect 11287 13345 11299 13379
rect 11624 13379 11759 13385
rect 11624 13372 11713 13379
rect 11241 13339 11299 13345
rect 11701 13345 11713 13372
rect 11747 13345 11759 13379
rect 11701 13339 11759 13345
rect 11974 13336 11980 13388
rect 12032 13336 12038 13388
rect 12268 13385 12296 13416
rect 12526 13404 12532 13416
rect 12584 13404 12590 13456
rect 13906 13404 13912 13456
rect 13964 13444 13970 13456
rect 13964 13416 17172 13444
rect 13964 13404 13970 13416
rect 14844 13385 14872 13416
rect 12253 13379 12311 13385
rect 12253 13345 12265 13379
rect 12299 13345 12311 13379
rect 14829 13379 14887 13385
rect 12253 13339 12311 13345
rect 12360 13348 12943 13376
rect 9824 13280 10640 13308
rect 9824 13268 9830 13280
rect 10778 13268 10784 13320
rect 10836 13308 10842 13320
rect 12360 13308 12388 13348
rect 10836 13280 12388 13308
rect 10836 13268 10842 13280
rect 12434 13268 12440 13320
rect 12492 13268 12498 13320
rect 12915 13317 12943 13348
rect 14829 13345 14841 13379
rect 14875 13345 14887 13379
rect 14829 13339 14887 13345
rect 15381 13379 15439 13385
rect 15381 13345 15393 13379
rect 15427 13376 15439 13379
rect 15470 13376 15476 13388
rect 15427 13348 15476 13376
rect 15427 13345 15439 13348
rect 15381 13339 15439 13345
rect 15470 13336 15476 13348
rect 15528 13376 15534 13388
rect 15746 13376 15752 13388
rect 15528 13348 15752 13376
rect 15528 13336 15534 13348
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 15933 13379 15991 13385
rect 15933 13345 15945 13379
rect 15979 13376 15991 13379
rect 16022 13376 16028 13388
rect 15979 13348 16028 13376
rect 15979 13345 15991 13348
rect 15933 13339 15991 13345
rect 12900 13311 12958 13317
rect 12900 13277 12912 13311
rect 12946 13277 12958 13311
rect 12900 13271 12958 13277
rect 12986 13268 12992 13320
rect 13044 13308 13050 13320
rect 13173 13311 13231 13317
rect 13173 13308 13185 13311
rect 13044 13280 13185 13308
rect 13044 13268 13050 13280
rect 13173 13277 13185 13280
rect 13219 13277 13231 13311
rect 13173 13271 13231 13277
rect 13262 13268 13268 13320
rect 13320 13308 13326 13320
rect 13906 13308 13912 13320
rect 13320 13280 13912 13308
rect 13320 13268 13326 13280
rect 13906 13268 13912 13280
rect 13964 13268 13970 13320
rect 14918 13268 14924 13320
rect 14976 13308 14982 13320
rect 15013 13311 15071 13317
rect 15013 13308 15025 13311
rect 14976 13280 15025 13308
rect 14976 13268 14982 13280
rect 15013 13277 15025 13280
rect 15059 13277 15071 13311
rect 15013 13271 15071 13277
rect 9140 13212 10272 13240
rect 9033 13203 9091 13209
rect 10244 13184 10272 13212
rect 10410 13200 10416 13252
rect 10468 13240 10474 13252
rect 10597 13243 10655 13249
rect 10597 13240 10609 13243
rect 10468 13212 10609 13240
rect 10468 13200 10474 13212
rect 10597 13209 10609 13212
rect 10643 13209 10655 13243
rect 10597 13203 10655 13209
rect 10686 13200 10692 13252
rect 10744 13200 10750 13252
rect 11054 13200 11060 13252
rect 11112 13240 11118 13252
rect 11112 13212 11284 13240
rect 11112 13200 11118 13212
rect 9306 13172 9312 13184
rect 8956 13144 9312 13172
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 9490 13132 9496 13184
rect 9548 13172 9554 13184
rect 10045 13175 10103 13181
rect 10045 13172 10057 13175
rect 9548 13144 10057 13172
rect 9548 13132 9554 13144
rect 10045 13141 10057 13144
rect 10091 13141 10103 13175
rect 10045 13135 10103 13141
rect 10226 13132 10232 13184
rect 10284 13132 10290 13184
rect 10321 13175 10379 13181
rect 10321 13141 10333 13175
rect 10367 13172 10379 13175
rect 10502 13172 10508 13184
rect 10367 13144 10508 13172
rect 10367 13141 10379 13144
rect 10321 13135 10379 13141
rect 10502 13132 10508 13144
rect 10560 13132 10566 13184
rect 10704 13172 10732 13200
rect 11149 13175 11207 13181
rect 11149 13172 11161 13175
rect 10704 13144 11161 13172
rect 11149 13141 11161 13144
rect 11195 13141 11207 13175
rect 11256 13172 11284 13212
rect 11514 13200 11520 13252
rect 11572 13200 11578 13252
rect 12069 13243 12127 13249
rect 12069 13240 12081 13243
rect 11624 13212 12081 13240
rect 11624 13172 11652 13212
rect 12069 13209 12081 13212
rect 12115 13209 12127 13243
rect 15565 13243 15623 13249
rect 15565 13240 15577 13243
rect 12069 13203 12127 13209
rect 14200 13212 15577 13240
rect 11256 13144 11652 13172
rect 11793 13175 11851 13181
rect 11149 13135 11207 13141
rect 11793 13141 11805 13175
rect 11839 13172 11851 13175
rect 11882 13172 11888 13184
rect 11839 13144 11888 13172
rect 11839 13141 11851 13144
rect 11793 13135 11851 13141
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 12250 13132 12256 13184
rect 12308 13172 12314 13184
rect 14200 13172 14228 13212
rect 15565 13209 15577 13212
rect 15611 13240 15623 13243
rect 15948 13240 15976 13339
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16114 13336 16120 13388
rect 16172 13336 16178 13388
rect 16482 13336 16488 13388
rect 16540 13336 16546 13388
rect 17034 13336 17040 13388
rect 17092 13336 17098 13388
rect 17144 13376 17172 13416
rect 18506 13404 18512 13456
rect 18564 13444 18570 13456
rect 21652 13444 21680 13475
rect 24228 13456 24256 13484
rect 24587 13481 24599 13484
rect 24633 13481 24645 13515
rect 24587 13475 24645 13481
rect 25314 13472 25320 13524
rect 25372 13512 25378 13524
rect 26326 13512 26332 13524
rect 25372 13484 26332 13512
rect 25372 13472 25378 13484
rect 26326 13472 26332 13484
rect 26384 13472 26390 13524
rect 26418 13472 26424 13524
rect 26476 13472 26482 13524
rect 26878 13472 26884 13524
rect 26936 13521 26942 13524
rect 26936 13512 26945 13521
rect 26936 13484 26981 13512
rect 26936 13475 26945 13484
rect 26936 13472 26942 13475
rect 27062 13472 27068 13524
rect 27120 13512 27126 13524
rect 27120 13484 27844 13512
rect 27120 13472 27126 13484
rect 18564 13416 18828 13444
rect 18564 13404 18570 13416
rect 17402 13376 17408 13388
rect 17144 13348 17408 13376
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 17773 13379 17831 13385
rect 17773 13345 17785 13379
rect 17819 13376 17831 13379
rect 18690 13376 18696 13388
rect 17819 13348 18696 13376
rect 17819 13345 17831 13348
rect 17773 13339 17831 13345
rect 18690 13336 18696 13348
rect 18748 13336 18754 13388
rect 18800 13376 18828 13416
rect 20364 13416 21588 13444
rect 21652 13416 21956 13444
rect 19797 13379 19855 13385
rect 19797 13376 19809 13379
rect 18800 13348 19809 13376
rect 19797 13345 19809 13348
rect 19843 13376 19855 13379
rect 19978 13376 19984 13388
rect 19843 13348 19984 13376
rect 19843 13345 19855 13348
rect 19797 13339 19855 13345
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 20254 13336 20260 13388
rect 20312 13376 20318 13388
rect 20364 13385 20392 13416
rect 20349 13379 20407 13385
rect 20349 13376 20361 13379
rect 20312 13348 20361 13376
rect 20312 13336 20318 13348
rect 20349 13345 20361 13348
rect 20395 13345 20407 13379
rect 20349 13339 20407 13345
rect 20530 13336 20536 13388
rect 20588 13376 20594 13388
rect 20625 13379 20683 13385
rect 20625 13376 20637 13379
rect 20588 13348 20637 13376
rect 20588 13336 20594 13348
rect 20625 13345 20637 13348
rect 20671 13376 20683 13379
rect 21560 13376 21588 13416
rect 21726 13376 21732 13388
rect 20671 13348 21496 13376
rect 21560 13348 21732 13376
rect 20671 13345 20683 13348
rect 20625 13339 20683 13345
rect 17533 13329 17591 13335
rect 17533 13326 17545 13329
rect 17512 13295 17545 13326
rect 17579 13308 17591 13329
rect 21266 13308 21272 13320
rect 17579 13295 21272 13308
rect 17512 13280 21272 13295
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 21468 13308 21496 13348
rect 21726 13336 21732 13348
rect 21784 13376 21790 13388
rect 21821 13379 21879 13385
rect 21821 13376 21833 13379
rect 21784 13348 21833 13376
rect 21784 13336 21790 13348
rect 21821 13345 21833 13348
rect 21867 13345 21879 13379
rect 21928 13376 21956 13416
rect 24026 13404 24032 13456
rect 24084 13404 24090 13456
rect 24210 13404 24216 13456
rect 24268 13404 24274 13456
rect 26436 13444 26464 13472
rect 25608 13416 26464 13444
rect 22649 13379 22707 13385
rect 22649 13376 22661 13379
rect 21928 13348 22661 13376
rect 21821 13339 21879 13345
rect 22649 13345 22661 13348
rect 22695 13345 22707 13379
rect 22649 13339 22707 13345
rect 23566 13336 23572 13388
rect 23624 13376 23630 13388
rect 24857 13379 24915 13385
rect 24857 13376 24869 13379
rect 23624 13348 24869 13376
rect 23624 13336 23630 13348
rect 24857 13345 24869 13348
rect 24903 13345 24915 13379
rect 24857 13339 24915 13345
rect 21634 13308 21640 13320
rect 21468 13280 21640 13308
rect 21634 13268 21640 13280
rect 21692 13268 21698 13320
rect 21913 13311 21971 13317
rect 21913 13277 21925 13311
rect 21959 13308 21971 13311
rect 22186 13308 22192 13320
rect 21959 13280 22192 13308
rect 21959 13277 21971 13280
rect 21913 13271 21971 13277
rect 22186 13268 22192 13280
rect 22244 13268 22250 13320
rect 22278 13268 22284 13320
rect 22336 13310 22342 13320
rect 22376 13311 22434 13317
rect 22376 13310 22388 13311
rect 22336 13282 22388 13310
rect 22336 13268 22342 13282
rect 22376 13277 22388 13282
rect 22422 13277 22434 13311
rect 22376 13271 22434 13277
rect 24118 13268 24124 13320
rect 24176 13308 24182 13320
rect 24394 13308 24400 13320
rect 24176 13280 24400 13308
rect 24176 13268 24182 13280
rect 24394 13268 24400 13280
rect 24452 13268 24458 13320
rect 24486 13268 24492 13320
rect 24544 13310 24550 13320
rect 24584 13313 24642 13319
rect 24584 13310 24596 13313
rect 24544 13282 24596 13310
rect 24544 13268 24550 13282
rect 24584 13279 24596 13282
rect 24630 13279 24642 13313
rect 24584 13273 24642 13279
rect 24670 13268 24676 13320
rect 24728 13308 24734 13320
rect 25608 13308 25636 13416
rect 26436 13385 26464 13416
rect 26421 13379 26479 13385
rect 26421 13345 26433 13379
rect 26467 13345 26479 13379
rect 26421 13339 26479 13345
rect 26510 13336 26516 13388
rect 26568 13376 26574 13388
rect 27157 13379 27215 13385
rect 27157 13376 27169 13379
rect 26568 13348 27169 13376
rect 26568 13336 26574 13348
rect 27157 13345 27169 13348
rect 27203 13345 27215 13379
rect 27157 13339 27215 13345
rect 27614 13336 27620 13388
rect 27672 13336 27678 13388
rect 27816 13376 27844 13484
rect 28258 13472 28264 13524
rect 28316 13472 28322 13524
rect 28166 13404 28172 13456
rect 28224 13444 28230 13456
rect 28626 13444 28632 13456
rect 28224 13416 28632 13444
rect 28224 13404 28230 13416
rect 28626 13404 28632 13416
rect 28684 13404 28690 13456
rect 28905 13379 28963 13385
rect 28905 13376 28917 13379
rect 27816 13348 28917 13376
rect 28905 13345 28917 13348
rect 28951 13345 28963 13379
rect 28905 13339 28963 13345
rect 26884 13311 26942 13317
rect 26884 13308 26896 13311
rect 24728 13280 25636 13308
rect 26444 13280 26896 13308
rect 24728 13268 24734 13280
rect 15611 13212 15976 13240
rect 15611 13209 15623 13212
rect 15565 13203 15623 13209
rect 16390 13200 16396 13252
rect 16448 13240 16454 13252
rect 19521 13243 19579 13249
rect 16448 13212 16804 13240
rect 16448 13200 16454 13212
rect 12308 13144 14228 13172
rect 12308 13132 12314 13144
rect 14274 13132 14280 13184
rect 14332 13132 14338 13184
rect 15746 13132 15752 13184
rect 15804 13132 15810 13184
rect 15838 13132 15844 13184
rect 15896 13172 15902 13184
rect 16666 13172 16672 13184
rect 15896 13144 16672 13172
rect 15896 13132 15902 13144
rect 16666 13132 16672 13144
rect 16724 13132 16730 13184
rect 16776 13172 16804 13212
rect 19521 13209 19533 13243
rect 19567 13240 19579 13243
rect 20070 13240 20076 13252
rect 19567 13212 20076 13240
rect 19567 13209 19579 13212
rect 19521 13203 19579 13209
rect 20070 13200 20076 13212
rect 20128 13200 20134 13252
rect 20165 13243 20223 13249
rect 20165 13209 20177 13243
rect 20211 13240 20223 13243
rect 26145 13243 26203 13249
rect 20211 13212 21956 13240
rect 20211 13209 20223 13212
rect 20165 13203 20223 13209
rect 21928 13184 21956 13212
rect 26145 13209 26157 13243
rect 26191 13240 26203 13243
rect 26444 13240 26472 13280
rect 26884 13277 26896 13280
rect 26930 13277 26942 13311
rect 27632 13308 27660 13336
rect 28629 13311 28687 13317
rect 28629 13308 28641 13311
rect 27632 13280 28641 13308
rect 26884 13271 26942 13277
rect 28629 13277 28641 13280
rect 28675 13277 28687 13311
rect 28629 13271 28687 13277
rect 26191 13212 26472 13240
rect 26191 13209 26203 13212
rect 26145 13203 26203 13209
rect 19334 13172 19340 13184
rect 16776 13144 19340 13172
rect 19334 13132 19340 13144
rect 19392 13132 19398 13184
rect 19978 13132 19984 13184
rect 20036 13172 20042 13184
rect 20346 13172 20352 13184
rect 20036 13144 20352 13172
rect 20036 13132 20042 13144
rect 20346 13132 20352 13144
rect 20404 13132 20410 13184
rect 20441 13175 20499 13181
rect 20441 13141 20453 13175
rect 20487 13172 20499 13175
rect 21818 13172 21824 13184
rect 20487 13144 21824 13172
rect 20487 13141 20499 13144
rect 20441 13135 20499 13141
rect 21818 13132 21824 13144
rect 21876 13132 21882 13184
rect 21910 13132 21916 13184
rect 21968 13132 21974 13184
rect 23750 13132 23756 13184
rect 23808 13172 23814 13184
rect 27522 13172 27528 13184
rect 23808 13144 27528 13172
rect 23808 13132 23814 13144
rect 27522 13132 27528 13144
rect 27580 13132 27586 13184
rect 28810 13132 28816 13184
rect 28868 13172 28874 13184
rect 30009 13175 30067 13181
rect 30009 13172 30021 13175
rect 28868 13144 30021 13172
rect 28868 13132 28874 13144
rect 30009 13141 30021 13144
rect 30055 13141 30067 13175
rect 30009 13135 30067 13141
rect 552 13082 30912 13104
rect 552 13030 4193 13082
rect 4245 13030 4257 13082
rect 4309 13030 4321 13082
rect 4373 13030 4385 13082
rect 4437 13030 4449 13082
rect 4501 13030 11783 13082
rect 11835 13030 11847 13082
rect 11899 13030 11911 13082
rect 11963 13030 11975 13082
rect 12027 13030 12039 13082
rect 12091 13030 19373 13082
rect 19425 13030 19437 13082
rect 19489 13030 19501 13082
rect 19553 13030 19565 13082
rect 19617 13030 19629 13082
rect 19681 13030 26963 13082
rect 27015 13030 27027 13082
rect 27079 13030 27091 13082
rect 27143 13030 27155 13082
rect 27207 13030 27219 13082
rect 27271 13030 30912 13082
rect 552 13008 30912 13030
rect 1670 12928 1676 12980
rect 1728 12968 1734 12980
rect 3142 12968 3148 12980
rect 1728 12940 3148 12968
rect 1728 12928 1734 12940
rect 3142 12928 3148 12940
rect 3200 12928 3206 12980
rect 3510 12928 3516 12980
rect 3568 12968 3574 12980
rect 3878 12968 3884 12980
rect 3568 12940 3884 12968
rect 3568 12928 3574 12940
rect 3878 12928 3884 12940
rect 3936 12928 3942 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 7282 12968 7288 12980
rect 5951 12940 7288 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 7282 12928 7288 12940
rect 7340 12928 7346 12980
rect 7650 12928 7656 12980
rect 7708 12968 7714 12980
rect 9306 12968 9312 12980
rect 7708 12940 9312 12968
rect 7708 12928 7714 12940
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 10100 12940 12173 12968
rect 10100 12928 10106 12940
rect 12161 12937 12173 12940
rect 12207 12937 12219 12971
rect 12161 12931 12219 12937
rect 12342 12928 12348 12980
rect 12400 12968 12406 12980
rect 12710 12968 12716 12980
rect 12400 12940 12716 12968
rect 12400 12928 12406 12940
rect 9033 12903 9091 12909
rect 9033 12900 9045 12903
rect 3344 12872 3883 12900
rect 3344 12844 3372 12872
rect 937 12835 995 12841
rect 937 12801 949 12835
rect 983 12832 995 12835
rect 1302 12832 1308 12844
rect 983 12804 1308 12832
rect 983 12801 995 12804
rect 937 12795 995 12801
rect 1302 12792 1308 12804
rect 1360 12792 1366 12844
rect 1443 12835 1501 12841
rect 1443 12801 1455 12835
rect 1489 12832 1501 12835
rect 1489 12804 2774 12832
rect 1489 12801 1501 12804
rect 1443 12795 1501 12801
rect 1673 12767 1731 12773
rect 1673 12733 1685 12767
rect 1719 12764 1731 12767
rect 2130 12764 2136 12776
rect 1719 12736 2136 12764
rect 1719 12733 1731 12736
rect 1673 12727 1731 12733
rect 2130 12724 2136 12736
rect 2188 12724 2194 12776
rect 2746 12764 2774 12804
rect 3050 12792 3056 12844
rect 3108 12792 3114 12844
rect 3326 12792 3332 12844
rect 3384 12792 3390 12844
rect 3418 12792 3424 12844
rect 3476 12832 3482 12844
rect 3855 12841 3883 12872
rect 8864 12872 9045 12900
rect 3855 12835 3929 12841
rect 3476 12804 3746 12832
rect 3855 12804 3883 12835
rect 3476 12792 3482 12804
rect 3718 12780 3746 12804
rect 3871 12801 3883 12804
rect 3917 12801 3929 12835
rect 3871 12795 3929 12801
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4344 12835 4402 12841
rect 4344 12832 4356 12835
rect 4304 12804 4356 12832
rect 4304 12792 4310 12804
rect 4344 12801 4356 12804
rect 4390 12801 4402 12835
rect 4344 12795 4402 12801
rect 5350 12792 5356 12844
rect 5408 12832 5414 12844
rect 6552 12835 6610 12841
rect 6552 12832 6564 12835
rect 5408 12804 6564 12832
rect 5408 12792 5414 12804
rect 6552 12801 6564 12804
rect 6598 12801 6610 12835
rect 6552 12795 6610 12801
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 8864 12832 8892 12872
rect 9033 12869 9045 12872
rect 9079 12869 9091 12903
rect 9033 12863 9091 12869
rect 11238 12860 11244 12912
rect 11296 12900 11302 12912
rect 11885 12903 11943 12909
rect 11885 12900 11897 12903
rect 11296 12872 11897 12900
rect 11296 12860 11302 12872
rect 11885 12869 11897 12872
rect 11931 12869 11943 12903
rect 11885 12863 11943 12869
rect 12066 12860 12072 12912
rect 12124 12900 12130 12912
rect 12636 12900 12664 12940
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 12802 12928 12808 12980
rect 12860 12968 12866 12980
rect 12986 12968 12992 12980
rect 12860 12940 12992 12968
rect 12860 12928 12866 12940
rect 12986 12928 12992 12940
rect 13044 12928 13050 12980
rect 13170 12928 13176 12980
rect 13228 12968 13234 12980
rect 13630 12968 13636 12980
rect 13228 12940 13636 12968
rect 13228 12928 13234 12940
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 14090 12928 14096 12980
rect 14148 12968 14154 12980
rect 14148 12940 16712 12968
rect 14148 12928 14154 12940
rect 12897 12903 12955 12909
rect 12124 12872 12572 12900
rect 12636 12872 12848 12900
rect 12124 12860 12130 12872
rect 6871 12804 8892 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 10042 12792 10048 12844
rect 10100 12832 10106 12844
rect 10140 12835 10198 12841
rect 10140 12832 10152 12835
rect 10100 12804 10152 12832
rect 10100 12792 10106 12804
rect 10140 12801 10152 12804
rect 10186 12801 10198 12835
rect 10140 12795 10198 12801
rect 10410 12792 10416 12844
rect 10468 12792 10474 12844
rect 10502 12792 10508 12844
rect 10560 12832 10566 12844
rect 12250 12832 12256 12844
rect 10560 12804 12256 12832
rect 10560 12792 10566 12804
rect 12250 12792 12256 12804
rect 12308 12792 12314 12844
rect 12544 12780 12572 12872
rect 12820 12832 12848 12872
rect 12897 12869 12909 12903
rect 12943 12900 12955 12903
rect 14366 12900 14372 12912
rect 12943 12872 14372 12900
rect 12943 12869 12955 12872
rect 12897 12863 12955 12869
rect 14366 12860 14372 12872
rect 14424 12860 14430 12912
rect 16684 12900 16712 12940
rect 16758 12928 16764 12980
rect 16816 12928 16822 12980
rect 16850 12928 16856 12980
rect 16908 12968 16914 12980
rect 20073 12971 20131 12977
rect 16908 12940 19196 12968
rect 16908 12928 16914 12940
rect 16684 12872 18920 12900
rect 12820 12804 13400 12832
rect 3510 12764 3516 12776
rect 2746 12736 3516 12764
rect 3510 12724 3516 12736
rect 3568 12724 3574 12776
rect 3718 12773 3832 12780
rect 3718 12767 3847 12773
rect 3718 12752 3801 12767
rect 3789 12733 3801 12752
rect 3835 12733 3847 12767
rect 3789 12727 3847 12733
rect 4614 12724 4620 12776
rect 4672 12724 4678 12776
rect 5626 12724 5632 12776
rect 5684 12764 5690 12776
rect 6089 12767 6147 12773
rect 6089 12764 6101 12767
rect 5684 12736 6101 12764
rect 5684 12724 5690 12736
rect 6089 12733 6101 12736
rect 6135 12764 6147 12767
rect 6178 12764 6184 12776
rect 6135 12736 6184 12764
rect 6135 12733 6147 12736
rect 6089 12727 6147 12733
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 6416 12767 6474 12773
rect 6416 12733 6428 12767
rect 6462 12764 6474 12767
rect 7190 12764 7196 12776
rect 6462 12736 7196 12764
rect 6462 12733 6474 12736
rect 6416 12727 6474 12733
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 8754 12764 8760 12776
rect 8220 12736 8760 12764
rect 8220 12705 8248 12736
rect 8754 12724 8760 12736
rect 8812 12724 8818 12776
rect 9122 12724 9128 12776
rect 9180 12764 9186 12776
rect 9217 12767 9275 12773
rect 9217 12764 9229 12767
rect 9180 12736 9229 12764
rect 9180 12724 9186 12736
rect 9217 12733 9229 12736
rect 9263 12733 9275 12767
rect 9217 12727 9275 12733
rect 8205 12699 8263 12705
rect 2746 12668 3648 12696
rect 1403 12631 1461 12637
rect 1403 12597 1415 12631
rect 1449 12628 1461 12631
rect 1670 12628 1676 12640
rect 1449 12600 1676 12628
rect 1449 12597 1461 12600
rect 1403 12591 1461 12597
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 2590 12588 2596 12640
rect 2648 12628 2654 12640
rect 2746 12628 2774 12668
rect 3620 12637 3648 12668
rect 8205 12665 8217 12699
rect 8251 12665 8263 12699
rect 8205 12659 8263 12665
rect 8478 12656 8484 12708
rect 8536 12656 8542 12708
rect 9232 12696 9260 12727
rect 9306 12724 9312 12776
rect 9364 12724 9370 12776
rect 9674 12724 9680 12776
rect 9732 12724 9738 12776
rect 11606 12764 11612 12776
rect 9784 12736 11612 12764
rect 9784 12696 9812 12736
rect 11606 12724 11612 12736
rect 11664 12724 11670 12776
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 12069 12767 12127 12773
rect 12069 12764 12081 12767
rect 12032 12736 12081 12764
rect 12032 12724 12038 12736
rect 12069 12733 12081 12736
rect 12115 12733 12127 12767
rect 12069 12727 12127 12733
rect 12342 12724 12348 12776
rect 12400 12773 12406 12776
rect 12400 12764 12411 12773
rect 12400 12736 12445 12764
rect 12544 12752 12664 12780
rect 12400 12727 12411 12736
rect 12400 12724 12406 12727
rect 9232 12668 9812 12696
rect 11146 12656 11152 12708
rect 11204 12696 11210 12708
rect 11992 12696 12020 12724
rect 11204 12668 12020 12696
rect 12636 12696 12664 12752
rect 12805 12767 12863 12773
rect 12805 12733 12817 12767
rect 12851 12760 12863 12767
rect 13081 12767 13139 12773
rect 12851 12733 12940 12760
rect 12805 12732 12940 12733
rect 12805 12727 12863 12732
rect 12912 12696 12940 12732
rect 13081 12733 13093 12767
rect 13127 12764 13139 12767
rect 13170 12764 13176 12776
rect 13127 12736 13176 12764
rect 13127 12733 13139 12736
rect 13081 12727 13139 12733
rect 13170 12724 13176 12736
rect 13228 12724 13234 12776
rect 13372 12773 13400 12804
rect 13630 12792 13636 12844
rect 13688 12832 13694 12844
rect 13725 12835 13783 12841
rect 13725 12832 13737 12835
rect 13688 12804 13737 12832
rect 13688 12792 13694 12804
rect 13725 12801 13737 12804
rect 13771 12832 13783 12835
rect 13906 12832 13912 12844
rect 13771 12804 13912 12832
rect 13771 12801 13783 12804
rect 13725 12795 13783 12801
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 14550 12792 14556 12844
rect 14608 12792 14614 12844
rect 14918 12841 14924 12844
rect 14880 12835 14924 12841
rect 14880 12801 14892 12835
rect 14880 12795 14924 12801
rect 14918 12792 14924 12795
rect 14976 12792 14982 12844
rect 15059 12835 15117 12841
rect 15059 12801 15071 12835
rect 15105 12832 15117 12835
rect 15289 12835 15347 12841
rect 15105 12804 15240 12832
rect 15105 12801 15117 12804
rect 15059 12795 15117 12801
rect 13357 12767 13415 12773
rect 13357 12733 13369 12767
rect 13403 12733 13415 12767
rect 13357 12727 13415 12733
rect 13541 12767 13599 12773
rect 13541 12733 13553 12767
rect 13587 12764 13599 12767
rect 13814 12764 13820 12776
rect 13587 12736 13820 12764
rect 13587 12733 13599 12736
rect 13541 12727 13599 12733
rect 13814 12724 13820 12736
rect 13872 12724 13878 12776
rect 15212 12764 15240 12804
rect 15289 12801 15301 12835
rect 15335 12832 15347 12835
rect 15746 12832 15752 12844
rect 15335 12804 15752 12832
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 18230 12832 18236 12844
rect 15856 12804 18236 12832
rect 15856 12764 15884 12804
rect 18230 12792 18236 12804
rect 18288 12792 18294 12844
rect 15212 12736 15884 12764
rect 16298 12724 16304 12776
rect 16356 12764 16362 12776
rect 18892 12773 18920 12872
rect 19168 12773 19196 12940
rect 20073 12937 20085 12971
rect 20119 12968 20131 12971
rect 20622 12968 20628 12980
rect 20119 12940 20628 12968
rect 20119 12937 20131 12940
rect 20073 12931 20131 12937
rect 20622 12928 20628 12940
rect 20680 12928 20686 12980
rect 23566 12928 23572 12980
rect 23624 12968 23630 12980
rect 24486 12968 24492 12980
rect 23624 12940 24492 12968
rect 23624 12928 23630 12940
rect 24486 12928 24492 12940
rect 24544 12928 24550 12980
rect 25682 12928 25688 12980
rect 25740 12928 25746 12980
rect 26602 12928 26608 12980
rect 26660 12968 26666 12980
rect 28721 12971 28779 12977
rect 26660 12940 28396 12968
rect 26660 12928 26666 12940
rect 22833 12903 22891 12909
rect 22833 12869 22845 12903
rect 22879 12900 22891 12903
rect 22922 12900 22928 12912
rect 22879 12872 22928 12900
rect 22879 12869 22891 12872
rect 22833 12863 22891 12869
rect 22922 12860 22928 12872
rect 22980 12860 22986 12912
rect 23201 12903 23259 12909
rect 23201 12869 23213 12903
rect 23247 12900 23259 12903
rect 23750 12900 23756 12912
rect 23247 12872 23756 12900
rect 23247 12869 23259 12872
rect 23201 12863 23259 12869
rect 23750 12860 23756 12872
rect 23808 12860 23814 12912
rect 19886 12792 19892 12844
rect 19944 12832 19950 12844
rect 20806 12832 20812 12844
rect 19944 12804 20392 12832
rect 20770 12804 20812 12832
rect 19944 12792 19950 12804
rect 20364 12776 20392 12804
rect 20806 12792 20812 12804
rect 20864 12792 20870 12844
rect 22002 12832 22008 12844
rect 21008 12804 22008 12832
rect 16945 12767 17003 12773
rect 16945 12764 16957 12767
rect 16356 12736 16957 12764
rect 16356 12724 16362 12736
rect 16945 12733 16957 12736
rect 16991 12733 17003 12767
rect 16945 12727 17003 12733
rect 18877 12767 18935 12773
rect 18877 12733 18889 12767
rect 18923 12733 18935 12767
rect 18877 12727 18935 12733
rect 19153 12767 19211 12773
rect 19153 12733 19165 12767
rect 19199 12764 19211 12767
rect 19794 12764 19800 12776
rect 19199 12736 19800 12764
rect 19199 12733 19211 12736
rect 19153 12727 19211 12733
rect 12636 12668 13308 12696
rect 11204 12656 11210 12668
rect 2648 12600 2774 12628
rect 3605 12631 3663 12637
rect 2648 12588 2654 12600
rect 3605 12597 3617 12631
rect 3651 12597 3663 12631
rect 3605 12591 3663 12597
rect 3970 12588 3976 12640
rect 4028 12628 4034 12640
rect 4347 12631 4405 12637
rect 4347 12628 4359 12631
rect 4028 12600 4359 12628
rect 4028 12588 4034 12600
rect 4347 12597 4359 12600
rect 4393 12597 4405 12631
rect 4347 12591 4405 12597
rect 4890 12588 4896 12640
rect 4948 12628 4954 12640
rect 7466 12628 7472 12640
rect 4948 12600 7472 12628
rect 4948 12588 4954 12600
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 8570 12588 8576 12640
rect 8628 12588 8634 12640
rect 9030 12588 9036 12640
rect 9088 12628 9094 12640
rect 9582 12628 9588 12640
rect 9088 12600 9588 12628
rect 9088 12588 9094 12600
rect 9582 12588 9588 12600
rect 9640 12628 9646 12640
rect 10143 12631 10201 12637
rect 10143 12628 10155 12631
rect 9640 12600 10155 12628
rect 9640 12588 9646 12600
rect 10143 12597 10155 12600
rect 10189 12597 10201 12631
rect 10143 12591 10201 12597
rect 11701 12631 11759 12637
rect 11701 12597 11713 12631
rect 11747 12628 11759 12631
rect 12250 12628 12256 12640
rect 11747 12600 12256 12628
rect 11747 12597 11759 12600
rect 11701 12591 11759 12597
rect 12250 12588 12256 12600
rect 12308 12588 12314 12640
rect 12342 12588 12348 12640
rect 12400 12628 12406 12640
rect 12621 12631 12679 12637
rect 12621 12628 12633 12631
rect 12400 12600 12633 12628
rect 12400 12588 12406 12600
rect 12621 12597 12633 12600
rect 12667 12597 12679 12631
rect 12621 12591 12679 12597
rect 13170 12588 13176 12640
rect 13228 12588 13234 12640
rect 13280 12628 13308 12668
rect 13998 12656 14004 12708
rect 14056 12696 14062 12708
rect 14185 12699 14243 12705
rect 14185 12696 14197 12699
rect 14056 12668 14197 12696
rect 14056 12656 14062 12668
rect 14185 12665 14197 12668
rect 14231 12665 14243 12699
rect 14185 12659 14243 12665
rect 17957 12699 18015 12705
rect 17957 12665 17969 12699
rect 18003 12696 18015 12699
rect 18046 12696 18052 12708
rect 18003 12668 18052 12696
rect 18003 12665 18015 12668
rect 17957 12659 18015 12665
rect 18046 12656 18052 12668
rect 18104 12656 18110 12708
rect 18322 12656 18328 12708
rect 18380 12656 18386 12708
rect 18892 12696 18920 12727
rect 19794 12724 19800 12736
rect 19852 12764 19858 12776
rect 19981 12767 20039 12773
rect 19981 12764 19993 12767
rect 19852 12736 19993 12764
rect 19852 12724 19858 12736
rect 19981 12733 19993 12736
rect 20027 12733 20039 12767
rect 19981 12727 20039 12733
rect 20254 12724 20260 12776
rect 20312 12724 20318 12776
rect 20346 12724 20352 12776
rect 20404 12724 20410 12776
rect 20676 12767 20734 12773
rect 20676 12733 20688 12767
rect 20722 12764 20734 12767
rect 20898 12764 20904 12776
rect 20722 12736 20904 12764
rect 20722 12733 20734 12736
rect 20676 12727 20734 12733
rect 20898 12724 20904 12736
rect 20956 12764 20962 12776
rect 21008 12764 21036 12804
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 22186 12792 22192 12844
rect 22244 12832 22250 12844
rect 23842 12832 23848 12844
rect 22244 12804 23848 12832
rect 22244 12792 22250 12804
rect 23842 12792 23848 12804
rect 23900 12832 23906 12844
rect 24118 12832 24124 12844
rect 23900 12804 24124 12832
rect 23900 12792 23906 12804
rect 24118 12792 24124 12804
rect 24176 12792 24182 12844
rect 24308 12817 24366 12823
rect 24308 12814 24320 12817
rect 24228 12786 24320 12814
rect 20956 12736 21036 12764
rect 20956 12724 20962 12736
rect 21082 12724 21088 12776
rect 21140 12724 21146 12776
rect 22830 12764 22836 12776
rect 22066 12736 22836 12764
rect 20272 12696 20300 12724
rect 18892 12668 20300 12696
rect 14277 12631 14335 12637
rect 14277 12628 14289 12631
rect 13280 12600 14289 12628
rect 14277 12597 14289 12600
rect 14323 12628 14335 12631
rect 14550 12628 14556 12640
rect 14323 12600 14556 12628
rect 14323 12597 14335 12600
rect 14277 12591 14335 12597
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 14826 12588 14832 12640
rect 14884 12628 14890 12640
rect 16393 12631 16451 12637
rect 16393 12628 16405 12631
rect 14884 12600 16405 12628
rect 14884 12588 14890 12600
rect 16393 12597 16405 12600
rect 16439 12597 16451 12631
rect 16393 12591 16451 12597
rect 16942 12588 16948 12640
rect 17000 12628 17006 12640
rect 17221 12631 17279 12637
rect 17221 12628 17233 12631
rect 17000 12600 17233 12628
rect 17000 12588 17006 12600
rect 17221 12597 17233 12600
rect 17267 12628 17279 12631
rect 17589 12631 17647 12637
rect 17589 12628 17601 12631
rect 17267 12600 17601 12628
rect 17267 12597 17279 12600
rect 17221 12591 17279 12597
rect 17589 12597 17601 12600
rect 17635 12597 17647 12631
rect 17589 12591 17647 12597
rect 18690 12588 18696 12640
rect 18748 12588 18754 12640
rect 18969 12631 19027 12637
rect 18969 12597 18981 12631
rect 19015 12628 19027 12631
rect 19702 12628 19708 12640
rect 19015 12600 19708 12628
rect 19015 12597 19027 12600
rect 18969 12591 19027 12597
rect 19702 12588 19708 12600
rect 19760 12588 19766 12640
rect 19797 12631 19855 12637
rect 19797 12597 19809 12631
rect 19843 12628 19855 12631
rect 21174 12628 21180 12640
rect 19843 12600 21180 12628
rect 19843 12597 19855 12600
rect 19797 12591 19855 12597
rect 21174 12588 21180 12600
rect 21232 12588 21238 12640
rect 21450 12588 21456 12640
rect 21508 12628 21514 12640
rect 22066 12628 22094 12736
rect 22830 12724 22836 12736
rect 22888 12764 22894 12776
rect 23017 12767 23075 12773
rect 23017 12764 23029 12767
rect 22888 12736 23029 12764
rect 22888 12724 22894 12736
rect 23017 12733 23029 12736
rect 23063 12733 23075 12767
rect 23017 12727 23075 12733
rect 23106 12724 23112 12776
rect 23164 12764 23170 12776
rect 23385 12767 23443 12773
rect 23385 12764 23397 12767
rect 23164 12736 23397 12764
rect 23164 12724 23170 12736
rect 23385 12733 23397 12736
rect 23431 12764 23443 12767
rect 23661 12767 23719 12773
rect 23661 12764 23673 12767
rect 23431 12736 23673 12764
rect 23431 12733 23443 12736
rect 23385 12727 23443 12733
rect 23661 12733 23673 12736
rect 23707 12764 23719 12767
rect 23750 12764 23756 12776
rect 23707 12736 23756 12764
rect 23707 12733 23719 12736
rect 23661 12727 23719 12733
rect 23750 12724 23756 12736
rect 23808 12724 23814 12776
rect 24228 12764 24256 12786
rect 24308 12783 24320 12786
rect 24354 12783 24366 12817
rect 24486 12792 24492 12844
rect 24544 12832 24550 12844
rect 26712 12841 26740 12940
rect 28368 12900 28396 12940
rect 28721 12937 28733 12971
rect 28767 12968 28779 12971
rect 28902 12968 28908 12980
rect 28767 12940 28908 12968
rect 28767 12937 28779 12940
rect 28721 12931 28779 12937
rect 28902 12928 28908 12940
rect 28960 12928 28966 12980
rect 29181 12971 29239 12977
rect 29181 12937 29193 12971
rect 29227 12937 29239 12971
rect 29181 12931 29239 12937
rect 29196 12900 29224 12931
rect 29822 12928 29828 12980
rect 29880 12928 29886 12980
rect 28368 12872 29224 12900
rect 24581 12835 24639 12841
rect 24581 12832 24593 12835
rect 24544 12804 24593 12832
rect 24544 12792 24550 12804
rect 24581 12801 24593 12804
rect 24627 12801 24639 12835
rect 24581 12795 24639 12801
rect 26697 12835 26755 12841
rect 26697 12801 26709 12835
rect 26743 12801 26755 12835
rect 27798 12832 27804 12844
rect 26697 12795 26755 12801
rect 27172 12817 27804 12832
rect 24308 12777 24366 12783
rect 23955 12736 24256 12764
rect 22465 12699 22523 12705
rect 22465 12665 22477 12699
rect 22511 12696 22523 12699
rect 23955 12696 23983 12736
rect 24394 12724 24400 12776
rect 24452 12764 24458 12776
rect 26145 12767 26203 12773
rect 26145 12764 26157 12767
rect 24452 12736 26157 12764
rect 24452 12724 24458 12736
rect 26145 12733 26157 12736
rect 26191 12764 26203 12767
rect 26418 12764 26424 12776
rect 26191 12736 26424 12764
rect 26191 12733 26203 12736
rect 26145 12727 26203 12733
rect 26418 12724 26424 12736
rect 26476 12764 26482 12776
rect 26712 12764 26740 12795
rect 27172 12786 27205 12817
rect 27193 12783 27205 12786
rect 27239 12804 27804 12817
rect 27239 12783 27251 12804
rect 27798 12792 27804 12804
rect 27856 12792 27862 12844
rect 29546 12792 29552 12844
rect 29604 12832 29610 12844
rect 29604 12804 29684 12832
rect 29604 12792 29610 12804
rect 27193 12777 27251 12783
rect 26476 12736 26740 12764
rect 27433 12767 27491 12773
rect 26476 12724 26482 12736
rect 27433 12733 27445 12767
rect 27479 12764 27491 12767
rect 29656 12764 29684 12804
rect 30006 12773 30012 12776
rect 29733 12767 29791 12773
rect 29733 12764 29745 12767
rect 27479 12736 29592 12764
rect 29656 12736 29745 12764
rect 27479 12733 27491 12736
rect 27433 12727 27491 12733
rect 22511 12668 23983 12696
rect 29089 12699 29147 12705
rect 22511 12665 22523 12668
rect 22465 12659 22523 12665
rect 29089 12665 29101 12699
rect 29135 12696 29147 12699
rect 29362 12696 29368 12708
rect 29135 12668 29368 12696
rect 29135 12665 29147 12668
rect 29089 12659 29147 12665
rect 29362 12656 29368 12668
rect 29420 12656 29426 12708
rect 21508 12600 22094 12628
rect 23477 12631 23535 12637
rect 21508 12588 21514 12600
rect 23477 12597 23489 12631
rect 23523 12628 23535 12631
rect 24118 12628 24124 12640
rect 23523 12600 24124 12628
rect 23523 12597 23535 12600
rect 23477 12591 23535 12597
rect 24118 12588 24124 12600
rect 24176 12588 24182 12640
rect 24210 12588 24216 12640
rect 24268 12628 24274 12640
rect 24311 12631 24369 12637
rect 24311 12628 24323 12631
rect 24268 12600 24323 12628
rect 24268 12588 24274 12600
rect 24311 12597 24323 12600
rect 24357 12628 24369 12631
rect 26142 12628 26148 12640
rect 24357 12600 26148 12628
rect 24357 12597 24369 12600
rect 24311 12591 24369 12597
rect 26142 12588 26148 12600
rect 26200 12588 26206 12640
rect 26421 12631 26479 12637
rect 26421 12597 26433 12631
rect 26467 12628 26479 12631
rect 26510 12628 26516 12640
rect 26467 12600 26516 12628
rect 26467 12597 26479 12600
rect 26421 12591 26479 12597
rect 26510 12588 26516 12600
rect 26568 12588 26574 12640
rect 27163 12631 27221 12637
rect 27163 12597 27175 12631
rect 27209 12628 27221 12631
rect 27430 12628 27436 12640
rect 27209 12600 27436 12628
rect 27209 12597 27221 12600
rect 27163 12591 27221 12597
rect 27430 12588 27436 12600
rect 27488 12588 27494 12640
rect 28074 12588 28080 12640
rect 28132 12628 28138 12640
rect 28626 12628 28632 12640
rect 28132 12600 28632 12628
rect 28132 12588 28138 12600
rect 28626 12588 28632 12600
rect 28684 12588 28690 12640
rect 29564 12637 29592 12736
rect 29733 12733 29745 12736
rect 29779 12733 29791 12767
rect 30001 12764 30012 12773
rect 29967 12736 30012 12764
rect 29733 12727 29791 12733
rect 30001 12727 30012 12736
rect 30006 12724 30012 12727
rect 30064 12724 30070 12776
rect 29549 12631 29607 12637
rect 29549 12597 29561 12631
rect 29595 12597 29607 12631
rect 29549 12591 29607 12597
rect 552 12538 31072 12560
rect 552 12486 7988 12538
rect 8040 12486 8052 12538
rect 8104 12486 8116 12538
rect 8168 12486 8180 12538
rect 8232 12486 8244 12538
rect 8296 12486 15578 12538
rect 15630 12486 15642 12538
rect 15694 12486 15706 12538
rect 15758 12486 15770 12538
rect 15822 12486 15834 12538
rect 15886 12486 23168 12538
rect 23220 12486 23232 12538
rect 23284 12486 23296 12538
rect 23348 12486 23360 12538
rect 23412 12486 23424 12538
rect 23476 12486 30758 12538
rect 30810 12486 30822 12538
rect 30874 12486 30886 12538
rect 30938 12486 30950 12538
rect 31002 12486 31014 12538
rect 31066 12486 31072 12538
rect 552 12464 31072 12486
rect 1026 12384 1032 12436
rect 1084 12424 1090 12436
rect 1946 12424 1952 12436
rect 1084 12396 1952 12424
rect 1084 12384 1090 12396
rect 1946 12384 1952 12396
rect 2004 12384 2010 12436
rect 3970 12384 3976 12436
rect 4028 12433 4034 12436
rect 4028 12424 4037 12433
rect 4028 12396 4073 12424
rect 4028 12387 4037 12396
rect 4028 12384 4034 12387
rect 5258 12384 5264 12436
rect 5316 12384 5322 12436
rect 5537 12427 5595 12433
rect 5537 12393 5549 12427
rect 5583 12424 5595 12427
rect 5718 12424 5724 12436
rect 5583 12396 5724 12424
rect 5583 12393 5595 12396
rect 5537 12387 5595 12393
rect 5718 12384 5724 12396
rect 5776 12384 5782 12436
rect 6086 12384 6092 12436
rect 6144 12424 6150 12436
rect 6144 12396 6595 12424
rect 6144 12384 6150 12396
rect 5276 12356 5304 12384
rect 5276 12328 6316 12356
rect 1213 12291 1271 12297
rect 1213 12257 1225 12291
rect 1259 12288 1271 12291
rect 2866 12288 2872 12300
rect 1259 12260 2872 12288
rect 1259 12257 1271 12260
rect 1213 12251 1271 12257
rect 2866 12248 2872 12260
rect 2924 12248 2930 12300
rect 3421 12291 3479 12297
rect 3421 12257 3433 12291
rect 3467 12288 3479 12291
rect 3467 12260 4022 12288
rect 3467 12257 3479 12260
rect 3421 12251 3479 12257
rect 1302 12180 1308 12232
rect 1360 12180 1366 12232
rect 1670 12229 1676 12232
rect 1632 12223 1676 12229
rect 1632 12189 1644 12223
rect 1632 12183 1676 12189
rect 1670 12180 1676 12183
rect 1728 12180 1734 12232
rect 1854 12229 1860 12232
rect 1811 12223 1860 12229
rect 1811 12189 1823 12223
rect 1857 12189 1860 12223
rect 1811 12183 1860 12189
rect 1854 12180 1860 12183
rect 1912 12180 1918 12232
rect 1946 12180 1952 12232
rect 2004 12220 2010 12232
rect 2041 12223 2099 12229
rect 2041 12220 2053 12223
rect 2004 12192 2053 12220
rect 2004 12180 2010 12192
rect 2041 12189 2053 12192
rect 2087 12189 2099 12223
rect 2041 12183 2099 12189
rect 3326 12180 3332 12232
rect 3384 12220 3390 12232
rect 3994 12231 4022 12260
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 6288 12297 6316 12328
rect 4249 12291 4307 12297
rect 4249 12288 4261 12291
rect 4212 12260 4261 12288
rect 4212 12248 4218 12260
rect 4249 12257 4261 12260
rect 4295 12257 4307 12291
rect 4249 12251 4307 12257
rect 5997 12291 6055 12297
rect 5997 12257 6009 12291
rect 6043 12288 6055 12291
rect 6273 12291 6331 12297
rect 6043 12260 6224 12288
rect 6043 12257 6055 12260
rect 5997 12251 6055 12257
rect 3513 12223 3571 12229
rect 3513 12220 3525 12223
rect 3384 12192 3525 12220
rect 3384 12180 3390 12192
rect 3513 12189 3525 12192
rect 3559 12189 3571 12223
rect 3513 12183 3571 12189
rect 3992 12225 4050 12231
rect 3992 12191 4004 12225
rect 4038 12191 4050 12225
rect 3992 12185 4050 12191
rect 5074 12180 5080 12232
rect 5132 12220 5138 12232
rect 5132 12192 5856 12220
rect 5132 12180 5138 12192
rect 5828 12161 5856 12192
rect 5813 12155 5871 12161
rect 5460 12124 5672 12152
rect 1029 12087 1087 12093
rect 1029 12053 1041 12087
rect 1075 12084 1087 12087
rect 1578 12084 1584 12096
rect 1075 12056 1584 12084
rect 1075 12053 1087 12056
rect 1029 12047 1087 12053
rect 1578 12044 1584 12056
rect 1636 12044 1642 12096
rect 1762 12044 1768 12096
rect 1820 12084 1826 12096
rect 5460 12084 5488 12124
rect 1820 12056 5488 12084
rect 5644 12084 5672 12124
rect 5813 12121 5825 12155
rect 5859 12121 5871 12155
rect 5813 12115 5871 12121
rect 5994 12084 6000 12096
rect 5644 12056 6000 12084
rect 1820 12044 1826 12056
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6086 12044 6092 12096
rect 6144 12044 6150 12096
rect 6196 12084 6224 12260
rect 6273 12257 6285 12291
rect 6319 12257 6331 12291
rect 6273 12251 6331 12257
rect 6362 12248 6368 12300
rect 6420 12288 6426 12300
rect 6457 12291 6515 12297
rect 6457 12288 6469 12291
rect 6420 12260 6469 12288
rect 6420 12248 6426 12260
rect 6457 12257 6469 12260
rect 6503 12257 6515 12291
rect 6567 12288 6595 12396
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 7190 12424 7196 12436
rect 6880 12396 7196 12424
rect 6880 12384 6886 12396
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 7466 12384 7472 12436
rect 7524 12424 7530 12436
rect 7926 12424 7932 12436
rect 7524 12396 7932 12424
rect 7524 12384 7530 12396
rect 7926 12384 7932 12396
rect 7984 12424 7990 12436
rect 8570 12424 8576 12436
rect 7984 12396 8576 12424
rect 7984 12384 7990 12396
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 8754 12384 8760 12436
rect 8812 12424 8818 12436
rect 10042 12424 10048 12436
rect 8812 12396 10048 12424
rect 8812 12384 8818 12396
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 10689 12427 10747 12433
rect 10689 12393 10701 12427
rect 10735 12424 10747 12427
rect 10778 12424 10784 12436
rect 10735 12396 10784 12424
rect 10735 12393 10747 12396
rect 10689 12387 10747 12393
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 11330 12384 11336 12436
rect 11388 12384 11394 12436
rect 11974 12424 11980 12436
rect 11716 12396 11980 12424
rect 11348 12356 11376 12384
rect 11606 12356 11612 12368
rect 11348 12328 11612 12356
rect 7193 12291 7251 12297
rect 7193 12288 7205 12291
rect 6567 12260 7205 12288
rect 6457 12251 6515 12257
rect 7193 12257 7205 12260
rect 7239 12257 7251 12291
rect 7193 12251 7251 12257
rect 8573 12291 8631 12297
rect 8573 12257 8585 12291
rect 8619 12288 8631 12291
rect 8619 12260 9171 12288
rect 8619 12257 8631 12260
rect 8573 12251 8631 12257
rect 6822 12229 6828 12232
rect 6784 12223 6828 12229
rect 6784 12189 6796 12223
rect 6784 12183 6828 12189
rect 6822 12180 6828 12183
rect 6880 12180 6886 12232
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 6972 12192 7017 12220
rect 6972 12180 6978 12192
rect 8662 12180 8668 12232
rect 8720 12180 8726 12232
rect 9030 12229 9036 12232
rect 8992 12223 9036 12229
rect 8992 12189 9004 12223
rect 8992 12183 9036 12189
rect 9030 12180 9036 12183
rect 9088 12180 9094 12232
rect 9143 12231 9171 12260
rect 10870 12248 10876 12300
rect 10928 12288 10934 12300
rect 11149 12291 11207 12297
rect 10928 12260 11100 12288
rect 10928 12248 10934 12260
rect 9128 12225 9186 12231
rect 9128 12191 9140 12225
rect 9174 12191 9186 12225
rect 9128 12185 9186 12191
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12220 9459 12223
rect 9447 12192 10364 12220
rect 9447 12189 9459 12192
rect 9401 12183 9459 12189
rect 6730 12084 6736 12096
rect 6196 12056 6736 12084
rect 6730 12044 6736 12056
rect 6788 12084 6794 12096
rect 8202 12084 8208 12096
rect 6788 12056 8208 12084
rect 6788 12044 6794 12056
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 10336 12084 10364 12192
rect 10410 12180 10416 12232
rect 10468 12220 10474 12232
rect 10468 12192 11008 12220
rect 10468 12180 10474 12192
rect 10980 12161 11008 12192
rect 10965 12155 11023 12161
rect 10965 12121 10977 12155
rect 11011 12121 11023 12155
rect 11072 12152 11100 12260
rect 11149 12257 11161 12291
rect 11195 12288 11207 12291
rect 11348 12288 11376 12328
rect 11606 12316 11612 12328
rect 11664 12316 11670 12368
rect 11716 12297 11744 12396
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12253 12427 12311 12433
rect 12253 12393 12265 12427
rect 12299 12424 12311 12427
rect 12802 12424 12808 12436
rect 12299 12396 12808 12424
rect 12299 12393 12311 12396
rect 12253 12387 12311 12393
rect 12802 12384 12808 12396
rect 12860 12384 12866 12436
rect 12995 12427 13053 12433
rect 12995 12393 13007 12427
rect 13041 12424 13053 12427
rect 13630 12424 13636 12436
rect 13041 12396 13636 12424
rect 13041 12393 13053 12396
rect 12995 12387 13053 12393
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 14918 12384 14924 12436
rect 14976 12384 14982 12436
rect 15286 12384 15292 12436
rect 15344 12384 15350 12436
rect 15378 12384 15384 12436
rect 15436 12424 15442 12436
rect 15749 12427 15807 12433
rect 15749 12424 15761 12427
rect 15436 12396 15761 12424
rect 15436 12384 15442 12396
rect 15749 12393 15761 12396
rect 15795 12393 15807 12427
rect 15749 12387 15807 12393
rect 16393 12427 16451 12433
rect 16393 12393 16405 12427
rect 16439 12393 16451 12427
rect 16393 12387 16451 12393
rect 16945 12427 17003 12433
rect 16945 12393 16957 12427
rect 16991 12424 17003 12427
rect 17034 12424 17040 12436
rect 16991 12396 17040 12424
rect 16991 12393 17003 12396
rect 16945 12387 17003 12393
rect 11790 12316 11796 12368
rect 11848 12356 11854 12368
rect 14936 12356 14964 12384
rect 16408 12356 16436 12387
rect 17034 12384 17040 12396
rect 17092 12384 17098 12436
rect 18515 12427 18573 12433
rect 18515 12424 18527 12427
rect 17788 12396 18527 12424
rect 17788 12365 17816 12396
rect 18515 12393 18527 12396
rect 18561 12424 18573 12427
rect 19150 12424 19156 12436
rect 18561 12396 19156 12424
rect 18561 12393 18573 12396
rect 18515 12387 18573 12393
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 20073 12427 20131 12433
rect 20073 12393 20085 12427
rect 20119 12424 20131 12427
rect 20162 12424 20168 12436
rect 20119 12396 20168 12424
rect 20119 12393 20131 12396
rect 20073 12387 20131 12393
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 20809 12427 20867 12433
rect 20809 12393 20821 12427
rect 20855 12424 20867 12427
rect 21082 12424 21088 12436
rect 20855 12396 21088 12424
rect 20855 12393 20867 12396
rect 20809 12387 20867 12393
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 21174 12384 21180 12436
rect 21232 12424 21238 12436
rect 21542 12424 21548 12436
rect 21232 12396 21548 12424
rect 21232 12384 21238 12396
rect 21542 12384 21548 12396
rect 21600 12384 21606 12436
rect 21735 12427 21793 12433
rect 21735 12393 21747 12427
rect 21781 12424 21793 12427
rect 22002 12424 22008 12436
rect 21781 12396 22008 12424
rect 21781 12393 21793 12396
rect 21735 12387 21793 12393
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 23293 12427 23351 12433
rect 23293 12393 23305 12427
rect 23339 12424 23351 12427
rect 23382 12424 23388 12436
rect 23339 12396 23388 12424
rect 23339 12393 23351 12396
rect 23293 12387 23351 12393
rect 23382 12384 23388 12396
rect 23440 12384 23446 12436
rect 23943 12427 24001 12433
rect 23943 12393 23955 12427
rect 23989 12424 24001 12427
rect 24210 12424 24216 12436
rect 23989 12396 24216 12424
rect 23989 12393 24001 12396
rect 23943 12387 24001 12393
rect 24210 12384 24216 12396
rect 24268 12384 24274 12436
rect 25501 12427 25559 12433
rect 25501 12393 25513 12427
rect 25547 12424 25559 12427
rect 25774 12424 25780 12436
rect 25547 12396 25780 12424
rect 25547 12393 25559 12396
rect 25501 12387 25559 12393
rect 25774 12384 25780 12396
rect 25832 12384 25838 12436
rect 26142 12384 26148 12436
rect 26200 12424 26206 12436
rect 26887 12427 26945 12433
rect 26887 12424 26899 12427
rect 26200 12396 26899 12424
rect 26200 12384 26206 12396
rect 26887 12393 26899 12396
rect 26933 12424 26945 12427
rect 27430 12424 27436 12436
rect 26933 12396 27436 12424
rect 26933 12393 26945 12396
rect 26887 12387 26945 12393
rect 27430 12384 27436 12396
rect 27488 12384 27494 12436
rect 27890 12384 27896 12436
rect 27948 12424 27954 12436
rect 28261 12427 28319 12433
rect 28261 12424 28273 12427
rect 27948 12396 28273 12424
rect 27948 12384 27954 12396
rect 28261 12393 28273 12396
rect 28307 12393 28319 12427
rect 28261 12387 28319 12393
rect 28994 12384 29000 12436
rect 29052 12424 29058 12436
rect 30377 12427 30435 12433
rect 30377 12424 30389 12427
rect 29052 12396 30389 12424
rect 29052 12384 29058 12396
rect 30377 12393 30389 12396
rect 30423 12393 30435 12427
rect 30377 12387 30435 12393
rect 11848 12328 12664 12356
rect 14936 12328 16436 12356
rect 17773 12359 17831 12365
rect 11848 12316 11854 12328
rect 11195 12260 11376 12288
rect 11425 12291 11483 12297
rect 11195 12257 11207 12260
rect 11149 12251 11207 12257
rect 11425 12257 11437 12291
rect 11471 12257 11483 12291
rect 11425 12251 11483 12257
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12257 11759 12291
rect 11701 12251 11759 12257
rect 11977 12291 12035 12297
rect 11977 12257 11989 12291
rect 12023 12288 12035 12291
rect 12066 12288 12072 12300
rect 12023 12260 12072 12288
rect 12023 12257 12035 12260
rect 11977 12251 12035 12257
rect 11440 12220 11468 12251
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 12437 12291 12495 12297
rect 12437 12257 12449 12291
rect 12483 12257 12495 12291
rect 12437 12251 12495 12257
rect 12452 12220 12480 12251
rect 12526 12248 12532 12300
rect 12584 12248 12590 12300
rect 11440 12192 12480 12220
rect 12636 12220 12664 12328
rect 17773 12325 17785 12359
rect 17819 12325 17831 12359
rect 17773 12319 17831 12325
rect 25976 12328 26559 12356
rect 25976 12300 26004 12328
rect 13170 12248 13176 12300
rect 13228 12288 13234 12300
rect 13265 12291 13323 12297
rect 13265 12288 13277 12291
rect 13228 12260 13277 12288
rect 13228 12248 13234 12260
rect 13265 12257 13277 12260
rect 13311 12257 13323 12291
rect 13265 12251 13323 12257
rect 13722 12248 13728 12300
rect 13780 12248 13786 12300
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 14921 12291 14979 12297
rect 14921 12288 14933 12291
rect 13964 12260 14933 12288
rect 13964 12248 13970 12260
rect 14921 12257 14933 12260
rect 14967 12288 14979 12291
rect 15102 12288 15108 12300
rect 14967 12260 15108 12288
rect 14967 12257 14979 12260
rect 14921 12251 14979 12257
rect 15102 12248 15108 12260
rect 15160 12248 15166 12300
rect 15194 12248 15200 12300
rect 15252 12248 15258 12300
rect 15473 12291 15531 12297
rect 15473 12257 15485 12291
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 15933 12291 15991 12297
rect 15933 12257 15945 12291
rect 15979 12257 15991 12291
rect 15933 12251 15991 12257
rect 12992 12223 13050 12229
rect 12992 12220 13004 12223
rect 12636 12192 13004 12220
rect 11793 12155 11851 12161
rect 11793 12152 11805 12155
rect 11072 12124 11805 12152
rect 10965 12115 11023 12121
rect 11793 12121 11805 12124
rect 11839 12121 11851 12155
rect 11793 12115 11851 12121
rect 11241 12087 11299 12093
rect 11241 12084 11253 12087
rect 10336 12056 11253 12084
rect 11241 12053 11253 12056
rect 11287 12053 11299 12087
rect 11241 12047 11299 12053
rect 11514 12044 11520 12096
rect 11572 12044 11578 12096
rect 12452 12084 12480 12192
rect 12992 12189 13004 12192
rect 13038 12189 13050 12223
rect 13740 12220 13768 12248
rect 15488 12220 15516 12251
rect 13740 12192 15516 12220
rect 15948 12220 15976 12251
rect 16022 12248 16028 12300
rect 16080 12288 16086 12300
rect 16301 12291 16359 12297
rect 16301 12288 16313 12291
rect 16080 12260 16313 12288
rect 16080 12248 16086 12260
rect 16301 12257 16313 12260
rect 16347 12257 16359 12291
rect 16301 12251 16359 12257
rect 16390 12248 16396 12300
rect 16448 12288 16454 12300
rect 16577 12291 16635 12297
rect 16577 12288 16589 12291
rect 16448 12260 16589 12288
rect 16448 12248 16454 12260
rect 16577 12257 16589 12260
rect 16623 12257 16635 12291
rect 16577 12251 16635 12257
rect 17218 12248 17224 12300
rect 17276 12248 17282 12300
rect 17497 12291 17555 12297
rect 17497 12257 17509 12291
rect 17543 12288 17555 12291
rect 17586 12288 17592 12300
rect 17543 12260 17592 12288
rect 17543 12257 17555 12260
rect 17497 12251 17555 12257
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 17972 12260 18644 12288
rect 16408 12220 16436 12248
rect 15948 12192 16436 12220
rect 12992 12183 13050 12189
rect 12894 12084 12900 12096
rect 12452 12056 12900 12084
rect 12894 12044 12900 12056
rect 12952 12044 12958 12096
rect 13078 12044 13084 12096
rect 13136 12084 13142 12096
rect 13906 12084 13912 12096
rect 13136 12056 13912 12084
rect 13136 12044 13142 12056
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 14366 12044 14372 12096
rect 14424 12044 14430 12096
rect 14734 12044 14740 12096
rect 14792 12044 14798 12096
rect 15010 12044 15016 12096
rect 15068 12044 15074 12096
rect 15488 12084 15516 12192
rect 15562 12112 15568 12164
rect 15620 12152 15626 12164
rect 16117 12155 16175 12161
rect 16117 12152 16129 12155
rect 15620 12124 16129 12152
rect 15620 12112 15626 12124
rect 16117 12121 16129 12124
rect 16163 12121 16175 12155
rect 16117 12115 16175 12121
rect 16390 12112 16396 12164
rect 16448 12152 16454 12164
rect 17972 12152 18000 12260
rect 18046 12180 18052 12232
rect 18104 12180 18110 12232
rect 18506 12180 18512 12232
rect 18564 12180 18570 12232
rect 18616 12220 18644 12260
rect 18690 12248 18696 12300
rect 18748 12288 18754 12300
rect 18785 12291 18843 12297
rect 18785 12288 18797 12291
rect 18748 12260 18797 12288
rect 18748 12248 18754 12260
rect 18785 12257 18797 12260
rect 18831 12257 18843 12291
rect 18785 12251 18843 12257
rect 19242 12248 19248 12300
rect 19300 12288 19306 12300
rect 20993 12291 21051 12297
rect 20993 12288 21005 12291
rect 19300 12260 21005 12288
rect 19300 12248 19306 12260
rect 19812 12232 19840 12260
rect 20993 12257 21005 12260
rect 21039 12288 21051 12291
rect 21358 12288 21364 12300
rect 21039 12260 21364 12288
rect 21039 12257 21051 12260
rect 20993 12251 21051 12257
rect 21358 12248 21364 12260
rect 21416 12248 21422 12300
rect 21542 12248 21548 12300
rect 21600 12288 21606 12300
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 21600 12260 22017 12288
rect 21600 12248 21606 12260
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 23477 12291 23535 12297
rect 23477 12257 23489 12291
rect 23523 12288 23535 12291
rect 23842 12288 23848 12300
rect 23523 12260 23848 12288
rect 23523 12257 23535 12260
rect 23477 12251 23535 12257
rect 23842 12248 23848 12260
rect 23900 12248 23906 12300
rect 24118 12248 24124 12300
rect 24176 12288 24182 12300
rect 24213 12291 24271 12297
rect 24213 12288 24225 12291
rect 24176 12260 24225 12288
rect 24176 12248 24182 12260
rect 24213 12257 24225 12260
rect 24259 12257 24271 12291
rect 24213 12251 24271 12257
rect 25406 12248 25412 12300
rect 25464 12288 25470 12300
rect 25685 12291 25743 12297
rect 25685 12288 25697 12291
rect 25464 12260 25697 12288
rect 25464 12248 25470 12260
rect 25685 12257 25697 12260
rect 25731 12288 25743 12291
rect 25958 12288 25964 12300
rect 25731 12260 25964 12288
rect 25731 12257 25743 12260
rect 25685 12251 25743 12257
rect 25958 12248 25964 12260
rect 26016 12248 26022 12300
rect 26142 12248 26148 12300
rect 26200 12248 26206 12300
rect 26418 12248 26424 12300
rect 26476 12248 26482 12300
rect 26531 12288 26559 12328
rect 28534 12288 28540 12300
rect 26531 12260 28540 12288
rect 28534 12248 28540 12260
rect 28592 12248 28598 12300
rect 28629 12291 28687 12297
rect 28629 12257 28641 12291
rect 28675 12288 28687 12291
rect 28675 12260 29408 12288
rect 28675 12257 28687 12260
rect 28629 12251 28687 12257
rect 18616 12192 19472 12220
rect 16448 12124 18000 12152
rect 16448 12112 16454 12124
rect 16574 12084 16580 12096
rect 15488 12056 16580 12084
rect 16574 12044 16580 12056
rect 16632 12044 16638 12096
rect 17034 12044 17040 12096
rect 17092 12044 17098 12096
rect 18064 12084 18092 12180
rect 18874 12084 18880 12096
rect 18064 12056 18880 12084
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 19444 12084 19472 12192
rect 19794 12180 19800 12232
rect 19852 12180 19858 12232
rect 20346 12180 20352 12232
rect 20404 12220 20410 12232
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 20404 12192 21281 12220
rect 20404 12180 20410 12192
rect 21269 12189 21281 12192
rect 21315 12189 21327 12223
rect 21269 12183 21327 12189
rect 21174 12084 21180 12096
rect 19444 12056 21180 12084
rect 21174 12044 21180 12056
rect 21232 12044 21238 12096
rect 21284 12084 21312 12183
rect 21726 12180 21732 12232
rect 21784 12180 21790 12232
rect 21818 12180 21824 12232
rect 21876 12220 21882 12232
rect 23014 12220 23020 12232
rect 21876 12192 23020 12220
rect 21876 12180 21882 12192
rect 23014 12180 23020 12192
rect 23072 12180 23078 12232
rect 23934 12180 23940 12232
rect 23992 12180 23998 12232
rect 25869 12223 25927 12229
rect 25869 12189 25881 12223
rect 25915 12220 25927 12223
rect 26160 12220 26188 12248
rect 29380 12232 29408 12260
rect 30466 12248 30472 12300
rect 30524 12288 30530 12300
rect 30561 12291 30619 12297
rect 30561 12288 30573 12291
rect 30524 12260 30573 12288
rect 30524 12248 30530 12260
rect 30561 12257 30573 12260
rect 30607 12257 30619 12291
rect 30561 12251 30619 12257
rect 25915 12192 26188 12220
rect 25915 12189 25927 12192
rect 25869 12183 25927 12189
rect 26878 12180 26884 12232
rect 26936 12180 26942 12232
rect 27157 12223 27215 12229
rect 27157 12189 27169 12223
rect 27203 12220 27215 12223
rect 28074 12220 28080 12232
rect 27203 12192 28080 12220
rect 27203 12189 27215 12192
rect 27157 12183 27215 12189
rect 28074 12180 28080 12192
rect 28132 12180 28138 12232
rect 28905 12223 28963 12229
rect 28905 12220 28917 12223
rect 28644 12192 28917 12220
rect 21910 12084 21916 12096
rect 21284 12056 21916 12084
rect 21910 12044 21916 12056
rect 21968 12044 21974 12096
rect 22646 12044 22652 12096
rect 22704 12084 22710 12096
rect 28644 12084 28672 12192
rect 28905 12189 28917 12192
rect 28951 12189 28963 12223
rect 28905 12183 28963 12189
rect 29362 12180 29368 12232
rect 29420 12180 29426 12232
rect 22704 12056 28672 12084
rect 22704 12044 22710 12056
rect 28810 12044 28816 12096
rect 28868 12084 28874 12096
rect 30009 12087 30067 12093
rect 30009 12084 30021 12087
rect 28868 12056 30021 12084
rect 28868 12044 28874 12056
rect 30009 12053 30021 12056
rect 30055 12053 30067 12087
rect 30009 12047 30067 12053
rect 552 11994 30912 12016
rect 552 11942 4193 11994
rect 4245 11942 4257 11994
rect 4309 11942 4321 11994
rect 4373 11942 4385 11994
rect 4437 11942 4449 11994
rect 4501 11942 11783 11994
rect 11835 11942 11847 11994
rect 11899 11942 11911 11994
rect 11963 11942 11975 11994
rect 12027 11942 12039 11994
rect 12091 11942 19373 11994
rect 19425 11942 19437 11994
rect 19489 11942 19501 11994
rect 19553 11942 19565 11994
rect 19617 11942 19629 11994
rect 19681 11942 26963 11994
rect 27015 11942 27027 11994
rect 27079 11942 27091 11994
rect 27143 11942 27155 11994
rect 27207 11942 27219 11994
rect 27271 11942 30912 11994
rect 552 11920 30912 11942
rect 4430 11880 4436 11892
rect 3252 11852 4436 11880
rect 3252 11824 3280 11852
rect 4430 11840 4436 11852
rect 4488 11880 4494 11892
rect 4982 11880 4988 11892
rect 4488 11852 4988 11880
rect 4488 11840 4494 11852
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 5350 11840 5356 11892
rect 5408 11840 5414 11892
rect 6086 11880 6092 11892
rect 5552 11852 6092 11880
rect 3234 11772 3240 11824
rect 3292 11772 3298 11824
rect 1486 11753 1492 11756
rect 1443 11747 1492 11753
rect 1443 11713 1455 11747
rect 1489 11713 1492 11747
rect 1443 11707 1492 11713
rect 1486 11704 1492 11707
rect 1544 11704 1550 11756
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 3694 11744 3700 11756
rect 1719 11716 3700 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 3694 11704 3700 11716
rect 3752 11704 3758 11756
rect 3878 11753 3884 11756
rect 3835 11747 3884 11753
rect 3835 11713 3847 11747
rect 3881 11713 3884 11747
rect 3835 11707 3884 11713
rect 3878 11704 3884 11707
rect 3936 11704 3942 11756
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11744 4123 11747
rect 5552 11744 5580 11852
rect 6086 11840 6092 11852
rect 6144 11840 6150 11892
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 8021 11883 8079 11889
rect 8021 11880 8033 11883
rect 7616 11852 8033 11880
rect 7616 11840 7622 11852
rect 8021 11849 8033 11852
rect 8067 11849 8079 11883
rect 11514 11880 11520 11892
rect 8021 11843 8079 11849
rect 10612 11852 11520 11880
rect 7374 11772 7380 11824
rect 7432 11812 7438 11824
rect 7432 11784 8708 11812
rect 7432 11772 7438 11784
rect 4111 11716 5580 11744
rect 4111 11713 4123 11716
rect 4065 11707 4123 11713
rect 5902 11704 5908 11756
rect 5960 11744 5966 11756
rect 6000 11747 6058 11753
rect 6000 11744 6012 11747
rect 5960 11716 6012 11744
rect 5960 11704 5966 11716
rect 6000 11713 6012 11716
rect 6046 11713 6058 11747
rect 6000 11707 6058 11713
rect 6086 11704 6092 11756
rect 6144 11744 6150 11756
rect 6144 11716 8340 11744
rect 6144 11704 6150 11716
rect 937 11679 995 11685
rect 937 11645 949 11679
rect 983 11676 995 11679
rect 1210 11676 1216 11688
rect 983 11648 1216 11676
rect 983 11645 995 11648
rect 937 11639 995 11645
rect 1210 11636 1216 11648
rect 1268 11676 1274 11688
rect 1762 11676 1768 11688
rect 1268 11648 1768 11676
rect 1268 11636 1274 11648
rect 1762 11636 1768 11648
rect 1820 11636 1826 11688
rect 3326 11636 3332 11688
rect 3384 11676 3390 11688
rect 4798 11676 4804 11688
rect 3384 11648 4804 11676
rect 3384 11636 3390 11648
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 5537 11679 5595 11685
rect 5537 11645 5549 11679
rect 5583 11676 5595 11679
rect 5626 11676 5632 11688
rect 5583 11648 5632 11676
rect 5583 11645 5595 11648
rect 5537 11639 5595 11645
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 5810 11636 5816 11688
rect 5868 11676 5874 11688
rect 6273 11679 6331 11685
rect 6273 11676 6285 11679
rect 5868 11648 6285 11676
rect 5868 11636 5874 11648
rect 6273 11645 6285 11648
rect 6319 11645 6331 11679
rect 6273 11639 6331 11645
rect 7926 11636 7932 11688
rect 7984 11636 7990 11688
rect 8202 11636 8208 11688
rect 8260 11636 8266 11688
rect 3053 11611 3111 11617
rect 3053 11577 3065 11611
rect 3099 11608 3111 11611
rect 3418 11608 3424 11620
rect 3099 11580 3424 11608
rect 3099 11577 3111 11580
rect 3053 11571 3111 11577
rect 3418 11568 3424 11580
rect 3476 11568 3482 11620
rect 8312 11608 8340 11716
rect 8570 11636 8576 11688
rect 8628 11636 8634 11688
rect 8680 11685 8708 11784
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 9496 11747 9554 11753
rect 9496 11744 9508 11747
rect 8904 11716 9508 11744
rect 8904 11704 8910 11716
rect 9496 11713 9508 11716
rect 9542 11713 9554 11747
rect 9496 11707 9554 11713
rect 9769 11747 9827 11753
rect 9769 11713 9781 11747
rect 9815 11744 9827 11747
rect 10612 11744 10640 11852
rect 11514 11840 11520 11852
rect 11572 11840 11578 11892
rect 11606 11840 11612 11892
rect 11664 11880 11670 11892
rect 11664 11852 12664 11880
rect 11664 11840 11670 11852
rect 12636 11812 12664 11852
rect 12710 11840 12716 11892
rect 12768 11880 12774 11892
rect 15933 11883 15991 11889
rect 15933 11880 15945 11883
rect 12768 11852 15945 11880
rect 12768 11840 12774 11852
rect 15933 11849 15945 11852
rect 15979 11880 15991 11883
rect 16022 11880 16028 11892
rect 15979 11852 16028 11880
rect 15979 11849 15991 11852
rect 15933 11843 15991 11849
rect 16022 11840 16028 11852
rect 16080 11840 16086 11892
rect 18417 11883 18475 11889
rect 18417 11849 18429 11883
rect 18463 11880 18475 11883
rect 18506 11880 18512 11892
rect 18463 11852 18512 11880
rect 18463 11849 18475 11852
rect 18417 11843 18475 11849
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 20717 11883 20775 11889
rect 18708 11852 20668 11880
rect 13078 11812 13084 11824
rect 12636 11784 13084 11812
rect 13078 11772 13084 11784
rect 13136 11772 13142 11824
rect 13538 11812 13544 11824
rect 13372 11784 13544 11812
rect 9815 11716 10640 11744
rect 11149 11747 11207 11753
rect 9815 11713 9827 11716
rect 9769 11707 9827 11713
rect 11149 11713 11161 11747
rect 11195 11744 11207 11747
rect 11514 11744 11520 11756
rect 11195 11716 11520 11744
rect 11195 11713 11207 11716
rect 11149 11707 11207 11713
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 11977 11747 12035 11753
rect 11719 11735 11836 11744
rect 11704 11729 11836 11735
rect 11704 11695 11716 11729
rect 11750 11716 11836 11729
rect 11750 11695 11762 11716
rect 11704 11689 11762 11695
rect 11808 11688 11836 11716
rect 11977 11713 11989 11747
rect 12023 11744 12035 11747
rect 12342 11744 12348 11756
rect 12023 11716 12348 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 12434 11704 12440 11756
rect 12492 11744 12498 11756
rect 13372 11744 13400 11784
rect 13538 11772 13544 11784
rect 13596 11772 13602 11824
rect 15102 11772 15108 11824
rect 15160 11812 15166 11824
rect 16298 11812 16304 11824
rect 15160 11784 16304 11812
rect 15160 11772 15166 11784
rect 16298 11772 16304 11784
rect 16356 11772 16362 11824
rect 18708 11812 18736 11852
rect 18340 11784 18736 11812
rect 20640 11812 20668 11852
rect 20717 11849 20729 11883
rect 20763 11880 20775 11883
rect 21726 11880 21732 11892
rect 20763 11852 21732 11880
rect 20763 11849 20775 11852
rect 20717 11843 20775 11849
rect 21726 11840 21732 11852
rect 21784 11840 21790 11892
rect 21910 11840 21916 11892
rect 21968 11880 21974 11892
rect 23569 11883 23627 11889
rect 21968 11852 23152 11880
rect 21968 11840 21974 11852
rect 20990 11812 20996 11824
rect 20640 11784 20996 11812
rect 14047 11745 14105 11751
rect 14047 11744 14059 11745
rect 12492 11716 13400 11744
rect 13464 11716 14059 11744
rect 12492 11704 12498 11716
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 8754 11636 8760 11688
rect 8812 11676 8818 11688
rect 9033 11679 9091 11685
rect 9033 11676 9045 11679
rect 8812 11648 9045 11676
rect 8812 11636 8818 11648
rect 9033 11645 9045 11648
rect 9079 11645 9091 11679
rect 9033 11639 9091 11645
rect 9140 11648 10456 11676
rect 9140 11608 9168 11648
rect 8312 11580 9168 11608
rect 10428 11608 10456 11648
rect 11238 11636 11244 11688
rect 11296 11636 11302 11688
rect 11606 11676 11612 11688
rect 11348 11648 11612 11676
rect 11348 11608 11376 11648
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 11790 11636 11796 11688
rect 11848 11636 11854 11688
rect 11882 11636 11888 11688
rect 11940 11676 11946 11688
rect 13464 11676 13492 11716
rect 14047 11711 14059 11716
rect 14093 11711 14105 11745
rect 14047 11705 14105 11711
rect 14274 11704 14280 11756
rect 14332 11704 14338 11756
rect 16758 11744 16764 11756
rect 16316 11716 16764 11744
rect 11940 11648 13492 11676
rect 11940 11636 11946 11648
rect 13538 11636 13544 11688
rect 13596 11636 13602 11688
rect 13630 11636 13636 11688
rect 13688 11676 13694 11688
rect 13868 11679 13926 11685
rect 13868 11676 13880 11679
rect 13688 11648 13880 11676
rect 13688 11636 13694 11648
rect 13868 11645 13880 11648
rect 13914 11645 13926 11679
rect 13868 11639 13926 11645
rect 14550 11636 14556 11688
rect 14608 11676 14614 11688
rect 15102 11676 15108 11688
rect 14608 11648 15108 11676
rect 14608 11636 14614 11648
rect 15102 11636 15108 11648
rect 15160 11636 15166 11688
rect 16316 11685 16344 11716
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 16942 11751 16948 11756
rect 16899 11745 16948 11751
rect 16899 11711 16911 11745
rect 16945 11711 16948 11745
rect 16899 11705 16948 11711
rect 16942 11704 16948 11705
rect 17000 11704 17006 11756
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 17092 11716 17141 11744
rect 17092 11704 17098 11716
rect 17129 11713 17141 11716
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 18340 11688 18368 11784
rect 20990 11772 20996 11784
rect 21048 11772 21054 11824
rect 18874 11744 18880 11756
rect 18708 11716 18880 11744
rect 16301 11679 16359 11685
rect 16301 11645 16313 11679
rect 16347 11645 16359 11679
rect 16301 11639 16359 11645
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11676 16451 11679
rect 16666 11676 16672 11688
rect 16439 11648 16672 11676
rect 16439 11645 16451 11648
rect 16393 11639 16451 11645
rect 16666 11636 16672 11648
rect 16724 11676 16730 11688
rect 18322 11676 18328 11688
rect 16724 11648 18328 11676
rect 16724 11636 16730 11648
rect 18322 11636 18328 11648
rect 18380 11636 18386 11688
rect 18708 11685 18736 11716
rect 18874 11704 18880 11716
rect 18932 11704 18938 11756
rect 19156 11747 19214 11753
rect 19156 11744 19168 11747
rect 18984 11716 19168 11744
rect 18984 11688 19012 11716
rect 19156 11713 19168 11716
rect 19202 11713 19214 11747
rect 19156 11707 19214 11713
rect 19426 11704 19432 11756
rect 19484 11704 19490 11756
rect 21545 11747 21603 11753
rect 21545 11713 21557 11747
rect 21591 11744 21603 11747
rect 21910 11744 21916 11756
rect 21591 11716 21916 11744
rect 21591 11713 21603 11716
rect 21545 11707 21603 11713
rect 21910 11704 21916 11716
rect 21968 11704 21974 11756
rect 22051 11747 22109 11753
rect 22051 11713 22063 11747
rect 22097 11744 22109 11747
rect 22097 11716 22784 11744
rect 22097 11713 22109 11716
rect 22051 11707 22109 11713
rect 22756 11688 22784 11716
rect 18693 11679 18751 11685
rect 18693 11645 18705 11679
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 18966 11636 18972 11688
rect 19024 11636 19030 11688
rect 22278 11636 22284 11688
rect 22336 11636 22342 11688
rect 22738 11636 22744 11688
rect 22796 11636 22802 11688
rect 10428 11580 11376 11608
rect 13354 11568 13360 11620
rect 13412 11568 13418 11620
rect 1394 11500 1400 11552
rect 1452 11549 1458 11552
rect 1452 11540 1461 11549
rect 1762 11540 1768 11552
rect 1452 11512 1768 11540
rect 1452 11503 1461 11512
rect 1452 11500 1458 11503
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 3795 11543 3853 11549
rect 3795 11509 3807 11543
rect 3841 11540 3853 11543
rect 3970 11540 3976 11552
rect 3841 11512 3976 11540
rect 3841 11509 3853 11512
rect 3795 11503 3853 11509
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 4890 11500 4896 11552
rect 4948 11540 4954 11552
rect 5810 11540 5816 11552
rect 4948 11512 5816 11540
rect 4948 11500 4954 11512
rect 5810 11500 5816 11512
rect 5868 11500 5874 11552
rect 5994 11500 6000 11552
rect 6052 11549 6058 11552
rect 6052 11540 6061 11549
rect 6052 11512 6097 11540
rect 6052 11503 6061 11512
rect 6052 11500 6058 11503
rect 7006 11500 7012 11552
rect 7064 11540 7070 11552
rect 7377 11543 7435 11549
rect 7377 11540 7389 11543
rect 7064 11512 7389 11540
rect 7064 11500 7070 11512
rect 7377 11509 7389 11512
rect 7423 11509 7435 11543
rect 7377 11503 7435 11509
rect 7742 11500 7748 11552
rect 7800 11500 7806 11552
rect 8386 11500 8392 11552
rect 8444 11500 8450 11552
rect 8846 11500 8852 11552
rect 8904 11500 8910 11552
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 9398 11540 9404 11552
rect 9088 11512 9404 11540
rect 9088 11500 9094 11512
rect 9398 11500 9404 11512
rect 9456 11540 9462 11552
rect 9499 11543 9557 11549
rect 9499 11540 9511 11543
rect 9456 11512 9511 11540
rect 9456 11500 9462 11512
rect 9499 11509 9511 11512
rect 9545 11509 9557 11543
rect 9499 11503 9557 11509
rect 11707 11543 11765 11549
rect 11707 11509 11719 11543
rect 11753 11540 11765 11543
rect 12250 11540 12256 11552
rect 11753 11512 12256 11540
rect 11753 11509 11765 11512
rect 11707 11503 11765 11509
rect 12250 11500 12256 11512
rect 12308 11540 12314 11552
rect 13648 11540 13676 11636
rect 23124 11608 23152 11852
rect 23569 11849 23581 11883
rect 23615 11880 23627 11883
rect 23934 11880 23940 11892
rect 23615 11852 23940 11880
rect 23615 11849 23627 11852
rect 23569 11843 23627 11849
rect 23934 11840 23940 11852
rect 23992 11840 23998 11892
rect 24670 11840 24676 11892
rect 24728 11880 24734 11892
rect 26510 11880 26516 11892
rect 24728 11852 26516 11880
rect 24728 11840 24734 11852
rect 26510 11840 26516 11852
rect 26568 11840 26574 11892
rect 26697 11883 26755 11889
rect 26697 11849 26709 11883
rect 26743 11880 26755 11883
rect 26786 11880 26792 11892
rect 26743 11852 26792 11880
rect 26743 11849 26755 11852
rect 26697 11843 26755 11849
rect 26786 11840 26792 11852
rect 26844 11840 26850 11892
rect 27522 11840 27528 11892
rect 27580 11880 27586 11892
rect 27580 11852 27844 11880
rect 27580 11840 27586 11852
rect 23845 11815 23903 11821
rect 23845 11781 23857 11815
rect 23891 11812 23903 11815
rect 27816 11812 27844 11852
rect 28626 11840 28632 11892
rect 28684 11840 28690 11892
rect 28736 11852 29776 11880
rect 23891 11784 24660 11812
rect 27816 11784 28488 11812
rect 23891 11781 23903 11784
rect 23845 11775 23903 11781
rect 24118 11744 24124 11756
rect 24044 11716 24124 11744
rect 24044 11685 24072 11716
rect 24118 11704 24124 11716
rect 24176 11704 24182 11756
rect 24632 11744 24660 11784
rect 25179 11747 25237 11753
rect 24632 11716 24808 11744
rect 24029 11679 24087 11685
rect 24029 11645 24041 11679
rect 24075 11645 24087 11679
rect 24029 11639 24087 11645
rect 24213 11679 24271 11685
rect 24213 11645 24225 11679
rect 24259 11676 24271 11679
rect 24670 11676 24676 11688
rect 24259 11648 24676 11676
rect 24259 11645 24271 11648
rect 24213 11639 24271 11645
rect 24228 11608 24256 11639
rect 24670 11636 24676 11648
rect 24728 11636 24734 11688
rect 24780 11676 24808 11716
rect 25179 11713 25191 11747
rect 25225 11744 25237 11747
rect 25225 11716 25728 11744
rect 25225 11713 25237 11716
rect 25179 11707 25237 11713
rect 25700 11688 25728 11716
rect 26050 11704 26056 11756
rect 26108 11744 26114 11756
rect 26881 11747 26939 11753
rect 26881 11744 26893 11747
rect 26108 11716 26893 11744
rect 26108 11704 26114 11716
rect 26881 11713 26893 11716
rect 26927 11713 26939 11747
rect 26881 11707 26939 11713
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11744 27215 11747
rect 28166 11744 28172 11756
rect 27203 11716 28172 11744
rect 27203 11713 27215 11716
rect 27157 11707 27215 11713
rect 28166 11704 28172 11716
rect 28224 11704 28230 11756
rect 28460 11744 28488 11784
rect 28460 11742 28672 11744
rect 28736 11742 28764 11852
rect 29638 11812 29644 11824
rect 28460 11716 28764 11742
rect 28644 11714 28764 11716
rect 28828 11784 29644 11812
rect 25409 11679 25467 11685
rect 25409 11676 25421 11679
rect 24780 11648 25421 11676
rect 25409 11645 25421 11648
rect 25455 11645 25467 11679
rect 25409 11639 25467 11645
rect 25682 11636 25688 11688
rect 25740 11636 25746 11688
rect 27522 11676 27528 11688
rect 26068 11648 27528 11676
rect 23124 11580 24256 11608
rect 24394 11568 24400 11620
rect 24452 11608 24458 11620
rect 24581 11611 24639 11617
rect 24581 11608 24593 11611
rect 24452 11580 24593 11608
rect 24452 11568 24458 11580
rect 24581 11577 24593 11580
rect 24627 11608 24639 11611
rect 24762 11608 24768 11620
rect 24627 11580 24768 11608
rect 24627 11577 24639 11580
rect 24581 11571 24639 11577
rect 24762 11568 24768 11580
rect 24820 11568 24826 11620
rect 12308 11512 13676 11540
rect 12308 11500 12314 11512
rect 15010 11500 15016 11552
rect 15068 11540 15074 11552
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 15068 11512 15393 11540
rect 15068 11500 15074 11512
rect 15381 11509 15393 11512
rect 15427 11509 15439 11543
rect 15381 11503 15439 11509
rect 16114 11500 16120 11552
rect 16172 11500 16178 11552
rect 16859 11543 16917 11549
rect 16859 11509 16871 11543
rect 16905 11540 16917 11543
rect 17126 11540 17132 11552
rect 16905 11512 17132 11540
rect 16905 11509 16917 11512
rect 16859 11503 16917 11509
rect 17126 11500 17132 11512
rect 17184 11500 17190 11552
rect 19150 11500 19156 11552
rect 19208 11549 19214 11552
rect 19208 11540 19217 11549
rect 19208 11512 19253 11540
rect 19208 11503 19217 11512
rect 19208 11500 19214 11503
rect 22002 11500 22008 11552
rect 22060 11549 22066 11552
rect 22060 11540 22069 11549
rect 25139 11543 25197 11549
rect 25139 11540 25151 11543
rect 22060 11512 25151 11540
rect 22060 11503 22069 11512
rect 25139 11509 25151 11512
rect 25185 11540 25197 11543
rect 26068 11540 26096 11648
rect 27522 11636 27528 11648
rect 27580 11636 27586 11688
rect 27614 11636 27620 11688
rect 27672 11676 27678 11688
rect 28828 11685 28856 11784
rect 29638 11772 29644 11784
rect 29696 11772 29702 11824
rect 29748 11753 29776 11852
rect 29733 11747 29791 11753
rect 29733 11713 29745 11747
rect 29779 11713 29791 11747
rect 29733 11707 29791 11713
rect 28813 11679 28871 11685
rect 28813 11676 28825 11679
rect 27672 11648 28825 11676
rect 27672 11636 27678 11648
rect 28813 11645 28825 11648
rect 28859 11645 28871 11679
rect 29457 11679 29515 11685
rect 29457 11676 29469 11679
rect 28813 11639 28871 11645
rect 29012 11648 29469 11676
rect 29012 11608 29040 11648
rect 29457 11645 29469 11648
rect 29503 11676 29515 11679
rect 29549 11679 29607 11685
rect 29549 11676 29561 11679
rect 29503 11648 29561 11676
rect 29503 11645 29515 11648
rect 29457 11639 29515 11645
rect 29549 11645 29561 11648
rect 29595 11645 29607 11679
rect 29549 11639 29607 11645
rect 27816 11580 29040 11608
rect 29089 11611 29147 11617
rect 25185 11512 26096 11540
rect 25185 11509 25197 11512
rect 25139 11503 25197 11509
rect 22060 11500 22066 11503
rect 26602 11500 26608 11552
rect 26660 11540 26666 11552
rect 27816 11540 27844 11580
rect 29089 11577 29101 11611
rect 29135 11577 29147 11611
rect 29089 11571 29147 11577
rect 26660 11512 27844 11540
rect 26660 11500 26666 11512
rect 28258 11500 28264 11552
rect 28316 11500 28322 11552
rect 28534 11500 28540 11552
rect 28592 11540 28598 11552
rect 29104 11540 29132 11571
rect 28592 11512 29132 11540
rect 28592 11500 28598 11512
rect 552 11450 31072 11472
rect 552 11398 7988 11450
rect 8040 11398 8052 11450
rect 8104 11398 8116 11450
rect 8168 11398 8180 11450
rect 8232 11398 8244 11450
rect 8296 11398 15578 11450
rect 15630 11398 15642 11450
rect 15694 11398 15706 11450
rect 15758 11398 15770 11450
rect 15822 11398 15834 11450
rect 15886 11398 23168 11450
rect 23220 11398 23232 11450
rect 23284 11398 23296 11450
rect 23348 11398 23360 11450
rect 23412 11398 23424 11450
rect 23476 11398 30758 11450
rect 30810 11398 30822 11450
rect 30874 11398 30886 11450
rect 30938 11398 30950 11450
rect 31002 11398 31014 11450
rect 31066 11398 31072 11450
rect 552 11376 31072 11398
rect 934 11296 940 11348
rect 992 11336 998 11348
rect 2130 11336 2136 11348
rect 992 11308 2136 11336
rect 992 11296 998 11308
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 3513 11339 3571 11345
rect 3513 11305 3525 11339
rect 3559 11336 3571 11339
rect 4522 11336 4528 11348
rect 3559 11308 4528 11336
rect 3559 11305 3571 11308
rect 3513 11299 3571 11305
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 4798 11296 4804 11348
rect 4856 11336 4862 11348
rect 4856 11308 5580 11336
rect 4856 11296 4862 11308
rect 3878 11268 3884 11280
rect 3252 11240 3884 11268
rect 1213 11203 1271 11209
rect 1213 11169 1225 11203
rect 1259 11200 1271 11203
rect 1259 11172 2038 11200
rect 1259 11169 1271 11172
rect 1213 11163 1271 11169
rect 1394 11092 1400 11144
rect 1452 11132 1458 11144
rect 1489 11135 1547 11141
rect 1489 11132 1501 11135
rect 1452 11104 1501 11132
rect 1452 11092 1458 11104
rect 1489 11101 1501 11104
rect 1535 11101 1547 11135
rect 1489 11095 1547 11101
rect 1670 11092 1676 11144
rect 1728 11132 1734 11144
rect 2010 11141 2038 11172
rect 2130 11160 2136 11212
rect 2188 11200 2194 11212
rect 2225 11203 2283 11209
rect 2225 11200 2237 11203
rect 2188 11172 2237 11200
rect 2188 11160 2194 11172
rect 2225 11169 2237 11172
rect 2271 11169 2283 11203
rect 2225 11163 2283 11169
rect 1816 11135 1874 11141
rect 1816 11132 1828 11135
rect 1728 11104 1828 11132
rect 1728 11092 1734 11104
rect 1816 11101 1828 11104
rect 1862 11101 1874 11135
rect 1816 11095 1874 11101
rect 1995 11135 2053 11141
rect 1995 11101 2007 11135
rect 2041 11132 2053 11135
rect 3252 11132 3280 11240
rect 3878 11228 3884 11240
rect 3936 11228 3942 11280
rect 4430 11228 4436 11280
rect 4488 11268 4494 11280
rect 4488 11240 4568 11268
rect 4488 11228 4494 11240
rect 4540 11209 4568 11240
rect 4614 11228 4620 11280
rect 4672 11268 4678 11280
rect 4709 11271 4767 11277
rect 4709 11268 4721 11271
rect 4672 11240 4721 11268
rect 4672 11228 4678 11240
rect 4709 11237 4721 11240
rect 4755 11237 4767 11271
rect 4709 11231 4767 11237
rect 5074 11228 5080 11280
rect 5132 11268 5138 11280
rect 5445 11271 5503 11277
rect 5445 11268 5457 11271
rect 5132 11240 5457 11268
rect 5132 11228 5138 11240
rect 5445 11237 5457 11240
rect 5491 11237 5503 11271
rect 5552 11268 5580 11308
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 5776 11308 6868 11336
rect 5776 11296 5782 11308
rect 5905 11271 5963 11277
rect 5905 11268 5917 11271
rect 5552 11240 5917 11268
rect 5445 11231 5503 11237
rect 5905 11237 5917 11240
rect 5951 11237 5963 11271
rect 5905 11231 5963 11237
rect 6380 11240 6776 11268
rect 6380 11212 6408 11240
rect 6748 11212 6776 11240
rect 3697 11203 3755 11209
rect 3697 11169 3709 11203
rect 3743 11200 3755 11203
rect 4525 11203 4583 11209
rect 3743 11172 4476 11200
rect 3743 11169 3755 11172
rect 3697 11163 3755 11169
rect 2041 11104 3280 11132
rect 2041 11101 2053 11104
rect 1995 11095 2053 11101
rect 3970 11092 3976 11144
rect 4028 11092 4034 11144
rect 4448 11132 4476 11172
rect 4525 11169 4537 11203
rect 4571 11169 4583 11203
rect 5169 11203 5227 11209
rect 5169 11200 5181 11203
rect 4525 11163 4583 11169
rect 4632 11172 5181 11200
rect 4632 11132 4660 11172
rect 5169 11169 5181 11172
rect 5215 11200 5227 11203
rect 5350 11200 5356 11212
rect 5215 11172 5356 11200
rect 5215 11169 5227 11172
rect 5169 11163 5227 11169
rect 5350 11160 5356 11172
rect 5408 11160 5414 11212
rect 6362 11160 6368 11212
rect 6420 11160 6426 11212
rect 6454 11160 6460 11212
rect 6512 11200 6518 11212
rect 6549 11203 6607 11209
rect 6549 11200 6561 11203
rect 6512 11172 6561 11200
rect 6512 11160 6518 11172
rect 6549 11169 6561 11172
rect 6595 11169 6607 11203
rect 6549 11163 6607 11169
rect 6730 11160 6736 11212
rect 6788 11160 6794 11212
rect 6840 11200 6868 11308
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 8662 11336 8668 11348
rect 8260 11308 8668 11336
rect 8260 11296 8266 11308
rect 8662 11296 8668 11308
rect 8720 11336 8726 11348
rect 9582 11336 9588 11348
rect 8720 11308 9588 11336
rect 8720 11296 8726 11308
rect 9582 11296 9588 11308
rect 9640 11336 9646 11348
rect 9677 11339 9735 11345
rect 9677 11336 9689 11339
rect 9640 11308 9689 11336
rect 9640 11296 9646 11308
rect 9677 11305 9689 11308
rect 9723 11305 9735 11339
rect 11793 11339 11851 11345
rect 9677 11299 9735 11305
rect 10336 11308 11284 11336
rect 10336 11268 10364 11308
rect 11054 11268 11060 11280
rect 8588 11240 10364 11268
rect 10428 11240 11060 11268
rect 8588 11212 8616 11240
rect 7469 11203 7527 11209
rect 6840 11172 7239 11200
rect 4448 11104 4660 11132
rect 5994 11092 6000 11144
rect 6052 11132 6058 11144
rect 6914 11132 6920 11144
rect 6052 11104 6920 11132
rect 6052 11092 6058 11104
rect 6914 11092 6920 11104
rect 6972 11132 6978 11144
rect 7211 11143 7239 11172
rect 7469 11169 7481 11203
rect 7515 11200 7527 11203
rect 7742 11200 7748 11212
rect 7515 11172 7748 11200
rect 7515 11169 7527 11172
rect 7469 11163 7527 11169
rect 7742 11160 7748 11172
rect 7800 11160 7806 11212
rect 8570 11160 8576 11212
rect 8628 11160 8634 11212
rect 8938 11160 8944 11212
rect 8996 11160 9002 11212
rect 9490 11160 9496 11212
rect 9548 11200 9554 11212
rect 10428 11209 10456 11240
rect 11054 11228 11060 11240
rect 11112 11228 11118 11280
rect 9585 11203 9643 11209
rect 9585 11200 9597 11203
rect 9548 11172 9597 11200
rect 9548 11160 9554 11172
rect 9585 11169 9597 11172
rect 9631 11169 9643 11203
rect 9585 11163 9643 11169
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11169 10471 11203
rect 10413 11163 10471 11169
rect 10502 11160 10508 11212
rect 10560 11200 10566 11212
rect 10689 11203 10747 11209
rect 10689 11200 10701 11203
rect 10560 11172 10701 11200
rect 10560 11160 10566 11172
rect 10689 11169 10701 11172
rect 10735 11169 10747 11203
rect 10689 11163 10747 11169
rect 10778 11160 10784 11212
rect 10836 11200 10842 11212
rect 11256 11209 11284 11308
rect 11793 11305 11805 11339
rect 11839 11305 11851 11339
rect 11793 11299 11851 11305
rect 11808 11268 11836 11299
rect 12066 11296 12072 11348
rect 12124 11296 12130 11348
rect 12250 11296 12256 11348
rect 12308 11336 12314 11348
rect 12903 11339 12961 11345
rect 12903 11336 12915 11339
rect 12308 11308 12915 11336
rect 12308 11296 12314 11308
rect 12903 11305 12915 11308
rect 12949 11305 12961 11339
rect 12903 11299 12961 11305
rect 14734 11296 14740 11348
rect 14792 11296 14798 11348
rect 15102 11336 15108 11348
rect 14844 11308 15108 11336
rect 11440 11240 11836 11268
rect 11149 11203 11207 11209
rect 11149 11200 11161 11203
rect 10836 11172 11161 11200
rect 10836 11160 10842 11172
rect 11149 11169 11161 11172
rect 11195 11169 11207 11203
rect 11149 11163 11207 11169
rect 11241 11203 11299 11209
rect 11241 11169 11253 11203
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 7060 11135 7118 11141
rect 7060 11132 7072 11135
rect 6972 11104 7072 11132
rect 6972 11092 6978 11104
rect 7060 11101 7072 11104
rect 7106 11101 7118 11135
rect 7060 11095 7118 11101
rect 7196 11137 7254 11143
rect 7196 11103 7208 11137
rect 7242 11103 7254 11137
rect 7196 11097 7254 11103
rect 8849 11135 8907 11141
rect 8849 11101 8861 11135
rect 8895 11132 8907 11135
rect 9858 11132 9864 11144
rect 8895 11104 9864 11132
rect 8895 11101 8907 11104
rect 8849 11095 8907 11101
rect 9858 11092 9864 11104
rect 9916 11092 9922 11144
rect 11440 11132 11468 11240
rect 12342 11228 12348 11280
rect 12400 11228 12406 11280
rect 11517 11203 11575 11209
rect 11517 11169 11529 11203
rect 11563 11169 11575 11203
rect 11517 11163 11575 11169
rect 11977 11203 12035 11209
rect 11977 11169 11989 11203
rect 12023 11200 12035 11203
rect 12253 11203 12311 11209
rect 12253 11200 12265 11203
rect 12023 11172 12265 11200
rect 12023 11169 12035 11172
rect 11977 11163 12035 11169
rect 12253 11169 12265 11172
rect 12299 11169 12311 11203
rect 12360 11200 12388 11228
rect 13173 11203 13231 11209
rect 12360 11172 12943 11200
rect 12253 11163 12311 11169
rect 10060 11104 11468 11132
rect 11532 11134 11560 11163
rect 11532 11132 11652 11134
rect 12158 11132 12164 11144
rect 11532 11106 12164 11132
rect 11624 11104 12164 11106
rect 3234 11024 3240 11076
rect 3292 11064 3298 11076
rect 6089 11067 6147 11073
rect 6089 11064 6101 11067
rect 3292 11036 6101 11064
rect 3292 11024 3298 11036
rect 6089 11033 6101 11036
rect 6135 11033 6147 11067
rect 6089 11027 6147 11033
rect 6362 11024 6368 11076
rect 6420 11024 6426 11076
rect 10060 11064 10088 11104
rect 12158 11092 12164 11104
rect 12216 11092 12222 11144
rect 8128 11036 10088 11064
rect 1854 10956 1860 11008
rect 1912 10996 1918 11008
rect 3142 10996 3148 11008
rect 1912 10968 3148 10996
rect 1912 10956 1918 10968
rect 3142 10956 3148 10968
rect 3200 10956 3206 11008
rect 3786 10956 3792 11008
rect 3844 10996 3850 11008
rect 4062 10996 4068 11008
rect 3844 10968 4068 10996
rect 3844 10956 3850 10968
rect 4062 10956 4068 10968
rect 4120 10956 4126 11008
rect 4341 10999 4399 11005
rect 4341 10965 4353 10999
rect 4387 10996 4399 10999
rect 4614 10996 4620 11008
rect 4387 10968 4620 10996
rect 4387 10965 4399 10968
rect 4341 10959 4399 10965
rect 4614 10956 4620 10968
rect 4672 10956 4678 11008
rect 4798 10956 4804 11008
rect 4856 10996 4862 11008
rect 8128 10996 8156 11036
rect 10134 11024 10140 11076
rect 10192 11064 10198 11076
rect 10229 11067 10287 11073
rect 10229 11064 10241 11067
rect 10192 11036 10241 11064
rect 10192 11024 10198 11036
rect 10229 11033 10241 11036
rect 10275 11033 10287 11067
rect 10229 11027 10287 11033
rect 10502 11024 10508 11076
rect 10560 11024 10566 11076
rect 10962 11024 10968 11076
rect 11020 11024 11026 11076
rect 11054 11024 11060 11076
rect 11112 11064 11118 11076
rect 12268 11064 12296 11163
rect 12434 11132 12440 11144
rect 12406 11092 12440 11132
rect 12492 11132 12498 11144
rect 12915 11141 12943 11172
rect 13173 11169 13185 11203
rect 13219 11200 13231 11203
rect 14752 11200 14780 11296
rect 14844 11209 14872 11308
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 16114 11296 16120 11348
rect 16172 11296 16178 11348
rect 16298 11296 16304 11348
rect 16356 11336 16362 11348
rect 16669 11339 16727 11345
rect 16669 11336 16681 11339
rect 16356 11308 16681 11336
rect 16356 11296 16362 11308
rect 16669 11305 16681 11308
rect 16715 11305 16727 11339
rect 16669 11299 16727 11305
rect 17126 11296 17132 11348
rect 17184 11336 17190 11348
rect 17319 11339 17377 11345
rect 17319 11336 17331 11339
rect 17184 11308 17331 11336
rect 17184 11296 17190 11308
rect 17319 11305 17331 11308
rect 17365 11336 17377 11339
rect 18877 11339 18935 11345
rect 17365 11308 18828 11336
rect 17365 11305 17377 11308
rect 17319 11299 17377 11305
rect 15378 11268 15384 11280
rect 15120 11240 15384 11268
rect 15120 11209 15148 11240
rect 15378 11228 15384 11240
rect 15436 11268 15442 11280
rect 15436 11240 16068 11268
rect 15436 11228 15442 11240
rect 16040 11212 16068 11240
rect 13219 11172 14780 11200
rect 14829 11203 14887 11209
rect 13219 11169 13231 11172
rect 13173 11163 13231 11169
rect 14829 11169 14841 11203
rect 14875 11169 14887 11203
rect 14829 11163 14887 11169
rect 15105 11203 15163 11209
rect 15105 11169 15117 11203
rect 15151 11169 15163 11203
rect 15105 11163 15163 11169
rect 15470 11160 15476 11212
rect 15528 11160 15534 11212
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11169 15807 11203
rect 15749 11163 15807 11169
rect 12900 11135 12958 11141
rect 12492 11104 12537 11132
rect 12492 11092 12498 11104
rect 12900 11101 12912 11135
rect 12946 11101 12958 11135
rect 12900 11095 12958 11101
rect 13538 11092 13544 11144
rect 13596 11132 13602 11144
rect 15764 11132 15792 11163
rect 16022 11160 16028 11212
rect 16080 11160 16086 11212
rect 16132 11200 16160 11296
rect 18800 11268 18828 11308
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 18966 11336 18972 11348
rect 18923 11308 18972 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 21637 11339 21695 11345
rect 21637 11305 21649 11339
rect 21683 11336 21695 11339
rect 22278 11336 22284 11348
rect 21683 11308 22284 11336
rect 21683 11305 21695 11308
rect 21637 11299 21695 11305
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 22462 11296 22468 11348
rect 22520 11336 22526 11348
rect 24587 11339 24645 11345
rect 24587 11336 24599 11339
rect 22520 11308 24599 11336
rect 22520 11296 22526 11308
rect 24587 11305 24599 11308
rect 24633 11336 24645 11339
rect 24633 11308 25544 11336
rect 24633 11305 24645 11308
rect 24587 11299 24645 11305
rect 19337 11271 19395 11277
rect 19337 11268 19349 11271
rect 18800 11240 19349 11268
rect 19337 11237 19349 11240
rect 19383 11268 19395 11271
rect 19383 11240 20484 11268
rect 19383 11237 19395 11240
rect 19337 11231 19395 11237
rect 17589 11203 17647 11209
rect 17589 11200 17601 11203
rect 16132 11172 17601 11200
rect 17589 11169 17601 11172
rect 17635 11169 17647 11203
rect 17589 11163 17647 11169
rect 18966 11160 18972 11212
rect 19024 11200 19030 11212
rect 19061 11203 19119 11209
rect 19061 11200 19073 11203
rect 19024 11172 19073 11200
rect 19024 11160 19030 11172
rect 19061 11169 19073 11172
rect 19107 11169 19119 11203
rect 19061 11163 19119 11169
rect 19518 11160 19524 11212
rect 19576 11200 19582 11212
rect 19794 11200 19800 11212
rect 19576 11172 19800 11200
rect 19576 11160 19582 11172
rect 19794 11160 19800 11172
rect 19852 11160 19858 11212
rect 20456 11200 20484 11240
rect 21082 11228 21088 11280
rect 21140 11268 21146 11280
rect 25516 11268 25544 11308
rect 25682 11296 25688 11348
rect 25740 11336 25746 11348
rect 25961 11339 26019 11345
rect 25961 11336 25973 11339
rect 25740 11308 25973 11336
rect 25740 11296 25746 11308
rect 25961 11305 25973 11308
rect 26007 11305 26019 11339
rect 26694 11336 26700 11348
rect 25961 11299 26019 11305
rect 26068 11308 26700 11336
rect 26068 11268 26096 11308
rect 26694 11296 26700 11308
rect 26752 11336 26758 11348
rect 26887 11339 26945 11345
rect 26887 11336 26899 11339
rect 26752 11308 26899 11336
rect 26752 11296 26758 11308
rect 26887 11305 26899 11308
rect 26933 11305 26945 11339
rect 26887 11299 26945 11305
rect 27430 11296 27436 11348
rect 27488 11336 27494 11348
rect 30377 11339 30435 11345
rect 30377 11336 30389 11339
rect 27488 11308 30389 11336
rect 27488 11296 27494 11308
rect 30377 11305 30389 11308
rect 30423 11305 30435 11339
rect 30377 11299 30435 11305
rect 21140 11240 21496 11268
rect 25516 11240 26096 11268
rect 21140 11228 21146 11240
rect 20898 11200 20904 11212
rect 20456 11172 20904 11200
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 21468 11209 21496 11240
rect 21453 11203 21511 11209
rect 21453 11169 21465 11203
rect 21499 11169 21511 11203
rect 21453 11163 21511 11169
rect 21818 11160 21824 11212
rect 21876 11160 21882 11212
rect 22002 11160 22008 11212
rect 22060 11200 22066 11212
rect 22240 11203 22298 11209
rect 22240 11200 22252 11203
rect 22060 11172 22252 11200
rect 22060 11160 22066 11172
rect 22240 11169 22252 11172
rect 22286 11169 22298 11203
rect 22240 11163 22298 11169
rect 24029 11203 24087 11209
rect 24029 11169 24041 11203
rect 24075 11200 24087 11203
rect 24075 11172 24532 11200
rect 24075 11169 24087 11172
rect 24029 11163 24087 11169
rect 13596 11104 15792 11132
rect 13596 11092 13602 11104
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 16853 11135 16911 11141
rect 16853 11132 16865 11135
rect 16724 11104 16865 11132
rect 16724 11092 16730 11104
rect 16853 11101 16865 11104
rect 16899 11101 16911 11135
rect 16853 11095 16911 11101
rect 17359 11135 17417 11141
rect 17359 11101 17371 11135
rect 17405 11132 17417 11135
rect 17405 11104 19012 11132
rect 17405 11101 17417 11104
rect 17359 11095 17417 11101
rect 12406 11076 12434 11092
rect 11112 11036 12296 11064
rect 11112 11024 11118 11036
rect 12342 11024 12348 11076
rect 12400 11036 12434 11076
rect 12400 11024 12406 11036
rect 14182 11024 14188 11076
rect 14240 11064 14246 11076
rect 14277 11067 14335 11073
rect 14277 11064 14289 11067
rect 14240 11036 14289 11064
rect 14240 11024 14246 11036
rect 14277 11033 14289 11036
rect 14323 11033 14335 11067
rect 14277 11027 14335 11033
rect 14458 11024 14464 11076
rect 14516 11064 14522 11076
rect 14516 11036 14872 11064
rect 14516 11024 14522 11036
rect 4856 10968 8156 10996
rect 4856 10956 4862 10968
rect 9122 10956 9128 11008
rect 9180 10956 9186 11008
rect 9490 10956 9496 11008
rect 9548 10996 9554 11008
rect 11238 10996 11244 11008
rect 9548 10968 11244 10996
rect 9548 10956 9554 10968
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 11422 10956 11428 11008
rect 11480 10956 11486 11008
rect 11514 10956 11520 11008
rect 11572 10996 11578 11008
rect 11701 10999 11759 11005
rect 11701 10996 11713 10999
rect 11572 10968 11713 10996
rect 11572 10956 11578 10968
rect 11701 10965 11713 10968
rect 11747 10965 11759 10999
rect 11701 10959 11759 10965
rect 14642 10956 14648 11008
rect 14700 10956 14706 11008
rect 14844 10996 14872 11036
rect 14918 11024 14924 11076
rect 14976 11024 14982 11076
rect 18984 11064 19012 11104
rect 20806 11092 20812 11144
rect 20864 11092 20870 11144
rect 20990 11092 20996 11144
rect 21048 11132 21054 11144
rect 21913 11135 21971 11141
rect 21913 11132 21925 11135
rect 21048 11104 21925 11132
rect 21048 11092 21054 11104
rect 21913 11101 21925 11104
rect 21959 11101 21971 11135
rect 21913 11095 21971 11101
rect 22419 11135 22477 11141
rect 22419 11101 22431 11135
rect 22465 11132 22477 11135
rect 22554 11132 22560 11144
rect 22465 11104 22560 11132
rect 22465 11101 22477 11104
rect 22419 11095 22477 11101
rect 22554 11092 22560 11104
rect 22612 11092 22618 11144
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 24121 11135 24179 11141
rect 24121 11101 24133 11135
rect 24167 11132 24179 11135
rect 24394 11132 24400 11144
rect 24167 11104 24400 11132
rect 24167 11101 24179 11104
rect 24121 11095 24179 11101
rect 20824 11064 20852 11092
rect 24136 11064 24164 11095
rect 24394 11092 24400 11104
rect 24452 11092 24458 11144
rect 24504 11134 24532 11172
rect 24762 11160 24768 11212
rect 24820 11200 24826 11212
rect 24820 11172 24992 11200
rect 24820 11160 24826 11172
rect 24584 11137 24642 11143
rect 24584 11134 24596 11137
rect 24504 11106 24596 11134
rect 24584 11103 24596 11106
rect 24630 11103 24642 11137
rect 24584 11097 24642 11103
rect 24854 11092 24860 11144
rect 24912 11092 24918 11144
rect 24964 11132 24992 11172
rect 26326 11160 26332 11212
rect 26384 11200 26390 11212
rect 27157 11203 27215 11209
rect 27157 11200 27169 11203
rect 26384 11172 27169 11200
rect 26384 11160 26390 11172
rect 27157 11169 27169 11172
rect 27203 11169 27215 11203
rect 27157 11163 27215 11169
rect 28902 11160 28908 11212
rect 28960 11160 28966 11212
rect 29362 11160 29368 11212
rect 29420 11160 29426 11212
rect 30282 11160 30288 11212
rect 30340 11200 30346 11212
rect 30561 11203 30619 11209
rect 30561 11200 30573 11203
rect 30340 11172 30573 11200
rect 30340 11160 30346 11172
rect 30561 11169 30573 11172
rect 30607 11169 30619 11203
rect 30561 11163 30619 11169
rect 26418 11132 26424 11144
rect 24964 11104 26424 11132
rect 26418 11092 26424 11104
rect 26476 11092 26482 11144
rect 26878 11092 26884 11144
rect 26936 11092 26942 11144
rect 28534 11092 28540 11144
rect 28592 11132 28598 11144
rect 28629 11135 28687 11141
rect 28629 11132 28641 11135
rect 28592 11104 28641 11132
rect 28592 11092 28598 11104
rect 28629 11101 28641 11104
rect 28675 11132 28687 11135
rect 29380 11132 29408 11160
rect 28675 11104 29408 11132
rect 28675 11101 28687 11104
rect 28629 11095 28687 11101
rect 18984 11036 20852 11064
rect 23308 11036 24164 11064
rect 16301 10999 16359 11005
rect 16301 10996 16313 10999
rect 14844 10968 16313 10996
rect 16301 10965 16313 10968
rect 16347 10965 16359 10999
rect 16301 10959 16359 10965
rect 17034 10956 17040 11008
rect 17092 10996 17098 11008
rect 19518 10996 19524 11008
rect 17092 10968 19524 10996
rect 17092 10956 17098 10968
rect 19518 10956 19524 10968
rect 19576 10956 19582 11008
rect 19613 10999 19671 11005
rect 19613 10965 19625 10999
rect 19659 10996 19671 10999
rect 19702 10996 19708 11008
rect 19659 10968 19708 10996
rect 19659 10965 19671 10968
rect 19613 10959 19671 10965
rect 19702 10956 19708 10968
rect 19760 10956 19766 11008
rect 21269 10999 21327 11005
rect 21269 10965 21281 10999
rect 21315 10996 21327 10999
rect 21542 10996 21548 11008
rect 21315 10968 21548 10996
rect 21315 10965 21327 10968
rect 21269 10959 21327 10965
rect 21542 10956 21548 10968
rect 21600 10956 21606 11008
rect 22278 10956 22284 11008
rect 22336 10996 22342 11008
rect 23308 10996 23336 11036
rect 28074 11024 28080 11076
rect 28132 11064 28138 11076
rect 28261 11067 28319 11073
rect 28261 11064 28273 11067
rect 28132 11036 28273 11064
rect 28132 11024 28138 11036
rect 28261 11033 28273 11036
rect 28307 11033 28319 11067
rect 28261 11027 28319 11033
rect 30006 11024 30012 11076
rect 30064 11024 30070 11076
rect 22336 10968 23336 10996
rect 22336 10956 22342 10968
rect 24026 10956 24032 11008
rect 24084 10996 24090 11008
rect 29270 10996 29276 11008
rect 24084 10968 29276 10996
rect 24084 10956 24090 10968
rect 29270 10956 29276 10968
rect 29328 10956 29334 11008
rect 552 10906 30912 10928
rect 552 10854 4193 10906
rect 4245 10854 4257 10906
rect 4309 10854 4321 10906
rect 4373 10854 4385 10906
rect 4437 10854 4449 10906
rect 4501 10854 11783 10906
rect 11835 10854 11847 10906
rect 11899 10854 11911 10906
rect 11963 10854 11975 10906
rect 12027 10854 12039 10906
rect 12091 10854 19373 10906
rect 19425 10854 19437 10906
rect 19489 10854 19501 10906
rect 19553 10854 19565 10906
rect 19617 10854 19629 10906
rect 19681 10854 26963 10906
rect 27015 10854 27027 10906
rect 27079 10854 27091 10906
rect 27143 10854 27155 10906
rect 27207 10854 27219 10906
rect 27271 10854 30912 10906
rect 552 10832 30912 10854
rect 4614 10792 4620 10804
rect 2746 10764 4620 10792
rect 937 10659 995 10665
rect 937 10625 949 10659
rect 983 10656 995 10659
rect 1302 10656 1308 10668
rect 983 10628 1308 10656
rect 983 10625 995 10628
rect 937 10619 995 10625
rect 1302 10616 1308 10628
rect 1360 10616 1366 10668
rect 1443 10659 1501 10665
rect 1443 10625 1455 10659
rect 1489 10656 1501 10659
rect 2130 10656 2136 10668
rect 1489 10628 2136 10656
rect 1489 10625 1501 10628
rect 1443 10619 1501 10625
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 2746 10588 2774 10764
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 4724 10764 11652 10792
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 3200 10628 3372 10656
rect 3200 10616 3206 10628
rect 1719 10560 2774 10588
rect 3237 10591 3295 10597
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 3237 10557 3249 10591
rect 3283 10557 3295 10591
rect 3344 10588 3372 10628
rect 3694 10616 3700 10668
rect 3752 10663 3758 10668
rect 3752 10657 3801 10663
rect 3752 10623 3755 10657
rect 3789 10623 3801 10657
rect 4724 10656 4752 10764
rect 8021 10727 8079 10733
rect 8021 10724 8033 10727
rect 6932 10696 8033 10724
rect 3752 10617 3801 10623
rect 3896 10628 4752 10656
rect 3752 10616 3758 10617
rect 3896 10588 3924 10628
rect 5534 10616 5540 10668
rect 5592 10616 5598 10668
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 6000 10659 6058 10665
rect 6000 10656 6012 10659
rect 5868 10628 6012 10656
rect 5868 10616 5874 10628
rect 6000 10625 6012 10628
rect 6046 10625 6058 10659
rect 6000 10619 6058 10625
rect 6730 10616 6736 10668
rect 6788 10656 6794 10668
rect 6932 10656 6960 10696
rect 8021 10693 8033 10696
rect 8067 10693 8079 10727
rect 9674 10724 9680 10736
rect 8021 10687 8079 10693
rect 8404 10696 9680 10724
rect 6788 10628 6960 10656
rect 7653 10659 7711 10665
rect 6788 10616 6794 10628
rect 7653 10625 7665 10659
rect 7699 10656 7711 10659
rect 7834 10656 7840 10668
rect 7699 10628 7840 10656
rect 7699 10625 7711 10628
rect 7653 10619 7711 10625
rect 7834 10616 7840 10628
rect 7892 10616 7898 10668
rect 3344 10560 3924 10588
rect 3973 10591 4031 10597
rect 3237 10551 3295 10557
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 4062 10588 4068 10600
rect 4019 10560 4068 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 1403 10455 1461 10461
rect 1403 10421 1415 10455
rect 1449 10452 1461 10455
rect 1670 10452 1676 10464
rect 1449 10424 1676 10452
rect 1449 10421 1461 10424
rect 1403 10415 1461 10421
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 2958 10412 2964 10464
rect 3016 10412 3022 10464
rect 3252 10452 3280 10551
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 5552 10588 5580 10616
rect 6086 10588 6092 10600
rect 4672 10560 5580 10588
rect 5644 10560 6092 10588
rect 4672 10548 4678 10560
rect 5353 10523 5411 10529
rect 5353 10489 5365 10523
rect 5399 10520 5411 10523
rect 5644 10520 5672 10560
rect 6086 10548 6092 10560
rect 6144 10548 6150 10600
rect 6270 10548 6276 10600
rect 6328 10548 6334 10600
rect 6914 10548 6920 10600
rect 6972 10588 6978 10600
rect 8404 10597 8432 10696
rect 9674 10684 9680 10696
rect 9732 10684 9738 10736
rect 11624 10724 11652 10764
rect 11698 10752 11704 10804
rect 11756 10752 11762 10804
rect 12986 10792 12992 10804
rect 12176 10764 12992 10792
rect 12176 10724 12204 10764
rect 12986 10752 12992 10764
rect 13044 10792 13050 10804
rect 15194 10792 15200 10804
rect 13044 10764 15200 10792
rect 13044 10752 13050 10764
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 16301 10795 16359 10801
rect 16301 10761 16313 10795
rect 16347 10792 16359 10795
rect 16390 10792 16396 10804
rect 16347 10764 16396 10792
rect 16347 10761 16359 10764
rect 16301 10755 16359 10761
rect 16390 10752 16396 10764
rect 16448 10752 16454 10804
rect 16942 10752 16948 10804
rect 17000 10792 17006 10804
rect 17862 10792 17868 10804
rect 17000 10764 17868 10792
rect 17000 10752 17006 10764
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 20530 10792 20536 10804
rect 18432 10764 20536 10792
rect 11624 10696 12204 10724
rect 12253 10727 12311 10733
rect 12253 10693 12265 10727
rect 12299 10724 12311 10727
rect 12342 10724 12348 10736
rect 12299 10696 12348 10724
rect 12299 10693 12311 10696
rect 12253 10687 12311 10693
rect 9582 10616 9588 10668
rect 9640 10616 9646 10668
rect 9858 10616 9864 10668
rect 9916 10656 9922 10668
rect 10140 10659 10198 10665
rect 10140 10656 10152 10659
rect 9916 10628 10152 10656
rect 9916 10616 9922 10628
rect 10140 10625 10152 10628
rect 10186 10625 10198 10659
rect 10140 10619 10198 10625
rect 10413 10659 10471 10665
rect 10413 10625 10425 10659
rect 10459 10656 10471 10659
rect 10870 10656 10876 10668
rect 10459 10628 10876 10656
rect 10459 10625 10471 10628
rect 10413 10619 10471 10625
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 11238 10616 11244 10668
rect 11296 10656 11302 10668
rect 12268 10656 12296 10687
rect 12342 10684 12348 10696
rect 12400 10684 12406 10736
rect 12437 10727 12495 10733
rect 12437 10693 12449 10727
rect 12483 10693 12495 10727
rect 12437 10687 12495 10693
rect 11296 10628 12296 10656
rect 11296 10616 11302 10628
rect 8389 10591 8447 10597
rect 6972 10560 8340 10588
rect 6972 10548 6978 10560
rect 5399 10492 5672 10520
rect 5399 10489 5411 10492
rect 5353 10483 5411 10489
rect 7374 10480 7380 10532
rect 7432 10520 7438 10532
rect 7837 10523 7895 10529
rect 7837 10520 7849 10523
rect 7432 10492 7849 10520
rect 7432 10480 7438 10492
rect 7837 10489 7849 10492
rect 7883 10520 7895 10523
rect 8202 10520 8208 10532
rect 7883 10492 8208 10520
rect 7883 10489 7895 10492
rect 7837 10483 7895 10489
rect 8202 10480 8208 10492
rect 8260 10480 8266 10532
rect 8312 10520 8340 10560
rect 8389 10557 8401 10591
rect 8435 10557 8447 10591
rect 8389 10551 8447 10557
rect 8938 10548 8944 10600
rect 8996 10548 9002 10600
rect 9600 10588 9628 10616
rect 9677 10591 9735 10597
rect 9677 10588 9689 10591
rect 9600 10560 9689 10588
rect 9677 10557 9689 10560
rect 9723 10557 9735 10591
rect 10004 10591 10062 10597
rect 10004 10588 10016 10591
rect 9677 10551 9735 10557
rect 9784 10560 10016 10588
rect 9217 10523 9275 10529
rect 9217 10520 9229 10523
rect 8312 10492 9229 10520
rect 9217 10489 9229 10492
rect 9263 10520 9275 10523
rect 9398 10520 9404 10532
rect 9263 10492 9404 10520
rect 9263 10489 9275 10492
rect 9217 10483 9275 10489
rect 9398 10480 9404 10492
rect 9456 10520 9462 10532
rect 9784 10520 9812 10560
rect 10004 10557 10016 10560
rect 10050 10557 10062 10591
rect 10004 10551 10062 10557
rect 10226 10548 10232 10600
rect 10284 10588 10290 10600
rect 12452 10588 12480 10687
rect 13170 10684 13176 10736
rect 13228 10684 13234 10736
rect 13354 10684 13360 10736
rect 13412 10684 13418 10736
rect 18432 10733 18460 10764
rect 20530 10752 20536 10764
rect 20588 10752 20594 10804
rect 20714 10752 20720 10804
rect 20772 10752 20778 10804
rect 22278 10792 22284 10804
rect 20916 10764 22284 10792
rect 18417 10727 18475 10733
rect 18417 10693 18429 10727
rect 18463 10693 18475 10727
rect 18417 10687 18475 10693
rect 12544 10628 12756 10656
rect 12544 10600 12572 10628
rect 10284 10560 12480 10588
rect 10284 10548 10290 10560
rect 12526 10548 12532 10600
rect 12584 10548 12590 10600
rect 12618 10548 12624 10600
rect 12676 10548 12682 10600
rect 12728 10597 12756 10628
rect 12713 10591 12771 10597
rect 12713 10557 12725 10591
rect 12759 10557 12771 10591
rect 13188 10588 13216 10684
rect 13372 10656 13400 10684
rect 14004 10659 14062 10665
rect 14004 10656 14016 10659
rect 13372 10628 14016 10656
rect 14004 10625 14016 10628
rect 14050 10625 14062 10659
rect 14004 10619 14062 10625
rect 14277 10659 14335 10665
rect 14277 10625 14289 10659
rect 14323 10656 14335 10659
rect 14642 10656 14648 10668
rect 14323 10628 14648 10656
rect 14323 10625 14335 10628
rect 14277 10619 14335 10625
rect 14642 10616 14648 10628
rect 14700 10616 14706 10668
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 16856 10659 16914 10665
rect 16856 10656 16868 10659
rect 16632 10628 16868 10656
rect 16632 10616 16638 10628
rect 16856 10625 16868 10628
rect 16902 10625 16914 10659
rect 18138 10656 18144 10668
rect 16856 10619 16914 10625
rect 17052 10628 18144 10656
rect 13357 10591 13415 10597
rect 13357 10588 13369 10591
rect 13188 10560 13369 10588
rect 12713 10551 12771 10557
rect 13357 10557 13369 10560
rect 13403 10557 13415 10591
rect 13357 10551 13415 10557
rect 13538 10548 13544 10600
rect 13596 10548 13602 10600
rect 13814 10548 13820 10600
rect 13872 10588 13878 10600
rect 15194 10588 15200 10600
rect 13872 10560 15200 10588
rect 13872 10548 13878 10560
rect 15194 10548 15200 10560
rect 15252 10548 15258 10600
rect 16393 10591 16451 10597
rect 16393 10557 16405 10591
rect 16439 10588 16451 10591
rect 17052 10588 17080 10628
rect 18138 10616 18144 10628
rect 18196 10616 18202 10668
rect 18693 10659 18751 10665
rect 18693 10625 18705 10659
rect 18739 10656 18751 10659
rect 18874 10656 18880 10668
rect 18739 10628 18880 10656
rect 18739 10625 18751 10628
rect 18693 10619 18751 10625
rect 18874 10616 18880 10628
rect 18932 10616 18938 10668
rect 19172 10641 19230 10647
rect 19172 10607 19184 10641
rect 19218 10607 19230 10641
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 20916 10665 20944 10764
rect 22278 10752 22284 10764
rect 22336 10752 22342 10804
rect 22646 10752 22652 10804
rect 22704 10792 22710 10804
rect 23109 10795 23167 10801
rect 23109 10792 23121 10795
rect 22704 10764 23121 10792
rect 22704 10752 22710 10764
rect 23109 10761 23121 10764
rect 23155 10761 23167 10795
rect 23109 10755 23167 10761
rect 23845 10795 23903 10801
rect 23845 10761 23857 10795
rect 23891 10792 23903 10795
rect 24854 10792 24860 10804
rect 23891 10764 24860 10792
rect 23891 10761 23903 10764
rect 23845 10755 23903 10761
rect 24854 10752 24860 10764
rect 24912 10752 24918 10804
rect 25130 10752 25136 10804
rect 25188 10792 25194 10804
rect 25682 10792 25688 10804
rect 25188 10764 25688 10792
rect 25188 10752 25194 10764
rect 25682 10752 25688 10764
rect 25740 10792 25746 10804
rect 29914 10792 29920 10804
rect 25740 10764 29920 10792
rect 25740 10752 25746 10764
rect 22738 10684 22744 10736
rect 22796 10684 22802 10736
rect 20901 10659 20959 10665
rect 20901 10656 20913 10659
rect 19392 10628 20913 10656
rect 19392 10616 19398 10628
rect 20901 10625 20913 10628
rect 20947 10625 20959 10659
rect 20901 10619 20959 10625
rect 21379 10641 21772 10656
rect 21379 10610 21409 10641
rect 19172 10604 19230 10607
rect 21397 10607 21409 10610
rect 21443 10628 21772 10641
rect 21443 10607 21455 10628
rect 19172 10601 19288 10604
rect 21397 10601 21455 10607
rect 19174 10600 19288 10601
rect 16439 10560 17080 10588
rect 17129 10591 17187 10597
rect 16439 10557 16451 10560
rect 16393 10551 16451 10557
rect 17129 10557 17141 10591
rect 17175 10588 17187 10591
rect 18598 10588 18604 10600
rect 17175 10560 18604 10588
rect 17175 10557 17187 10560
rect 17129 10551 17187 10557
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 19174 10576 19248 10600
rect 19242 10548 19248 10576
rect 19300 10548 19306 10600
rect 19429 10591 19487 10597
rect 19429 10557 19441 10591
rect 19475 10588 19487 10591
rect 19702 10588 19708 10600
rect 19475 10560 19708 10588
rect 19475 10557 19487 10560
rect 19429 10551 19487 10557
rect 19702 10548 19708 10560
rect 19760 10548 19766 10600
rect 21542 10548 21548 10600
rect 21600 10588 21606 10600
rect 21637 10591 21695 10597
rect 21637 10588 21649 10591
rect 21600 10560 21649 10588
rect 21600 10548 21606 10560
rect 21637 10557 21649 10560
rect 21683 10557 21695 10591
rect 21744 10588 21772 10628
rect 21818 10616 21824 10668
rect 21876 10656 21882 10668
rect 25087 10659 25145 10665
rect 21876 10628 23336 10656
rect 21876 10616 21882 10628
rect 23308 10597 23336 10628
rect 25087 10625 25099 10659
rect 25133 10656 25145 10659
rect 27065 10659 27123 10665
rect 25133 10628 25728 10656
rect 25133 10625 25145 10628
rect 25087 10619 25145 10625
rect 25700 10600 25728 10628
rect 27065 10625 27077 10659
rect 27111 10656 27123 10659
rect 28258 10656 28264 10668
rect 27111 10628 28264 10656
rect 27111 10625 27123 10628
rect 27065 10619 27123 10625
rect 28258 10616 28264 10628
rect 28316 10616 28322 10668
rect 23293 10591 23351 10597
rect 21744 10560 22692 10588
rect 21637 10551 21695 10557
rect 9456 10492 9812 10520
rect 11977 10523 12035 10529
rect 9456 10480 9462 10492
rect 11977 10489 11989 10523
rect 12023 10520 12035 10523
rect 13556 10520 13584 10548
rect 12023 10492 13584 10520
rect 12023 10489 12035 10492
rect 11977 10483 12035 10489
rect 3510 10452 3516 10464
rect 3252 10424 3516 10452
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 3703 10455 3761 10461
rect 3703 10421 3715 10455
rect 3749 10452 3761 10455
rect 5626 10452 5632 10464
rect 3749 10424 5632 10452
rect 3749 10421 3761 10424
rect 3703 10415 3761 10421
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 5994 10412 6000 10464
rect 6052 10461 6058 10464
rect 6052 10452 6061 10461
rect 6052 10424 6097 10452
rect 6052 10415 6061 10424
rect 6052 10412 6058 10415
rect 7650 10412 7656 10464
rect 7708 10452 7714 10464
rect 8573 10455 8631 10461
rect 8573 10452 8585 10455
rect 7708 10424 8585 10452
rect 7708 10412 7714 10424
rect 8573 10421 8585 10424
rect 8619 10452 8631 10455
rect 10134 10452 10140 10464
rect 8619 10424 10140 10452
rect 8619 10421 8631 10424
rect 8573 10415 8631 10421
rect 10134 10412 10140 10424
rect 10192 10412 10198 10464
rect 10870 10412 10876 10464
rect 10928 10452 10934 10464
rect 11992 10452 12020 10483
rect 22664 10464 22692 10560
rect 23293 10557 23305 10591
rect 23339 10588 23351 10591
rect 24026 10588 24032 10600
rect 23339 10560 24032 10588
rect 23339 10557 23351 10560
rect 23293 10551 23351 10557
rect 24026 10548 24032 10560
rect 24084 10548 24090 10600
rect 24581 10591 24639 10597
rect 24581 10588 24593 10591
rect 24136 10560 24593 10588
rect 24136 10464 24164 10560
rect 24581 10557 24593 10560
rect 24627 10557 24639 10591
rect 24581 10551 24639 10557
rect 25314 10548 25320 10600
rect 25372 10548 25378 10600
rect 25682 10548 25688 10600
rect 25740 10548 25746 10600
rect 26789 10591 26847 10597
rect 26789 10557 26801 10591
rect 26835 10588 26847 10591
rect 28534 10588 28540 10600
rect 26835 10560 28540 10588
rect 26835 10557 26847 10560
rect 26789 10551 26847 10557
rect 28534 10548 28540 10560
rect 28592 10548 28598 10600
rect 29104 10597 29132 10764
rect 29914 10752 29920 10764
rect 29972 10752 29978 10804
rect 30282 10684 30288 10736
rect 30340 10684 30346 10736
rect 29362 10616 29368 10668
rect 29420 10656 29426 10668
rect 30300 10656 30328 10684
rect 29420 10628 30328 10656
rect 29420 10616 29426 10628
rect 29089 10591 29147 10597
rect 29089 10557 29101 10591
rect 29135 10557 29147 10591
rect 29089 10551 29147 10557
rect 29454 10548 29460 10600
rect 29512 10588 29518 10600
rect 30101 10591 30159 10597
rect 30101 10588 30113 10591
rect 29512 10560 30113 10588
rect 29512 10548 29518 10560
rect 30101 10557 30113 10560
rect 30147 10557 30159 10591
rect 30101 10551 30159 10557
rect 26050 10480 26056 10532
rect 26108 10520 26114 10532
rect 26697 10523 26755 10529
rect 26108 10492 26372 10520
rect 26108 10480 26114 10492
rect 10928 10424 12020 10452
rect 10928 10412 10934 10424
rect 12158 10412 12164 10464
rect 12216 10452 12222 10464
rect 12526 10452 12532 10464
rect 12216 10424 12532 10452
rect 12216 10412 12222 10424
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 12894 10412 12900 10464
rect 12952 10412 12958 10464
rect 13173 10455 13231 10461
rect 13173 10421 13185 10455
rect 13219 10452 13231 10455
rect 13814 10452 13820 10464
rect 13219 10424 13820 10452
rect 13219 10421 13231 10424
rect 13173 10415 13231 10421
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 14007 10455 14065 10461
rect 14007 10452 14019 10455
rect 13964 10424 14019 10452
rect 13964 10412 13970 10424
rect 14007 10421 14019 10424
rect 14053 10421 14065 10455
rect 14007 10415 14065 10421
rect 15378 10412 15384 10464
rect 15436 10412 15442 10464
rect 16859 10455 16917 10461
rect 16859 10421 16871 10455
rect 16905 10452 16917 10455
rect 18782 10452 18788 10464
rect 16905 10424 18788 10452
rect 16905 10421 16917 10424
rect 16859 10415 16917 10421
rect 18782 10412 18788 10424
rect 18840 10412 18846 10464
rect 19150 10412 19156 10464
rect 19208 10461 19214 10464
rect 19208 10452 19217 10461
rect 21367 10455 21425 10461
rect 21367 10452 21379 10455
rect 19208 10424 21379 10452
rect 19208 10415 19217 10424
rect 21367 10421 21379 10424
rect 21413 10452 21425 10455
rect 22462 10452 22468 10464
rect 21413 10424 22468 10452
rect 21413 10421 21425 10424
rect 21367 10415 21425 10421
rect 19208 10412 19214 10415
rect 22462 10412 22468 10424
rect 22520 10412 22526 10464
rect 22646 10412 22652 10464
rect 22704 10412 22710 10464
rect 24118 10412 24124 10464
rect 24176 10412 24182 10464
rect 24486 10412 24492 10464
rect 24544 10452 24550 10464
rect 25047 10455 25105 10461
rect 25047 10452 25059 10455
rect 24544 10424 25059 10452
rect 24544 10412 24550 10424
rect 25047 10421 25059 10424
rect 25093 10452 25105 10455
rect 26234 10452 26240 10464
rect 25093 10424 26240 10452
rect 25093 10421 25105 10424
rect 25047 10415 25105 10421
rect 26234 10412 26240 10424
rect 26292 10412 26298 10464
rect 26344 10452 26372 10492
rect 26697 10489 26709 10523
rect 26743 10520 26755 10523
rect 26878 10520 26884 10532
rect 26743 10492 26884 10520
rect 26743 10489 26755 10492
rect 26697 10483 26755 10489
rect 26878 10480 26884 10492
rect 26936 10480 26942 10532
rect 29641 10523 29699 10529
rect 29641 10489 29653 10523
rect 29687 10520 29699 10523
rect 30466 10520 30472 10532
rect 29687 10492 30472 10520
rect 29687 10489 29699 10492
rect 29641 10483 29699 10489
rect 30466 10480 30472 10492
rect 30524 10480 30530 10532
rect 28169 10455 28227 10461
rect 28169 10452 28181 10455
rect 26344 10424 28181 10452
rect 28169 10421 28181 10424
rect 28215 10421 28227 10455
rect 28169 10415 28227 10421
rect 28994 10412 29000 10464
rect 29052 10452 29058 10464
rect 29181 10455 29239 10461
rect 29181 10452 29193 10455
rect 29052 10424 29193 10452
rect 29052 10412 29058 10424
rect 29181 10421 29193 10424
rect 29227 10421 29239 10455
rect 29181 10415 29239 10421
rect 29730 10412 29736 10464
rect 29788 10412 29794 10464
rect 552 10362 31072 10384
rect 552 10310 7988 10362
rect 8040 10310 8052 10362
rect 8104 10310 8116 10362
rect 8168 10310 8180 10362
rect 8232 10310 8244 10362
rect 8296 10310 15578 10362
rect 15630 10310 15642 10362
rect 15694 10310 15706 10362
rect 15758 10310 15770 10362
rect 15822 10310 15834 10362
rect 15886 10310 23168 10362
rect 23220 10310 23232 10362
rect 23284 10310 23296 10362
rect 23348 10310 23360 10362
rect 23412 10310 23424 10362
rect 23476 10310 30758 10362
rect 30810 10310 30822 10362
rect 30874 10310 30886 10362
rect 30938 10310 30950 10362
rect 31002 10310 31014 10362
rect 31066 10310 31072 10362
rect 552 10288 31072 10310
rect 1302 10248 1308 10260
rect 1044 10220 1308 10248
rect 934 10072 940 10124
rect 992 10112 998 10124
rect 1044 10121 1072 10220
rect 1302 10208 1308 10220
rect 1360 10208 1366 10260
rect 1394 10208 1400 10260
rect 1452 10248 1458 10260
rect 1495 10251 1553 10257
rect 1495 10248 1507 10251
rect 1452 10220 1507 10248
rect 1452 10208 1458 10220
rect 1495 10217 1507 10220
rect 1541 10248 1553 10251
rect 1670 10248 1676 10260
rect 1541 10220 1676 10248
rect 1541 10217 1553 10220
rect 1495 10211 1553 10217
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 3234 10208 3240 10260
rect 3292 10248 3298 10260
rect 3703 10251 3761 10257
rect 3703 10248 3715 10251
rect 3292 10220 3715 10248
rect 3292 10208 3298 10220
rect 3703 10217 3715 10220
rect 3749 10217 3761 10251
rect 3703 10211 3761 10217
rect 3878 10208 3884 10260
rect 3936 10248 3942 10260
rect 5166 10248 5172 10260
rect 3936 10220 5172 10248
rect 3936 10208 3942 10220
rect 5166 10208 5172 10220
rect 5224 10208 5230 10260
rect 6914 10208 6920 10260
rect 6972 10257 6978 10260
rect 6972 10248 6981 10257
rect 6972 10220 7017 10248
rect 6972 10211 6981 10220
rect 6972 10208 6978 10211
rect 8938 10208 8944 10260
rect 8996 10248 9002 10260
rect 8996 10220 12434 10248
rect 8996 10208 9002 10220
rect 5350 10140 5356 10192
rect 5408 10180 5414 10192
rect 6546 10180 6552 10192
rect 5408 10152 6552 10180
rect 5408 10140 5414 10152
rect 5920 10121 5948 10152
rect 6546 10140 6552 10152
rect 6604 10140 6610 10192
rect 10134 10140 10140 10192
rect 10192 10180 10198 10192
rect 11054 10180 11060 10192
rect 10192 10152 11060 10180
rect 10192 10140 10198 10152
rect 11054 10140 11060 10152
rect 11112 10140 11118 10192
rect 12406 10180 12434 10220
rect 12618 10208 12624 10260
rect 12676 10248 12682 10260
rect 16482 10248 16488 10260
rect 12676 10220 16488 10248
rect 12676 10208 12682 10220
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 17126 10208 17132 10260
rect 17184 10248 17190 10260
rect 17687 10251 17745 10257
rect 17687 10248 17699 10251
rect 17184 10220 17699 10248
rect 17184 10208 17190 10220
rect 17687 10217 17699 10220
rect 17733 10217 17745 10251
rect 17687 10211 17745 10217
rect 18782 10208 18788 10260
rect 18840 10208 18846 10260
rect 19242 10208 19248 10260
rect 19300 10208 19306 10260
rect 20898 10208 20904 10260
rect 20956 10248 20962 10260
rect 21735 10251 21793 10257
rect 21735 10248 21747 10251
rect 20956 10220 21747 10248
rect 20956 10208 20962 10220
rect 21735 10217 21747 10220
rect 21781 10248 21793 10251
rect 22002 10248 22008 10260
rect 21781 10220 22008 10248
rect 21781 10217 21793 10220
rect 21735 10211 21793 10217
rect 22002 10208 22008 10220
rect 22060 10208 22066 10260
rect 22646 10208 22652 10260
rect 22704 10248 22710 10260
rect 23109 10251 23167 10257
rect 23109 10248 23121 10251
rect 22704 10220 23121 10248
rect 22704 10208 22710 10220
rect 23109 10217 23121 10220
rect 23155 10217 23167 10251
rect 23109 10211 23167 10217
rect 24026 10208 24032 10260
rect 24084 10248 24090 10260
rect 24762 10248 24768 10260
rect 24084 10220 24768 10248
rect 24084 10208 24090 10220
rect 24762 10208 24768 10220
rect 24820 10208 24826 10260
rect 26694 10208 26700 10260
rect 26752 10248 26758 10260
rect 26878 10248 26884 10260
rect 26936 10257 26942 10260
rect 26752 10220 26884 10248
rect 26752 10208 26758 10220
rect 26878 10208 26884 10220
rect 26936 10211 26945 10257
rect 26936 10208 26942 10211
rect 29914 10208 29920 10260
rect 29972 10208 29978 10260
rect 12406 10152 12940 10180
rect 1029 10115 1087 10121
rect 1029 10112 1041 10115
rect 992 10084 1041 10112
rect 992 10072 998 10084
rect 1029 10081 1041 10084
rect 1075 10081 1087 10115
rect 1029 10075 1087 10081
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10112 5687 10115
rect 5905 10115 5963 10121
rect 5675 10084 5856 10112
rect 5675 10081 5687 10084
rect 5629 10075 5687 10081
rect 1525 10065 1583 10071
rect 1525 10031 1537 10065
rect 1571 10044 1583 10065
rect 1670 10044 1676 10056
rect 1571 10031 1676 10044
rect 1525 10025 1676 10031
rect 1550 10016 1676 10025
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 1762 10004 1768 10056
rect 1820 10004 1826 10056
rect 2958 10004 2964 10056
rect 3016 10004 3022 10056
rect 3234 10004 3240 10056
rect 3292 10004 3298 10056
rect 3694 10004 3700 10056
rect 3752 10044 3758 10056
rect 3973 10047 4031 10053
rect 3752 10016 3797 10044
rect 3752 10004 3758 10016
rect 3973 10013 3985 10047
rect 4019 10044 4031 10047
rect 4154 10044 4160 10056
rect 4019 10016 4160 10044
rect 4019 10013 4031 10016
rect 3973 10007 4031 10013
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 5353 10047 5411 10053
rect 5353 10013 5365 10047
rect 5399 10044 5411 10047
rect 5718 10044 5724 10056
rect 5399 10016 5724 10044
rect 5399 10013 5411 10016
rect 5353 10007 5411 10013
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 2976 9976 3004 10004
rect 5828 9976 5856 10084
rect 5905 10081 5917 10115
rect 5951 10081 5963 10115
rect 5905 10075 5963 10081
rect 6457 10115 6515 10121
rect 6457 10081 6469 10115
rect 6503 10112 6515 10115
rect 7282 10112 7288 10124
rect 6503 10084 7288 10112
rect 6503 10081 6515 10084
rect 6457 10075 6515 10081
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 8573 10115 8631 10121
rect 8573 10081 8585 10115
rect 8619 10112 8631 10115
rect 9401 10115 9459 10121
rect 8619 10084 9171 10112
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 5994 10004 6000 10056
rect 6052 10044 6058 10056
rect 6089 10047 6147 10053
rect 6089 10044 6101 10047
rect 6052 10016 6101 10044
rect 6052 10004 6058 10016
rect 6089 10013 6101 10016
rect 6135 10013 6147 10047
rect 6822 10044 6828 10056
rect 6089 10007 6147 10013
rect 6196 10016 6828 10044
rect 6196 9976 6224 10016
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 6963 10047 7021 10053
rect 6963 10013 6975 10047
rect 7009 10044 7021 10047
rect 7098 10044 7104 10056
rect 7009 10016 7104 10044
rect 7009 10013 7021 10016
rect 6963 10007 7021 10013
rect 7098 10004 7104 10016
rect 7156 10004 7162 10056
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10044 7251 10047
rect 7558 10044 7564 10056
rect 7239 10016 7564 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 9030 10053 9036 10056
rect 8665 10047 8723 10053
rect 8665 10013 8677 10047
rect 8711 10013 8723 10047
rect 8665 10007 8723 10013
rect 8992 10047 9036 10053
rect 8992 10013 9004 10047
rect 8992 10007 9036 10013
rect 2976 9948 3280 9976
rect 5828 9948 6224 9976
rect 3050 9868 3056 9920
rect 3108 9868 3114 9920
rect 3252 9908 3280 9948
rect 3694 9908 3700 9920
rect 3252 9880 3700 9908
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 5445 9911 5503 9917
rect 5445 9877 5457 9911
rect 5491 9908 5503 9911
rect 8478 9908 8484 9920
rect 5491 9880 8484 9908
rect 5491 9877 5503 9880
rect 5445 9871 5503 9877
rect 8478 9868 8484 9880
rect 8536 9868 8542 9920
rect 8570 9868 8576 9920
rect 8628 9908 8634 9920
rect 8680 9908 8708 10007
rect 9030 10004 9036 10007
rect 9088 10004 9094 10056
rect 9143 10055 9171 10084
rect 9401 10081 9413 10115
rect 9447 10112 9459 10115
rect 10502 10112 10508 10124
rect 9447 10084 10508 10112
rect 9447 10081 9459 10084
rect 9401 10075 9459 10081
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 10744 10084 11471 10112
rect 10744 10072 10750 10084
rect 9128 10049 9186 10055
rect 9128 10015 9140 10049
rect 9174 10015 9186 10049
rect 9128 10009 9186 10015
rect 10870 10004 10876 10056
rect 10928 10044 10934 10056
rect 11330 10053 11336 10056
rect 10965 10047 11023 10053
rect 10965 10044 10977 10047
rect 10928 10016 10977 10044
rect 10928 10004 10934 10016
rect 10965 10013 10977 10016
rect 11011 10013 11023 10047
rect 10965 10007 11023 10013
rect 11292 10047 11336 10053
rect 11292 10013 11304 10047
rect 11292 10007 11336 10013
rect 11330 10004 11336 10007
rect 11388 10004 11394 10056
rect 11443 10053 11471 10084
rect 11428 10047 11486 10053
rect 11428 10013 11440 10047
rect 11474 10013 11486 10047
rect 11428 10007 11486 10013
rect 11698 10004 11704 10056
rect 11756 10004 11762 10056
rect 12912 9920 12940 10152
rect 13262 10140 13268 10192
rect 13320 10140 13326 10192
rect 16390 10140 16396 10192
rect 16448 10140 16454 10192
rect 17310 10180 17316 10192
rect 16868 10152 17316 10180
rect 13538 10072 13544 10124
rect 13596 10072 13602 10124
rect 14366 10112 14372 10124
rect 14200 10084 14372 10112
rect 13906 10053 13912 10056
rect 13868 10047 13912 10053
rect 13868 10013 13880 10047
rect 13868 10007 13912 10013
rect 13906 10004 13912 10007
rect 13964 10004 13970 10056
rect 14047 10047 14105 10053
rect 14047 10013 14059 10047
rect 14093 10044 14105 10047
rect 14200 10044 14228 10084
rect 14366 10072 14372 10084
rect 14424 10072 14430 10124
rect 15194 10072 15200 10124
rect 15252 10112 15258 10124
rect 15933 10115 15991 10121
rect 15933 10112 15945 10115
rect 15252 10084 15945 10112
rect 15252 10072 15258 10084
rect 15933 10081 15945 10084
rect 15979 10081 15991 10115
rect 15933 10075 15991 10081
rect 16301 10115 16359 10121
rect 16301 10081 16313 10115
rect 16347 10112 16359 10115
rect 16408 10112 16436 10140
rect 16347 10084 16436 10112
rect 16347 10081 16359 10084
rect 16301 10075 16359 10081
rect 16666 10072 16672 10124
rect 16724 10072 16730 10124
rect 16868 10121 16896 10152
rect 17310 10140 17316 10152
rect 17368 10140 17374 10192
rect 18800 10180 18828 10208
rect 19978 10180 19984 10192
rect 18800 10152 19984 10180
rect 19978 10140 19984 10152
rect 20036 10140 20042 10192
rect 20717 10183 20775 10189
rect 20717 10149 20729 10183
rect 20763 10180 20775 10183
rect 20990 10180 20996 10192
rect 20763 10152 20996 10180
rect 20763 10149 20775 10152
rect 20717 10143 20775 10149
rect 20990 10140 20996 10152
rect 21048 10180 21054 10192
rect 21266 10180 21272 10192
rect 21048 10152 21272 10180
rect 21048 10140 21054 10152
rect 21266 10140 21272 10152
rect 21324 10140 21330 10192
rect 23676 10152 24256 10180
rect 16853 10115 16911 10121
rect 16853 10081 16865 10115
rect 16899 10081 16911 10115
rect 16853 10075 16911 10081
rect 17034 10072 17040 10124
rect 17092 10112 17098 10124
rect 17129 10115 17187 10121
rect 17129 10112 17141 10115
rect 17092 10084 17141 10112
rect 17092 10072 17098 10084
rect 17129 10081 17141 10084
rect 17175 10081 17187 10115
rect 20165 10115 20223 10121
rect 17129 10075 17187 10081
rect 17880 10084 18092 10112
rect 14093 10016 14228 10044
rect 14277 10047 14335 10053
rect 14093 10013 14105 10016
rect 14047 10007 14105 10013
rect 14277 10013 14289 10047
rect 14323 10044 14335 10047
rect 16684 10044 16712 10072
rect 17221 10047 17279 10053
rect 17221 10044 17233 10047
rect 14323 10016 15792 10044
rect 16684 10016 17233 10044
rect 14323 10013 14335 10016
rect 14277 10007 14335 10013
rect 15764 9985 15792 10016
rect 17221 10013 17233 10016
rect 17267 10013 17279 10047
rect 17221 10007 17279 10013
rect 17727 10047 17785 10053
rect 17727 10013 17739 10047
rect 17773 10044 17785 10047
rect 17880 10044 17908 10084
rect 18064 10056 18092 10084
rect 20165 10081 20177 10115
rect 20211 10112 20223 10115
rect 20254 10112 20260 10124
rect 20211 10084 20260 10112
rect 20211 10081 20223 10084
rect 20165 10075 20223 10081
rect 20254 10072 20260 10084
rect 20312 10112 20318 10124
rect 21082 10112 21088 10124
rect 20312 10084 21088 10112
rect 20312 10072 20318 10084
rect 21082 10072 21088 10084
rect 21140 10072 21146 10124
rect 22005 10115 22063 10121
rect 22005 10112 22017 10115
rect 21192 10084 22017 10112
rect 17773 10016 17908 10044
rect 17773 10013 17785 10016
rect 17727 10007 17785 10013
rect 17954 10004 17960 10056
rect 18012 10004 18018 10056
rect 18046 10004 18052 10056
rect 18104 10004 18110 10056
rect 15749 9979 15807 9985
rect 15749 9945 15761 9979
rect 15795 9945 15807 9979
rect 15749 9939 15807 9945
rect 16669 9979 16727 9985
rect 16669 9945 16681 9979
rect 16715 9976 16727 9979
rect 17126 9976 17132 9988
rect 16715 9948 17132 9976
rect 16715 9945 16727 9948
rect 16669 9939 16727 9945
rect 17126 9936 17132 9948
rect 17184 9936 17190 9988
rect 19981 9979 20039 9985
rect 19981 9945 19993 9979
rect 20027 9976 20039 9979
rect 21192 9976 21220 10084
rect 22005 10081 22017 10084
rect 22051 10081 22063 10115
rect 22005 10075 22063 10081
rect 21266 10004 21272 10056
rect 21324 10004 21330 10056
rect 21726 10004 21732 10056
rect 21784 10004 21790 10056
rect 21910 10004 21916 10056
rect 21968 10044 21974 10056
rect 23676 10044 23704 10152
rect 23750 10072 23756 10124
rect 23808 10112 23814 10124
rect 24029 10115 24087 10121
rect 24029 10112 24041 10115
rect 23808 10084 24041 10112
rect 23808 10072 23814 10084
rect 24029 10081 24041 10084
rect 24075 10081 24087 10115
rect 24228 10112 24256 10152
rect 24486 10121 24492 10124
rect 24448 10115 24492 10121
rect 24448 10112 24460 10115
rect 24228 10084 24460 10112
rect 24029 10075 24087 10081
rect 24448 10081 24460 10084
rect 24448 10075 24492 10081
rect 24486 10072 24492 10075
rect 24544 10072 24550 10124
rect 24946 10112 24952 10124
rect 24599 10084 24952 10112
rect 24118 10044 24124 10056
rect 21968 10016 23704 10044
rect 23768 10016 24124 10044
rect 21968 10004 21974 10016
rect 20027 9948 21220 9976
rect 20027 9945 20039 9948
rect 19981 9939 20039 9945
rect 9490 9908 9496 9920
rect 8628 9880 9496 9908
rect 8628 9868 8634 9880
rect 9490 9868 9496 9880
rect 9548 9868 9554 9920
rect 10689 9911 10747 9917
rect 10689 9877 10701 9911
rect 10735 9908 10747 9911
rect 11146 9908 11152 9920
rect 10735 9880 11152 9908
rect 10735 9877 10747 9880
rect 10689 9871 10747 9877
rect 11146 9868 11152 9880
rect 11204 9868 11210 9920
rect 12342 9868 12348 9920
rect 12400 9908 12406 9920
rect 12805 9911 12863 9917
rect 12805 9908 12817 9911
rect 12400 9880 12817 9908
rect 12400 9868 12406 9880
rect 12805 9877 12817 9880
rect 12851 9877 12863 9911
rect 12805 9871 12863 9877
rect 12894 9868 12900 9920
rect 12952 9908 12958 9920
rect 13357 9911 13415 9917
rect 13357 9908 13369 9911
rect 12952 9880 13369 9908
rect 12952 9868 12958 9880
rect 13357 9877 13369 9880
rect 13403 9877 13415 9911
rect 13357 9871 13415 9877
rect 15286 9868 15292 9920
rect 15344 9908 15350 9920
rect 15381 9911 15439 9917
rect 15381 9908 15393 9911
rect 15344 9880 15393 9908
rect 15344 9868 15350 9880
rect 15381 9877 15393 9880
rect 15427 9877 15439 9911
rect 15381 9871 15439 9877
rect 15470 9868 15476 9920
rect 15528 9908 15534 9920
rect 16117 9911 16175 9917
rect 16117 9908 16129 9911
rect 15528 9880 16129 9908
rect 15528 9868 15534 9880
rect 16117 9877 16129 9880
rect 16163 9877 16175 9911
rect 16117 9871 16175 9877
rect 16945 9911 17003 9917
rect 16945 9877 16957 9911
rect 16991 9908 17003 9911
rect 17954 9908 17960 9920
rect 16991 9880 17960 9908
rect 16991 9877 17003 9880
rect 16945 9871 17003 9877
rect 17954 9868 17960 9880
rect 18012 9868 18018 9920
rect 20990 9868 20996 9920
rect 21048 9868 21054 9920
rect 21284 9908 21312 10004
rect 23768 9908 23796 10016
rect 24118 10004 24124 10016
rect 24176 10004 24182 10056
rect 24599 10053 24627 10084
rect 24946 10072 24952 10084
rect 25004 10072 25010 10124
rect 26237 10115 26295 10121
rect 26237 10081 26249 10115
rect 26283 10112 26295 10115
rect 28629 10115 28687 10121
rect 26283 10084 26924 10112
rect 26283 10081 26295 10084
rect 26237 10075 26295 10081
rect 24584 10047 24642 10053
rect 24584 10013 24596 10047
rect 24630 10013 24642 10047
rect 24584 10007 24642 10013
rect 24670 10004 24676 10056
rect 24728 10044 24734 10056
rect 24857 10047 24915 10053
rect 24857 10044 24869 10047
rect 24728 10016 24869 10044
rect 24728 10004 24734 10016
rect 24857 10013 24869 10016
rect 24903 10013 24915 10047
rect 24857 10007 24915 10013
rect 26418 10004 26424 10056
rect 26476 10004 26482 10056
rect 26896 10053 26924 10084
rect 28629 10081 28641 10115
rect 28675 10112 28687 10115
rect 29178 10112 29184 10124
rect 28675 10084 29184 10112
rect 28675 10081 28687 10084
rect 28629 10075 28687 10081
rect 29178 10072 29184 10084
rect 29236 10072 29242 10124
rect 29932 10112 29960 10208
rect 30561 10115 30619 10121
rect 30561 10112 30573 10115
rect 29932 10084 30573 10112
rect 30561 10081 30573 10084
rect 30607 10081 30619 10115
rect 30561 10075 30619 10081
rect 26884 10047 26942 10053
rect 26884 10013 26896 10047
rect 26930 10013 26942 10047
rect 26884 10007 26942 10013
rect 27157 10047 27215 10053
rect 27157 10013 27169 10047
rect 27203 10044 27215 10047
rect 28258 10044 28264 10056
rect 27203 10016 28264 10044
rect 27203 10013 27215 10016
rect 27157 10007 27215 10013
rect 28258 10004 28264 10016
rect 28316 10004 28322 10056
rect 28810 10004 28816 10056
rect 28868 10044 28874 10056
rect 28905 10047 28963 10053
rect 28905 10044 28917 10047
rect 28868 10016 28917 10044
rect 28868 10004 28874 10016
rect 28905 10013 28917 10016
rect 28951 10013 28963 10047
rect 28905 10007 28963 10013
rect 21284 9880 23796 9908
rect 23845 9911 23903 9917
rect 23845 9877 23857 9911
rect 23891 9908 23903 9911
rect 24670 9908 24676 9920
rect 23891 9880 24676 9908
rect 23891 9877 23903 9880
rect 23845 9871 23903 9877
rect 24670 9868 24676 9880
rect 24728 9868 24734 9920
rect 28442 9868 28448 9920
rect 28500 9868 28506 9920
rect 30006 9868 30012 9920
rect 30064 9868 30070 9920
rect 30098 9868 30104 9920
rect 30156 9908 30162 9920
rect 30377 9911 30435 9917
rect 30377 9908 30389 9911
rect 30156 9880 30389 9908
rect 30156 9868 30162 9880
rect 30377 9877 30389 9880
rect 30423 9877 30435 9911
rect 30377 9871 30435 9877
rect 552 9818 30912 9840
rect 552 9766 4193 9818
rect 4245 9766 4257 9818
rect 4309 9766 4321 9818
rect 4373 9766 4385 9818
rect 4437 9766 4449 9818
rect 4501 9766 11783 9818
rect 11835 9766 11847 9818
rect 11899 9766 11911 9818
rect 11963 9766 11975 9818
rect 12027 9766 12039 9818
rect 12091 9766 19373 9818
rect 19425 9766 19437 9818
rect 19489 9766 19501 9818
rect 19553 9766 19565 9818
rect 19617 9766 19629 9818
rect 19681 9766 26963 9818
rect 27015 9766 27027 9818
rect 27079 9766 27091 9818
rect 27143 9766 27155 9818
rect 27207 9766 27219 9818
rect 27271 9766 30912 9818
rect 552 9744 30912 9766
rect 1118 9664 1124 9716
rect 1176 9704 1182 9716
rect 1762 9704 1768 9716
rect 1176 9676 1768 9704
rect 1176 9664 1182 9676
rect 1762 9664 1768 9676
rect 1820 9664 1826 9716
rect 1854 9664 1860 9716
rect 1912 9704 1918 9716
rect 5442 9704 5448 9716
rect 1912 9676 5448 9704
rect 1912 9664 1918 9676
rect 5442 9664 5448 9676
rect 5500 9664 5506 9716
rect 5810 9704 5816 9716
rect 5736 9676 5816 9704
rect 5353 9639 5411 9645
rect 5353 9605 5365 9639
rect 5399 9636 5411 9639
rect 5736 9636 5764 9676
rect 5810 9664 5816 9676
rect 5868 9664 5874 9716
rect 7282 9704 7288 9716
rect 6104 9676 7288 9704
rect 5399 9608 5764 9636
rect 5399 9605 5411 9608
rect 5353 9599 5411 9605
rect 934 9528 940 9580
rect 992 9528 998 9580
rect 1458 9559 2360 9568
rect 1433 9553 2360 9559
rect 1433 9519 1445 9553
rect 1479 9540 2360 9553
rect 1479 9519 1491 9540
rect 1433 9513 1491 9519
rect 1578 9460 1584 9512
rect 1636 9500 1642 9512
rect 1673 9503 1731 9509
rect 1673 9500 1685 9503
rect 1636 9472 1685 9500
rect 1636 9460 1642 9472
rect 1673 9469 1685 9472
rect 1719 9469 1731 9503
rect 1673 9463 1731 9469
rect 1394 9324 1400 9376
rect 1452 9373 1458 9376
rect 1452 9327 1461 9373
rect 2332 9364 2360 9540
rect 3050 9528 3056 9580
rect 3108 9568 3114 9580
rect 3792 9571 3850 9577
rect 3792 9568 3804 9571
rect 3108 9540 3804 9568
rect 3108 9528 3114 9540
rect 3792 9537 3804 9540
rect 3838 9537 3850 9571
rect 3792 9531 3850 9537
rect 3878 9528 3884 9580
rect 3936 9568 3942 9580
rect 4706 9568 4712 9580
rect 3936 9540 4712 9568
rect 3936 9528 3942 9540
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 6104 9577 6132 9676
rect 7282 9664 7288 9676
rect 7340 9664 7346 9716
rect 8478 9664 8484 9716
rect 8536 9704 8542 9716
rect 8754 9704 8760 9716
rect 8536 9676 8760 9704
rect 8536 9664 8542 9676
rect 8754 9664 8760 9676
rect 8812 9664 8818 9716
rect 10686 9664 10692 9716
rect 10744 9664 10750 9716
rect 10962 9664 10968 9716
rect 11020 9704 11026 9716
rect 11698 9704 11704 9716
rect 11020 9676 11704 9704
rect 11020 9664 11026 9676
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 11882 9664 11888 9716
rect 11940 9704 11946 9716
rect 17218 9704 17224 9716
rect 11940 9676 12388 9704
rect 11940 9664 11946 9676
rect 10597 9639 10655 9645
rect 10597 9605 10609 9639
rect 10643 9636 10655 9639
rect 10704 9636 10732 9664
rect 10643 9608 10732 9636
rect 12360 9636 12388 9676
rect 16316 9676 17224 9704
rect 13173 9639 13231 9645
rect 13173 9636 13185 9639
rect 12360 9608 13185 9636
rect 10643 9605 10655 9608
rect 10597 9599 10655 9605
rect 13173 9605 13185 9608
rect 13219 9605 13231 9639
rect 13173 9599 13231 9605
rect 6089 9571 6147 9577
rect 5316 9540 6040 9568
rect 5316 9528 5322 9540
rect 3234 9460 3240 9512
rect 3292 9500 3298 9512
rect 3329 9503 3387 9509
rect 3329 9500 3341 9503
rect 3292 9472 3341 9500
rect 3292 9460 3298 9472
rect 3329 9469 3341 9472
rect 3375 9469 3387 9503
rect 3329 9463 3387 9469
rect 3602 9460 3608 9512
rect 3660 9500 3666 9512
rect 6012 9509 6040 9540
rect 6089 9537 6101 9571
rect 6135 9537 6147 9571
rect 6089 9531 6147 9537
rect 6546 9528 6552 9580
rect 6604 9568 6610 9580
rect 6604 9540 6649 9568
rect 6604 9528 6610 9540
rect 8386 9528 8392 9580
rect 8444 9528 8450 9580
rect 8570 9528 8576 9580
rect 8628 9528 8634 9580
rect 9079 9571 9137 9577
rect 9079 9537 9091 9571
rect 9125 9568 9137 9571
rect 9125 9540 9444 9568
rect 9125 9537 9137 9540
rect 9079 9531 9137 9537
rect 4065 9503 4123 9509
rect 4065 9500 4077 9503
rect 3660 9472 4077 9500
rect 3660 9460 3666 9472
rect 4065 9469 4077 9472
rect 4111 9469 4123 9503
rect 5721 9503 5779 9509
rect 5721 9500 5733 9503
rect 4065 9463 4123 9469
rect 4724 9472 5733 9500
rect 2746 9404 3096 9432
rect 2746 9364 2774 9404
rect 2332 9336 2774 9364
rect 1452 9324 1458 9327
rect 2958 9324 2964 9376
rect 3016 9324 3022 9376
rect 3068 9364 3096 9404
rect 4724 9376 4752 9472
rect 5721 9469 5733 9472
rect 5767 9500 5779 9503
rect 5997 9503 6055 9509
rect 5767 9472 5948 9500
rect 5767 9469 5779 9472
rect 5721 9463 5779 9469
rect 4982 9392 4988 9444
rect 5040 9432 5046 9444
rect 5040 9404 5856 9432
rect 5040 9392 5046 9404
rect 3694 9364 3700 9376
rect 3068 9336 3700 9364
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 3795 9367 3853 9373
rect 3795 9333 3807 9367
rect 3841 9364 3853 9367
rect 3970 9364 3976 9376
rect 3841 9336 3976 9364
rect 3841 9333 3853 9336
rect 3795 9327 3853 9333
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 4706 9324 4712 9376
rect 4764 9324 4770 9376
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 5626 9364 5632 9376
rect 5583 9336 5632 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 5828 9373 5856 9404
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9333 5871 9367
rect 5920 9364 5948 9472
rect 5997 9469 6009 9503
rect 6043 9500 6055 9503
rect 6730 9500 6736 9512
rect 6043 9472 6736 9500
rect 6043 9469 6055 9472
rect 5997 9463 6055 9469
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9496 6883 9503
rect 7024 9500 7236 9516
rect 8404 9500 8432 9528
rect 9416 9512 9444 9540
rect 10778 9528 10784 9580
rect 10836 9528 10842 9580
rect 11108 9571 11166 9577
rect 11108 9537 11120 9571
rect 11154 9568 11166 9571
rect 11154 9537 11192 9568
rect 11108 9531 11192 9537
rect 6932 9496 8432 9500
rect 6871 9488 8432 9496
rect 6871 9472 7052 9488
rect 7208 9472 8432 9488
rect 6871 9469 6960 9472
rect 6825 9468 6960 9469
rect 6825 9463 6883 9468
rect 9306 9460 9312 9512
rect 9364 9460 9370 9512
rect 9398 9460 9404 9512
rect 9456 9460 9462 9512
rect 11164 9500 11192 9531
rect 11238 9528 11244 9580
rect 11296 9528 11302 9580
rect 11330 9528 11336 9580
rect 11388 9568 11394 9580
rect 13078 9568 13084 9580
rect 11388 9540 13084 9568
rect 11388 9528 11394 9540
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 13538 9528 13544 9580
rect 13596 9528 13602 9580
rect 13814 9528 13820 9580
rect 13872 9528 13878 9580
rect 14047 9571 14105 9577
rect 14047 9537 14059 9571
rect 14093 9568 14105 9571
rect 15010 9568 15016 9580
rect 14093 9540 15016 9568
rect 14093 9537 14105 9540
rect 14047 9531 14105 9537
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 11348 9500 11376 9528
rect 11164 9472 11376 9500
rect 11514 9460 11520 9512
rect 11572 9460 11578 9512
rect 11606 9460 11612 9512
rect 11664 9500 11670 9512
rect 12989 9503 13047 9509
rect 12989 9500 13001 9503
rect 11664 9472 13001 9500
rect 11664 9460 11670 9472
rect 12989 9469 13001 9472
rect 13035 9469 13047 9503
rect 13832 9500 13860 9528
rect 16316 9509 16344 9676
rect 17218 9664 17224 9676
rect 17276 9704 17282 9716
rect 17586 9704 17592 9716
rect 17276 9676 17592 9704
rect 17276 9664 17282 9676
rect 17586 9664 17592 9676
rect 17644 9664 17650 9716
rect 18046 9664 18052 9716
rect 18104 9704 18110 9716
rect 18233 9707 18291 9713
rect 18233 9704 18245 9707
rect 18104 9676 18245 9704
rect 18104 9664 18110 9676
rect 18233 9673 18245 9676
rect 18279 9673 18291 9707
rect 18233 9667 18291 9673
rect 18598 9664 18604 9716
rect 18656 9704 18662 9716
rect 24026 9704 24032 9716
rect 18656 9676 24032 9704
rect 18656 9664 18662 9676
rect 24026 9664 24032 9676
rect 24084 9664 24090 9716
rect 24118 9664 24124 9716
rect 24176 9704 24182 9716
rect 24176 9676 25268 9704
rect 24176 9664 24182 9676
rect 22554 9596 22560 9648
rect 22612 9636 22618 9648
rect 22741 9639 22799 9645
rect 22741 9636 22753 9639
rect 22612 9608 22753 9636
rect 22612 9596 22618 9608
rect 22741 9605 22753 9608
rect 22787 9605 22799 9639
rect 22741 9599 22799 9605
rect 19242 9575 19248 9580
rect 16899 9569 16957 9575
rect 16899 9535 16911 9569
rect 16945 9535 16957 9569
rect 16899 9529 16957 9535
rect 19199 9569 19248 9575
rect 19199 9535 19211 9569
rect 19245 9535 19248 9569
rect 19199 9529 19248 9535
rect 16758 9509 16764 9512
rect 14277 9503 14335 9509
rect 14277 9500 14289 9503
rect 13832 9472 14289 9500
rect 12989 9463 13047 9469
rect 14277 9469 14289 9472
rect 14323 9469 14335 9503
rect 14277 9463 14335 9469
rect 16301 9503 16359 9509
rect 16301 9469 16313 9503
rect 16347 9469 16359 9503
rect 16301 9463 16359 9469
rect 16393 9503 16451 9509
rect 16393 9469 16405 9503
rect 16439 9469 16451 9503
rect 16393 9463 16451 9469
rect 16720 9503 16764 9509
rect 16720 9469 16732 9503
rect 16720 9463 16764 9469
rect 16025 9435 16083 9441
rect 16025 9401 16037 9435
rect 16071 9432 16083 9435
rect 16071 9404 16344 9432
rect 16071 9401 16083 9404
rect 16025 9395 16083 9401
rect 16316 9376 16344 9404
rect 6454 9364 6460 9376
rect 5920 9336 6460 9364
rect 5813 9327 5871 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6555 9367 6613 9373
rect 6555 9333 6567 9367
rect 6601 9364 6613 9367
rect 6914 9364 6920 9376
rect 6601 9336 6920 9364
rect 6601 9333 6613 9336
rect 6555 9327 6613 9333
rect 6914 9324 6920 9336
rect 6972 9364 6978 9376
rect 7742 9364 7748 9376
rect 6972 9336 7748 9364
rect 6972 9324 6978 9336
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 8113 9367 8171 9373
rect 8113 9333 8125 9367
rect 8159 9364 8171 9367
rect 8938 9364 8944 9376
rect 8159 9336 8944 9364
rect 8159 9333 8171 9336
rect 8113 9327 8171 9333
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 9030 9324 9036 9376
rect 9088 9373 9094 9376
rect 9088 9364 9097 9373
rect 9582 9364 9588 9376
rect 9088 9336 9588 9364
rect 9088 9327 9097 9336
rect 9088 9324 9094 9327
rect 9582 9324 9588 9336
rect 9640 9364 9646 9376
rect 10778 9364 10784 9376
rect 9640 9336 10784 9364
rect 9640 9324 9646 9336
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 12621 9367 12679 9373
rect 12621 9364 12633 9367
rect 12492 9336 12633 9364
rect 12492 9324 12498 9336
rect 12621 9333 12633 9336
rect 12667 9333 12679 9367
rect 12621 9327 12679 9333
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14007 9367 14065 9373
rect 14007 9364 14019 9367
rect 13964 9336 14019 9364
rect 13964 9324 13970 9336
rect 14007 9333 14019 9336
rect 14053 9333 14065 9367
rect 14007 9327 14065 9333
rect 15010 9324 15016 9376
rect 15068 9364 15074 9376
rect 15381 9367 15439 9373
rect 15381 9364 15393 9367
rect 15068 9336 15393 9364
rect 15068 9324 15074 9336
rect 15381 9333 15393 9336
rect 15427 9333 15439 9367
rect 15381 9327 15439 9333
rect 16114 9324 16120 9376
rect 16172 9324 16178 9376
rect 16298 9324 16304 9376
rect 16356 9324 16362 9376
rect 16408 9364 16436 9463
rect 16758 9460 16764 9463
rect 16816 9460 16822 9512
rect 16914 9500 16942 9529
rect 19242 9528 19248 9529
rect 19300 9528 19306 9580
rect 19426 9528 19432 9580
rect 19484 9528 19490 9580
rect 20806 9528 20812 9580
rect 20864 9528 20870 9580
rect 21726 9568 21732 9580
rect 21379 9553 21732 9568
rect 21379 9522 21409 9553
rect 21397 9519 21409 9522
rect 21443 9540 21732 9553
rect 21443 9519 21455 9540
rect 21726 9528 21732 9540
rect 21784 9528 21790 9580
rect 23768 9540 23980 9568
rect 21397 9513 21455 9519
rect 23768 9512 23796 9540
rect 17034 9500 17040 9512
rect 16914 9472 17040 9500
rect 17034 9460 17040 9472
rect 17092 9460 17098 9512
rect 17126 9460 17132 9512
rect 17184 9460 17190 9512
rect 18690 9460 18696 9512
rect 18748 9500 18754 9512
rect 20901 9503 20959 9509
rect 20901 9500 20913 9503
rect 18748 9472 20913 9500
rect 18748 9460 18754 9472
rect 20901 9469 20913 9472
rect 20947 9500 20959 9503
rect 20990 9500 20996 9512
rect 20947 9472 20996 9500
rect 20947 9469 20959 9472
rect 20901 9463 20959 9469
rect 20990 9460 20996 9472
rect 21048 9460 21054 9512
rect 21634 9460 21640 9512
rect 21692 9460 21698 9512
rect 21910 9460 21916 9512
rect 21968 9500 21974 9512
rect 23569 9503 23627 9509
rect 23569 9500 23581 9503
rect 21968 9472 23581 9500
rect 21968 9460 21974 9472
rect 23569 9469 23581 9472
rect 23615 9500 23627 9503
rect 23750 9500 23756 9512
rect 23615 9472 23756 9500
rect 23615 9469 23627 9472
rect 23569 9463 23627 9469
rect 23750 9460 23756 9472
rect 23808 9460 23814 9512
rect 23845 9503 23903 9509
rect 23845 9469 23857 9503
rect 23891 9469 23903 9503
rect 23952 9500 23980 9540
rect 24118 9528 24124 9580
rect 24176 9568 24182 9580
rect 24308 9571 24366 9577
rect 24308 9568 24320 9571
rect 24176 9540 24320 9568
rect 24176 9528 24182 9540
rect 24308 9537 24320 9540
rect 24354 9537 24366 9571
rect 25240 9568 25268 9676
rect 25682 9664 25688 9716
rect 25740 9664 25746 9716
rect 28258 9664 28264 9716
rect 28316 9664 28322 9716
rect 28810 9636 28816 9648
rect 27448 9608 28816 9636
rect 26053 9571 26111 9577
rect 26053 9568 26065 9571
rect 25240 9540 26065 9568
rect 24308 9531 24366 9537
rect 26053 9537 26065 9540
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 26234 9528 26240 9580
rect 26292 9568 26298 9580
rect 26380 9571 26438 9577
rect 26380 9568 26392 9571
rect 26292 9540 26392 9568
rect 26292 9528 26298 9540
rect 26380 9537 26392 9540
rect 26426 9537 26438 9571
rect 26380 9531 26438 9537
rect 26516 9569 26574 9575
rect 26516 9535 26528 9569
rect 26562 9535 26574 9569
rect 26516 9529 26574 9535
rect 24486 9500 24492 9512
rect 23952 9472 24492 9500
rect 23845 9463 23903 9469
rect 23860 9432 23888 9463
rect 24486 9460 24492 9472
rect 24544 9460 24550 9512
rect 24581 9503 24639 9509
rect 24581 9469 24593 9503
rect 24627 9500 24639 9503
rect 25682 9500 25688 9512
rect 24627 9472 25688 9500
rect 24627 9469 24639 9472
rect 24581 9463 24639 9469
rect 25682 9460 25688 9472
rect 25740 9460 25746 9512
rect 25884 9496 26472 9500
rect 26531 9496 26559 9529
rect 26694 9528 26700 9580
rect 26752 9568 26758 9580
rect 27448 9568 27476 9608
rect 28810 9596 28816 9608
rect 28868 9636 28874 9648
rect 29730 9636 29736 9648
rect 28868 9608 29736 9636
rect 28868 9596 28874 9608
rect 28994 9568 29000 9580
rect 26752 9540 27476 9568
rect 28460 9540 29000 9568
rect 26752 9528 26758 9540
rect 25884 9472 26559 9496
rect 25884 9444 25912 9472
rect 26444 9468 26559 9472
rect 26786 9460 26792 9512
rect 26844 9460 26850 9512
rect 28460 9509 28488 9540
rect 28994 9528 29000 9540
rect 29052 9528 29058 9580
rect 28445 9503 28503 9509
rect 28445 9500 28457 9503
rect 27448 9472 28457 9500
rect 23934 9432 23940 9444
rect 23032 9404 23796 9432
rect 23860 9404 23940 9432
rect 23032 9376 23060 9404
rect 16666 9364 16672 9376
rect 16408 9336 16672 9364
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 16850 9324 16856 9376
rect 16908 9364 16914 9376
rect 17586 9364 17592 9376
rect 16908 9336 17592 9364
rect 16908 9324 16914 9336
rect 17586 9324 17592 9336
rect 17644 9324 17650 9376
rect 17770 9324 17776 9376
rect 17828 9364 17834 9376
rect 19058 9364 19064 9376
rect 17828 9336 19064 9364
rect 17828 9324 17834 9336
rect 19058 9324 19064 9336
rect 19116 9364 19122 9376
rect 19159 9367 19217 9373
rect 19159 9364 19171 9367
rect 19116 9336 19171 9364
rect 19116 9324 19122 9336
rect 19159 9333 19171 9336
rect 19205 9364 19217 9367
rect 21367 9367 21425 9373
rect 21367 9364 21379 9367
rect 19205 9336 21379 9364
rect 19205 9333 19217 9336
rect 19159 9327 19217 9333
rect 21367 9333 21379 9336
rect 21413 9364 21425 9367
rect 23014 9364 23020 9376
rect 21413 9336 23020 9364
rect 21413 9333 21425 9336
rect 21367 9327 21425 9333
rect 23014 9324 23020 9336
rect 23072 9324 23078 9376
rect 23385 9367 23443 9373
rect 23385 9333 23397 9367
rect 23431 9364 23443 9367
rect 23658 9364 23664 9376
rect 23431 9336 23664 9364
rect 23431 9333 23443 9336
rect 23385 9327 23443 9333
rect 23658 9324 23664 9336
rect 23716 9324 23722 9376
rect 23768 9364 23796 9404
rect 23934 9392 23940 9404
rect 23992 9392 23998 9444
rect 25866 9392 25872 9444
rect 25924 9392 25930 9444
rect 24210 9364 24216 9376
rect 23768 9336 24216 9364
rect 24210 9324 24216 9336
rect 24268 9364 24274 9376
rect 24311 9367 24369 9373
rect 24311 9364 24323 9367
rect 24268 9336 24323 9364
rect 24268 9324 24274 9336
rect 24311 9333 24323 9336
rect 24357 9333 24369 9367
rect 24311 9327 24369 9333
rect 24486 9324 24492 9376
rect 24544 9364 24550 9376
rect 27448 9364 27476 9472
rect 28445 9469 28457 9472
rect 28491 9469 28503 9503
rect 28445 9463 28503 9469
rect 28721 9503 28779 9509
rect 28721 9469 28733 9503
rect 28767 9500 28779 9503
rect 29104 9500 29132 9608
rect 29730 9596 29736 9608
rect 29788 9596 29794 9648
rect 29178 9500 29184 9512
rect 28767 9472 29184 9500
rect 28767 9469 28779 9472
rect 28721 9463 28779 9469
rect 29178 9460 29184 9472
rect 29236 9460 29242 9512
rect 30466 9460 30472 9512
rect 30524 9460 30530 9512
rect 24544 9336 27476 9364
rect 24544 9324 24550 9336
rect 27890 9324 27896 9376
rect 27948 9324 27954 9376
rect 28534 9324 28540 9376
rect 28592 9324 28598 9376
rect 30282 9324 30288 9376
rect 30340 9324 30346 9376
rect 552 9274 31072 9296
rect 552 9222 7988 9274
rect 8040 9222 8052 9274
rect 8104 9222 8116 9274
rect 8168 9222 8180 9274
rect 8232 9222 8244 9274
rect 8296 9222 15578 9274
rect 15630 9222 15642 9274
rect 15694 9222 15706 9274
rect 15758 9222 15770 9274
rect 15822 9222 15834 9274
rect 15886 9222 23168 9274
rect 23220 9222 23232 9274
rect 23284 9222 23296 9274
rect 23348 9222 23360 9274
rect 23412 9222 23424 9274
rect 23476 9222 30758 9274
rect 30810 9222 30822 9274
rect 30874 9222 30886 9274
rect 30938 9222 30950 9274
rect 31002 9222 31014 9274
rect 31066 9222 31072 9274
rect 552 9200 31072 9222
rect 2958 9120 2964 9172
rect 3016 9120 3022 9172
rect 3703 9163 3761 9169
rect 3703 9129 3715 9163
rect 3749 9160 3761 9163
rect 3970 9160 3976 9172
rect 3749 9132 3976 9160
rect 3749 9129 3761 9132
rect 3703 9123 3761 9129
rect 3970 9120 3976 9132
rect 4028 9120 4034 9172
rect 5276 9132 6040 9160
rect 2976 9024 3004 9120
rect 5276 9104 5304 9132
rect 5258 9052 5264 9104
rect 5316 9052 5322 9104
rect 5353 9095 5411 9101
rect 5353 9061 5365 9095
rect 5399 9092 5411 9095
rect 5902 9092 5908 9104
rect 5399 9064 5908 9092
rect 5399 9061 5411 9064
rect 5353 9055 5411 9061
rect 5902 9052 5908 9064
rect 5960 9052 5966 9104
rect 6012 9092 6040 9132
rect 6730 9120 6736 9172
rect 6788 9160 6794 9172
rect 7190 9160 7196 9172
rect 6788 9132 7196 9160
rect 6788 9120 6794 9132
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 7285 9163 7343 9169
rect 7285 9129 7297 9163
rect 7331 9160 7343 9163
rect 7331 9132 7604 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 6012 9064 7328 9092
rect 6012 9033 6040 9064
rect 7300 9036 7328 9064
rect 5629 9027 5687 9033
rect 1688 8996 2774 9024
rect 2976 8996 3372 9024
rect 1525 8977 1583 8983
rect 842 8916 848 8968
rect 900 8956 906 8968
rect 1394 8965 1400 8968
rect 1029 8959 1087 8965
rect 1029 8956 1041 8959
rect 900 8928 1041 8956
rect 900 8916 906 8928
rect 1029 8925 1041 8928
rect 1075 8925 1087 8959
rect 1029 8919 1087 8925
rect 1356 8959 1400 8965
rect 1356 8925 1368 8959
rect 1356 8919 1400 8925
rect 1394 8916 1400 8919
rect 1452 8916 1458 8968
rect 1525 8943 1537 8977
rect 1571 8956 1583 8977
rect 1688 8956 1716 8996
rect 1571 8943 1716 8956
rect 1525 8937 1716 8943
rect 1550 8928 1716 8937
rect 1762 8916 1768 8968
rect 1820 8916 1826 8968
rect 934 8780 940 8832
rect 992 8820 998 8832
rect 2406 8820 2412 8832
rect 992 8792 2412 8820
rect 992 8780 998 8792
rect 2406 8780 2412 8792
rect 2464 8780 2470 8832
rect 2746 8820 2774 8996
rect 3142 8916 3148 8968
rect 3200 8916 3206 8968
rect 3234 8916 3240 8968
rect 3292 8916 3298 8968
rect 3344 8956 3372 8996
rect 5629 8993 5641 9027
rect 5675 9024 5687 9027
rect 5997 9027 6055 9033
rect 5675 9008 5907 9024
rect 5675 8996 5948 9008
rect 5675 8993 5687 8996
rect 5629 8987 5687 8993
rect 3700 8977 3758 8983
rect 5879 8980 5948 8996
rect 5997 8993 6009 9027
rect 6043 8993 6055 9027
rect 5997 8987 6055 8993
rect 6178 8984 6184 9036
rect 6236 9024 6242 9036
rect 6362 9024 6368 9036
rect 6236 8996 6368 9024
rect 6236 8984 6242 8996
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 6454 8984 6460 9036
rect 6512 9024 6518 9036
rect 6641 9028 6699 9033
rect 6567 9027 6699 9028
rect 6567 9024 6653 9027
rect 6512 9000 6653 9024
rect 6512 8996 6595 9000
rect 6512 8984 6518 8996
rect 6641 8993 6653 9000
rect 6687 8993 6699 9027
rect 6641 8987 6699 8993
rect 6730 8984 6736 9036
rect 6788 8984 6794 9036
rect 7282 8984 7288 9036
rect 7340 8984 7346 9036
rect 7466 8984 7472 9036
rect 7524 8984 7530 9036
rect 7576 9024 7604 9132
rect 9306 9120 9312 9172
rect 9364 9120 9370 9172
rect 9398 9120 9404 9172
rect 9456 9120 9462 9172
rect 9769 9163 9827 9169
rect 9769 9129 9781 9163
rect 9815 9129 9827 9163
rect 9769 9123 9827 9129
rect 9324 9092 9352 9120
rect 9784 9092 9812 9123
rect 10318 9120 10324 9172
rect 10376 9120 10382 9172
rect 10597 9163 10655 9169
rect 10597 9129 10609 9163
rect 10643 9160 10655 9163
rect 11514 9160 11520 9172
rect 10643 9132 11520 9160
rect 10643 9129 10655 9132
rect 10597 9123 10655 9129
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 14734 9120 14740 9172
rect 14792 9160 14798 9172
rect 15749 9163 15807 9169
rect 15749 9160 15761 9163
rect 14792 9132 15761 9160
rect 14792 9120 14798 9132
rect 15749 9129 15761 9132
rect 15795 9129 15807 9163
rect 15749 9123 15807 9129
rect 16577 9163 16635 9169
rect 16577 9129 16589 9163
rect 16623 9160 16635 9163
rect 16850 9160 16856 9172
rect 16623 9132 16856 9160
rect 16623 9129 16635 9132
rect 16577 9123 16635 9129
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 17586 9120 17592 9172
rect 17644 9160 17650 9172
rect 19426 9160 19432 9172
rect 17644 9132 19432 9160
rect 17644 9120 17650 9132
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 21269 9163 21327 9169
rect 21269 9129 21281 9163
rect 21315 9160 21327 9163
rect 21634 9160 21640 9172
rect 21315 9132 21640 9160
rect 21315 9129 21327 9132
rect 21269 9123 21327 9129
rect 21634 9120 21640 9132
rect 21692 9120 21698 9172
rect 23934 9160 23940 9172
rect 21744 9132 23940 9160
rect 9324 9064 9812 9092
rect 12710 9052 12716 9104
rect 12768 9092 12774 9104
rect 13265 9095 13323 9101
rect 13265 9092 13277 9095
rect 12768 9064 13277 9092
rect 12768 9052 12774 9064
rect 13265 9061 13277 9064
rect 13311 9061 13323 9095
rect 13265 9055 13323 9061
rect 15194 9052 15200 9104
rect 15252 9092 15258 9104
rect 15562 9092 15568 9104
rect 15252 9064 15568 9092
rect 15252 9052 15258 9064
rect 15562 9052 15568 9064
rect 15620 9052 15626 9104
rect 15856 9064 16344 9092
rect 8297 9027 8355 9033
rect 8297 9024 8309 9027
rect 7576 8996 8309 9024
rect 8297 8993 8309 8996
rect 8343 8993 8355 9027
rect 8297 8987 8355 8993
rect 9953 9027 10011 9033
rect 9953 8993 9965 9027
rect 9999 9024 10011 9027
rect 10229 9027 10287 9033
rect 10229 9024 10241 9027
rect 9999 8996 10241 9024
rect 9999 8993 10011 8996
rect 9953 8987 10011 8993
rect 10229 8993 10241 8996
rect 10275 9024 10287 9027
rect 10410 9024 10416 9036
rect 10275 8996 10416 9024
rect 10275 8993 10287 8996
rect 10229 8987 10287 8993
rect 10410 8984 10416 8996
rect 10468 8984 10474 9036
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 9024 10563 9027
rect 10594 9024 10600 9036
rect 10551 8996 10600 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 10594 8984 10600 8996
rect 10652 8984 10658 9036
rect 11330 9033 11336 9036
rect 10781 9027 10839 9033
rect 10781 8993 10793 9027
rect 10827 8993 10839 9027
rect 10781 8987 10839 8993
rect 11292 9027 11336 9033
rect 11292 8993 11304 9027
rect 11292 8987 11336 8993
rect 3700 8956 3712 8977
rect 3344 8943 3712 8956
rect 3746 8943 3758 8977
rect 3344 8937 3758 8943
rect 3973 8959 4031 8965
rect 3344 8928 3743 8937
rect 3973 8925 3985 8959
rect 4019 8956 4031 8959
rect 5920 8956 5948 8980
rect 6822 8956 6828 8968
rect 4019 8928 5856 8956
rect 5920 8928 6828 8956
rect 4019 8925 4031 8928
rect 3973 8919 4031 8925
rect 5258 8848 5264 8900
rect 5316 8888 5322 8900
rect 5828 8897 5856 8928
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 6914 8916 6920 8968
rect 6972 8916 6978 8968
rect 7374 8916 7380 8968
rect 7432 8956 7438 8968
rect 7561 8959 7619 8965
rect 7561 8956 7573 8959
rect 7432 8928 7573 8956
rect 7432 8916 7438 8928
rect 7561 8925 7573 8928
rect 7607 8925 7619 8959
rect 7561 8919 7619 8925
rect 7742 8916 7748 8968
rect 7800 8956 7806 8968
rect 7888 8959 7946 8965
rect 7888 8956 7900 8959
rect 7800 8928 7900 8956
rect 7800 8916 7806 8928
rect 7888 8925 7900 8928
rect 7934 8925 7946 8959
rect 7888 8919 7946 8925
rect 8018 8916 8024 8968
rect 8076 8956 8082 8968
rect 8076 8928 8121 8956
rect 8076 8916 8082 8928
rect 8202 8916 8208 8968
rect 8260 8956 8266 8968
rect 10042 8956 10048 8968
rect 8260 8928 10048 8956
rect 8260 8916 8266 8928
rect 10042 8916 10048 8928
rect 10100 8956 10106 8968
rect 10318 8956 10324 8968
rect 10100 8928 10324 8956
rect 10100 8916 10106 8928
rect 10318 8916 10324 8928
rect 10376 8956 10382 8968
rect 10796 8956 10824 8987
rect 11330 8984 11336 8987
rect 11388 8984 11394 9036
rect 11606 8984 11612 9036
rect 11664 9024 11670 9036
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 11664 8996 11713 9024
rect 11664 8984 11670 8996
rect 11701 8993 11713 8996
rect 11747 8993 11759 9027
rect 11701 8987 11759 8993
rect 13078 8984 13084 9036
rect 13136 9024 13142 9036
rect 13906 9033 13912 9036
rect 13868 9027 13912 9033
rect 13868 9024 13880 9027
rect 13136 8996 13880 9024
rect 13136 8984 13142 8996
rect 13868 8993 13880 8996
rect 13868 8987 13912 8993
rect 13906 8984 13912 8987
rect 13964 8984 13970 9036
rect 14277 9027 14335 9033
rect 14277 8993 14289 9027
rect 14323 9024 14335 9027
rect 14918 9024 14924 9036
rect 14323 8996 14924 9024
rect 14323 8993 14335 8996
rect 14277 8987 14335 8993
rect 14918 8984 14924 8996
rect 14976 8984 14982 9036
rect 14037 8977 14095 8983
rect 14037 8974 14049 8977
rect 10376 8928 10824 8956
rect 10965 8959 11023 8965
rect 10376 8916 10382 8928
rect 10965 8925 10977 8959
rect 11011 8956 11023 8959
rect 11146 8956 11152 8968
rect 11011 8928 11152 8956
rect 11011 8925 11023 8928
rect 10965 8919 11023 8925
rect 11146 8916 11152 8928
rect 11204 8916 11210 8968
rect 11428 8961 11486 8967
rect 11428 8927 11440 8961
rect 11474 8956 11486 8961
rect 11514 8956 11520 8968
rect 11474 8928 11520 8956
rect 11474 8927 11486 8928
rect 11428 8921 11486 8927
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 13538 8916 13544 8968
rect 13596 8916 13602 8968
rect 14016 8943 14049 8974
rect 14083 8968 14095 8977
rect 15856 8968 15884 9064
rect 16316 9033 16344 9064
rect 16666 9052 16672 9104
rect 16724 9092 16730 9104
rect 16724 9064 16896 9092
rect 16724 9052 16730 9064
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 8993 15991 9027
rect 15933 8987 15991 8993
rect 16301 9027 16359 9033
rect 16301 8993 16313 9027
rect 16347 8993 16359 9027
rect 16301 8987 16359 8993
rect 14083 8943 14096 8968
rect 14016 8928 14096 8943
rect 14090 8916 14096 8928
rect 14148 8916 14154 8968
rect 15838 8916 15844 8968
rect 15896 8916 15902 8968
rect 15948 8956 15976 8987
rect 16758 8984 16764 9036
rect 16816 8984 16822 9036
rect 16868 9033 16896 9064
rect 19058 9052 19064 9104
rect 19116 9092 19122 9104
rect 20533 9095 20591 9101
rect 20533 9092 20545 9095
rect 19116 9064 20545 9092
rect 19116 9052 19122 9064
rect 20533 9061 20545 9064
rect 20579 9061 20591 9095
rect 20533 9055 20591 9061
rect 20990 9052 20996 9104
rect 21048 9092 21054 9104
rect 21744 9092 21772 9132
rect 21048 9064 21772 9092
rect 21048 9052 21054 9064
rect 21818 9052 21824 9104
rect 21876 9052 21882 9104
rect 16853 9027 16911 9033
rect 16853 8993 16865 9027
rect 16899 9024 16911 9027
rect 17334 9024 17540 9028
rect 17954 9024 17960 9036
rect 16899 9000 17960 9024
rect 16899 8996 17362 9000
rect 17512 8996 17960 9000
rect 16899 8993 16911 8996
rect 16853 8987 16911 8993
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 19242 8984 19248 9036
rect 19300 9024 19306 9036
rect 20162 9024 20168 9036
rect 19300 8996 20168 9024
rect 19300 8984 19306 8996
rect 20162 8984 20168 8996
rect 20220 8984 20226 9036
rect 20257 9027 20315 9033
rect 20257 8993 20269 9027
rect 20303 8993 20315 9027
rect 20257 8987 20315 8993
rect 16482 8956 16488 8968
rect 15948 8928 16488 8956
rect 16482 8916 16488 8928
rect 16540 8916 16546 8968
rect 17126 8916 17132 8968
rect 17184 8965 17190 8968
rect 17402 8965 17408 8968
rect 17184 8959 17238 8965
rect 17184 8925 17192 8959
rect 17226 8925 17238 8959
rect 17184 8919 17238 8925
rect 17359 8959 17408 8965
rect 17359 8925 17371 8959
rect 17405 8925 17408 8959
rect 17359 8919 17408 8925
rect 17184 8916 17190 8919
rect 17402 8916 17408 8919
rect 17460 8916 17466 8968
rect 17589 8959 17647 8965
rect 17589 8925 17601 8959
rect 17635 8956 17647 8959
rect 17770 8956 17776 8968
rect 17635 8928 17776 8956
rect 17635 8925 17647 8928
rect 17589 8919 17647 8925
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 18414 8916 18420 8968
rect 18472 8956 18478 8968
rect 19794 8956 19800 8968
rect 18472 8928 19800 8956
rect 18472 8916 18478 8928
rect 19794 8916 19800 8928
rect 19852 8916 19858 8968
rect 5813 8891 5871 8897
rect 5316 8860 5764 8888
rect 5316 8848 5322 8860
rect 5350 8820 5356 8832
rect 2746 8792 5356 8820
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 5442 8780 5448 8832
rect 5500 8780 5506 8832
rect 5736 8820 5764 8860
rect 5813 8857 5825 8891
rect 5859 8857 5871 8891
rect 10226 8888 10232 8900
rect 5813 8851 5871 8857
rect 6104 8860 7420 8888
rect 6104 8820 6132 8860
rect 5736 8792 6132 8820
rect 6178 8780 6184 8832
rect 6236 8780 6242 8832
rect 6454 8780 6460 8832
rect 6512 8780 6518 8832
rect 7392 8820 7420 8860
rect 9968 8860 10232 8888
rect 9968 8820 9996 8860
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 10468 8860 11008 8888
rect 10468 8848 10474 8860
rect 7392 8792 9996 8820
rect 10045 8823 10103 8829
rect 10045 8789 10057 8823
rect 10091 8820 10103 8823
rect 10870 8820 10876 8832
rect 10091 8792 10876 8820
rect 10091 8789 10103 8792
rect 10045 8783 10103 8789
rect 10870 8780 10876 8792
rect 10928 8780 10934 8832
rect 10980 8820 11008 8860
rect 15120 8860 16712 8888
rect 11330 8820 11336 8832
rect 10980 8792 11336 8820
rect 11330 8780 11336 8792
rect 11388 8780 11394 8832
rect 12802 8780 12808 8832
rect 12860 8780 12866 8832
rect 13354 8780 13360 8832
rect 13412 8780 13418 8832
rect 13722 8780 13728 8832
rect 13780 8820 13786 8832
rect 15120 8820 15148 8860
rect 16684 8832 16712 8860
rect 18322 8848 18328 8900
rect 18380 8888 18386 8900
rect 18966 8888 18972 8900
rect 18380 8860 18972 8888
rect 18380 8848 18386 8860
rect 18966 8848 18972 8860
rect 19024 8888 19030 8900
rect 20272 8888 20300 8987
rect 20898 8984 20904 9036
rect 20956 9024 20962 9036
rect 21453 9027 21511 9033
rect 21453 9024 21465 9027
rect 20956 8996 21465 9024
rect 20956 8984 20962 8996
rect 21453 8993 21465 8996
rect 21499 9024 21511 9027
rect 21836 9024 21864 9052
rect 21499 8996 21864 9024
rect 22189 9027 22247 9033
rect 21499 8993 21511 8996
rect 21453 8987 21511 8993
rect 22189 8993 22201 9027
rect 22235 9024 22247 9027
rect 22830 9024 22836 9036
rect 22235 8996 22836 9024
rect 22235 8993 22247 8996
rect 22189 8987 22247 8993
rect 22830 8984 22836 8996
rect 22888 8984 22894 9036
rect 22940 9033 22968 9132
rect 23934 9120 23940 9132
rect 23992 9120 23998 9172
rect 25682 9120 25688 9172
rect 25740 9120 25746 9172
rect 25961 9163 26019 9169
rect 25961 9129 25973 9163
rect 26007 9160 26019 9163
rect 26786 9160 26792 9172
rect 26007 9132 26792 9160
rect 26007 9129 26019 9132
rect 25961 9123 26019 9129
rect 26786 9120 26792 9132
rect 26844 9120 26850 9172
rect 26878 9120 26884 9172
rect 26936 9169 26942 9172
rect 26936 9160 26945 9169
rect 26936 9132 26981 9160
rect 26936 9123 26945 9132
rect 26936 9120 26942 9123
rect 27890 9120 27896 9172
rect 27948 9120 27954 9172
rect 28534 9120 28540 9172
rect 28592 9120 28598 9172
rect 30193 9163 30251 9169
rect 30193 9129 30205 9163
rect 30239 9160 30251 9163
rect 31110 9160 31116 9172
rect 30239 9132 31116 9160
rect 30239 9129 30251 9132
rect 30193 9123 30251 9129
rect 31110 9120 31116 9132
rect 31168 9120 31174 9172
rect 23014 9052 23020 9104
rect 23072 9052 23078 9104
rect 24854 9052 24860 9104
rect 24912 9092 24918 9104
rect 25225 9095 25283 9101
rect 25225 9092 25237 9095
rect 24912 9064 25237 9092
rect 24912 9052 24918 9064
rect 25225 9061 25237 9064
rect 25271 9061 25283 9095
rect 25225 9055 25283 9061
rect 22925 9027 22983 9033
rect 22925 8993 22937 9027
rect 22971 8993 22983 9027
rect 23032 9024 23060 9052
rect 23252 9027 23310 9033
rect 23252 9024 23264 9027
rect 23032 8996 23264 9024
rect 22925 8987 22983 8993
rect 23252 8993 23264 8996
rect 23298 8993 23310 9027
rect 23252 8987 23310 8993
rect 23658 8984 23664 9036
rect 23716 8984 23722 9036
rect 23750 8984 23756 9036
rect 23808 9024 23814 9036
rect 25774 9024 25780 9036
rect 23808 8996 25780 9024
rect 23808 8984 23814 8996
rect 25774 8984 25780 8996
rect 25832 8984 25838 9036
rect 25869 9027 25927 9033
rect 25869 8993 25881 9027
rect 25915 9024 25927 9027
rect 25958 9024 25964 9036
rect 25915 8996 25964 9024
rect 25915 8993 25927 8996
rect 25869 8987 25927 8993
rect 25958 8984 25964 8996
rect 26016 8984 26022 9036
rect 26142 8984 26148 9036
rect 26200 8984 26206 9036
rect 26418 8984 26424 9036
rect 26476 8984 26482 9036
rect 26694 8984 26700 9036
rect 26752 8984 26758 9036
rect 27908 9024 27936 9120
rect 27080 8996 27936 9024
rect 20530 8916 20536 8968
rect 20588 8956 20594 8968
rect 22738 8956 22744 8968
rect 20588 8928 22744 8956
rect 20588 8916 20594 8928
rect 22738 8916 22744 8928
rect 22796 8916 22802 8968
rect 23431 8959 23489 8965
rect 23431 8925 23443 8959
rect 23477 8956 23489 8959
rect 23566 8956 23572 8968
rect 23477 8928 23572 8956
rect 23477 8925 23489 8928
rect 23431 8919 23489 8925
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 23842 8916 23848 8968
rect 23900 8956 23906 8968
rect 25501 8959 25559 8965
rect 25501 8956 25513 8959
rect 23900 8928 25513 8956
rect 23900 8916 23906 8928
rect 25501 8925 25513 8928
rect 25547 8925 25559 8959
rect 26160 8956 26188 8984
rect 26712 8956 26740 8984
rect 26160 8928 26740 8956
rect 26927 8959 26985 8965
rect 25501 8919 25559 8925
rect 26927 8925 26939 8959
rect 26973 8956 26985 8959
rect 27080 8956 27108 8996
rect 26973 8928 27108 8956
rect 27157 8959 27215 8965
rect 26973 8925 26985 8928
rect 26927 8919 26985 8925
rect 27157 8925 27169 8959
rect 27203 8956 27215 8959
rect 28552 8956 28580 9120
rect 28629 9027 28687 9033
rect 28629 8993 28641 9027
rect 28675 8993 28687 9027
rect 28629 8987 28687 8993
rect 28905 9027 28963 9033
rect 28905 8993 28917 9027
rect 28951 9024 28963 9027
rect 30006 9024 30012 9036
rect 28951 8996 30012 9024
rect 28951 8993 28963 8996
rect 28905 8987 28963 8993
rect 27203 8928 28580 8956
rect 27203 8925 27215 8928
rect 27157 8919 27215 8925
rect 19024 8860 20300 8888
rect 19024 8848 19030 8860
rect 28166 8848 28172 8900
rect 28224 8888 28230 8900
rect 28644 8888 28672 8987
rect 30006 8984 30012 8996
rect 30064 8984 30070 9036
rect 28224 8860 28672 8888
rect 28224 8848 28230 8860
rect 13780 8792 15148 8820
rect 13780 8780 13786 8792
rect 15194 8780 15200 8832
rect 15252 8820 15258 8832
rect 15381 8823 15439 8829
rect 15381 8820 15393 8823
rect 15252 8792 15393 8820
rect 15252 8780 15258 8792
rect 15381 8789 15393 8792
rect 15427 8789 15439 8823
rect 15381 8783 15439 8789
rect 16114 8780 16120 8832
rect 16172 8780 16178 8832
rect 16666 8780 16672 8832
rect 16724 8780 16730 8832
rect 17770 8780 17776 8832
rect 17828 8820 17834 8832
rect 18693 8823 18751 8829
rect 18693 8820 18705 8823
rect 17828 8792 18705 8820
rect 17828 8780 17834 8792
rect 18693 8789 18705 8792
rect 18739 8789 18751 8823
rect 18693 8783 18751 8789
rect 18782 8780 18788 8832
rect 18840 8820 18846 8832
rect 19061 8823 19119 8829
rect 19061 8820 19073 8823
rect 18840 8792 19073 8820
rect 18840 8780 18846 8792
rect 19061 8789 19073 8792
rect 19107 8789 19119 8823
rect 19061 8783 19119 8789
rect 22005 8823 22063 8829
rect 22005 8789 22017 8823
rect 22051 8820 22063 8823
rect 22186 8820 22192 8832
rect 22051 8792 22192 8820
rect 22051 8789 22063 8792
rect 22005 8783 22063 8789
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 22649 8823 22707 8829
rect 22649 8789 22661 8823
rect 22695 8820 22707 8823
rect 24486 8820 24492 8832
rect 22695 8792 24492 8820
rect 22695 8789 22707 8792
rect 22649 8783 22707 8789
rect 24486 8780 24492 8792
rect 24544 8780 24550 8832
rect 24946 8780 24952 8832
rect 25004 8780 25010 8832
rect 26878 8780 26884 8832
rect 26936 8820 26942 8832
rect 27522 8820 27528 8832
rect 26936 8792 27528 8820
rect 26936 8780 26942 8792
rect 27522 8780 27528 8792
rect 27580 8820 27586 8832
rect 27890 8820 27896 8832
rect 27580 8792 27896 8820
rect 27580 8780 27586 8792
rect 27890 8780 27896 8792
rect 27948 8780 27954 8832
rect 28258 8780 28264 8832
rect 28316 8780 28322 8832
rect 552 8730 30912 8752
rect 552 8678 4193 8730
rect 4245 8678 4257 8730
rect 4309 8678 4321 8730
rect 4373 8678 4385 8730
rect 4437 8678 4449 8730
rect 4501 8678 11783 8730
rect 11835 8678 11847 8730
rect 11899 8678 11911 8730
rect 11963 8678 11975 8730
rect 12027 8678 12039 8730
rect 12091 8678 19373 8730
rect 19425 8678 19437 8730
rect 19489 8678 19501 8730
rect 19553 8678 19565 8730
rect 19617 8678 19629 8730
rect 19681 8678 26963 8730
rect 27015 8678 27027 8730
rect 27079 8678 27091 8730
rect 27143 8678 27155 8730
rect 27207 8678 27219 8730
rect 27271 8678 30912 8730
rect 552 8656 30912 8678
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 2777 8619 2835 8625
rect 2777 8616 2789 8619
rect 2096 8588 2789 8616
rect 2096 8576 2102 8588
rect 2777 8585 2789 8588
rect 2823 8585 2835 8619
rect 2777 8579 2835 8585
rect 2958 8576 2964 8628
rect 3016 8616 3022 8628
rect 3016 8588 6960 8616
rect 3016 8576 3022 8588
rect 2406 8508 2412 8560
rect 2464 8548 2470 8560
rect 2464 8520 3372 8548
rect 2464 8508 2470 8520
rect 3344 8492 3372 8520
rect 5166 8508 5172 8560
rect 5224 8508 5230 8560
rect 6932 8548 6960 8588
rect 7098 8576 7104 8628
rect 7156 8616 7162 8628
rect 7377 8619 7435 8625
rect 7377 8616 7389 8619
rect 7156 8588 7389 8616
rect 7156 8576 7162 8588
rect 7377 8585 7389 8588
rect 7423 8585 7435 8619
rect 7377 8579 7435 8585
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 7745 8619 7803 8625
rect 7745 8616 7757 8619
rect 7616 8588 7757 8616
rect 7616 8576 7622 8588
rect 7745 8585 7757 8588
rect 7791 8585 7803 8619
rect 7745 8579 7803 8585
rect 8938 8576 8944 8628
rect 8996 8616 9002 8628
rect 8996 8588 9260 8616
rect 8996 8576 9002 8588
rect 9125 8551 9183 8557
rect 9125 8548 9137 8551
rect 6932 8520 9137 8548
rect 9125 8517 9137 8520
rect 9171 8517 9183 8551
rect 9125 8511 9183 8517
rect 1443 8483 1501 8489
rect 1443 8449 1455 8483
rect 1489 8480 1501 8483
rect 3142 8480 3148 8492
rect 1489 8452 3148 8480
rect 1489 8449 1501 8452
rect 1443 8443 1501 8449
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 3326 8440 3332 8492
rect 3384 8440 3390 8492
rect 3835 8483 3893 8489
rect 3835 8449 3847 8483
rect 3881 8480 3893 8483
rect 3970 8480 3976 8492
rect 3881 8452 3976 8480
rect 3881 8449 3893 8452
rect 3835 8443 3893 8449
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8480 4123 8483
rect 5258 8480 5264 8492
rect 4111 8452 5264 8480
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 5718 8440 5724 8492
rect 5776 8480 5782 8492
rect 6000 8483 6058 8489
rect 6000 8480 6012 8483
rect 5776 8452 6012 8480
rect 5776 8440 5782 8452
rect 6000 8449 6012 8452
rect 6046 8449 6058 8483
rect 6000 8443 6058 8449
rect 6362 8440 6368 8492
rect 6420 8440 6426 8492
rect 7006 8440 7012 8492
rect 7064 8480 7070 8492
rect 9232 8480 9260 8588
rect 11514 8576 11520 8628
rect 11572 8576 11578 8628
rect 11606 8576 11612 8628
rect 11664 8616 11670 8628
rect 18138 8616 18144 8628
rect 11664 8588 12020 8616
rect 11664 8576 11670 8588
rect 11992 8548 12020 8588
rect 16408 8588 18144 8616
rect 12805 8551 12863 8557
rect 12805 8548 12817 8551
rect 11992 8520 12817 8548
rect 12805 8517 12817 8520
rect 12851 8517 12863 8551
rect 12805 8511 12863 8517
rect 9956 8483 10014 8489
rect 9956 8480 9968 8483
rect 7064 8452 8156 8480
rect 9232 8452 9968 8480
rect 7064 8440 7070 8452
rect 842 8372 848 8424
rect 900 8412 906 8424
rect 937 8415 995 8421
rect 937 8412 949 8415
rect 900 8384 949 8412
rect 900 8372 906 8384
rect 937 8381 949 8384
rect 983 8381 995 8415
rect 937 8375 995 8381
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 2958 8412 2964 8424
rect 1719 8384 2964 8412
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 2958 8372 2964 8384
rect 3016 8372 3022 8424
rect 3602 8412 3608 8424
rect 3436 8384 3608 8412
rect 2774 8304 2780 8356
rect 2832 8344 2838 8356
rect 3436 8344 3464 8384
rect 3602 8372 3608 8384
rect 3660 8421 3666 8424
rect 3660 8415 3714 8421
rect 3660 8381 3668 8415
rect 3702 8381 3714 8415
rect 6273 8415 6331 8421
rect 6273 8412 6285 8415
rect 3660 8375 3714 8381
rect 5644 8384 6285 8412
rect 3660 8372 3666 8375
rect 2832 8316 3464 8344
rect 2832 8304 2838 8316
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 5644 8344 5672 8384
rect 6273 8381 6285 8384
rect 6319 8381 6331 8415
rect 6380 8412 6408 8440
rect 6380 8384 6960 8412
rect 6273 8375 6331 8381
rect 5500 8316 5672 8344
rect 6932 8344 6960 8384
rect 7098 8372 7104 8424
rect 7156 8412 7162 8424
rect 7650 8412 7656 8424
rect 7156 8384 7656 8412
rect 7156 8372 7162 8384
rect 7650 8372 7656 8384
rect 7708 8412 7714 8424
rect 7929 8415 7987 8421
rect 7929 8412 7941 8415
rect 7708 8384 7941 8412
rect 7708 8372 7714 8384
rect 7929 8381 7941 8384
rect 7975 8381 7987 8415
rect 8128 8412 8156 8452
rect 9956 8449 9968 8452
rect 10002 8449 10014 8483
rect 9956 8443 10014 8449
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10686 8480 10692 8492
rect 10275 8452 10692 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10686 8440 10692 8452
rect 10744 8440 10750 8492
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 12069 8483 12127 8489
rect 12069 8480 12081 8483
rect 11204 8452 12081 8480
rect 11204 8440 11210 8452
rect 12069 8449 12081 8452
rect 12115 8480 12127 8483
rect 13538 8480 13544 8492
rect 12115 8452 13544 8480
rect 12115 8449 12127 8452
rect 12069 8443 12127 8449
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 14047 8483 14105 8489
rect 14047 8449 14059 8483
rect 14093 8480 14105 8483
rect 14182 8480 14188 8492
rect 14093 8452 14188 8480
rect 14093 8449 14105 8452
rect 14047 8443 14105 8449
rect 14182 8440 14188 8452
rect 14240 8440 14246 8492
rect 14277 8483 14335 8489
rect 14277 8449 14289 8483
rect 14323 8480 14335 8483
rect 15470 8480 15476 8492
rect 14323 8452 15476 8480
rect 14323 8449 14335 8452
rect 14277 8443 14335 8449
rect 15470 8440 15476 8452
rect 15528 8440 15534 8492
rect 16408 8480 16436 8588
rect 18138 8576 18144 8588
rect 18196 8576 18202 8628
rect 18230 8576 18236 8628
rect 18288 8576 18294 8628
rect 20717 8619 20775 8625
rect 20717 8585 20729 8619
rect 20763 8616 20775 8619
rect 21542 8616 21548 8628
rect 20763 8588 21548 8616
rect 20763 8585 20775 8588
rect 20717 8579 20775 8585
rect 21542 8576 21548 8588
rect 21600 8576 21606 8628
rect 21726 8576 21732 8628
rect 21784 8616 21790 8628
rect 22741 8619 22799 8625
rect 22741 8616 22753 8619
rect 21784 8588 22753 8616
rect 21784 8576 21790 8588
rect 22741 8585 22753 8588
rect 22787 8585 22799 8619
rect 22741 8579 22799 8585
rect 22830 8576 22836 8628
rect 22888 8616 22894 8628
rect 22888 8588 25268 8616
rect 22888 8576 22894 8588
rect 23750 8548 23756 8560
rect 23676 8520 23756 8548
rect 16720 8483 16778 8489
rect 16720 8480 16732 8483
rect 16408 8452 16732 8480
rect 16720 8449 16732 8452
rect 16766 8449 16778 8483
rect 16720 8443 16778 8449
rect 16868 8465 17908 8480
rect 16868 8434 16901 8465
rect 16889 8431 16901 8434
rect 16935 8452 17908 8465
rect 16935 8431 16947 8452
rect 16889 8425 16947 8431
rect 8202 8412 8208 8424
rect 8128 8384 8208 8412
rect 7929 8375 7987 8381
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 8662 8412 8668 8424
rect 8312 8384 8668 8412
rect 6932 8316 7052 8344
rect 5500 8304 5506 8316
rect 1394 8236 1400 8288
rect 1452 8285 1458 8288
rect 1452 8276 1461 8285
rect 1452 8248 1497 8276
rect 1452 8239 1461 8248
rect 1452 8236 1458 8239
rect 5994 8236 6000 8288
rect 6052 8285 6058 8288
rect 6052 8239 6061 8285
rect 6052 8236 6058 8239
rect 6362 8236 6368 8288
rect 6420 8276 6426 8288
rect 6914 8276 6920 8288
rect 6420 8248 6920 8276
rect 6420 8236 6426 8248
rect 6914 8236 6920 8248
rect 6972 8236 6978 8288
rect 7024 8276 7052 8316
rect 7282 8304 7288 8356
rect 7340 8344 7346 8356
rect 7834 8344 7840 8356
rect 7340 8316 7840 8344
rect 7340 8304 7346 8316
rect 7834 8304 7840 8316
rect 7892 8344 7898 8356
rect 8312 8344 8340 8384
rect 8662 8372 8668 8384
rect 8720 8412 8726 8424
rect 8849 8415 8907 8421
rect 8849 8412 8861 8415
rect 8720 8384 8861 8412
rect 8720 8372 8726 8384
rect 8849 8381 8861 8384
rect 8895 8381 8907 8415
rect 8849 8375 8907 8381
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8412 9367 8415
rect 9398 8412 9404 8424
rect 9355 8384 9404 8412
rect 9355 8381 9367 8384
rect 9309 8375 9367 8381
rect 9398 8372 9404 8384
rect 9456 8372 9462 8424
rect 9490 8372 9496 8424
rect 9548 8372 9554 8424
rect 9582 8372 9588 8424
rect 9640 8412 9646 8424
rect 9820 8415 9878 8421
rect 9820 8412 9832 8415
rect 9640 8384 9832 8412
rect 9640 8372 9646 8384
rect 9820 8381 9832 8384
rect 9866 8381 9878 8415
rect 9820 8375 9878 8381
rect 10594 8372 10600 8424
rect 10652 8412 10658 8424
rect 12529 8415 12587 8421
rect 12529 8412 12541 8415
rect 10652 8384 12541 8412
rect 10652 8372 10658 8384
rect 10980 8356 11008 8384
rect 12529 8381 12541 8384
rect 12575 8381 12587 8415
rect 12529 8375 12587 8381
rect 12618 8372 12624 8424
rect 12676 8372 12682 8424
rect 12710 8372 12716 8424
rect 12768 8412 12774 8424
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12768 8384 12909 8412
rect 12768 8372 12774 8384
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 13078 8372 13084 8424
rect 13136 8412 13142 8424
rect 13173 8415 13231 8421
rect 13173 8412 13185 8415
rect 13136 8384 13185 8412
rect 13136 8372 13142 8384
rect 13173 8381 13185 8384
rect 13219 8412 13231 8415
rect 13868 8415 13926 8421
rect 13868 8412 13880 8415
rect 13219 8384 13880 8412
rect 13219 8381 13231 8384
rect 13173 8375 13231 8381
rect 13868 8381 13880 8384
rect 13914 8381 13926 8415
rect 13868 8375 13926 8381
rect 15562 8372 15568 8424
rect 15620 8412 15626 8424
rect 15841 8415 15899 8421
rect 15841 8412 15853 8415
rect 15620 8384 15853 8412
rect 15620 8372 15626 8384
rect 15841 8381 15853 8384
rect 15887 8381 15899 8415
rect 15841 8375 15899 8381
rect 16393 8415 16451 8421
rect 16393 8381 16405 8415
rect 16439 8412 16451 8415
rect 17129 8415 17187 8421
rect 16439 8384 16528 8412
rect 16439 8381 16451 8384
rect 16393 8375 16451 8381
rect 7892 8316 8340 8344
rect 8481 8347 8539 8353
rect 7892 8304 7898 8316
rect 8481 8313 8493 8347
rect 8527 8344 8539 8347
rect 8527 8316 9628 8344
rect 8527 8313 8539 8316
rect 8481 8307 8539 8313
rect 7098 8276 7104 8288
rect 7024 8248 7104 8276
rect 7098 8236 7104 8248
rect 7156 8236 7162 8288
rect 8021 8279 8079 8285
rect 8021 8245 8033 8279
rect 8067 8276 8079 8279
rect 9122 8276 9128 8288
rect 8067 8248 9128 8276
rect 8067 8245 8079 8248
rect 8021 8239 8079 8245
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 9600 8276 9628 8316
rect 10962 8304 10968 8356
rect 11020 8304 11026 8356
rect 11238 8304 11244 8356
rect 11296 8344 11302 8356
rect 11793 8347 11851 8353
rect 11793 8344 11805 8347
rect 11296 8316 11805 8344
rect 11296 8304 11302 8316
rect 11793 8313 11805 8316
rect 11839 8313 11851 8347
rect 12158 8344 12164 8356
rect 11793 8307 11851 8313
rect 11900 8316 12164 8344
rect 11900 8276 11928 8316
rect 12158 8304 12164 8316
rect 12216 8344 12222 8356
rect 12309 8347 12367 8353
rect 12309 8344 12321 8347
rect 12216 8316 12321 8344
rect 12216 8304 12222 8316
rect 12309 8313 12321 8316
rect 12355 8313 12367 8347
rect 12309 8307 12367 8313
rect 9600 8248 11928 8276
rect 13814 8236 13820 8288
rect 13872 8276 13878 8288
rect 15381 8279 15439 8285
rect 15381 8276 15393 8279
rect 13872 8248 15393 8276
rect 13872 8236 13878 8248
rect 15381 8245 15393 8248
rect 15427 8245 15439 8279
rect 15381 8239 15439 8245
rect 15838 8236 15844 8288
rect 15896 8276 15902 8288
rect 16117 8279 16175 8285
rect 16117 8276 16129 8279
rect 15896 8248 16129 8276
rect 15896 8236 15902 8248
rect 16117 8245 16129 8248
rect 16163 8276 16175 8279
rect 16206 8276 16212 8288
rect 16163 8248 16212 8276
rect 16163 8245 16175 8248
rect 16117 8239 16175 8245
rect 16206 8236 16212 8248
rect 16264 8236 16270 8288
rect 16500 8276 16528 8384
rect 17129 8381 17141 8415
rect 17175 8412 17187 8415
rect 17218 8412 17224 8424
rect 17175 8384 17224 8412
rect 17175 8381 17187 8384
rect 17129 8375 17187 8381
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 17770 8276 17776 8288
rect 16500 8248 17776 8276
rect 17770 8236 17776 8248
rect 17828 8236 17834 8288
rect 17880 8276 17908 8452
rect 17954 8440 17960 8492
rect 18012 8480 18018 8492
rect 18690 8480 18696 8492
rect 18012 8452 18696 8480
rect 18012 8440 18018 8452
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 19058 8489 19064 8492
rect 19020 8483 19064 8489
rect 19020 8449 19032 8483
rect 19020 8443 19064 8449
rect 19058 8440 19064 8443
rect 19116 8440 19122 8492
rect 19199 8483 19257 8489
rect 19199 8449 19211 8483
rect 19245 8480 19257 8483
rect 21228 8483 21286 8489
rect 21228 8480 21240 8483
rect 19245 8452 19748 8480
rect 19245 8449 19257 8452
rect 19199 8443 19257 8449
rect 19720 8424 19748 8452
rect 20732 8452 21240 8480
rect 20732 8424 20760 8452
rect 21228 8449 21240 8452
rect 21274 8449 21286 8483
rect 21228 8443 21286 8449
rect 21407 8483 21465 8489
rect 21407 8449 21419 8483
rect 21453 8480 21465 8483
rect 23676 8480 23704 8520
rect 23750 8508 23756 8520
rect 23808 8508 23814 8560
rect 24308 8483 24366 8489
rect 24308 8480 24320 8483
rect 21453 8452 23704 8480
rect 23768 8452 24320 8480
rect 21453 8449 21465 8452
rect 21407 8443 21465 8449
rect 18782 8372 18788 8424
rect 18840 8412 18846 8424
rect 19429 8415 19487 8421
rect 19429 8412 19441 8415
rect 18840 8384 19441 8412
rect 18840 8372 18846 8384
rect 19429 8381 19441 8384
rect 19475 8381 19487 8415
rect 19429 8375 19487 8381
rect 19702 8372 19708 8424
rect 19760 8372 19766 8424
rect 20714 8372 20720 8424
rect 20772 8372 20778 8424
rect 20806 8372 20812 8424
rect 20864 8412 20870 8424
rect 20901 8415 20959 8421
rect 20901 8412 20913 8415
rect 20864 8384 20913 8412
rect 20864 8372 20870 8384
rect 20901 8381 20913 8384
rect 20947 8381 20959 8415
rect 21637 8415 21695 8421
rect 21637 8412 21649 8415
rect 20901 8375 20959 8381
rect 21008 8384 21649 8412
rect 20438 8304 20444 8356
rect 20496 8344 20502 8356
rect 21008 8344 21036 8384
rect 21637 8381 21649 8384
rect 21683 8381 21695 8415
rect 21637 8375 21695 8381
rect 21726 8372 21732 8424
rect 21784 8412 21790 8424
rect 23201 8415 23259 8421
rect 23201 8412 23213 8415
rect 21784 8384 23213 8412
rect 21784 8372 21790 8384
rect 23201 8381 23213 8384
rect 23247 8381 23259 8415
rect 23201 8375 23259 8381
rect 23768 8356 23796 8452
rect 24308 8449 24320 8452
rect 24354 8449 24366 8483
rect 24308 8443 24366 8449
rect 24486 8440 24492 8492
rect 24544 8480 24550 8492
rect 24581 8483 24639 8489
rect 24581 8480 24593 8483
rect 24544 8452 24593 8480
rect 24544 8440 24550 8452
rect 24581 8449 24593 8452
rect 24627 8449 24639 8483
rect 25240 8480 25268 8588
rect 25314 8576 25320 8628
rect 25372 8616 25378 8628
rect 26053 8619 26111 8625
rect 26053 8616 26065 8619
rect 25372 8588 26065 8616
rect 25372 8576 25378 8588
rect 26053 8585 26065 8588
rect 26099 8585 26111 8619
rect 26053 8579 26111 8585
rect 26326 8576 26332 8628
rect 26384 8576 26390 8628
rect 26510 8576 26516 8628
rect 26568 8616 26574 8628
rect 27614 8616 27620 8628
rect 26568 8588 27620 8616
rect 26568 8576 26574 8588
rect 27614 8576 27620 8588
rect 27672 8576 27678 8628
rect 27798 8576 27804 8628
rect 27856 8616 27862 8628
rect 28537 8619 28595 8625
rect 28537 8616 28549 8619
rect 27856 8588 28549 8616
rect 27856 8576 27862 8588
rect 28537 8585 28549 8588
rect 28583 8585 28595 8619
rect 28537 8579 28595 8585
rect 28626 8576 28632 8628
rect 28684 8616 28690 8628
rect 29181 8619 29239 8625
rect 29181 8616 29193 8619
rect 28684 8588 29193 8616
rect 28684 8576 28690 8588
rect 29181 8585 29193 8588
rect 29227 8585 29239 8619
rect 29181 8579 29239 8585
rect 29270 8576 29276 8628
rect 29328 8616 29334 8628
rect 30190 8616 30196 8628
rect 29328 8588 30196 8616
rect 29328 8576 29334 8588
rect 30190 8576 30196 8588
rect 30248 8616 30254 8628
rect 30285 8619 30343 8625
rect 30285 8616 30297 8619
rect 30248 8588 30297 8616
rect 30248 8576 30254 8588
rect 30285 8585 30297 8588
rect 30331 8585 30343 8619
rect 30285 8579 30343 8585
rect 25866 8508 25872 8560
rect 25924 8508 25930 8560
rect 26528 8480 26556 8576
rect 29638 8508 29644 8560
rect 29696 8548 29702 8560
rect 29696 8520 30236 8548
rect 29696 8508 29702 8520
rect 26697 8483 26755 8489
rect 26697 8480 26709 8483
rect 25240 8452 26464 8480
rect 26528 8452 26709 8480
rect 24581 8443 24639 8449
rect 23845 8415 23903 8421
rect 23845 8381 23857 8415
rect 23891 8412 23903 8415
rect 23934 8412 23940 8424
rect 23891 8384 23940 8412
rect 23891 8381 23903 8384
rect 23845 8375 23903 8381
rect 23934 8372 23940 8384
rect 23992 8372 23998 8424
rect 24210 8421 24216 8424
rect 24172 8415 24216 8421
rect 24172 8381 24184 8415
rect 24172 8375 24216 8381
rect 24210 8372 24216 8375
rect 24268 8372 24274 8424
rect 24670 8372 24676 8424
rect 24728 8412 24734 8424
rect 25958 8412 25964 8424
rect 24728 8384 25964 8412
rect 24728 8372 24734 8384
rect 25958 8372 25964 8384
rect 26016 8412 26022 8424
rect 26237 8415 26295 8421
rect 26237 8412 26249 8415
rect 26016 8384 26249 8412
rect 26016 8372 26022 8384
rect 26237 8381 26249 8384
rect 26283 8381 26295 8415
rect 26237 8375 26295 8381
rect 23569 8347 23627 8353
rect 20496 8316 21036 8344
rect 23216 8316 23428 8344
rect 20496 8304 20502 8316
rect 23216 8276 23244 8316
rect 17880 8248 23244 8276
rect 23400 8276 23428 8316
rect 23569 8313 23581 8347
rect 23615 8344 23627 8347
rect 23658 8344 23664 8356
rect 23615 8316 23664 8344
rect 23615 8313 23627 8316
rect 23569 8307 23627 8313
rect 23658 8304 23664 8316
rect 23716 8304 23722 8356
rect 23750 8304 23756 8356
rect 23808 8304 23814 8356
rect 25866 8276 25872 8288
rect 23400 8248 25872 8276
rect 25866 8236 25872 8248
rect 25924 8236 25930 8288
rect 26252 8276 26280 8375
rect 26436 8356 26464 8452
rect 26697 8449 26709 8452
rect 26743 8449 26755 8483
rect 26697 8443 26755 8449
rect 26878 8440 26884 8492
rect 26936 8480 26942 8492
rect 27024 8483 27082 8489
rect 27024 8480 27036 8483
rect 26936 8452 27036 8480
rect 26936 8440 26942 8452
rect 27024 8449 27036 8452
rect 27070 8449 27082 8483
rect 27024 8443 27082 8449
rect 27203 8483 27261 8489
rect 27203 8449 27215 8483
rect 27249 8480 27261 8483
rect 28074 8480 28080 8492
rect 27249 8452 28080 8480
rect 27249 8449 27261 8452
rect 27203 8443 27261 8449
rect 28074 8440 28080 8452
rect 28132 8440 28138 8492
rect 29362 8480 29368 8492
rect 28176 8452 29368 8480
rect 26513 8415 26571 8421
rect 26513 8381 26525 8415
rect 26559 8381 26571 8415
rect 26513 8375 26571 8381
rect 26418 8304 26424 8356
rect 26476 8304 26482 8356
rect 26528 8276 26556 8375
rect 27430 8372 27436 8424
rect 27488 8372 27494 8424
rect 28176 8276 28204 8452
rect 29362 8440 29368 8452
rect 29420 8440 29426 8492
rect 28350 8372 28356 8424
rect 28408 8372 28414 8424
rect 29086 8372 29092 8424
rect 29144 8372 29150 8424
rect 30208 8421 30236 8520
rect 30193 8415 30251 8421
rect 30193 8381 30205 8415
rect 30239 8381 30251 8415
rect 30193 8375 30251 8381
rect 28368 8344 28396 8372
rect 29641 8347 29699 8353
rect 29641 8344 29653 8347
rect 28368 8316 29653 8344
rect 29641 8313 29653 8316
rect 29687 8313 29699 8347
rect 29641 8307 29699 8313
rect 26252 8248 28204 8276
rect 29086 8236 29092 8288
rect 29144 8276 29150 8288
rect 29733 8279 29791 8285
rect 29733 8276 29745 8279
rect 29144 8248 29745 8276
rect 29144 8236 29150 8248
rect 29733 8245 29745 8248
rect 29779 8245 29791 8279
rect 29733 8239 29791 8245
rect 552 8186 31072 8208
rect 552 8134 7988 8186
rect 8040 8134 8052 8186
rect 8104 8134 8116 8186
rect 8168 8134 8180 8186
rect 8232 8134 8244 8186
rect 8296 8134 15578 8186
rect 15630 8134 15642 8186
rect 15694 8134 15706 8186
rect 15758 8134 15770 8186
rect 15822 8134 15834 8186
rect 15886 8134 23168 8186
rect 23220 8134 23232 8186
rect 23284 8134 23296 8186
rect 23348 8134 23360 8186
rect 23412 8134 23424 8186
rect 23476 8134 30758 8186
rect 30810 8134 30822 8186
rect 30874 8134 30886 8186
rect 30938 8134 30950 8186
rect 31002 8134 31014 8186
rect 31066 8134 31072 8186
rect 552 8112 31072 8134
rect 5166 8032 5172 8084
rect 5224 8032 5230 8084
rect 5442 8032 5448 8084
rect 5500 8032 5506 8084
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 5813 8075 5871 8081
rect 5813 8072 5825 8075
rect 5776 8044 5825 8072
rect 5776 8032 5782 8044
rect 5813 8041 5825 8044
rect 5859 8041 5871 8075
rect 8021 8075 8079 8081
rect 8021 8072 8033 8075
rect 5813 8035 5871 8041
rect 6294 8044 8033 8072
rect 3237 7939 3295 7945
rect 3237 7905 3249 7939
rect 3283 7936 3295 7939
rect 3326 7936 3332 7948
rect 3283 7908 3332 7936
rect 3283 7905 3295 7908
rect 3237 7899 3295 7905
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 3973 7939 4031 7945
rect 3436 7908 3740 7936
rect 3436 7880 3464 7908
rect 3712 7895 3740 7908
rect 3973 7905 3985 7939
rect 4019 7936 4031 7939
rect 4798 7936 4804 7948
rect 4019 7908 4804 7936
rect 4019 7905 4031 7908
rect 3973 7899 4031 7905
rect 4798 7896 4804 7908
rect 4856 7896 4862 7948
rect 5184 7936 5212 8032
rect 5350 7964 5356 8016
rect 5408 8004 5414 8016
rect 6294 8004 6322 8044
rect 8021 8041 8033 8044
rect 8067 8041 8079 8075
rect 12250 8072 12256 8084
rect 8021 8035 8079 8041
rect 8404 8044 11100 8072
rect 5408 7976 6322 8004
rect 5408 7964 5414 7976
rect 8404 7948 8432 8044
rect 10502 7964 10508 8016
rect 10560 8004 10566 8016
rect 11072 8013 11100 8044
rect 11624 8044 12256 8072
rect 11057 8007 11115 8013
rect 10560 7976 10824 8004
rect 10560 7964 10566 7976
rect 5629 7939 5687 7945
rect 5629 7936 5641 7939
rect 5184 7908 5641 7936
rect 5629 7905 5641 7908
rect 5675 7936 5687 7939
rect 5902 7936 5908 7948
rect 5675 7908 5908 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 5902 7896 5908 7908
rect 5960 7896 5966 7948
rect 5994 7896 6000 7948
rect 6052 7896 6058 7948
rect 8386 7936 8392 7948
rect 6196 7908 8392 7936
rect 3712 7889 3774 7895
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1394 7877 1400 7880
rect 1029 7871 1087 7877
rect 1029 7868 1041 7871
rect 900 7840 1041 7868
rect 900 7828 906 7840
rect 1029 7837 1041 7840
rect 1075 7837 1087 7871
rect 1029 7831 1087 7837
rect 1356 7871 1400 7877
rect 1356 7837 1368 7871
rect 1356 7831 1400 7837
rect 1394 7828 1400 7831
rect 1452 7828 1458 7880
rect 1535 7871 1593 7877
rect 1535 7837 1547 7871
rect 1581 7868 1593 7871
rect 1670 7868 1676 7880
rect 1581 7840 1676 7868
rect 1581 7837 1593 7840
rect 1535 7831 1593 7837
rect 1670 7828 1676 7840
rect 1728 7828 1734 7880
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7868 1823 7871
rect 2590 7868 2596 7880
rect 1811 7840 2596 7868
rect 1811 7837 1823 7840
rect 1765 7831 1823 7837
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 3418 7828 3424 7880
rect 3476 7828 3482 7880
rect 3602 7877 3608 7880
rect 3564 7871 3608 7877
rect 3564 7837 3576 7871
rect 3564 7831 3608 7837
rect 3602 7828 3608 7831
rect 3660 7828 3666 7880
rect 3712 7858 3728 7889
rect 3716 7855 3728 7858
rect 3762 7855 3774 7889
rect 6196 7877 6224 7908
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 10796 7945 10824 7976
rect 11057 7973 11069 8007
rect 11103 7973 11115 8007
rect 11057 7967 11115 7973
rect 10781 7939 10839 7945
rect 9048 7908 10732 7936
rect 3716 7849 3774 7855
rect 6181 7871 6239 7877
rect 6181 7837 6193 7871
rect 6227 7837 6239 7871
rect 6181 7831 6239 7837
rect 5902 7760 5908 7812
rect 5960 7800 5966 7812
rect 6196 7800 6224 7831
rect 6362 7828 6368 7880
rect 6420 7868 6426 7880
rect 6730 7879 6736 7880
rect 6508 7871 6566 7877
rect 6508 7868 6520 7871
rect 6420 7840 6520 7868
rect 6420 7828 6426 7840
rect 6508 7837 6520 7840
rect 6554 7837 6566 7871
rect 6508 7831 6566 7837
rect 6687 7873 6736 7879
rect 6687 7839 6699 7873
rect 6733 7839 6736 7873
rect 6687 7833 6736 7839
rect 6730 7828 6736 7833
rect 6788 7828 6794 7880
rect 6914 7828 6920 7880
rect 6972 7828 6978 7880
rect 8754 7877 8760 7880
rect 8716 7871 8760 7877
rect 8716 7837 8728 7871
rect 8716 7831 8760 7837
rect 8754 7828 8760 7831
rect 8812 7828 8818 7880
rect 8895 7871 8953 7877
rect 8895 7837 8907 7871
rect 8941 7868 8953 7871
rect 9048 7868 9076 7908
rect 8941 7840 9076 7868
rect 9125 7871 9183 7877
rect 8941 7837 8953 7840
rect 8895 7831 8953 7837
rect 9125 7837 9137 7871
rect 9171 7868 9183 7871
rect 9306 7868 9312 7880
rect 9171 7840 9312 7868
rect 9171 7837 9183 7840
rect 9125 7831 9183 7837
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 5960 7772 6224 7800
rect 5960 7760 5966 7772
rect 10594 7760 10600 7812
rect 10652 7760 10658 7812
rect 10704 7800 10732 7908
rect 10781 7905 10793 7939
rect 10827 7905 10839 7939
rect 10781 7899 10839 7905
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 11624 7877 11652 8044
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 13446 8032 13452 8084
rect 13504 8032 13510 8084
rect 13814 8032 13820 8084
rect 13872 8032 13878 8084
rect 14090 8032 14096 8084
rect 14148 8072 14154 8084
rect 14283 8075 14341 8081
rect 14283 8072 14295 8075
rect 14148 8044 14295 8072
rect 14148 8032 14154 8044
rect 14283 8041 14295 8044
rect 14329 8041 14341 8075
rect 14283 8035 14341 8041
rect 14550 8032 14556 8084
rect 14608 8072 14614 8084
rect 16114 8072 16120 8084
rect 14608 8044 16120 8072
rect 14608 8032 14614 8044
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 16206 8032 16212 8084
rect 16264 8072 16270 8084
rect 16264 8044 17632 8072
rect 16264 8032 16270 8044
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 11936 7939 11994 7945
rect 11936 7936 11948 7939
rect 11756 7908 11948 7936
rect 11756 7896 11762 7908
rect 11936 7905 11948 7908
rect 11982 7905 11994 7939
rect 13832 7936 13860 8032
rect 16022 7964 16028 8016
rect 16080 8004 16086 8016
rect 16945 8007 17003 8013
rect 16945 8004 16957 8007
rect 16080 7976 16957 8004
rect 16080 7964 16086 7976
rect 16945 7973 16957 7976
rect 16991 7973 17003 8007
rect 16945 7967 17003 7973
rect 17494 7964 17500 8016
rect 17552 7964 17558 8016
rect 17604 7948 17632 8044
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 18515 8075 18573 8081
rect 18515 8072 18527 8075
rect 18196 8044 18527 8072
rect 18196 8032 18202 8044
rect 18515 8041 18527 8044
rect 18561 8041 18573 8075
rect 18515 8035 18573 8041
rect 19886 8032 19892 8084
rect 19944 8032 19950 8084
rect 20438 8032 20444 8084
rect 20496 8032 20502 8084
rect 21269 8075 21327 8081
rect 21269 8041 21281 8075
rect 21315 8072 21327 8075
rect 21450 8072 21456 8084
rect 21315 8044 21456 8072
rect 21315 8041 21327 8044
rect 21269 8035 21327 8041
rect 21450 8032 21456 8044
rect 21508 8032 21514 8084
rect 21560 8044 23520 8072
rect 21560 8004 21588 8044
rect 20548 7976 21588 8004
rect 23492 8004 23520 8044
rect 23566 8032 23572 8084
rect 23624 8032 23630 8084
rect 25961 8075 26019 8081
rect 25961 8072 25973 8075
rect 23676 8044 25973 8072
rect 23676 8004 23704 8044
rect 25961 8041 25973 8044
rect 26007 8041 26019 8075
rect 28166 8072 28172 8084
rect 25961 8035 26019 8041
rect 27724 8044 28172 8072
rect 23492 7976 23704 8004
rect 11936 7899 11994 7905
rect 12268 7908 13860 7936
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 11296 7840 11345 7868
rect 11296 7828 11302 7840
rect 11333 7837 11345 7840
rect 11379 7868 11391 7871
rect 11609 7871 11667 7877
rect 11609 7868 11621 7871
rect 11379 7840 11621 7868
rect 11379 7837 11391 7840
rect 11333 7831 11391 7837
rect 11609 7837 11621 7840
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 12115 7871 12173 7877
rect 12115 7837 12127 7871
rect 12161 7868 12173 7871
rect 12268 7868 12296 7908
rect 14550 7896 14556 7948
rect 14608 7896 14614 7948
rect 16390 7896 16396 7948
rect 16448 7896 16454 7948
rect 17586 7896 17592 7948
rect 17644 7896 17650 7948
rect 17770 7896 17776 7948
rect 17828 7936 17834 7948
rect 18049 7939 18107 7945
rect 18049 7936 18061 7939
rect 17828 7908 18061 7936
rect 17828 7896 17834 7908
rect 18049 7905 18061 7908
rect 18095 7905 18107 7939
rect 20548 7936 20576 7976
rect 18049 7899 18107 7905
rect 18708 7908 20576 7936
rect 20625 7939 20683 7945
rect 12161 7840 12296 7868
rect 12345 7871 12403 7877
rect 12161 7837 12173 7840
rect 12115 7831 12173 7837
rect 12345 7837 12357 7871
rect 12391 7868 12403 7871
rect 12391 7840 13768 7868
rect 12391 7837 12403 7840
rect 12345 7831 12403 7837
rect 10704 7772 11284 7800
rect 2869 7735 2927 7741
rect 2869 7701 2881 7735
rect 2915 7732 2927 7735
rect 2958 7732 2964 7744
rect 2915 7704 2964 7732
rect 2915 7701 2927 7704
rect 2869 7695 2927 7701
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 5077 7735 5135 7741
rect 5077 7701 5089 7735
rect 5123 7732 5135 7735
rect 5166 7732 5172 7744
rect 5123 7704 5172 7732
rect 5123 7701 5135 7704
rect 5077 7695 5135 7701
rect 5166 7692 5172 7704
rect 5224 7692 5230 7744
rect 6546 7692 6552 7744
rect 6604 7732 6610 7744
rect 9766 7732 9772 7744
rect 6604 7704 9772 7732
rect 6604 7692 6610 7704
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 10226 7692 10232 7744
rect 10284 7692 10290 7744
rect 11256 7732 11284 7772
rect 13170 7732 13176 7744
rect 11256 7704 13176 7732
rect 13170 7692 13176 7704
rect 13228 7692 13234 7744
rect 13740 7732 13768 7840
rect 13814 7828 13820 7880
rect 13872 7828 13878 7880
rect 14323 7871 14381 7877
rect 14323 7837 14335 7871
rect 14369 7868 14381 7871
rect 15286 7868 15292 7880
rect 14369 7840 15292 7868
rect 14369 7837 14381 7840
rect 14323 7831 14381 7837
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 16758 7828 16764 7880
rect 16816 7868 16822 7880
rect 17954 7868 17960 7880
rect 16816 7840 17960 7868
rect 16816 7828 16822 7840
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 18555 7873 18613 7879
rect 18555 7839 18567 7873
rect 18601 7868 18613 7873
rect 18708 7868 18736 7908
rect 20625 7905 20637 7939
rect 20671 7936 20683 7939
rect 20898 7936 20904 7948
rect 20671 7908 20904 7936
rect 20671 7905 20683 7908
rect 20625 7899 20683 7905
rect 20898 7896 20904 7908
rect 20956 7896 20962 7948
rect 21450 7945 21456 7948
rect 21085 7939 21143 7945
rect 21085 7905 21097 7939
rect 21131 7905 21143 7939
rect 21085 7899 21143 7905
rect 21429 7939 21456 7945
rect 21429 7905 21441 7939
rect 21429 7899 21456 7905
rect 18601 7840 18736 7868
rect 18601 7839 18613 7840
rect 18555 7833 18613 7839
rect 18782 7828 18788 7880
rect 18840 7828 18846 7880
rect 16114 7800 16120 7812
rect 15212 7772 16120 7800
rect 15212 7732 15240 7772
rect 16114 7760 16120 7772
rect 16172 7760 16178 7812
rect 17681 7803 17739 7809
rect 17681 7800 17693 7803
rect 16500 7772 17693 7800
rect 16500 7744 16528 7772
rect 17681 7769 17693 7772
rect 17727 7769 17739 7803
rect 21100 7800 21128 7899
rect 21450 7896 21456 7899
rect 21508 7896 21514 7948
rect 21634 7896 21640 7948
rect 21692 7936 21698 7948
rect 22281 7939 22339 7945
rect 22281 7936 22293 7939
rect 21692 7908 22293 7936
rect 21692 7896 21698 7908
rect 22281 7905 22293 7908
rect 22327 7905 22339 7939
rect 22281 7899 22339 7905
rect 22554 7896 22560 7948
rect 22612 7936 22618 7948
rect 26421 7939 26479 7945
rect 22612 7908 24627 7936
rect 22612 7896 22618 7908
rect 21545 7871 21603 7877
rect 21545 7837 21557 7871
rect 21591 7868 21603 7871
rect 21726 7868 21732 7880
rect 21591 7840 21732 7868
rect 21591 7837 21603 7840
rect 21545 7831 21603 7837
rect 21174 7800 21180 7812
rect 21100 7772 21180 7800
rect 17681 7763 17739 7769
rect 21174 7760 21180 7772
rect 21232 7760 21238 7812
rect 21450 7760 21456 7812
rect 21508 7800 21514 7812
rect 21560 7800 21588 7831
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 21910 7877 21916 7880
rect 21872 7871 21916 7877
rect 21872 7837 21884 7871
rect 21872 7831 21916 7837
rect 21910 7828 21916 7831
rect 21968 7828 21974 7880
rect 22002 7828 22008 7880
rect 22060 7877 22066 7880
rect 22060 7871 22109 7877
rect 22060 7837 22063 7871
rect 22097 7868 22109 7871
rect 22097 7840 22153 7868
rect 22097 7837 22109 7840
rect 22060 7831 22109 7837
rect 22060 7828 22066 7831
rect 23658 7828 23664 7880
rect 23716 7868 23722 7880
rect 24486 7877 24492 7880
rect 24121 7871 24179 7877
rect 24121 7868 24133 7871
rect 23716 7840 24133 7868
rect 23716 7828 23722 7840
rect 24121 7837 24133 7840
rect 24167 7837 24179 7871
rect 24121 7831 24179 7837
rect 24448 7871 24492 7877
rect 24448 7837 24460 7871
rect 24448 7831 24492 7837
rect 24486 7828 24492 7831
rect 24544 7828 24550 7880
rect 24599 7879 24627 7908
rect 26421 7905 26433 7939
rect 26467 7936 26479 7939
rect 26602 7936 26608 7948
rect 26467 7908 26608 7936
rect 26467 7905 26479 7908
rect 26421 7899 26479 7905
rect 26602 7896 26608 7908
rect 26660 7896 26666 7948
rect 27614 7896 27620 7948
rect 27672 7896 27678 7948
rect 27724 7945 27752 8044
rect 28166 8032 28172 8044
rect 28224 8072 28230 8084
rect 28626 8072 28632 8084
rect 28224 8044 28632 8072
rect 28224 8032 28230 8044
rect 28626 8032 28632 8044
rect 28684 8032 28690 8084
rect 28902 8032 28908 8084
rect 28960 8072 28966 8084
rect 29641 8075 29699 8081
rect 29641 8072 29653 8075
rect 28960 8044 29653 8072
rect 28960 8032 28966 8044
rect 29641 8041 29653 8044
rect 29687 8041 29699 8075
rect 29641 8035 29699 8041
rect 30190 8032 30196 8084
rect 30248 8032 30254 8084
rect 27890 7964 27896 8016
rect 27948 7964 27954 8016
rect 27709 7939 27767 7945
rect 27709 7905 27721 7939
rect 27755 7905 27767 7939
rect 27908 7936 27936 7964
rect 28128 7939 28186 7945
rect 28128 7936 28140 7939
rect 27908 7908 28140 7936
rect 27709 7899 27767 7905
rect 28128 7905 28140 7908
rect 28174 7905 28186 7939
rect 28128 7899 28186 7905
rect 28442 7896 28448 7948
rect 28500 7896 28506 7948
rect 28537 7939 28595 7945
rect 28537 7905 28549 7939
rect 28583 7936 28595 7939
rect 30098 7936 30104 7948
rect 28583 7908 30104 7936
rect 28583 7905 28595 7908
rect 28537 7899 28595 7905
rect 30098 7896 30104 7908
rect 30156 7896 30162 7948
rect 30208 7936 30236 8032
rect 30285 7939 30343 7945
rect 30285 7936 30297 7939
rect 30208 7908 30297 7936
rect 30285 7905 30297 7908
rect 30331 7905 30343 7939
rect 30285 7899 30343 7905
rect 30561 7939 30619 7945
rect 30561 7905 30573 7939
rect 30607 7905 30619 7939
rect 30561 7899 30619 7905
rect 24584 7873 24642 7879
rect 24584 7839 24596 7873
rect 24630 7839 24642 7873
rect 24584 7833 24642 7839
rect 24857 7871 24915 7877
rect 24857 7837 24869 7871
rect 24903 7868 24915 7871
rect 26697 7871 26755 7877
rect 24903 7840 26559 7868
rect 24903 7837 24915 7840
rect 24857 7831 24915 7837
rect 21508 7772 21588 7800
rect 26531 7800 26559 7840
rect 26697 7837 26709 7871
rect 26743 7868 26755 7871
rect 26786 7868 26792 7880
rect 26743 7840 26792 7868
rect 26743 7837 26755 7840
rect 26697 7831 26755 7837
rect 26786 7828 26792 7840
rect 26844 7828 26850 7880
rect 27632 7868 27660 7896
rect 27798 7868 27804 7880
rect 27632 7840 27804 7868
rect 27798 7828 27804 7840
rect 27856 7828 27862 7880
rect 28307 7871 28365 7877
rect 28307 7837 28319 7871
rect 28353 7868 28365 7871
rect 28460 7868 28488 7896
rect 28353 7840 28488 7868
rect 28353 7837 28365 7840
rect 28307 7831 28365 7837
rect 28994 7828 29000 7880
rect 29052 7868 29058 7880
rect 29546 7868 29552 7880
rect 29052 7840 29552 7868
rect 29052 7828 29058 7840
rect 29546 7828 29552 7840
rect 29604 7868 29610 7880
rect 30576 7868 30604 7899
rect 29604 7840 30604 7868
rect 29604 7828 29610 7840
rect 30377 7803 30435 7809
rect 30377 7800 30389 7803
rect 26531 7772 27844 7800
rect 21508 7760 21514 7772
rect 13740 7704 15240 7732
rect 15286 7692 15292 7744
rect 15344 7732 15350 7744
rect 15657 7735 15715 7741
rect 15657 7732 15669 7735
rect 15344 7704 15669 7732
rect 15344 7692 15350 7704
rect 15657 7701 15669 7704
rect 15703 7701 15715 7735
rect 15657 7695 15715 7701
rect 16482 7692 16488 7744
rect 16540 7692 16546 7744
rect 16669 7735 16727 7741
rect 16669 7701 16681 7735
rect 16715 7732 16727 7735
rect 16758 7732 16764 7744
rect 16715 7704 16764 7732
rect 16715 7701 16727 7704
rect 16669 7695 16727 7701
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 16942 7692 16948 7744
rect 17000 7732 17006 7744
rect 17037 7735 17095 7741
rect 17037 7732 17049 7735
rect 17000 7704 17049 7732
rect 17000 7692 17006 7704
rect 17037 7701 17049 7704
rect 17083 7701 17095 7735
rect 17037 7695 17095 7701
rect 18598 7692 18604 7744
rect 18656 7732 18662 7744
rect 20806 7732 20812 7744
rect 18656 7704 20812 7732
rect 18656 7692 18662 7704
rect 20806 7692 20812 7704
rect 20864 7692 20870 7744
rect 20901 7735 20959 7741
rect 20901 7701 20913 7735
rect 20947 7732 20959 7735
rect 21542 7732 21548 7744
rect 20947 7704 21548 7732
rect 20947 7701 20959 7704
rect 20901 7695 20959 7701
rect 21542 7692 21548 7704
rect 21600 7692 21606 7744
rect 21726 7692 21732 7744
rect 21784 7732 21790 7744
rect 24670 7732 24676 7744
rect 21784 7704 24676 7732
rect 21784 7692 21790 7704
rect 24670 7692 24676 7704
rect 24728 7692 24734 7744
rect 24762 7692 24768 7744
rect 24820 7732 24826 7744
rect 27430 7732 27436 7744
rect 24820 7704 27436 7732
rect 24820 7692 24826 7704
rect 27430 7692 27436 7704
rect 27488 7692 27494 7744
rect 27522 7692 27528 7744
rect 27580 7692 27586 7744
rect 27816 7732 27844 7772
rect 29196 7772 30389 7800
rect 28442 7732 28448 7744
rect 27816 7704 28448 7732
rect 28442 7692 28448 7704
rect 28500 7692 28506 7744
rect 28626 7692 28632 7744
rect 28684 7732 28690 7744
rect 29196 7732 29224 7772
rect 30377 7769 30389 7772
rect 30423 7769 30435 7803
rect 30377 7763 30435 7769
rect 28684 7704 29224 7732
rect 28684 7692 28690 7704
rect 30098 7692 30104 7744
rect 30156 7692 30162 7744
rect 552 7642 30912 7664
rect 552 7590 4193 7642
rect 4245 7590 4257 7642
rect 4309 7590 4321 7642
rect 4373 7590 4385 7642
rect 4437 7590 4449 7642
rect 4501 7590 11783 7642
rect 11835 7590 11847 7642
rect 11899 7590 11911 7642
rect 11963 7590 11975 7642
rect 12027 7590 12039 7642
rect 12091 7590 19373 7642
rect 19425 7590 19437 7642
rect 19489 7590 19501 7642
rect 19553 7590 19565 7642
rect 19617 7590 19629 7642
rect 19681 7590 26963 7642
rect 27015 7590 27027 7642
rect 27079 7590 27091 7642
rect 27143 7590 27155 7642
rect 27207 7590 27219 7642
rect 27271 7590 30912 7642
rect 552 7568 30912 7590
rect 4706 7528 4712 7540
rect 3528 7500 4712 7528
rect 3528 7401 3556 7500
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 6454 7528 6460 7540
rect 4908 7500 6460 7528
rect 4062 7401 4068 7404
rect 1443 7395 1501 7401
rect 1443 7361 1455 7395
rect 1489 7392 1501 7395
rect 3513 7395 3571 7401
rect 1489 7364 2774 7392
rect 1489 7361 1501 7364
rect 1443 7355 1501 7361
rect 842 7284 848 7336
rect 900 7324 906 7336
rect 937 7327 995 7333
rect 937 7324 949 7327
rect 900 7296 949 7324
rect 900 7284 906 7296
rect 937 7293 949 7296
rect 983 7293 995 7327
rect 937 7287 995 7293
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 2406 7324 2412 7336
rect 1719 7296 2412 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 2746 7256 2774 7364
rect 3513 7361 3525 7395
rect 3559 7361 3571 7395
rect 3513 7355 3571 7361
rect 4019 7395 4068 7401
rect 4019 7361 4031 7395
rect 4065 7361 4068 7395
rect 4019 7355 4068 7361
rect 4062 7352 4068 7355
rect 4120 7352 4126 7404
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7392 4307 7395
rect 4908 7392 4936 7500
rect 6454 7488 6460 7500
rect 6512 7488 6518 7540
rect 6914 7488 6920 7540
rect 6972 7528 6978 7540
rect 7929 7531 7987 7537
rect 7929 7528 7941 7531
rect 6972 7500 7941 7528
rect 6972 7488 6978 7500
rect 7929 7497 7941 7500
rect 7975 7497 7987 7531
rect 13081 7531 13139 7537
rect 13081 7528 13093 7531
rect 7929 7491 7987 7497
rect 8036 7500 10364 7528
rect 5350 7420 5356 7472
rect 5408 7420 5414 7472
rect 7190 7420 7196 7472
rect 7248 7460 7254 7472
rect 7466 7460 7472 7472
rect 7248 7432 7472 7460
rect 7248 7420 7254 7432
rect 7466 7420 7472 7432
rect 7524 7420 7530 7472
rect 5902 7392 5908 7404
rect 4295 7364 4936 7392
rect 5736 7364 5908 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 5736 7336 5764 7364
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 6270 7399 6276 7404
rect 6227 7393 6276 7399
rect 6227 7359 6239 7393
rect 6273 7359 6276 7393
rect 6227 7353 6276 7359
rect 6270 7352 6276 7353
rect 6328 7352 6334 7404
rect 8036 7392 8064 7500
rect 10336 7469 10364 7500
rect 10704 7500 13093 7528
rect 10321 7463 10379 7469
rect 10321 7429 10333 7463
rect 10367 7429 10379 7463
rect 10321 7423 10379 7429
rect 6380 7364 8064 7392
rect 2866 7284 2872 7336
rect 2924 7324 2930 7336
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 2924 7296 3433 7324
rect 2924 7284 2930 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 3620 7296 4936 7324
rect 3620 7256 3648 7296
rect 2746 7228 3648 7256
rect 4908 7256 4936 7296
rect 5718 7284 5724 7336
rect 5776 7284 5782 7336
rect 6380 7324 6408 7364
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 8481 7395 8539 7401
rect 8481 7392 8493 7395
rect 8444 7364 8493 7392
rect 8444 7352 8450 7364
rect 8481 7361 8493 7364
rect 8527 7361 8539 7395
rect 8481 7355 8539 7361
rect 8987 7395 9045 7401
rect 8987 7361 8999 7395
rect 9033 7392 9045 7395
rect 10704 7392 10732 7500
rect 13081 7497 13093 7500
rect 13127 7497 13139 7531
rect 15102 7528 15108 7540
rect 13081 7491 13139 7497
rect 14016 7500 15108 7528
rect 10965 7463 11023 7469
rect 10965 7429 10977 7463
rect 11011 7429 11023 7463
rect 10965 7423 11023 7429
rect 9033 7364 10732 7392
rect 10980 7392 11008 7423
rect 14016 7404 14044 7500
rect 15102 7488 15108 7500
rect 15160 7528 15166 7540
rect 15160 7500 17264 7528
rect 15160 7488 15166 7500
rect 14093 7463 14151 7469
rect 14093 7429 14105 7463
rect 14139 7429 14151 7463
rect 14093 7423 14151 7429
rect 11747 7395 11805 7401
rect 10980 7364 11560 7392
rect 9033 7361 9045 7364
rect 8987 7355 9045 7361
rect 5828 7296 6408 7324
rect 5828 7256 5856 7296
rect 6454 7284 6460 7336
rect 6512 7284 6518 7336
rect 6822 7284 6828 7336
rect 6880 7324 6886 7336
rect 8110 7324 8116 7336
rect 6880 7296 8116 7324
rect 6880 7284 6886 7296
rect 8110 7284 8116 7296
rect 8168 7284 8174 7336
rect 8754 7324 8760 7336
rect 8588 7296 8760 7324
rect 8588 7256 8616 7296
rect 8754 7284 8760 7296
rect 8812 7333 8818 7336
rect 8812 7327 8866 7333
rect 8812 7293 8820 7327
rect 8854 7293 8866 7327
rect 8812 7287 8866 7293
rect 8812 7284 8818 7287
rect 9214 7284 9220 7336
rect 9272 7284 9278 7336
rect 10410 7284 10416 7336
rect 10468 7324 10474 7336
rect 10873 7327 10931 7333
rect 10873 7324 10885 7327
rect 10468 7296 10885 7324
rect 10468 7284 10474 7296
rect 10873 7293 10885 7296
rect 10919 7324 10931 7327
rect 10962 7324 10968 7336
rect 10919 7296 10968 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11149 7327 11207 7333
rect 11149 7293 11161 7327
rect 11195 7293 11207 7327
rect 11149 7287 11207 7293
rect 11164 7256 11192 7287
rect 11238 7284 11244 7336
rect 11296 7284 11302 7336
rect 11330 7284 11336 7336
rect 11388 7284 11394 7336
rect 11532 7324 11560 7364
rect 11747 7361 11759 7395
rect 11793 7392 11805 7395
rect 12342 7392 12348 7404
rect 11793 7364 12348 7392
rect 11793 7361 11805 7364
rect 11747 7355 11805 7361
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 13814 7392 13820 7404
rect 13464 7364 13820 7392
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11532 7296 11989 7324
rect 11977 7293 11989 7296
rect 12023 7293 12035 7327
rect 11977 7287 12035 7293
rect 12250 7284 12256 7336
rect 12308 7324 12314 7336
rect 13464 7324 13492 7364
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 13998 7352 14004 7404
rect 14056 7352 14062 7404
rect 14108 7392 14136 7423
rect 14875 7395 14933 7401
rect 14108 7364 14688 7392
rect 12308 7296 13492 7324
rect 13541 7327 13599 7333
rect 12308 7284 12314 7296
rect 13541 7293 13553 7327
rect 13587 7293 13599 7327
rect 13832 7324 13860 7352
rect 13832 7296 14228 7324
rect 13541 7287 13599 7293
rect 11348 7256 11376 7284
rect 4908 7228 5856 7256
rect 7484 7228 8616 7256
rect 9968 7228 11376 7256
rect 1394 7148 1400 7200
rect 1452 7197 1458 7200
rect 1452 7188 1461 7197
rect 1452 7160 1497 7188
rect 1452 7151 1461 7160
rect 1452 7148 1458 7151
rect 2130 7148 2136 7200
rect 2188 7188 2194 7200
rect 2777 7191 2835 7197
rect 2777 7188 2789 7191
rect 2188 7160 2789 7188
rect 2188 7148 2194 7160
rect 2777 7157 2789 7160
rect 2823 7157 2835 7191
rect 2777 7151 2835 7157
rect 3234 7148 3240 7200
rect 3292 7148 3298 7200
rect 3979 7191 4037 7197
rect 3979 7157 3991 7191
rect 4025 7188 4037 7191
rect 5994 7188 6000 7200
rect 4025 7160 6000 7188
rect 4025 7157 4037 7160
rect 3979 7151 4037 7157
rect 5994 7148 6000 7160
rect 6052 7188 6058 7200
rect 6187 7191 6245 7197
rect 6187 7188 6199 7191
rect 6052 7160 6199 7188
rect 6052 7148 6058 7160
rect 6187 7157 6199 7160
rect 6233 7188 6245 7191
rect 6362 7188 6368 7200
rect 6233 7160 6368 7188
rect 6233 7157 6245 7160
rect 6187 7151 6245 7157
rect 6362 7148 6368 7160
rect 6420 7188 6426 7200
rect 7484 7188 7512 7228
rect 6420 7160 7512 7188
rect 6420 7148 6426 7160
rect 7558 7148 7564 7200
rect 7616 7148 7622 7200
rect 8386 7148 8392 7200
rect 8444 7188 8450 7200
rect 9968 7188 9996 7228
rect 12710 7216 12716 7268
rect 12768 7256 12774 7268
rect 13556 7256 13584 7287
rect 12768 7228 13584 7256
rect 13817 7259 13875 7265
rect 12768 7216 12774 7228
rect 13817 7225 13829 7259
rect 13863 7225 13875 7259
rect 14200 7256 14228 7296
rect 14274 7284 14280 7336
rect 14332 7284 14338 7336
rect 14369 7327 14427 7333
rect 14369 7293 14381 7327
rect 14415 7293 14427 7327
rect 14660 7324 14688 7364
rect 14875 7361 14887 7395
rect 14921 7392 14933 7395
rect 15194 7392 15200 7404
rect 14921 7364 15200 7392
rect 14921 7361 14933 7364
rect 14875 7355 14933 7361
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 16574 7352 16580 7404
rect 16632 7392 16638 7404
rect 16632 7364 16896 7392
rect 16632 7352 16638 7364
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 14660 7296 15117 7324
rect 14369 7287 14427 7293
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 14384 7256 14412 7287
rect 16758 7284 16764 7336
rect 16816 7284 16822 7336
rect 16868 7333 16896 7364
rect 16853 7327 16911 7333
rect 16853 7293 16865 7327
rect 16899 7293 16911 7327
rect 17236 7324 17264 7500
rect 17770 7488 17776 7540
rect 17828 7528 17834 7540
rect 17865 7531 17923 7537
rect 17865 7528 17877 7531
rect 17828 7500 17877 7528
rect 17828 7488 17834 7500
rect 17865 7497 17877 7500
rect 17911 7528 17923 7531
rect 18598 7528 18604 7540
rect 17911 7500 18604 7528
rect 17911 7497 17923 7500
rect 17865 7491 17923 7497
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 19794 7488 19800 7540
rect 19852 7528 19858 7540
rect 20533 7531 20591 7537
rect 20533 7528 20545 7531
rect 19852 7500 20545 7528
rect 19852 7488 19858 7500
rect 20533 7497 20545 7500
rect 20579 7497 20591 7531
rect 20533 7491 20591 7497
rect 21358 7488 21364 7540
rect 21416 7528 21422 7540
rect 21818 7528 21824 7540
rect 21416 7500 21824 7528
rect 21416 7488 21422 7500
rect 21818 7488 21824 7500
rect 21876 7488 21882 7540
rect 23569 7531 23627 7537
rect 23569 7497 23581 7531
rect 23615 7528 23627 7531
rect 23750 7528 23756 7540
rect 23615 7500 23756 7528
rect 23615 7497 23627 7500
rect 23569 7491 23627 7497
rect 23750 7488 23756 7500
rect 23808 7488 23814 7540
rect 25130 7488 25136 7540
rect 25188 7528 25194 7540
rect 25188 7500 28120 7528
rect 25188 7488 25194 7500
rect 25866 7420 25872 7472
rect 25924 7420 25930 7472
rect 28092 7469 28120 7500
rect 28442 7488 28448 7540
rect 28500 7488 28506 7540
rect 28077 7463 28135 7469
rect 28077 7429 28089 7463
rect 28123 7429 28135 7463
rect 28077 7423 28135 7429
rect 28718 7420 28724 7472
rect 28776 7460 28782 7472
rect 29273 7463 29331 7469
rect 29273 7460 29285 7463
rect 28776 7432 29285 7460
rect 28776 7420 28782 7432
rect 29273 7429 29285 7432
rect 29319 7429 29331 7463
rect 29273 7423 29331 7429
rect 17494 7352 17500 7404
rect 17552 7392 17558 7404
rect 19199 7395 19257 7401
rect 17552 7364 18828 7392
rect 17552 7352 17558 7364
rect 17405 7327 17463 7333
rect 17405 7324 17417 7327
rect 17236 7296 17417 7324
rect 16853 7287 16911 7293
rect 17405 7293 17417 7296
rect 17451 7293 17463 7327
rect 17405 7287 17463 7293
rect 17589 7327 17647 7333
rect 17589 7293 17601 7327
rect 17635 7324 17647 7327
rect 17862 7324 17868 7336
rect 17635 7296 17868 7324
rect 17635 7293 17647 7296
rect 17589 7287 17647 7293
rect 17862 7284 17868 7296
rect 17920 7284 17926 7336
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 14200 7228 14412 7256
rect 16776 7256 16804 7284
rect 18064 7256 18092 7287
rect 18138 7284 18144 7336
rect 18196 7324 18202 7336
rect 18325 7327 18383 7333
rect 18325 7324 18337 7327
rect 18196 7296 18337 7324
rect 18196 7284 18202 7296
rect 18325 7293 18337 7296
rect 18371 7293 18383 7327
rect 18325 7287 18383 7293
rect 18230 7256 18236 7268
rect 16776 7228 17448 7256
rect 18064 7228 18236 7256
rect 13817 7219 13875 7225
rect 8444 7160 9996 7188
rect 10689 7191 10747 7197
rect 8444 7148 8450 7160
rect 10689 7157 10701 7191
rect 10735 7188 10747 7191
rect 11330 7188 11336 7200
rect 10735 7160 11336 7188
rect 10735 7157 10747 7160
rect 10689 7151 10747 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11698 7148 11704 7200
rect 11756 7197 11762 7200
rect 11756 7188 11765 7197
rect 13832 7188 13860 7219
rect 17420 7200 17448 7228
rect 18230 7216 18236 7228
rect 18288 7216 18294 7268
rect 14090 7188 14096 7200
rect 11756 7160 14096 7188
rect 11756 7151 11765 7160
rect 11756 7148 11762 7151
rect 14090 7148 14096 7160
rect 14148 7188 14154 7200
rect 14734 7188 14740 7200
rect 14148 7160 14740 7188
rect 14148 7148 14154 7160
rect 14734 7148 14740 7160
rect 14792 7188 14798 7200
rect 14835 7191 14893 7197
rect 14835 7188 14847 7191
rect 14792 7160 14847 7188
rect 14792 7148 14798 7160
rect 14835 7157 14847 7160
rect 14881 7157 14893 7191
rect 14835 7151 14893 7157
rect 15194 7148 15200 7200
rect 15252 7188 15258 7200
rect 16209 7191 16267 7197
rect 16209 7188 16221 7191
rect 15252 7160 16221 7188
rect 15252 7148 15258 7160
rect 16209 7157 16221 7160
rect 16255 7157 16267 7191
rect 16209 7151 16267 7157
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 16577 7191 16635 7197
rect 16577 7188 16589 7191
rect 16356 7160 16589 7188
rect 16356 7148 16362 7160
rect 16577 7157 16589 7160
rect 16623 7157 16635 7191
rect 16577 7151 16635 7157
rect 17034 7148 17040 7200
rect 17092 7148 17098 7200
rect 17126 7148 17132 7200
rect 17184 7188 17190 7200
rect 17221 7191 17279 7197
rect 17221 7188 17233 7191
rect 17184 7160 17233 7188
rect 17184 7148 17190 7160
rect 17221 7157 17233 7160
rect 17267 7157 17279 7191
rect 17221 7151 17279 7157
rect 17402 7148 17408 7200
rect 17460 7148 17466 7200
rect 18340 7188 18368 7287
rect 18598 7284 18604 7336
rect 18656 7324 18662 7336
rect 18693 7327 18751 7333
rect 18693 7324 18705 7327
rect 18656 7296 18705 7324
rect 18656 7284 18662 7296
rect 18693 7293 18705 7296
rect 18739 7293 18751 7327
rect 18800 7324 18828 7364
rect 19199 7361 19211 7395
rect 19245 7392 19257 7395
rect 21726 7392 21732 7404
rect 19245 7364 21732 7392
rect 19245 7361 19257 7364
rect 19199 7355 19257 7361
rect 21726 7352 21732 7364
rect 21784 7352 21790 7404
rect 22094 7399 22100 7404
rect 22051 7393 22100 7399
rect 22051 7359 22063 7393
rect 22097 7359 22100 7393
rect 22051 7353 22100 7359
rect 22094 7352 22100 7353
rect 22152 7352 22158 7404
rect 22186 7352 22192 7404
rect 22244 7392 22250 7404
rect 22281 7395 22339 7401
rect 22281 7392 22293 7395
rect 22244 7364 22293 7392
rect 22244 7352 22250 7364
rect 22281 7361 22293 7364
rect 22327 7361 22339 7395
rect 24492 7395 24550 7401
rect 24492 7392 24504 7395
rect 22281 7355 22339 7361
rect 23492 7364 24504 7392
rect 23492 7336 23520 7364
rect 24492 7361 24504 7364
rect 24538 7361 24550 7395
rect 24492 7355 24550 7361
rect 24578 7352 24584 7404
rect 24636 7352 24642 7404
rect 24670 7352 24676 7404
rect 24728 7392 24734 7404
rect 26700 7395 26758 7401
rect 26700 7392 26712 7395
rect 24728 7364 26712 7392
rect 24728 7352 24734 7364
rect 26700 7361 26712 7364
rect 26746 7361 26758 7395
rect 26700 7355 26758 7361
rect 19429 7327 19487 7333
rect 19429 7324 19441 7327
rect 18800 7296 19441 7324
rect 18693 7287 18751 7293
rect 19429 7293 19441 7296
rect 19475 7293 19487 7327
rect 19429 7287 19487 7293
rect 20806 7284 20812 7336
rect 20864 7324 20870 7336
rect 21450 7324 21456 7336
rect 20864 7296 21456 7324
rect 20864 7284 20870 7296
rect 21450 7284 21456 7296
rect 21508 7324 21514 7336
rect 21545 7327 21603 7333
rect 21545 7324 21557 7327
rect 21508 7296 21557 7324
rect 21508 7284 21514 7296
rect 21545 7293 21557 7296
rect 21591 7293 21603 7327
rect 21545 7287 21603 7293
rect 21652 7296 22968 7324
rect 20162 7216 20168 7268
rect 20220 7256 20226 7268
rect 21085 7259 21143 7265
rect 21085 7256 21097 7259
rect 20220 7228 21097 7256
rect 20220 7216 20226 7228
rect 21085 7225 21097 7228
rect 21131 7225 21143 7259
rect 21085 7219 21143 7225
rect 21174 7216 21180 7268
rect 21232 7256 21238 7268
rect 21652 7256 21680 7296
rect 21232 7228 21680 7256
rect 22940 7256 22968 7296
rect 23474 7284 23480 7336
rect 23532 7284 23538 7336
rect 23658 7284 23664 7336
rect 23716 7324 23722 7336
rect 24029 7327 24087 7333
rect 24029 7324 24041 7327
rect 23716 7296 24041 7324
rect 23716 7284 23722 7296
rect 24029 7293 24041 7296
rect 24075 7293 24087 7327
rect 24596 7324 24624 7352
rect 24029 7287 24087 7293
rect 24136 7296 24624 7324
rect 23566 7256 23572 7268
rect 22940 7228 23572 7256
rect 21232 7216 21238 7228
rect 23566 7216 23572 7228
rect 23624 7256 23630 7268
rect 24136 7256 24164 7296
rect 24762 7284 24768 7336
rect 24820 7284 24826 7336
rect 26234 7284 26240 7336
rect 26292 7284 26298 7336
rect 26564 7327 26622 7333
rect 26564 7324 26576 7327
rect 26344 7296 26576 7324
rect 23624 7228 24164 7256
rect 23624 7216 23630 7228
rect 19159 7191 19217 7197
rect 19159 7188 19171 7191
rect 18340 7160 19171 7188
rect 19159 7157 19171 7160
rect 19205 7188 19217 7191
rect 20714 7188 20720 7200
rect 19205 7160 20720 7188
rect 19205 7157 19217 7160
rect 19159 7151 19217 7157
rect 20714 7148 20720 7160
rect 20772 7188 20778 7200
rect 21910 7188 21916 7200
rect 20772 7160 21916 7188
rect 20772 7148 20778 7160
rect 21910 7148 21916 7160
rect 21968 7188 21974 7200
rect 22011 7191 22069 7197
rect 22011 7188 22023 7191
rect 21968 7160 22023 7188
rect 21968 7148 21974 7160
rect 22011 7157 22023 7160
rect 22057 7157 22069 7191
rect 22011 7151 22069 7157
rect 24486 7148 24492 7200
rect 24544 7197 24550 7200
rect 24544 7188 24553 7197
rect 26344 7188 26372 7296
rect 26564 7293 26576 7296
rect 26610 7324 26622 7327
rect 26786 7324 26792 7336
rect 26610 7296 26792 7324
rect 26610 7293 26622 7296
rect 26564 7287 26622 7293
rect 26786 7284 26792 7296
rect 26844 7284 26850 7336
rect 26970 7284 26976 7336
rect 27028 7284 27034 7336
rect 27430 7284 27436 7336
rect 27488 7324 27494 7336
rect 28629 7327 28687 7333
rect 27488 7296 27660 7324
rect 27488 7284 27494 7296
rect 27632 7256 27660 7296
rect 28629 7293 28641 7327
rect 28675 7324 28687 7327
rect 29086 7324 29092 7336
rect 28675 7296 29092 7324
rect 28675 7293 28687 7296
rect 28629 7287 28687 7293
rect 29086 7284 29092 7296
rect 29144 7284 29150 7336
rect 29178 7284 29184 7336
rect 29236 7284 29242 7336
rect 29362 7284 29368 7336
rect 29420 7324 29426 7336
rect 29457 7327 29515 7333
rect 29457 7324 29469 7327
rect 29420 7296 29469 7324
rect 29420 7284 29426 7296
rect 29457 7293 29469 7296
rect 29503 7293 29515 7327
rect 29457 7287 29515 7293
rect 27632 7228 29776 7256
rect 29748 7200 29776 7228
rect 24544 7160 26372 7188
rect 24544 7151 24553 7160
rect 24544 7148 24550 7151
rect 28994 7148 29000 7200
rect 29052 7148 29058 7200
rect 29730 7148 29736 7200
rect 29788 7148 29794 7200
rect 552 7098 31072 7120
rect 552 7046 7988 7098
rect 8040 7046 8052 7098
rect 8104 7046 8116 7098
rect 8168 7046 8180 7098
rect 8232 7046 8244 7098
rect 8296 7046 15578 7098
rect 15630 7046 15642 7098
rect 15694 7046 15706 7098
rect 15758 7046 15770 7098
rect 15822 7046 15834 7098
rect 15886 7046 23168 7098
rect 23220 7046 23232 7098
rect 23284 7046 23296 7098
rect 23348 7046 23360 7098
rect 23412 7046 23424 7098
rect 23476 7046 30758 7098
rect 30810 7046 30822 7098
rect 30874 7046 30886 7098
rect 30938 7046 30950 7098
rect 31002 7046 31014 7098
rect 31066 7046 31072 7098
rect 552 7024 31072 7046
rect 1044 6956 2774 6984
rect 842 6740 848 6792
rect 900 6780 906 6792
rect 1044 6789 1072 6956
rect 2746 6848 2774 6956
rect 3234 6944 3240 6996
rect 3292 6984 3298 6996
rect 4890 6984 4896 6996
rect 3292 6956 4896 6984
rect 3292 6944 3298 6956
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 6270 6944 6276 6996
rect 6328 6984 6334 6996
rect 9398 6984 9404 6996
rect 6328 6956 9404 6984
rect 6328 6944 6334 6956
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 10318 6944 10324 6996
rect 10376 6984 10382 6996
rect 10376 6956 11284 6984
rect 10376 6944 10382 6956
rect 4798 6876 4804 6928
rect 4856 6916 4862 6928
rect 8386 6916 8392 6928
rect 4856 6888 5672 6916
rect 4856 6876 4862 6888
rect 5350 6848 5356 6860
rect 1550 6820 2176 6848
rect 2746 6820 3280 6848
rect 1394 6789 1400 6792
rect 1029 6783 1087 6789
rect 1029 6780 1041 6783
rect 900 6752 1041 6780
rect 900 6740 906 6752
rect 1029 6749 1041 6752
rect 1075 6749 1087 6783
rect 1029 6743 1087 6749
rect 1356 6783 1400 6789
rect 1356 6749 1368 6783
rect 1356 6743 1400 6749
rect 1394 6740 1400 6743
rect 1452 6740 1458 6792
rect 1550 6789 1578 6820
rect 1535 6783 1593 6789
rect 1535 6749 1547 6783
rect 1581 6749 1593 6783
rect 1535 6743 1593 6749
rect 1762 6740 1768 6792
rect 1820 6740 1826 6792
rect 2148 6780 2176 6820
rect 3252 6792 3280 6820
rect 3896 6820 5356 6848
rect 2148 6752 3188 6780
rect 1762 6604 1768 6656
rect 1820 6644 1826 6656
rect 2498 6644 2504 6656
rect 1820 6616 2504 6644
rect 1820 6604 1826 6616
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 2866 6604 2872 6656
rect 2924 6604 2930 6656
rect 3160 6644 3188 6752
rect 3234 6740 3240 6792
rect 3292 6740 3298 6792
rect 3602 6789 3608 6792
rect 3564 6783 3608 6789
rect 3564 6749 3576 6783
rect 3564 6743 3608 6749
rect 3602 6740 3608 6743
rect 3660 6740 3666 6792
rect 3743 6783 3801 6789
rect 3743 6749 3755 6783
rect 3789 6780 3801 6783
rect 3896 6780 3924 6820
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 5644 6857 5672 6888
rect 8220 6888 8392 6916
rect 8220 6857 8248 6888
rect 8386 6876 8392 6888
rect 8444 6876 8450 6928
rect 10704 6888 10916 6916
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6817 5687 6851
rect 8205 6851 8263 6857
rect 5629 6811 5687 6817
rect 5736 6820 7604 6848
rect 3789 6752 3924 6780
rect 3789 6749 3801 6752
rect 3743 6743 3801 6749
rect 3970 6740 3976 6792
rect 4028 6740 4034 6792
rect 5736 6780 5764 6820
rect 7576 6792 7604 6820
rect 8205 6817 8217 6851
rect 8251 6817 8263 6851
rect 8478 6848 8484 6860
rect 8205 6811 8263 6817
rect 8404 6820 8484 6848
rect 4632 6752 5764 6780
rect 5813 6783 5871 6789
rect 4632 6644 4660 6752
rect 5813 6749 5825 6783
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 4706 6672 4712 6724
rect 4764 6712 4770 6724
rect 5718 6712 5724 6724
rect 4764 6684 5724 6712
rect 4764 6672 4770 6684
rect 5718 6672 5724 6684
rect 5776 6712 5782 6724
rect 5828 6712 5856 6743
rect 5994 6740 6000 6792
rect 6052 6780 6058 6792
rect 6362 6789 6368 6792
rect 6140 6783 6198 6789
rect 6140 6780 6152 6783
rect 6052 6752 6152 6780
rect 6052 6740 6058 6752
rect 6140 6749 6152 6752
rect 6186 6749 6198 6783
rect 6140 6743 6198 6749
rect 6319 6783 6368 6789
rect 6319 6749 6331 6783
rect 6365 6749 6368 6783
rect 6319 6743 6368 6749
rect 6362 6740 6368 6743
rect 6420 6740 6426 6792
rect 6546 6740 6552 6792
rect 6604 6740 6610 6792
rect 7558 6740 7564 6792
rect 7616 6740 7622 6792
rect 8404 6789 8432 6820
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 9054 6848 9260 6852
rect 10704 6848 10732 6888
rect 8910 6824 10732 6848
rect 8910 6820 9082 6824
rect 9232 6820 10732 6824
rect 10781 6851 10839 6857
rect 8754 6789 8760 6792
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 8716 6783 8760 6789
rect 8716 6749 8728 6783
rect 8716 6743 8760 6749
rect 8754 6740 8760 6743
rect 8812 6740 8818 6792
rect 8910 6791 8938 6820
rect 10781 6817 10793 6851
rect 10827 6817 10839 6851
rect 10781 6811 10839 6817
rect 8895 6785 8953 6791
rect 8895 6751 8907 6785
rect 8941 6751 8953 6785
rect 8895 6745 8953 6751
rect 9122 6740 9128 6792
rect 9180 6740 9186 6792
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 10226 6780 10232 6792
rect 9548 6752 10232 6780
rect 9548 6740 9554 6752
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 10796 6712 10824 6811
rect 10888 6780 10916 6888
rect 11256 6857 11284 6956
rect 11330 6944 11336 6996
rect 11388 6984 11394 6996
rect 12066 6984 12072 6996
rect 11388 6956 12072 6984
rect 11388 6944 11394 6956
rect 12066 6944 12072 6956
rect 12124 6944 12130 6996
rect 13170 6944 13176 6996
rect 13228 6944 13234 6996
rect 14090 6944 14096 6996
rect 14148 6984 14154 6996
rect 14283 6987 14341 6993
rect 14283 6984 14295 6987
rect 14148 6956 14295 6984
rect 14148 6944 14154 6956
rect 14283 6953 14295 6956
rect 14329 6953 14341 6987
rect 14283 6947 14341 6953
rect 14642 6944 14648 6996
rect 14700 6984 14706 6996
rect 14700 6956 16068 6984
rect 14700 6944 14706 6956
rect 11698 6857 11704 6860
rect 11241 6851 11299 6857
rect 11241 6817 11253 6851
rect 11287 6848 11299 6851
rect 11660 6851 11704 6857
rect 11287 6820 11560 6848
rect 11287 6817 11299 6820
rect 11241 6811 11299 6817
rect 11532 6792 11560 6820
rect 11660 6817 11672 6851
rect 11660 6811 11704 6817
rect 11698 6808 11704 6811
rect 11756 6808 11762 6860
rect 11992 6820 12434 6848
rect 11146 6780 11152 6792
rect 10888 6752 11152 6780
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 11333 6783 11391 6789
rect 11333 6780 11345 6783
rect 11256 6752 11345 6780
rect 11256 6724 11284 6752
rect 11333 6749 11345 6752
rect 11379 6749 11391 6783
rect 11333 6743 11391 6749
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 11839 6783 11897 6789
rect 11839 6749 11851 6783
rect 11885 6780 11897 6783
rect 11992 6780 12020 6820
rect 11885 6752 12020 6780
rect 11885 6749 11897 6752
rect 11839 6743 11897 6749
rect 12066 6740 12072 6792
rect 12124 6740 12130 6792
rect 12406 6780 12434 6820
rect 13538 6808 13544 6860
rect 13596 6808 13602 6860
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 15933 6851 15991 6857
rect 15933 6848 15945 6851
rect 13780 6820 15945 6848
rect 13780 6808 13786 6820
rect 15933 6817 15945 6820
rect 15979 6817 15991 6851
rect 16040 6848 16068 6956
rect 16114 6944 16120 6996
rect 16172 6944 16178 6996
rect 17494 6944 17500 6996
rect 17552 6944 17558 6996
rect 17770 6944 17776 6996
rect 17828 6984 17834 6996
rect 17828 6956 18092 6984
rect 17828 6944 17834 6956
rect 17052 6888 17264 6916
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 16040 6820 16313 6848
rect 15933 6811 15991 6817
rect 16301 6817 16313 6820
rect 16347 6848 16359 6851
rect 16393 6851 16451 6857
rect 16393 6848 16405 6851
rect 16347 6820 16405 6848
rect 16347 6817 16359 6820
rect 16301 6811 16359 6817
rect 16393 6817 16405 6820
rect 16439 6848 16451 6851
rect 16482 6848 16488 6860
rect 16439 6820 16488 6848
rect 16439 6817 16451 6820
rect 16393 6811 16451 6817
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 16669 6851 16727 6857
rect 16669 6848 16681 6851
rect 16632 6820 16681 6848
rect 16632 6808 16638 6820
rect 16669 6817 16681 6820
rect 16715 6817 16727 6851
rect 16669 6811 16727 6817
rect 16758 6808 16764 6860
rect 16816 6848 16822 6860
rect 16945 6851 17003 6857
rect 16945 6848 16957 6851
rect 16816 6820 16957 6848
rect 16816 6808 16822 6820
rect 16945 6817 16957 6820
rect 16991 6848 17003 6851
rect 17052 6848 17080 6888
rect 16991 6820 17080 6848
rect 16991 6817 17003 6820
rect 16945 6811 17003 6817
rect 17126 6808 17132 6860
rect 17184 6808 17190 6860
rect 12802 6780 12808 6792
rect 12406 6752 12808 6780
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 13814 6740 13820 6792
rect 13872 6740 13878 6792
rect 14323 6783 14381 6789
rect 14323 6749 14335 6783
rect 14369 6780 14381 6783
rect 14458 6780 14464 6792
rect 14369 6752 14464 6780
rect 14369 6749 14381 6752
rect 14323 6743 14381 6749
rect 14458 6740 14464 6752
rect 14516 6740 14522 6792
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 17144 6780 17172 6808
rect 14599 6752 17172 6780
rect 17236 6780 17264 6888
rect 17696 6888 17908 6916
rect 17310 6808 17316 6860
rect 17368 6848 17374 6860
rect 17696 6857 17724 6888
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 17368 6820 17417 6848
rect 17368 6808 17374 6820
rect 17405 6817 17417 6820
rect 17451 6817 17463 6851
rect 17405 6811 17463 6817
rect 17681 6851 17739 6857
rect 17681 6817 17693 6851
rect 17727 6817 17739 6851
rect 17681 6811 17739 6817
rect 17773 6851 17831 6857
rect 17773 6817 17785 6851
rect 17819 6817 17831 6851
rect 17773 6811 17831 6817
rect 17788 6780 17816 6811
rect 17880 6792 17908 6888
rect 18064 6857 18092 6956
rect 18138 6944 18144 6996
rect 18196 6984 18202 6996
rect 18515 6987 18573 6993
rect 18515 6984 18527 6987
rect 18196 6956 18527 6984
rect 18196 6944 18202 6956
rect 18515 6953 18527 6956
rect 18561 6953 18573 6987
rect 18515 6947 18573 6953
rect 20898 6944 20904 6996
rect 20956 6984 20962 6996
rect 22002 6984 22008 6996
rect 20956 6956 22008 6984
rect 20956 6944 20962 6956
rect 22002 6944 22008 6956
rect 22060 6944 22066 6996
rect 23658 6944 23664 6996
rect 23716 6984 23722 6996
rect 26234 6984 26240 6996
rect 23716 6956 26240 6984
rect 23716 6944 23722 6956
rect 26234 6944 26240 6956
rect 26292 6944 26298 6996
rect 26421 6987 26479 6993
rect 26421 6953 26433 6987
rect 26467 6984 26479 6987
rect 26970 6984 26976 6996
rect 26467 6956 26976 6984
rect 26467 6953 26479 6956
rect 26421 6947 26479 6953
rect 26970 6944 26976 6956
rect 27028 6944 27034 6996
rect 27890 6944 27896 6996
rect 27948 6984 27954 6996
rect 28267 6987 28325 6993
rect 28267 6984 28279 6987
rect 27948 6956 28279 6984
rect 27948 6944 27954 6956
rect 28267 6953 28279 6956
rect 28313 6953 28325 6987
rect 28267 6947 28325 6953
rect 26252 6916 26280 6944
rect 26694 6916 26700 6928
rect 20640 6888 21128 6916
rect 26252 6888 26700 6916
rect 18049 6851 18107 6857
rect 18049 6817 18061 6851
rect 18095 6817 18107 6851
rect 18524 6848 18736 6852
rect 19242 6848 19248 6860
rect 18049 6811 18107 6817
rect 18340 6824 19248 6848
rect 18340 6820 18552 6824
rect 18708 6820 19248 6824
rect 17236 6752 17816 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 17862 6740 17868 6792
rect 17920 6740 17926 6792
rect 18230 6740 18236 6792
rect 18288 6780 18294 6792
rect 18340 6780 18368 6820
rect 19242 6808 19248 6820
rect 19300 6848 19306 6860
rect 20441 6851 20499 6857
rect 20441 6848 20453 6851
rect 19300 6820 20453 6848
rect 19300 6808 19306 6820
rect 20441 6817 20453 6820
rect 20487 6848 20499 6851
rect 20640 6848 20668 6888
rect 20487 6820 20668 6848
rect 20717 6851 20775 6857
rect 20487 6817 20499 6820
rect 20441 6811 20499 6817
rect 20717 6817 20729 6851
rect 20763 6848 20775 6851
rect 20993 6851 21051 6857
rect 20993 6848 21005 6851
rect 20763 6820 21005 6848
rect 20763 6817 20775 6820
rect 20717 6811 20775 6817
rect 20993 6817 21005 6820
rect 21039 6817 21051 6851
rect 21100 6848 21128 6888
rect 26694 6876 26700 6888
rect 26752 6916 26758 6928
rect 27341 6919 27399 6925
rect 27341 6916 27353 6919
rect 26752 6888 27353 6916
rect 26752 6876 26758 6888
rect 27341 6885 27353 6888
rect 27387 6916 27399 6919
rect 27430 6916 27436 6928
rect 27387 6888 27436 6916
rect 27387 6885 27399 6888
rect 27341 6879 27399 6885
rect 27430 6876 27436 6888
rect 27488 6876 27494 6928
rect 21266 6848 21272 6860
rect 21100 6820 21272 6848
rect 20993 6811 21051 6817
rect 18598 6791 18604 6792
rect 18288 6752 18368 6780
rect 18555 6785 18604 6791
rect 18288 6740 18294 6752
rect 18555 6751 18567 6785
rect 18601 6751 18604 6785
rect 18555 6745 18604 6751
rect 18598 6740 18604 6745
rect 18656 6740 18662 6792
rect 18690 6740 18696 6792
rect 18748 6780 18754 6792
rect 18785 6783 18843 6789
rect 18785 6780 18797 6783
rect 18748 6752 18797 6780
rect 18748 6740 18754 6752
rect 18785 6749 18797 6752
rect 18831 6749 18843 6783
rect 18785 6743 18843 6749
rect 5776 6684 5856 6712
rect 9784 6684 10824 6712
rect 5776 6672 5782 6684
rect 3160 6616 4660 6644
rect 5074 6604 5080 6656
rect 5132 6604 5138 6656
rect 5442 6604 5448 6656
rect 5500 6604 5506 6656
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 6270 6644 6276 6656
rect 5868 6616 6276 6644
rect 5868 6604 5874 6616
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 7650 6604 7656 6656
rect 7708 6604 7714 6656
rect 8021 6647 8079 6653
rect 8021 6613 8033 6647
rect 8067 6644 8079 6647
rect 9214 6644 9220 6656
rect 8067 6616 9220 6644
rect 8067 6613 8079 6616
rect 8021 6607 8079 6613
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 9582 6604 9588 6656
rect 9640 6644 9646 6656
rect 9784 6644 9812 6684
rect 11238 6672 11244 6724
rect 11296 6672 11302 6724
rect 15470 6672 15476 6724
rect 15528 6672 15534 6724
rect 19702 6672 19708 6724
rect 19760 6712 19766 6724
rect 19889 6715 19947 6721
rect 19889 6712 19901 6715
rect 19760 6684 19901 6712
rect 19760 6672 19766 6684
rect 19889 6681 19901 6684
rect 19935 6681 19947 6715
rect 20732 6712 20760 6811
rect 21008 6780 21036 6811
rect 21266 6808 21272 6820
rect 21324 6848 21330 6860
rect 21453 6851 21511 6857
rect 21453 6848 21465 6851
rect 21324 6820 21465 6848
rect 21324 6808 21330 6820
rect 21453 6817 21465 6820
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 21542 6808 21548 6860
rect 21600 6848 21606 6860
rect 22465 6851 22523 6857
rect 22465 6848 22477 6851
rect 21600 6820 22477 6848
rect 21600 6808 21606 6820
rect 22465 6817 22477 6820
rect 22511 6817 22523 6851
rect 22465 6811 22523 6817
rect 23845 6851 23903 6857
rect 23845 6817 23857 6851
rect 23891 6848 23903 6851
rect 24118 6848 24124 6860
rect 23891 6820 24124 6848
rect 23891 6817 23903 6820
rect 23845 6811 23903 6817
rect 24118 6808 24124 6820
rect 24176 6808 24182 6860
rect 24356 6851 24414 6857
rect 24356 6817 24368 6851
rect 24402 6848 24414 6851
rect 26605 6851 26663 6857
rect 24402 6820 24716 6848
rect 24402 6817 24414 6820
rect 24356 6811 24414 6817
rect 24688 6792 24716 6820
rect 26605 6817 26617 6851
rect 26651 6817 26663 6851
rect 28537 6851 28595 6857
rect 26605 6811 26663 6817
rect 27448 6820 28028 6848
rect 21174 6780 21180 6792
rect 21008 6752 21180 6780
rect 21174 6740 21180 6752
rect 21232 6740 21238 6792
rect 21358 6740 21364 6792
rect 21416 6780 21422 6792
rect 21729 6783 21787 6789
rect 21729 6780 21741 6783
rect 21416 6752 21741 6780
rect 21416 6740 21422 6752
rect 21729 6749 21741 6752
rect 21775 6749 21787 6783
rect 21729 6743 21787 6749
rect 21910 6740 21916 6792
rect 21968 6780 21974 6792
rect 22056 6783 22114 6789
rect 22056 6780 22068 6783
rect 21968 6752 22068 6780
rect 21968 6740 21974 6752
rect 22056 6749 22068 6752
rect 22102 6749 22114 6783
rect 22056 6743 22114 6749
rect 22235 6783 22293 6789
rect 22235 6749 22247 6783
rect 22281 6780 22293 6783
rect 23382 6780 23388 6792
rect 22281 6752 23388 6780
rect 22281 6749 22293 6752
rect 22235 6743 22293 6749
rect 23382 6740 23388 6752
rect 23440 6740 23446 6792
rect 24026 6740 24032 6792
rect 24084 6789 24090 6792
rect 24084 6780 24095 6789
rect 24084 6752 24129 6780
rect 24084 6743 24095 6752
rect 24084 6740 24090 6743
rect 24486 6740 24492 6792
rect 24544 6740 24550 6792
rect 24670 6740 24676 6792
rect 24728 6740 24734 6792
rect 24765 6783 24823 6789
rect 24765 6749 24777 6783
rect 24811 6780 24823 6783
rect 25958 6780 25964 6792
rect 24811 6752 25964 6780
rect 24811 6749 24823 6752
rect 24765 6743 24823 6749
rect 25958 6740 25964 6752
rect 26016 6740 26022 6792
rect 26620 6780 26648 6811
rect 27448 6780 27476 6820
rect 28000 6792 28028 6820
rect 28537 6817 28549 6851
rect 28583 6848 28595 6851
rect 30282 6848 30288 6860
rect 28583 6820 30288 6848
rect 28583 6817 28595 6820
rect 28537 6811 28595 6817
rect 30282 6808 30288 6820
rect 30340 6808 30346 6860
rect 26620 6752 27476 6780
rect 27798 6740 27804 6792
rect 27856 6740 27862 6792
rect 27982 6740 27988 6792
rect 28040 6740 28046 6792
rect 28258 6740 28264 6792
rect 28316 6780 28322 6792
rect 28316 6752 28361 6780
rect 28316 6740 28322 6752
rect 19889 6675 19947 6681
rect 20180 6684 20760 6712
rect 25884 6684 26188 6712
rect 9640 6616 9812 6644
rect 9640 6604 9646 6616
rect 9858 6604 9864 6656
rect 9916 6644 9922 6656
rect 10229 6647 10287 6653
rect 10229 6644 10241 6647
rect 9916 6616 10241 6644
rect 9916 6604 9922 6616
rect 10229 6613 10241 6616
rect 10275 6613 10287 6647
rect 10229 6607 10287 6613
rect 10594 6604 10600 6656
rect 10652 6604 10658 6656
rect 11054 6604 11060 6656
rect 11112 6604 11118 6656
rect 11330 6604 11336 6656
rect 11388 6644 11394 6656
rect 13354 6644 13360 6656
rect 11388 6616 13360 6644
rect 11388 6604 11394 6616
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 13722 6604 13728 6656
rect 13780 6604 13786 6656
rect 14458 6604 14464 6656
rect 14516 6644 14522 6656
rect 15488 6644 15516 6672
rect 14516 6616 15516 6644
rect 14516 6604 14522 6616
rect 16574 6604 16580 6656
rect 16632 6604 16638 6656
rect 16666 6604 16672 6656
rect 16724 6644 16730 6656
rect 16853 6647 16911 6653
rect 16853 6644 16865 6647
rect 16724 6616 16865 6644
rect 16724 6604 16730 6616
rect 16853 6613 16865 6616
rect 16899 6613 16911 6647
rect 16853 6607 16911 6613
rect 17126 6604 17132 6656
rect 17184 6604 17190 6656
rect 17218 6604 17224 6656
rect 17276 6604 17282 6656
rect 17770 6604 17776 6656
rect 17828 6644 17834 6656
rect 17957 6647 18015 6653
rect 17957 6644 17969 6647
rect 17828 6616 17969 6644
rect 17828 6604 17834 6616
rect 17957 6613 17969 6616
rect 18003 6613 18015 6647
rect 17957 6607 18015 6613
rect 18598 6604 18604 6656
rect 18656 6644 18662 6656
rect 20180 6644 20208 6684
rect 25884 6656 25912 6684
rect 18656 6616 20208 6644
rect 18656 6604 18662 6616
rect 20254 6604 20260 6656
rect 20312 6604 20318 6656
rect 20530 6604 20536 6656
rect 20588 6604 20594 6656
rect 20809 6647 20867 6653
rect 20809 6613 20821 6647
rect 20855 6644 20867 6647
rect 21174 6644 21180 6656
rect 20855 6616 21180 6644
rect 20855 6613 20867 6616
rect 20809 6607 20867 6613
rect 21174 6604 21180 6616
rect 21232 6604 21238 6656
rect 21269 6647 21327 6653
rect 21269 6613 21281 6647
rect 21315 6644 21327 6647
rect 21542 6644 21548 6656
rect 21315 6616 21548 6644
rect 21315 6613 21327 6616
rect 21269 6607 21327 6613
rect 21542 6604 21548 6616
rect 21600 6604 21606 6656
rect 21726 6604 21732 6656
rect 21784 6644 21790 6656
rect 25222 6644 25228 6656
rect 21784 6616 25228 6644
rect 21784 6604 21790 6616
rect 25222 6604 25228 6616
rect 25280 6604 25286 6656
rect 25866 6604 25872 6656
rect 25924 6604 25930 6656
rect 26050 6604 26056 6656
rect 26108 6604 26114 6656
rect 26160 6644 26188 6684
rect 27338 6672 27344 6724
rect 27396 6712 27402 6724
rect 29641 6715 29699 6721
rect 27396 6684 27568 6712
rect 27396 6672 27402 6684
rect 27433 6647 27491 6653
rect 27433 6644 27445 6647
rect 26160 6616 27445 6644
rect 27433 6613 27445 6616
rect 27479 6613 27491 6647
rect 27540 6644 27568 6684
rect 29641 6681 29653 6715
rect 29687 6681 29699 6715
rect 29641 6675 29699 6681
rect 29656 6644 29684 6675
rect 27540 6616 29684 6644
rect 27433 6607 27491 6613
rect 552 6554 30912 6576
rect 552 6502 4193 6554
rect 4245 6502 4257 6554
rect 4309 6502 4321 6554
rect 4373 6502 4385 6554
rect 4437 6502 4449 6554
rect 4501 6502 11783 6554
rect 11835 6502 11847 6554
rect 11899 6502 11911 6554
rect 11963 6502 11975 6554
rect 12027 6502 12039 6554
rect 12091 6502 19373 6554
rect 19425 6502 19437 6554
rect 19489 6502 19501 6554
rect 19553 6502 19565 6554
rect 19617 6502 19629 6554
rect 19681 6502 26963 6554
rect 27015 6502 27027 6554
rect 27079 6502 27091 6554
rect 27143 6502 27155 6554
rect 27207 6502 27219 6554
rect 27271 6502 30912 6554
rect 552 6480 30912 6502
rect 5074 6400 5080 6452
rect 5132 6400 5138 6452
rect 5350 6400 5356 6452
rect 5408 6440 5414 6452
rect 10597 6443 10655 6449
rect 10597 6440 10609 6443
rect 5408 6412 10609 6440
rect 5408 6400 5414 6412
rect 10597 6409 10609 6412
rect 10643 6409 10655 6443
rect 10597 6403 10655 6409
rect 11054 6400 11060 6452
rect 11112 6400 11118 6452
rect 11146 6400 11152 6452
rect 11204 6440 11210 6452
rect 13081 6443 13139 6449
rect 13081 6440 13093 6443
rect 11204 6412 13093 6440
rect 11204 6400 11210 6412
rect 13081 6409 13093 6412
rect 13127 6409 13139 6443
rect 13081 6403 13139 6409
rect 13817 6443 13875 6449
rect 13817 6409 13829 6443
rect 13863 6440 13875 6443
rect 14550 6440 14556 6452
rect 13863 6412 14556 6440
rect 13863 6409 13875 6412
rect 13817 6403 13875 6409
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 16206 6400 16212 6452
rect 16264 6400 16270 6452
rect 18049 6443 18107 6449
rect 17420 6412 17908 6440
rect 1443 6307 1501 6313
rect 1443 6273 1455 6307
rect 1489 6304 1501 6307
rect 2590 6304 2596 6316
rect 1489 6276 2596 6304
rect 1489 6273 1501 6276
rect 1443 6267 1501 6273
rect 2590 6264 2596 6276
rect 2648 6264 2654 6316
rect 3564 6307 3622 6313
rect 3564 6304 3576 6307
rect 2746 6276 3576 6304
rect 842 6196 848 6248
rect 900 6236 906 6248
rect 937 6239 995 6245
rect 937 6236 949 6239
rect 900 6208 949 6236
rect 900 6196 906 6208
rect 937 6205 949 6208
rect 983 6205 995 6239
rect 937 6199 995 6205
rect 1670 6196 1676 6248
rect 1728 6196 1734 6248
rect 2038 6196 2044 6248
rect 2096 6236 2102 6248
rect 2746 6236 2774 6276
rect 3564 6273 3576 6276
rect 3610 6273 3622 6307
rect 3564 6267 3622 6273
rect 3743 6307 3801 6313
rect 3743 6273 3755 6307
rect 3789 6304 3801 6307
rect 5092 6304 5120 6400
rect 7374 6332 7380 6384
rect 7432 6332 7438 6384
rect 8113 6375 8171 6381
rect 8113 6341 8125 6375
rect 8159 6372 8171 6375
rect 8386 6372 8392 6384
rect 8159 6344 8392 6372
rect 8159 6341 8171 6344
rect 8113 6335 8171 6341
rect 8386 6332 8392 6344
rect 8444 6332 8450 6384
rect 10873 6375 10931 6381
rect 10873 6341 10885 6375
rect 10919 6341 10931 6375
rect 10873 6335 10931 6341
rect 3789 6276 5120 6304
rect 3789 6273 3801 6276
rect 3743 6267 3801 6273
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 5902 6313 5908 6316
rect 5864 6307 5908 6313
rect 5864 6273 5876 6307
rect 5864 6267 5908 6273
rect 5902 6264 5908 6267
rect 5960 6264 5966 6316
rect 6086 6313 6092 6316
rect 6043 6307 6092 6313
rect 6043 6273 6055 6307
rect 6089 6273 6092 6307
rect 6043 6267 6092 6273
rect 6086 6264 6092 6267
rect 6144 6264 6150 6316
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 6273 6307 6331 6313
rect 6273 6304 6285 6307
rect 6236 6276 6285 6304
rect 6236 6264 6242 6276
rect 6273 6273 6285 6276
rect 6319 6273 6331 6307
rect 6273 6267 6331 6273
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 8852 6307 8910 6313
rect 8852 6304 8864 6307
rect 8628 6276 8864 6304
rect 8628 6264 8634 6276
rect 8852 6273 8864 6276
rect 8898 6273 8910 6307
rect 8852 6267 8910 6273
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 10888 6304 10916 6335
rect 9088 6276 10916 6304
rect 11072 6304 11100 6400
rect 11606 6313 11612 6316
rect 11568 6307 11612 6313
rect 11072 6276 11468 6304
rect 9088 6264 9094 6276
rect 2096 6208 2774 6236
rect 2096 6196 2102 6208
rect 3142 6196 3148 6248
rect 3200 6236 3206 6248
rect 3237 6239 3295 6245
rect 3237 6236 3249 6239
rect 3200 6208 3249 6236
rect 3200 6196 3206 6208
rect 3237 6205 3249 6208
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 3878 6196 3884 6248
rect 3936 6236 3942 6248
rect 3973 6239 4031 6245
rect 3973 6236 3985 6239
rect 3936 6208 3985 6236
rect 3936 6196 3942 6208
rect 3973 6205 3985 6208
rect 4019 6205 4031 6239
rect 3973 6199 4031 6205
rect 5537 6239 5595 6245
rect 5537 6205 5549 6239
rect 5583 6236 5595 6239
rect 5736 6236 5764 6264
rect 5583 6208 5764 6236
rect 5583 6205 5595 6208
rect 5537 6199 5595 6205
rect 8386 6196 8392 6248
rect 8444 6196 8450 6248
rect 8478 6196 8484 6248
rect 8536 6236 8542 6248
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 8536 6208 9137 6236
rect 8536 6196 8542 6208
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 9125 6199 9183 6205
rect 9784 6208 10793 6236
rect 7837 6171 7895 6177
rect 7837 6168 7849 6171
rect 4632 6140 5212 6168
rect 1394 6060 1400 6112
rect 1452 6109 1458 6112
rect 1452 6100 1461 6109
rect 1452 6072 1497 6100
rect 1452 6063 1461 6072
rect 1452 6060 1458 6063
rect 2774 6060 2780 6112
rect 2832 6060 2838 6112
rect 3234 6060 3240 6112
rect 3292 6100 3298 6112
rect 3694 6100 3700 6112
rect 3292 6072 3700 6100
rect 3292 6060 3298 6072
rect 3694 6060 3700 6072
rect 3752 6100 3758 6112
rect 4632 6100 4660 6140
rect 3752 6072 4660 6100
rect 3752 6060 3758 6072
rect 5074 6060 5080 6112
rect 5132 6060 5138 6112
rect 5184 6100 5212 6140
rect 6932 6140 7849 6168
rect 6932 6100 6960 6140
rect 7837 6137 7849 6140
rect 7883 6137 7895 6171
rect 7837 6131 7895 6137
rect 5184 6072 6960 6100
rect 8662 6060 8668 6112
rect 8720 6100 8726 6112
rect 8855 6103 8913 6109
rect 8855 6100 8867 6103
rect 8720 6072 8867 6100
rect 8720 6060 8726 6072
rect 8855 6069 8867 6072
rect 8901 6069 8913 6103
rect 8855 6063 8913 6069
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 9784 6100 9812 6208
rect 10781 6205 10793 6208
rect 10827 6236 10839 6239
rect 10870 6236 10876 6248
rect 10827 6208 10876 6236
rect 10827 6205 10839 6208
rect 10781 6199 10839 6205
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 11054 6196 11060 6248
rect 11112 6196 11118 6248
rect 11238 6196 11244 6248
rect 11296 6196 11302 6248
rect 11440 6236 11468 6276
rect 11568 6273 11580 6307
rect 11568 6267 11612 6273
rect 11606 6264 11612 6267
rect 11664 6264 11670 6316
rect 11747 6307 11805 6313
rect 11747 6273 11759 6307
rect 11793 6304 11805 6307
rect 12434 6304 12440 6316
rect 11793 6276 12440 6304
rect 11793 6273 11805 6276
rect 11747 6267 11805 6273
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 13814 6264 13820 6316
rect 13872 6304 13878 6316
rect 14734 6313 14740 6316
rect 14369 6307 14427 6313
rect 14369 6304 14381 6307
rect 13872 6276 14381 6304
rect 13872 6264 13878 6276
rect 14369 6273 14381 6276
rect 14415 6273 14427 6307
rect 14369 6267 14427 6273
rect 14696 6307 14740 6313
rect 14696 6273 14708 6307
rect 14696 6267 14740 6273
rect 14734 6264 14740 6267
rect 14792 6264 14798 6316
rect 14875 6307 14933 6313
rect 14875 6273 14887 6307
rect 14921 6304 14933 6307
rect 15010 6304 15016 6316
rect 14921 6276 15016 6304
rect 14921 6273 14933 6276
rect 14875 6267 14933 6273
rect 15010 6264 15016 6276
rect 15068 6264 15074 6316
rect 15105 6307 15163 6313
rect 15105 6273 15117 6307
rect 15151 6304 15163 6307
rect 16298 6304 16304 6316
rect 15151 6276 16304 6304
rect 15151 6273 15163 6276
rect 15105 6267 15163 6273
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 11977 6239 12035 6245
rect 11977 6236 11989 6239
rect 11440 6208 11989 6236
rect 11977 6205 11989 6208
rect 12023 6205 12035 6239
rect 11977 6199 12035 6205
rect 13354 6196 13360 6248
rect 13412 6236 13418 6248
rect 13725 6239 13783 6245
rect 13725 6236 13737 6239
rect 13412 6208 13737 6236
rect 13412 6196 13418 6208
rect 13725 6205 13737 6208
rect 13771 6236 13783 6239
rect 14001 6239 14059 6245
rect 14001 6236 14013 6239
rect 13771 6208 14013 6236
rect 13771 6205 13783 6208
rect 13725 6199 13783 6205
rect 14001 6205 14013 6208
rect 14047 6205 14059 6239
rect 14001 6199 14059 6205
rect 14090 6196 14096 6248
rect 14148 6236 14154 6248
rect 14277 6239 14335 6245
rect 14277 6236 14289 6239
rect 14148 6208 14289 6236
rect 14148 6196 14154 6208
rect 14277 6205 14289 6208
rect 14323 6205 14335 6239
rect 16666 6236 16672 6248
rect 14277 6199 14335 6205
rect 14384 6208 16672 6236
rect 9640 6072 9812 6100
rect 9640 6060 9646 6072
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 10229 6103 10287 6109
rect 10229 6100 10241 6103
rect 10100 6072 10241 6100
rect 10100 6060 10106 6072
rect 10229 6069 10241 6072
rect 10275 6069 10287 6103
rect 11072 6100 11100 6196
rect 13630 6128 13636 6180
rect 13688 6168 13694 6180
rect 14384 6168 14412 6208
rect 16666 6196 16672 6208
rect 16724 6196 16730 6248
rect 17420 6245 17448 6412
rect 17773 6375 17831 6381
rect 17773 6341 17785 6375
rect 17819 6341 17831 6375
rect 17880 6372 17908 6412
rect 18049 6409 18061 6443
rect 18095 6440 18107 6443
rect 18690 6440 18696 6452
rect 18095 6412 18696 6440
rect 18095 6409 18107 6412
rect 18049 6403 18107 6409
rect 18690 6400 18696 6412
rect 18748 6400 18754 6452
rect 20254 6400 20260 6452
rect 20312 6400 20318 6452
rect 21266 6400 21272 6452
rect 21324 6440 21330 6452
rect 23477 6443 23535 6449
rect 21324 6412 23428 6440
rect 21324 6400 21330 6412
rect 18230 6372 18236 6384
rect 17880 6344 18236 6372
rect 17773 6335 17831 6341
rect 17788 6304 17816 6335
rect 18230 6332 18236 6344
rect 18288 6332 18294 6384
rect 19156 6307 19214 6313
rect 19156 6304 19168 6307
rect 17788 6276 18828 6304
rect 18800 6248 18828 6276
rect 18984 6276 19168 6304
rect 18984 6248 19012 6276
rect 19156 6273 19168 6276
rect 19202 6273 19214 6307
rect 19156 6267 19214 6273
rect 19429 6307 19487 6313
rect 19429 6273 19441 6307
rect 19475 6304 19487 6307
rect 20272 6304 20300 6400
rect 23400 6372 23428 6412
rect 23477 6409 23489 6443
rect 23523 6440 23535 6443
rect 24762 6440 24768 6452
rect 23523 6412 24768 6440
rect 23523 6409 23535 6412
rect 23477 6403 23535 6409
rect 24762 6400 24768 6412
rect 24820 6400 24826 6452
rect 25222 6400 25228 6452
rect 25280 6440 25286 6452
rect 28537 6443 28595 6449
rect 28537 6440 28549 6443
rect 25280 6412 28549 6440
rect 25280 6400 25286 6412
rect 28537 6409 28549 6412
rect 28583 6409 28595 6443
rect 28537 6403 28595 6409
rect 29638 6400 29644 6452
rect 29696 6400 29702 6452
rect 23566 6372 23572 6384
rect 23400 6344 23572 6372
rect 23566 6332 23572 6344
rect 23624 6332 23630 6384
rect 19475 6276 20300 6304
rect 20809 6307 20867 6313
rect 19475 6273 19487 6276
rect 19429 6267 19487 6273
rect 20809 6273 20821 6307
rect 20855 6304 20867 6307
rect 21364 6307 21422 6313
rect 21364 6304 21376 6307
rect 20855 6276 21376 6304
rect 20855 6273 20867 6276
rect 20809 6267 20867 6273
rect 21364 6273 21376 6276
rect 21410 6273 21422 6307
rect 21364 6267 21422 6273
rect 21542 6264 21548 6316
rect 21600 6304 21606 6316
rect 21637 6307 21695 6313
rect 21637 6304 21649 6307
rect 21600 6276 21649 6304
rect 21600 6264 21606 6276
rect 21637 6273 21649 6276
rect 21683 6273 21695 6307
rect 21637 6267 21695 6273
rect 23474 6264 23480 6316
rect 23532 6264 23538 6316
rect 24535 6307 24593 6313
rect 24535 6273 24547 6307
rect 24581 6304 24593 6307
rect 24581 6276 24900 6304
rect 24581 6273 24593 6276
rect 24535 6267 24593 6273
rect 16853 6239 16911 6245
rect 16853 6205 16865 6239
rect 16899 6236 16911 6239
rect 17129 6239 17187 6245
rect 16899 6208 17080 6236
rect 16899 6205 16911 6208
rect 16853 6199 16911 6205
rect 13688 6140 14412 6168
rect 13688 6128 13694 6140
rect 17052 6112 17080 6208
rect 17129 6205 17141 6239
rect 17175 6205 17187 6239
rect 17129 6199 17187 6205
rect 17405 6239 17463 6245
rect 17405 6205 17417 6239
rect 17451 6205 17463 6239
rect 17405 6199 17463 6205
rect 17497 6239 17555 6245
rect 17497 6205 17509 6239
rect 17543 6236 17555 6239
rect 17586 6236 17592 6248
rect 17543 6208 17592 6236
rect 17543 6205 17555 6208
rect 17497 6199 17555 6205
rect 17144 6168 17172 6199
rect 17586 6196 17592 6208
rect 17644 6196 17650 6248
rect 17954 6196 17960 6248
rect 18012 6196 18018 6248
rect 18230 6196 18236 6248
rect 18288 6196 18294 6248
rect 18322 6196 18328 6248
rect 18380 6196 18386 6248
rect 18690 6196 18696 6248
rect 18748 6196 18754 6248
rect 18782 6196 18788 6248
rect 18840 6196 18846 6248
rect 18966 6196 18972 6248
rect 19024 6196 19030 6248
rect 20901 6239 20959 6245
rect 20901 6205 20913 6239
rect 20947 6236 20959 6239
rect 21266 6236 21272 6248
rect 20947 6208 21272 6236
rect 20947 6205 20959 6208
rect 20901 6199 20959 6205
rect 21266 6196 21272 6208
rect 21324 6196 21330 6248
rect 23293 6239 23351 6245
rect 23293 6205 23305 6239
rect 23339 6236 23351 6239
rect 23492 6236 23520 6264
rect 24872 6248 24900 6276
rect 26326 6264 26332 6316
rect 26384 6304 26390 6316
rect 27160 6307 27218 6313
rect 27160 6304 27172 6307
rect 26384 6276 27172 6304
rect 26384 6264 26390 6276
rect 27160 6273 27172 6276
rect 27206 6273 27218 6307
rect 27160 6267 27218 6273
rect 27433 6307 27491 6313
rect 27433 6273 27445 6307
rect 27479 6304 27491 6307
rect 27522 6304 27528 6316
rect 27479 6276 27528 6304
rect 27479 6273 27491 6276
rect 27433 6267 27491 6273
rect 27522 6264 27528 6276
rect 27580 6264 27586 6316
rect 28074 6264 28080 6316
rect 28132 6304 28138 6316
rect 29656 6304 29684 6400
rect 28132 6276 29684 6304
rect 28132 6264 28138 6276
rect 23339 6208 23520 6236
rect 23661 6239 23719 6245
rect 23339 6205 23351 6208
rect 23293 6199 23351 6205
rect 23661 6205 23673 6239
rect 23707 6236 23719 6239
rect 23750 6236 23756 6248
rect 23707 6208 23756 6236
rect 23707 6205 23719 6208
rect 23661 6199 23719 6205
rect 23750 6196 23756 6208
rect 23808 6196 23814 6248
rect 23934 6196 23940 6248
rect 23992 6236 23998 6248
rect 24029 6239 24087 6245
rect 24029 6236 24041 6239
rect 23992 6208 24041 6236
rect 23992 6196 23998 6208
rect 24029 6205 24041 6208
rect 24075 6205 24087 6239
rect 24029 6199 24087 6205
rect 24670 6196 24676 6248
rect 24728 6236 24734 6248
rect 24765 6239 24823 6245
rect 24765 6236 24777 6239
rect 24728 6208 24777 6236
rect 24728 6196 24734 6208
rect 24765 6205 24777 6208
rect 24811 6205 24823 6239
rect 24765 6199 24823 6205
rect 24854 6196 24860 6248
rect 24912 6196 24918 6248
rect 26605 6239 26663 6245
rect 26605 6205 26617 6239
rect 26651 6205 26663 6239
rect 26605 6199 26663 6205
rect 18598 6168 18604 6180
rect 17144 6140 18604 6168
rect 18598 6128 18604 6140
rect 18656 6128 18662 6180
rect 23017 6171 23075 6177
rect 23017 6137 23029 6171
rect 23063 6168 23075 6171
rect 24118 6168 24124 6180
rect 23063 6140 24124 6168
rect 23063 6137 23075 6140
rect 23017 6131 23075 6137
rect 24118 6128 24124 6140
rect 24176 6128 24182 6180
rect 26142 6128 26148 6180
rect 26200 6128 26206 6180
rect 26510 6128 26516 6180
rect 26568 6168 26574 6180
rect 26620 6168 26648 6199
rect 26694 6196 26700 6248
rect 26752 6196 26758 6248
rect 26786 6196 26792 6248
rect 26844 6236 26850 6248
rect 27024 6239 27082 6245
rect 27024 6236 27036 6239
rect 26844 6208 27036 6236
rect 26844 6196 26850 6208
rect 27024 6205 27036 6208
rect 27070 6236 27082 6239
rect 29181 6239 29239 6245
rect 27070 6208 28396 6236
rect 27070 6205 27082 6208
rect 27024 6199 27082 6205
rect 28368 6180 28396 6208
rect 29181 6205 29193 6239
rect 29227 6236 29239 6239
rect 29270 6236 29276 6248
rect 29227 6208 29276 6236
rect 29227 6205 29239 6208
rect 29181 6199 29239 6205
rect 29270 6196 29276 6208
rect 29328 6196 29334 6248
rect 26568 6140 26832 6168
rect 26568 6128 26574 6140
rect 13446 6100 13452 6112
rect 11072 6072 13452 6100
rect 10229 6063 10287 6069
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 13538 6060 13544 6112
rect 13596 6060 13602 6112
rect 14093 6103 14151 6109
rect 14093 6069 14105 6103
rect 14139 6100 14151 6103
rect 14458 6100 14464 6112
rect 14139 6072 14464 6100
rect 14139 6069 14151 6072
rect 14093 6063 14151 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 16669 6103 16727 6109
rect 16669 6069 16681 6103
rect 16715 6100 16727 6103
rect 16850 6100 16856 6112
rect 16715 6072 16856 6100
rect 16715 6069 16727 6072
rect 16669 6063 16727 6069
rect 16850 6060 16856 6072
rect 16908 6060 16914 6112
rect 16942 6060 16948 6112
rect 17000 6060 17006 6112
rect 17034 6060 17040 6112
rect 17092 6060 17098 6112
rect 17218 6060 17224 6112
rect 17276 6060 17282 6112
rect 17678 6060 17684 6112
rect 17736 6060 17742 6112
rect 18506 6060 18512 6112
rect 18564 6060 18570 6112
rect 18782 6060 18788 6112
rect 18840 6100 18846 6112
rect 19159 6103 19217 6109
rect 19159 6100 19171 6103
rect 18840 6072 19171 6100
rect 18840 6060 18846 6072
rect 19159 6069 19171 6072
rect 19205 6069 19217 6103
rect 19159 6063 19217 6069
rect 21367 6103 21425 6109
rect 21367 6069 21379 6103
rect 21413 6100 21425 6103
rect 21542 6100 21548 6112
rect 21413 6072 21548 6100
rect 21413 6069 21425 6072
rect 21367 6063 21425 6069
rect 21542 6060 21548 6072
rect 21600 6060 21606 6112
rect 22922 6060 22928 6112
rect 22980 6100 22986 6112
rect 23109 6103 23167 6109
rect 23109 6100 23121 6103
rect 22980 6072 23121 6100
rect 22980 6060 22986 6072
rect 23109 6069 23121 6072
rect 23155 6069 23167 6103
rect 23109 6063 23167 6069
rect 24495 6103 24553 6109
rect 24495 6069 24507 6103
rect 24541 6100 24553 6103
rect 24762 6100 24768 6112
rect 24541 6072 24768 6100
rect 24541 6069 24553 6072
rect 24495 6063 24553 6069
rect 24762 6060 24768 6072
rect 24820 6060 24826 6112
rect 26421 6103 26479 6109
rect 26421 6069 26433 6103
rect 26467 6100 26479 6103
rect 26694 6100 26700 6112
rect 26467 6072 26700 6100
rect 26467 6069 26479 6072
rect 26421 6063 26479 6069
rect 26694 6060 26700 6072
rect 26752 6060 26758 6112
rect 26804 6100 26832 6140
rect 28350 6128 28356 6180
rect 28408 6128 28414 6180
rect 27246 6100 27252 6112
rect 26804 6072 27252 6100
rect 27246 6060 27252 6072
rect 27304 6060 27310 6112
rect 27338 6060 27344 6112
rect 27396 6100 27402 6112
rect 28997 6103 29055 6109
rect 28997 6100 29009 6103
rect 27396 6072 29009 6100
rect 27396 6060 27402 6072
rect 28997 6069 29009 6072
rect 29043 6069 29055 6103
rect 28997 6063 29055 6069
rect 552 6010 31072 6032
rect 552 5958 7988 6010
rect 8040 5958 8052 6010
rect 8104 5958 8116 6010
rect 8168 5958 8180 6010
rect 8232 5958 8244 6010
rect 8296 5958 15578 6010
rect 15630 5958 15642 6010
rect 15694 5958 15706 6010
rect 15758 5958 15770 6010
rect 15822 5958 15834 6010
rect 15886 5958 23168 6010
rect 23220 5958 23232 6010
rect 23284 5958 23296 6010
rect 23348 5958 23360 6010
rect 23412 5958 23424 6010
rect 23476 5958 30758 6010
rect 30810 5958 30822 6010
rect 30874 5958 30886 6010
rect 30938 5958 30950 6010
rect 31002 5958 31014 6010
rect 31066 5958 31072 6010
rect 552 5936 31072 5958
rect 1210 5856 1216 5908
rect 1268 5856 1274 5908
rect 1578 5856 1584 5908
rect 1636 5896 1642 5908
rect 1771 5899 1829 5905
rect 1771 5896 1783 5899
rect 1636 5868 1783 5896
rect 1636 5856 1642 5868
rect 1771 5865 1783 5868
rect 1817 5896 1829 5899
rect 2038 5896 2044 5908
rect 1817 5868 2044 5896
rect 1817 5865 1829 5868
rect 1771 5859 1829 5865
rect 2038 5856 2044 5868
rect 2096 5856 2102 5908
rect 2866 5896 2872 5908
rect 2746 5868 2872 5896
rect 1228 5828 1256 5856
rect 1228 5800 1348 5828
rect 1320 5772 1348 5800
rect 1026 5720 1032 5772
rect 1084 5760 1090 5772
rect 1210 5760 1216 5772
rect 1084 5732 1216 5760
rect 1084 5720 1090 5732
rect 1210 5720 1216 5732
rect 1268 5720 1274 5772
rect 1302 5720 1308 5772
rect 1360 5720 1366 5772
rect 2746 5760 2774 5868
rect 2866 5856 2872 5868
rect 2924 5856 2930 5908
rect 3786 5856 3792 5908
rect 3844 5896 3850 5908
rect 3979 5899 4037 5905
rect 3979 5896 3991 5899
rect 3844 5868 3991 5896
rect 3844 5856 3850 5868
rect 3979 5865 3991 5868
rect 4025 5865 4037 5899
rect 3979 5859 4037 5865
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 6454 5896 6460 5908
rect 5592 5868 6460 5896
rect 5592 5856 5598 5868
rect 6454 5856 6460 5868
rect 6512 5856 6518 5908
rect 8487 5899 8545 5905
rect 8487 5865 8499 5899
rect 8533 5896 8545 5899
rect 8662 5896 8668 5908
rect 8533 5868 8668 5896
rect 8533 5865 8545 5868
rect 8487 5859 8545 5865
rect 8662 5856 8668 5868
rect 8720 5856 8726 5908
rect 11057 5899 11115 5905
rect 11057 5865 11069 5899
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 3421 5831 3479 5837
rect 3421 5797 3433 5831
rect 3467 5828 3479 5831
rect 3510 5828 3516 5840
rect 3467 5800 3516 5828
rect 3467 5797 3479 5800
rect 3421 5791 3479 5797
rect 3510 5788 3516 5800
rect 3568 5788 3574 5840
rect 5350 5788 5356 5840
rect 5408 5788 5414 5840
rect 11072 5828 11100 5859
rect 13446 5856 13452 5908
rect 13504 5896 13510 5908
rect 16758 5896 16764 5908
rect 13504 5868 16764 5896
rect 13504 5856 13510 5868
rect 16758 5856 16764 5868
rect 16816 5856 16822 5908
rect 17034 5856 17040 5908
rect 17092 5896 17098 5908
rect 20898 5896 20904 5908
rect 17092 5868 20904 5896
rect 17092 5856 17098 5868
rect 20898 5856 20904 5868
rect 20956 5856 20962 5908
rect 21542 5856 21548 5908
rect 21600 5896 21606 5908
rect 21735 5899 21793 5905
rect 21735 5896 21747 5899
rect 21600 5868 21747 5896
rect 21600 5856 21606 5868
rect 21735 5865 21747 5868
rect 21781 5865 21793 5899
rect 21735 5859 21793 5865
rect 23934 5856 23940 5908
rect 23992 5905 23998 5908
rect 23992 5896 24001 5905
rect 23992 5868 24037 5896
rect 23992 5859 24001 5868
rect 23992 5856 23998 5859
rect 24854 5856 24860 5908
rect 24912 5896 24918 5908
rect 25317 5899 25375 5905
rect 25317 5896 25329 5899
rect 24912 5868 25329 5896
rect 24912 5856 24918 5868
rect 25317 5865 25329 5868
rect 25363 5865 25375 5899
rect 25317 5859 25375 5865
rect 25958 5856 25964 5908
rect 26016 5856 26022 5908
rect 26887 5899 26945 5905
rect 26887 5896 26899 5899
rect 26068 5868 26899 5896
rect 5460 5800 5948 5828
rect 11072 5800 11744 5828
rect 1964 5732 2774 5760
rect 1801 5713 1859 5719
rect 1801 5710 1813 5713
rect 1780 5679 1813 5710
rect 1847 5692 1859 5713
rect 1964 5692 1992 5732
rect 2866 5720 2872 5772
rect 2924 5760 2930 5772
rect 4249 5763 4307 5769
rect 2924 5732 4200 5760
rect 2924 5720 2930 5732
rect 1847 5679 1992 5692
rect 1780 5664 1992 5679
rect 2038 5652 2044 5704
rect 2096 5652 2102 5704
rect 3326 5652 3332 5704
rect 3384 5692 3390 5704
rect 4062 5701 4068 5704
rect 3513 5695 3571 5701
rect 3513 5692 3525 5695
rect 3384 5664 3525 5692
rect 3384 5652 3390 5664
rect 3513 5661 3525 5664
rect 3559 5661 3571 5695
rect 3513 5655 3571 5661
rect 4019 5695 4068 5701
rect 4019 5661 4031 5695
rect 4065 5661 4068 5695
rect 4019 5655 4068 5661
rect 4062 5652 4068 5655
rect 4120 5652 4126 5704
rect 4172 5692 4200 5732
rect 4249 5729 4261 5763
rect 4295 5760 4307 5763
rect 5368 5760 5396 5788
rect 5460 5772 5488 5800
rect 4295 5732 5396 5760
rect 4295 5729 4307 5732
rect 4249 5723 4307 5729
rect 5442 5720 5448 5772
rect 5500 5720 5506 5772
rect 5920 5760 5948 5800
rect 6549 5763 6607 5769
rect 6549 5760 6561 5763
rect 5920 5732 6561 5760
rect 6549 5729 6561 5732
rect 6595 5729 6607 5763
rect 6549 5723 6607 5729
rect 7834 5720 7840 5772
rect 7892 5760 7898 5772
rect 7892 5732 8432 5760
rect 7892 5720 7898 5732
rect 8404 5710 8432 5732
rect 10410 5720 10416 5772
rect 10468 5769 10474 5772
rect 10468 5760 10479 5769
rect 10781 5763 10839 5769
rect 10468 5732 10513 5760
rect 10468 5723 10479 5732
rect 10781 5729 10793 5763
rect 10827 5729 10839 5763
rect 10781 5723 10839 5729
rect 10468 5720 10474 5723
rect 8484 5713 8542 5719
rect 8484 5710 8496 5713
rect 4172 5664 5672 5692
rect 2746 5596 3556 5624
rect 1029 5559 1087 5565
rect 1029 5525 1041 5559
rect 1075 5556 1087 5559
rect 2746 5556 2774 5596
rect 1075 5528 2774 5556
rect 3528 5556 3556 5596
rect 5442 5584 5448 5636
rect 5500 5584 5506 5636
rect 5460 5556 5488 5584
rect 3528 5528 5488 5556
rect 1075 5525 1087 5528
rect 1029 5519 1087 5525
rect 5534 5516 5540 5568
rect 5592 5516 5598 5568
rect 5644 5556 5672 5664
rect 5810 5652 5816 5704
rect 5868 5652 5874 5704
rect 6178 5701 6184 5704
rect 6140 5695 6184 5701
rect 6140 5661 6152 5695
rect 6140 5655 6184 5661
rect 6178 5652 6184 5655
rect 6236 5652 6242 5704
rect 6270 5652 6276 5704
rect 6328 5652 6334 5704
rect 6454 5652 6460 5704
rect 6512 5692 6518 5704
rect 8021 5695 8079 5701
rect 8021 5692 8033 5695
rect 6512 5664 8033 5692
rect 6512 5652 6518 5664
rect 8021 5661 8033 5664
rect 8067 5692 8079 5695
rect 8294 5692 8300 5704
rect 8067 5664 8300 5692
rect 8067 5661 8079 5664
rect 8021 5655 8079 5661
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8404 5682 8496 5710
rect 8484 5679 8496 5682
rect 8530 5679 8542 5713
rect 8484 5673 8542 5679
rect 8754 5652 8760 5704
rect 8812 5652 8818 5704
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5692 10195 5695
rect 10318 5692 10324 5704
rect 10183 5664 10324 5692
rect 10183 5661 10195 5664
rect 10137 5655 10195 5661
rect 10318 5652 10324 5664
rect 10376 5652 10382 5704
rect 10796 5692 10824 5723
rect 11238 5720 11244 5772
rect 11296 5720 11302 5772
rect 11517 5763 11575 5769
rect 11517 5729 11529 5763
rect 11563 5729 11575 5763
rect 11716 5760 11744 5800
rect 12345 5763 12403 5769
rect 12345 5760 12357 5763
rect 11716 5732 12357 5760
rect 11517 5723 11575 5729
rect 12345 5729 12357 5732
rect 12391 5729 12403 5763
rect 12345 5723 12403 5729
rect 11532 5692 11560 5723
rect 14458 5720 14464 5772
rect 14516 5760 14522 5772
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 14516 5732 14565 5760
rect 14516 5720 14522 5732
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 15933 5763 15991 5769
rect 15933 5729 15945 5763
rect 15979 5760 15991 5763
rect 15979 5732 16715 5760
rect 15979 5729 15991 5732
rect 15933 5723 15991 5729
rect 10796 5664 11560 5692
rect 11238 5624 11244 5636
rect 7208 5596 7788 5624
rect 7208 5556 7236 5596
rect 5644 5528 7236 5556
rect 7650 5516 7656 5568
rect 7708 5516 7714 5568
rect 7760 5556 7788 5596
rect 9600 5596 11244 5624
rect 8754 5556 8760 5568
rect 7760 5528 8760 5556
rect 8754 5516 8760 5528
rect 8812 5516 8818 5568
rect 8938 5516 8944 5568
rect 8996 5556 9002 5568
rect 9600 5556 9628 5596
rect 11238 5584 11244 5596
rect 11296 5584 11302 5636
rect 11532 5624 11560 5664
rect 11606 5652 11612 5704
rect 11664 5652 11670 5704
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 12158 5701 12164 5704
rect 11936 5695 11994 5701
rect 11936 5692 11948 5695
rect 11848 5664 11948 5692
rect 11848 5652 11854 5664
rect 11936 5661 11948 5664
rect 11982 5661 11994 5695
rect 11936 5655 11994 5661
rect 12115 5695 12164 5701
rect 12115 5661 12127 5695
rect 12161 5661 12164 5695
rect 12115 5655 12164 5661
rect 12158 5652 12164 5655
rect 12216 5652 12222 5704
rect 13817 5695 13875 5701
rect 13817 5661 13829 5695
rect 13863 5692 13875 5695
rect 13998 5692 14004 5704
rect 13863 5664 14004 5692
rect 13863 5661 13875 5664
rect 13817 5655 13875 5661
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 14182 5701 14188 5704
rect 14144 5695 14188 5701
rect 14144 5661 14156 5695
rect 14144 5655 14188 5661
rect 14182 5652 14188 5655
rect 14240 5652 14246 5704
rect 14274 5652 14280 5704
rect 14332 5652 14338 5704
rect 16206 5652 16212 5704
rect 16264 5652 16270 5704
rect 16574 5701 16580 5704
rect 16536 5695 16580 5701
rect 16536 5661 16548 5695
rect 16536 5655 16580 5661
rect 16574 5652 16580 5655
rect 16632 5652 16638 5704
rect 16687 5703 16715 5732
rect 16850 5720 16856 5772
rect 16908 5760 16914 5772
rect 16945 5763 17003 5769
rect 16945 5760 16957 5763
rect 16908 5732 16957 5760
rect 16908 5720 16914 5732
rect 16945 5729 16957 5732
rect 16991 5729 17003 5763
rect 16945 5723 17003 5729
rect 18325 5763 18383 5769
rect 18325 5729 18337 5763
rect 18371 5760 18383 5763
rect 20809 5763 20867 5769
rect 18371 5732 18923 5760
rect 18371 5729 18383 5732
rect 18325 5723 18383 5729
rect 16672 5697 16730 5703
rect 18782 5701 18788 5704
rect 16672 5663 16684 5697
rect 16718 5663 16730 5697
rect 16672 5657 16730 5663
rect 18417 5695 18475 5701
rect 18417 5661 18429 5695
rect 18463 5661 18475 5695
rect 18417 5655 18475 5661
rect 18744 5695 18788 5701
rect 18744 5661 18756 5695
rect 18744 5655 18788 5661
rect 13722 5624 13728 5636
rect 11532 5596 11652 5624
rect 8996 5528 9628 5556
rect 8996 5516 9002 5528
rect 10226 5516 10232 5568
rect 10284 5516 10290 5568
rect 10597 5559 10655 5565
rect 10597 5525 10609 5559
rect 10643 5556 10655 5559
rect 10778 5556 10784 5568
rect 10643 5528 10784 5556
rect 10643 5525 10655 5528
rect 10597 5519 10655 5525
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 11333 5559 11391 5565
rect 11333 5556 11345 5559
rect 11204 5528 11345 5556
rect 11204 5516 11210 5528
rect 11333 5525 11345 5528
rect 11379 5525 11391 5559
rect 11624 5556 11652 5596
rect 13556 5596 13728 5624
rect 13556 5556 13584 5596
rect 13722 5584 13728 5596
rect 13780 5584 13786 5636
rect 11624 5528 13584 5556
rect 13633 5559 13691 5565
rect 11333 5519 11391 5525
rect 13633 5525 13645 5559
rect 13679 5556 13691 5559
rect 14274 5556 14280 5568
rect 13679 5528 14280 5556
rect 13679 5525 13691 5528
rect 13633 5519 13691 5525
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 15378 5516 15384 5568
rect 15436 5556 15442 5568
rect 17126 5556 17132 5568
rect 15436 5528 17132 5556
rect 15436 5516 15442 5528
rect 17126 5516 17132 5528
rect 17184 5516 17190 5568
rect 18432 5556 18460 5655
rect 18782 5652 18788 5655
rect 18840 5652 18846 5704
rect 18895 5703 18923 5732
rect 20809 5729 20821 5763
rect 20855 5760 20867 5763
rect 20916 5760 20944 5856
rect 26068 5828 26096 5868
rect 26887 5865 26899 5868
rect 26933 5865 26945 5899
rect 26887 5859 26945 5865
rect 27246 5856 27252 5908
rect 27304 5896 27310 5908
rect 27304 5868 29040 5896
rect 27304 5856 27310 5868
rect 26510 5828 26516 5840
rect 24964 5800 26096 5828
rect 26160 5800 26516 5828
rect 24964 5772 24992 5800
rect 21085 5763 21143 5769
rect 21085 5760 21097 5763
rect 20855 5732 21097 5760
rect 20855 5729 20867 5732
rect 20809 5723 20867 5729
rect 21085 5729 21097 5732
rect 21131 5729 21143 5763
rect 22005 5763 22063 5769
rect 22005 5760 22017 5763
rect 21085 5723 21143 5729
rect 21192 5732 22017 5760
rect 18880 5697 18938 5703
rect 18880 5663 18892 5697
rect 18926 5663 18938 5697
rect 18880 5657 18938 5663
rect 19153 5695 19211 5701
rect 19153 5661 19165 5695
rect 19199 5692 19211 5695
rect 19199 5664 20668 5692
rect 19199 5661 19211 5664
rect 19153 5655 19211 5661
rect 20640 5633 20668 5664
rect 20625 5627 20683 5633
rect 20625 5593 20637 5627
rect 20671 5593 20683 5627
rect 20625 5587 20683 5593
rect 20901 5627 20959 5633
rect 20901 5593 20913 5627
rect 20947 5624 20959 5627
rect 21192 5624 21220 5732
rect 22005 5729 22017 5732
rect 22051 5729 22063 5763
rect 22005 5723 22063 5729
rect 23385 5763 23443 5769
rect 23385 5729 23397 5763
rect 23431 5760 23443 5763
rect 23431 5732 23980 5760
rect 23431 5729 23443 5732
rect 23385 5723 23443 5729
rect 21266 5652 21272 5704
rect 21324 5652 21330 5704
rect 21726 5652 21732 5704
rect 21784 5692 21790 5704
rect 23477 5695 23535 5701
rect 21784 5664 21829 5692
rect 21784 5652 21790 5664
rect 23477 5661 23489 5695
rect 23523 5692 23535 5695
rect 23658 5692 23664 5704
rect 23523 5664 23664 5692
rect 23523 5661 23535 5664
rect 23477 5655 23535 5661
rect 23658 5652 23664 5664
rect 23716 5652 23722 5704
rect 23952 5701 23980 5732
rect 24670 5720 24676 5772
rect 24728 5720 24734 5772
rect 24946 5720 24952 5772
rect 25004 5720 25010 5772
rect 25682 5720 25688 5772
rect 25740 5760 25746 5772
rect 26160 5769 26188 5800
rect 26510 5788 26516 5800
rect 26568 5788 26574 5840
rect 29012 5828 29040 5868
rect 29454 5856 29460 5908
rect 29512 5856 29518 5908
rect 29472 5828 29500 5856
rect 29012 5800 29500 5828
rect 25869 5763 25927 5769
rect 25740 5732 25802 5760
rect 25740 5720 25746 5732
rect 23940 5695 23998 5701
rect 23940 5661 23952 5695
rect 23986 5661 23998 5695
rect 23940 5655 23998 5661
rect 24210 5652 24216 5704
rect 24268 5652 24274 5704
rect 24688 5692 24716 5720
rect 24688 5664 25728 5692
rect 25700 5633 25728 5664
rect 20947 5596 21220 5624
rect 25685 5627 25743 5633
rect 20947 5593 20959 5596
rect 20901 5587 20959 5593
rect 25685 5593 25697 5627
rect 25731 5593 25743 5627
rect 25774 5624 25802 5732
rect 25869 5729 25881 5763
rect 25915 5760 25927 5763
rect 26145 5763 26203 5769
rect 25915 5732 26004 5760
rect 25915 5729 25927 5732
rect 25869 5723 25927 5729
rect 25976 5704 26004 5732
rect 26145 5729 26157 5763
rect 26191 5729 26203 5763
rect 26145 5723 26203 5729
rect 26234 5720 26240 5772
rect 26292 5760 26298 5772
rect 27157 5763 27215 5769
rect 27157 5760 27169 5763
rect 26292 5732 27169 5760
rect 26292 5720 26298 5732
rect 27157 5729 27169 5732
rect 27203 5729 27215 5763
rect 27157 5723 27215 5729
rect 27982 5720 27988 5772
rect 28040 5760 28046 5772
rect 29012 5769 29040 5800
rect 28629 5763 28687 5769
rect 28629 5760 28641 5763
rect 28040 5732 28641 5760
rect 28040 5720 28046 5732
rect 28629 5729 28641 5732
rect 28675 5729 28687 5763
rect 28629 5723 28687 5729
rect 28997 5763 29055 5769
rect 28997 5729 29009 5763
rect 29043 5729 29055 5763
rect 28997 5723 29055 5729
rect 29273 5763 29331 5769
rect 29273 5729 29285 5763
rect 29319 5729 29331 5763
rect 29273 5723 29331 5729
rect 25958 5652 25964 5704
rect 26016 5652 26022 5704
rect 26421 5695 26479 5701
rect 26421 5661 26433 5695
rect 26467 5661 26479 5695
rect 26421 5655 26479 5661
rect 26439 5624 26467 5655
rect 26878 5652 26884 5704
rect 26936 5652 26942 5704
rect 28644 5692 28672 5723
rect 29288 5692 29316 5723
rect 28644 5664 29316 5692
rect 25774 5596 26467 5624
rect 25685 5587 25743 5593
rect 27890 5584 27896 5636
rect 27948 5624 27954 5636
rect 28813 5627 28871 5633
rect 28813 5624 28825 5627
rect 27948 5596 28825 5624
rect 27948 5584 27954 5596
rect 28813 5593 28825 5596
rect 28859 5593 28871 5627
rect 28813 5587 28871 5593
rect 18690 5556 18696 5568
rect 18432 5528 18696 5556
rect 18690 5516 18696 5528
rect 18748 5516 18754 5568
rect 20441 5559 20499 5565
rect 20441 5525 20453 5559
rect 20487 5556 20499 5559
rect 21726 5556 21732 5568
rect 20487 5528 21732 5556
rect 20487 5525 20499 5528
rect 20441 5519 20499 5525
rect 21726 5516 21732 5528
rect 21784 5516 21790 5568
rect 23382 5516 23388 5568
rect 23440 5556 23446 5568
rect 24210 5556 24216 5568
rect 23440 5528 24216 5556
rect 23440 5516 23446 5528
rect 24210 5516 24216 5528
rect 24268 5516 24274 5568
rect 27798 5516 27804 5568
rect 27856 5556 27862 5568
rect 28261 5559 28319 5565
rect 28261 5556 28273 5559
rect 27856 5528 28273 5556
rect 27856 5516 27862 5528
rect 28261 5525 28273 5528
rect 28307 5525 28319 5559
rect 28261 5519 28319 5525
rect 29178 5516 29184 5568
rect 29236 5516 29242 5568
rect 29454 5516 29460 5568
rect 29512 5516 29518 5568
rect 552 5466 30912 5488
rect 552 5414 4193 5466
rect 4245 5414 4257 5466
rect 4309 5414 4321 5466
rect 4373 5414 4385 5466
rect 4437 5414 4449 5466
rect 4501 5414 11783 5466
rect 11835 5414 11847 5466
rect 11899 5414 11911 5466
rect 11963 5414 11975 5466
rect 12027 5414 12039 5466
rect 12091 5414 19373 5466
rect 19425 5414 19437 5466
rect 19489 5414 19501 5466
rect 19553 5414 19565 5466
rect 19617 5414 19629 5466
rect 19681 5414 26963 5466
rect 27015 5414 27027 5466
rect 27079 5414 27091 5466
rect 27143 5414 27155 5466
rect 27207 5414 27219 5466
rect 27271 5414 30912 5466
rect 552 5392 30912 5414
rect 1302 5352 1308 5364
rect 952 5324 1308 5352
rect 952 5228 980 5324
rect 1302 5312 1308 5324
rect 1360 5352 1366 5364
rect 2961 5355 3019 5361
rect 1360 5324 2774 5352
rect 1360 5312 1366 5324
rect 934 5176 940 5228
rect 992 5176 998 5228
rect 1443 5219 1501 5225
rect 1443 5185 1455 5219
rect 1489 5216 1501 5219
rect 2130 5216 2136 5228
rect 1489 5188 2136 5216
rect 1489 5185 1501 5188
rect 1443 5179 1501 5185
rect 2130 5176 2136 5188
rect 2188 5176 2194 5228
rect 2746 5216 2774 5324
rect 2961 5321 2973 5355
rect 3007 5352 3019 5355
rect 4062 5352 4068 5364
rect 3007 5324 4068 5352
rect 3007 5321 3019 5324
rect 2961 5315 3019 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 5905 5355 5963 5361
rect 5905 5321 5917 5355
rect 5951 5352 5963 5355
rect 6270 5352 6276 5364
rect 5951 5324 6276 5352
rect 5951 5321 5963 5324
rect 5905 5315 5963 5321
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 6362 5312 6368 5364
rect 6420 5352 6426 5364
rect 6638 5352 6644 5364
rect 6420 5324 6644 5352
rect 6420 5312 6426 5324
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 8389 5355 8447 5361
rect 8389 5321 8401 5355
rect 8435 5352 8447 5355
rect 9306 5352 9312 5364
rect 8435 5324 9312 5352
rect 8435 5321 8447 5324
rect 8389 5315 8447 5321
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 9398 5312 9404 5364
rect 9456 5352 9462 5364
rect 13265 5355 13323 5361
rect 9456 5324 13216 5352
rect 9456 5312 9462 5324
rect 3605 5287 3663 5293
rect 3605 5253 3617 5287
rect 3651 5284 3663 5287
rect 3694 5284 3700 5296
rect 3651 5256 3700 5284
rect 3651 5253 3663 5256
rect 3605 5247 3663 5253
rect 3694 5244 3700 5256
rect 3752 5244 3758 5296
rect 7558 5244 7564 5296
rect 7616 5284 7622 5296
rect 8665 5287 8723 5293
rect 8665 5284 8677 5287
rect 7616 5256 8677 5284
rect 7616 5244 7622 5256
rect 8665 5253 8677 5256
rect 8711 5253 8723 5287
rect 13188 5284 13216 5324
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 14366 5352 14372 5364
rect 13311 5324 14372 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 14366 5312 14372 5324
rect 14424 5312 14430 5364
rect 20622 5312 20628 5364
rect 20680 5352 20686 5364
rect 23106 5352 23112 5364
rect 20680 5324 23112 5352
rect 20680 5312 20686 5324
rect 23106 5312 23112 5324
rect 23164 5312 23170 5364
rect 24762 5312 24768 5364
rect 24820 5352 24826 5364
rect 25406 5352 25412 5364
rect 24820 5324 25412 5352
rect 24820 5312 24826 5324
rect 25406 5312 25412 5324
rect 25464 5312 25470 5364
rect 25869 5355 25927 5361
rect 25869 5321 25881 5355
rect 25915 5352 25927 5355
rect 26878 5352 26884 5364
rect 25915 5324 26884 5352
rect 25915 5321 25927 5324
rect 25869 5315 25927 5321
rect 26878 5312 26884 5324
rect 26936 5312 26942 5364
rect 27062 5312 27068 5364
rect 27120 5352 27126 5364
rect 28074 5352 28080 5364
rect 27120 5324 28080 5352
rect 27120 5312 27126 5324
rect 28074 5312 28080 5324
rect 28132 5312 28138 5364
rect 28534 5312 28540 5364
rect 28592 5312 28598 5364
rect 13906 5284 13912 5296
rect 13188 5256 13912 5284
rect 8665 5247 8723 5253
rect 13906 5244 13912 5256
rect 13964 5244 13970 5296
rect 23385 5287 23443 5293
rect 23385 5253 23397 5287
rect 23431 5253 23443 5287
rect 23385 5247 23443 5253
rect 3142 5216 3148 5228
rect 2746 5188 3148 5216
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 3881 5219 3939 5225
rect 3881 5216 3893 5219
rect 3384 5188 3893 5216
rect 3384 5176 3390 5188
rect 3881 5185 3893 5188
rect 3927 5185 3939 5219
rect 3881 5179 3939 5185
rect 4387 5219 4445 5225
rect 4387 5185 4399 5219
rect 4433 5216 4445 5219
rect 5074 5216 5080 5228
rect 4433 5188 5080 5216
rect 4433 5185 4445 5188
rect 4387 5179 4445 5185
rect 5074 5176 5080 5188
rect 5132 5176 5138 5228
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 6595 5219 6653 5225
rect 5684 5188 6224 5216
rect 5684 5176 5690 5188
rect 1264 5151 1322 5157
rect 1264 5117 1276 5151
rect 1310 5148 1322 5151
rect 1578 5148 1584 5160
rect 1310 5120 1584 5148
rect 1310 5117 1322 5120
rect 1264 5111 1322 5117
rect 1578 5108 1584 5120
rect 1636 5108 1642 5160
rect 1673 5151 1731 5157
rect 1673 5117 1685 5151
rect 1719 5148 1731 5151
rect 1946 5148 1952 5160
rect 1719 5120 1952 5148
rect 1719 5117 1731 5120
rect 1673 5111 1731 5117
rect 1946 5108 1952 5120
rect 2004 5108 2010 5160
rect 3786 5108 3792 5160
rect 3844 5148 3850 5160
rect 4208 5151 4266 5157
rect 4208 5148 4220 5151
rect 3844 5120 4220 5148
rect 3844 5108 3850 5120
rect 4208 5117 4220 5120
rect 4254 5117 4266 5151
rect 4208 5111 4266 5117
rect 4614 5108 4620 5160
rect 4672 5108 4678 5160
rect 6089 5151 6147 5157
rect 6089 5117 6101 5151
rect 6135 5117 6147 5151
rect 6196 5148 6224 5188
rect 6595 5185 6607 5219
rect 6641 5216 6653 5219
rect 7650 5216 7656 5228
rect 6641 5188 7656 5216
rect 6641 5185 6653 5188
rect 6595 5179 6653 5185
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 9398 5216 9404 5228
rect 7760 5188 9404 5216
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6196 5120 6837 5148
rect 6089 5111 6147 5117
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 3142 5040 3148 5092
rect 3200 5080 3206 5092
rect 3329 5083 3387 5089
rect 3329 5080 3341 5083
rect 3200 5052 3341 5080
rect 3200 5040 3206 5052
rect 3329 5049 3341 5052
rect 3375 5049 3387 5083
rect 3329 5043 3387 5049
rect 6104 5012 6132 5111
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 7760 5148 7788 5188
rect 9398 5176 9404 5188
rect 9456 5176 9462 5228
rect 9539 5219 9597 5225
rect 9539 5185 9551 5219
rect 9585 5216 9597 5219
rect 9674 5216 9680 5228
rect 9585 5188 9680 5216
rect 9585 5185 9597 5188
rect 9539 5179 9597 5185
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 9766 5174 9772 5226
rect 9824 5174 9830 5226
rect 11146 5176 11152 5228
rect 11204 5216 11210 5228
rect 11204 5188 11652 5216
rect 11204 5176 11210 5188
rect 6972 5120 7788 5148
rect 6972 5108 6978 5120
rect 7926 5108 7932 5160
rect 7984 5148 7990 5160
rect 8573 5151 8631 5157
rect 8573 5148 8585 5151
rect 7984 5120 8585 5148
rect 7984 5108 7990 5120
rect 8573 5117 8585 5120
rect 8619 5117 8631 5151
rect 8573 5111 8631 5117
rect 8849 5151 8907 5157
rect 8849 5117 8861 5151
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 8205 5083 8263 5089
rect 8205 5049 8217 5083
rect 8251 5080 8263 5083
rect 8754 5080 8760 5092
rect 8251 5052 8760 5080
rect 8251 5049 8263 5052
rect 8205 5043 8263 5049
rect 8754 5040 8760 5052
rect 8812 5040 8818 5092
rect 6454 5012 6460 5024
rect 6104 4984 6460 5012
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 6555 5015 6613 5021
rect 6555 4981 6567 5015
rect 6601 5012 6613 5015
rect 6822 5012 6828 5024
rect 6601 4984 6828 5012
rect 6601 4981 6613 4984
rect 6555 4975 6613 4981
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 7098 4972 7104 5024
rect 7156 5012 7162 5024
rect 8386 5012 8392 5024
rect 7156 4984 8392 5012
rect 7156 4972 7162 4984
rect 8386 4972 8392 4984
rect 8444 5012 8450 5024
rect 8864 5012 8892 5111
rect 8938 5108 8944 5160
rect 8996 5148 9002 5160
rect 9033 5151 9091 5157
rect 9033 5148 9045 5151
rect 8996 5120 9045 5148
rect 8996 5108 9002 5120
rect 9033 5117 9045 5120
rect 9079 5117 9091 5151
rect 9033 5111 9091 5117
rect 11241 5151 11299 5157
rect 11241 5117 11253 5151
rect 11287 5148 11299 5151
rect 11514 5148 11520 5160
rect 11287 5120 11520 5148
rect 11287 5117 11299 5120
rect 11241 5111 11299 5117
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 11624 5148 11652 5188
rect 11698 5176 11704 5228
rect 11756 5216 11762 5228
rect 11756 5188 11801 5216
rect 11756 5176 11762 5188
rect 11882 5176 11888 5228
rect 11940 5216 11946 5228
rect 11940 5188 12296 5216
rect 11940 5176 11946 5188
rect 12268 5160 12296 5188
rect 14182 5176 14188 5228
rect 14240 5216 14246 5228
rect 14328 5219 14386 5225
rect 14328 5216 14340 5219
rect 14240 5188 14340 5216
rect 14240 5176 14246 5188
rect 14328 5185 14340 5188
rect 14374 5185 14386 5219
rect 14328 5179 14386 5185
rect 14464 5217 14522 5223
rect 14464 5183 14476 5217
rect 14510 5183 14522 5217
rect 14464 5177 14522 5183
rect 11977 5151 12035 5157
rect 11977 5148 11989 5151
rect 11624 5120 11989 5148
rect 11977 5117 11989 5120
rect 12023 5117 12035 5151
rect 11977 5111 12035 5117
rect 12250 5108 12256 5160
rect 12308 5108 12314 5160
rect 13909 5151 13967 5157
rect 13909 5148 13921 5151
rect 13832 5120 13921 5148
rect 13832 5092 13860 5120
rect 13909 5117 13921 5120
rect 13955 5117 13967 5151
rect 13909 5111 13967 5117
rect 13998 5108 14004 5160
rect 14056 5108 14062 5160
rect 14479 5148 14507 5177
rect 14550 5176 14556 5228
rect 14608 5216 14614 5228
rect 14737 5219 14795 5225
rect 14737 5216 14749 5219
rect 14608 5188 14749 5216
rect 14608 5176 14614 5188
rect 14737 5185 14749 5188
rect 14783 5185 14795 5219
rect 14737 5179 14795 5185
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 16672 5219 16730 5225
rect 16672 5216 16684 5219
rect 16163 5188 16684 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 16672 5185 16684 5188
rect 16718 5185 16730 5219
rect 16672 5179 16730 5185
rect 16942 5176 16948 5228
rect 17000 5176 17006 5228
rect 18325 5219 18383 5225
rect 18325 5185 18337 5219
rect 18371 5216 18383 5219
rect 19156 5219 19214 5225
rect 19156 5216 19168 5219
rect 18371 5188 19168 5216
rect 18371 5185 18383 5188
rect 18325 5179 18383 5185
rect 19156 5185 19168 5188
rect 19202 5185 19214 5219
rect 19156 5179 19214 5185
rect 19429 5219 19487 5225
rect 19429 5185 19441 5219
rect 19475 5216 19487 5219
rect 20530 5216 20536 5228
rect 19475 5188 20536 5216
rect 19475 5185 19487 5188
rect 19429 5179 19487 5185
rect 20530 5176 20536 5188
rect 20588 5176 20594 5228
rect 20809 5219 20867 5225
rect 20809 5185 20821 5219
rect 20855 5216 20867 5219
rect 21364 5219 21422 5225
rect 21364 5216 21376 5219
rect 20855 5188 21376 5216
rect 20855 5185 20867 5188
rect 20809 5179 20867 5185
rect 21364 5185 21376 5188
rect 21410 5185 21422 5219
rect 21364 5179 21422 5185
rect 22002 5176 22008 5228
rect 22060 5216 22066 5228
rect 23400 5216 23428 5247
rect 22060 5176 22094 5216
rect 23400 5188 24072 5216
rect 14108 5120 14507 5148
rect 14108 5092 14136 5120
rect 16206 5108 16212 5160
rect 16264 5108 16270 5160
rect 16574 5157 16580 5160
rect 16536 5151 16580 5157
rect 16536 5117 16548 5151
rect 16536 5111 16580 5117
rect 16574 5108 16580 5111
rect 16632 5108 16638 5160
rect 18690 5108 18696 5160
rect 18748 5108 18754 5160
rect 20901 5151 20959 5157
rect 18800 5120 20760 5148
rect 13814 5080 13820 5092
rect 12636 5052 13820 5080
rect 8444 4984 8892 5012
rect 8444 4972 8450 4984
rect 9030 4972 9036 5024
rect 9088 5012 9094 5024
rect 9499 5015 9557 5021
rect 9499 5012 9511 5015
rect 9088 4984 9511 5012
rect 9088 4972 9094 4984
rect 9499 4981 9511 4984
rect 9545 4981 9557 5015
rect 9499 4975 9557 4981
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 10042 5012 10048 5024
rect 9732 4984 10048 5012
rect 9732 4972 9738 4984
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 11057 5015 11115 5021
rect 11057 4981 11069 5015
rect 11103 5012 11115 5015
rect 11514 5012 11520 5024
rect 11103 4984 11520 5012
rect 11103 4981 11115 4984
rect 11057 4975 11115 4981
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 11707 5015 11765 5021
rect 11707 4981 11719 5015
rect 11753 5012 11765 5015
rect 11882 5012 11888 5024
rect 11753 4984 11888 5012
rect 11753 4981 11765 4984
rect 11707 4975 11765 4981
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 12636 5012 12664 5052
rect 13814 5040 13820 5052
rect 13872 5040 13878 5092
rect 14090 5040 14096 5092
rect 14148 5040 14154 5092
rect 18800 5080 18828 5120
rect 17604 5052 18828 5080
rect 12032 4984 12664 5012
rect 12032 4972 12038 4984
rect 13722 4972 13728 5024
rect 13780 4972 13786 5024
rect 13906 4972 13912 5024
rect 13964 5012 13970 5024
rect 17604 5012 17632 5052
rect 20732 5024 20760 5120
rect 20901 5117 20913 5151
rect 20947 5117 20959 5151
rect 20901 5111 20959 5117
rect 20916 5024 20944 5111
rect 21174 5108 21180 5160
rect 21232 5148 21238 5160
rect 21637 5151 21695 5157
rect 21637 5148 21649 5151
rect 21232 5120 21649 5148
rect 21232 5108 21238 5120
rect 21637 5117 21649 5120
rect 21683 5117 21695 5151
rect 22066 5148 22094 5176
rect 23293 5151 23351 5157
rect 23293 5148 23305 5151
rect 22066 5120 23305 5148
rect 21637 5111 21695 5117
rect 23293 5117 23305 5120
rect 23339 5117 23351 5151
rect 23293 5111 23351 5117
rect 23382 5108 23388 5160
rect 23440 5108 23446 5160
rect 23566 5108 23572 5160
rect 23624 5108 23630 5160
rect 23658 5108 23664 5160
rect 23716 5148 23722 5160
rect 23845 5151 23903 5157
rect 23845 5148 23857 5151
rect 23716 5120 23857 5148
rect 23716 5108 23722 5120
rect 23845 5117 23857 5120
rect 23891 5117 23903 5151
rect 24044 5148 24072 5188
rect 24118 5176 24124 5228
rect 24176 5216 24182 5228
rect 24308 5219 24366 5225
rect 24308 5216 24320 5219
rect 24176 5188 24320 5216
rect 24176 5176 24182 5188
rect 24308 5185 24320 5188
rect 24354 5185 24366 5219
rect 24308 5179 24366 5185
rect 26418 5176 26424 5228
rect 26476 5216 26482 5228
rect 27160 5219 27218 5225
rect 27160 5216 27172 5219
rect 26476 5188 27172 5216
rect 26476 5176 26482 5188
rect 27160 5185 27172 5188
rect 27206 5185 27218 5219
rect 27160 5179 27218 5185
rect 27433 5219 27491 5225
rect 27433 5185 27445 5219
rect 27479 5216 27491 5219
rect 28994 5216 29000 5228
rect 27479 5188 29000 5216
rect 27479 5185 27491 5188
rect 27433 5179 27491 5185
rect 28994 5176 29000 5188
rect 29052 5176 29058 5228
rect 24581 5151 24639 5157
rect 24581 5148 24593 5151
rect 24044 5120 24593 5148
rect 23845 5111 23903 5117
rect 24581 5117 24593 5120
rect 24627 5117 24639 5151
rect 24581 5111 24639 5117
rect 13964 4984 17632 5012
rect 13964 4972 13970 4984
rect 18782 4972 18788 5024
rect 18840 5012 18846 5024
rect 19159 5015 19217 5021
rect 19159 5012 19171 5015
rect 18840 4984 19171 5012
rect 18840 4972 18846 4984
rect 19159 4981 19171 4984
rect 19205 4981 19217 5015
rect 19159 4975 19217 4981
rect 20714 4972 20720 5024
rect 20772 4972 20778 5024
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 21266 5012 21272 5024
rect 20956 4984 21272 5012
rect 20956 4972 20962 4984
rect 21266 4972 21272 4984
rect 21324 4972 21330 5024
rect 21367 5015 21425 5021
rect 21367 4981 21379 5015
rect 21413 5012 21425 5015
rect 21542 5012 21548 5024
rect 21413 4984 21548 5012
rect 21413 4981 21425 4984
rect 21367 4975 21425 4981
rect 21542 4972 21548 4984
rect 21600 4972 21606 5024
rect 22738 4972 22744 5024
rect 22796 4972 22802 5024
rect 23109 5015 23167 5021
rect 23109 4981 23121 5015
rect 23155 5012 23167 5015
rect 23400 5012 23428 5108
rect 23860 5024 23888 5111
rect 25958 5108 25964 5160
rect 26016 5148 26022 5160
rect 26513 5151 26571 5157
rect 26513 5148 26525 5151
rect 26016 5120 26525 5148
rect 26016 5108 26022 5120
rect 26513 5117 26525 5120
rect 26559 5117 26571 5151
rect 26513 5111 26571 5117
rect 26697 5151 26755 5157
rect 26697 5117 26709 5151
rect 26743 5148 26755 5151
rect 27522 5148 27528 5160
rect 26743 5120 27528 5148
rect 26743 5117 26755 5120
rect 26697 5111 26755 5117
rect 23934 5040 23940 5092
rect 23992 5040 23998 5092
rect 26528 5080 26556 5111
rect 27522 5108 27528 5120
rect 27580 5108 27586 5160
rect 26528 5052 26740 5080
rect 23155 4984 23428 5012
rect 23155 4981 23167 4984
rect 23109 4975 23167 4981
rect 23842 4972 23848 5024
rect 23900 4972 23906 5024
rect 23952 5012 23980 5040
rect 24118 5012 24124 5024
rect 23952 4984 24124 5012
rect 24118 4972 24124 4984
rect 24176 5012 24182 5024
rect 24311 5015 24369 5021
rect 24311 5012 24323 5015
rect 24176 4984 24323 5012
rect 24176 4972 24182 4984
rect 24311 4981 24323 4984
rect 24357 4981 24369 5015
rect 24311 4975 24369 4981
rect 26329 5015 26387 5021
rect 26329 4981 26341 5015
rect 26375 5012 26387 5015
rect 26602 5012 26608 5024
rect 26375 4984 26608 5012
rect 26375 4981 26387 4984
rect 26329 4975 26387 4981
rect 26602 4972 26608 4984
rect 26660 4972 26666 5024
rect 26712 5012 26740 5052
rect 27062 5012 27068 5024
rect 26712 4984 27068 5012
rect 27062 4972 27068 4984
rect 27120 4972 27126 5024
rect 27163 5015 27221 5021
rect 27163 4981 27175 5015
rect 27209 5012 27221 5015
rect 28350 5012 28356 5024
rect 27209 4984 28356 5012
rect 27209 4981 27221 4984
rect 27163 4975 27221 4981
rect 28350 4972 28356 4984
rect 28408 4972 28414 5024
rect 552 4922 31072 4944
rect 552 4870 7988 4922
rect 8040 4870 8052 4922
rect 8104 4870 8116 4922
rect 8168 4870 8180 4922
rect 8232 4870 8244 4922
rect 8296 4870 15578 4922
rect 15630 4870 15642 4922
rect 15694 4870 15706 4922
rect 15758 4870 15770 4922
rect 15822 4870 15834 4922
rect 15886 4870 23168 4922
rect 23220 4870 23232 4922
rect 23284 4870 23296 4922
rect 23348 4870 23360 4922
rect 23412 4870 23424 4922
rect 23476 4870 30758 4922
rect 30810 4870 30822 4922
rect 30874 4870 30886 4922
rect 30938 4870 30950 4922
rect 31002 4870 31014 4922
rect 31066 4870 31072 4922
rect 552 4848 31072 4870
rect 1486 4768 1492 4820
rect 1544 4808 1550 4820
rect 2685 4811 2743 4817
rect 2685 4808 2697 4811
rect 1544 4780 2697 4808
rect 1544 4768 1550 4780
rect 2685 4777 2697 4780
rect 2731 4777 2743 4811
rect 2685 4771 2743 4777
rect 3510 4768 3516 4820
rect 3568 4768 3574 4820
rect 3786 4768 3792 4820
rect 3844 4808 3850 4820
rect 3979 4811 4037 4817
rect 3979 4808 3991 4811
rect 3844 4780 3991 4808
rect 3844 4768 3850 4780
rect 3979 4777 3991 4780
rect 4025 4777 4037 4811
rect 3979 4771 4037 4777
rect 7834 4768 7840 4820
rect 7892 4768 7898 4820
rect 9490 4808 9496 4820
rect 8772 4780 9496 4808
rect 842 4632 848 4684
rect 900 4632 906 4684
rect 1854 4672 1860 4684
rect 1228 4644 1860 4672
rect 1228 4613 1256 4644
rect 1854 4632 1860 4644
rect 1912 4632 1918 4684
rect 3326 4632 3332 4684
rect 3384 4632 3390 4684
rect 3418 4632 3424 4684
rect 3476 4632 3482 4684
rect 3528 4672 3556 4768
rect 8772 4740 8800 4780
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 10965 4811 11023 4817
rect 10965 4808 10977 4811
rect 9824 4780 10977 4808
rect 9824 4768 9830 4780
rect 10965 4777 10977 4780
rect 11011 4777 11023 4811
rect 10965 4771 11023 4777
rect 11146 4768 11152 4820
rect 11204 4768 11210 4820
rect 11514 4768 11520 4820
rect 11572 4768 11578 4820
rect 12075 4811 12133 4817
rect 12075 4777 12087 4811
rect 12121 4808 12133 4811
rect 12250 4808 12256 4820
rect 12121 4780 12256 4808
rect 12121 4777 12133 4780
rect 12075 4771 12133 4777
rect 12250 4768 12256 4780
rect 12308 4768 12314 4820
rect 13633 4811 13691 4817
rect 13633 4777 13645 4811
rect 13679 4808 13691 4811
rect 14090 4808 14096 4820
rect 13679 4780 14096 4808
rect 13679 4777 13691 4780
rect 13633 4771 13691 4777
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 14182 4768 14188 4820
rect 14240 4808 14246 4820
rect 14283 4811 14341 4817
rect 14283 4808 14295 4811
rect 14240 4780 14295 4808
rect 14240 4768 14246 4780
rect 14283 4777 14295 4780
rect 14329 4777 14341 4811
rect 14283 4771 14341 4777
rect 16574 4768 16580 4820
rect 16632 4808 16638 4820
rect 16675 4811 16733 4817
rect 16675 4808 16687 4811
rect 16632 4780 16687 4808
rect 16632 4768 16638 4780
rect 16675 4777 16687 4780
rect 16721 4777 16733 4811
rect 16675 4771 16733 4777
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 19435 4811 19493 4817
rect 19435 4808 19447 4811
rect 19392 4780 19447 4808
rect 19392 4768 19398 4780
rect 19435 4777 19447 4780
rect 19481 4808 19493 4811
rect 19978 4808 19984 4820
rect 19481 4780 19984 4808
rect 19481 4777 19493 4780
rect 19435 4771 19493 4777
rect 19978 4768 19984 4780
rect 20036 4768 20042 4820
rect 20162 4768 20168 4820
rect 20220 4808 20226 4820
rect 24213 4811 24271 4817
rect 20220 4780 24164 4808
rect 20220 4768 20226 4780
rect 11164 4740 11192 4768
rect 8588 4712 8800 4740
rect 11072 4712 11192 4740
rect 4249 4675 4307 4681
rect 3528 4644 3648 4672
rect 1172 4607 1256 4613
rect 1172 4573 1184 4607
rect 1218 4576 1256 4607
rect 1351 4607 1409 4613
rect 1218 4573 1230 4576
rect 1172 4567 1230 4573
rect 1351 4573 1363 4607
rect 1397 4604 1409 4607
rect 1486 4604 1492 4616
rect 1397 4576 1492 4604
rect 1397 4573 1409 4576
rect 1351 4567 1409 4573
rect 1486 4564 1492 4576
rect 1544 4564 1550 4616
rect 1578 4564 1584 4616
rect 1636 4564 1642 4616
rect 3234 4604 3240 4616
rect 2746 4576 3240 4604
rect 1486 4428 1492 4480
rect 1544 4468 1550 4480
rect 2746 4468 2774 4576
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 3344 4604 3372 4632
rect 3513 4607 3571 4613
rect 3513 4604 3525 4607
rect 3344 4576 3525 4604
rect 3513 4573 3525 4576
rect 3559 4573 3571 4607
rect 3620 4604 3648 4644
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4982 4672 4988 4684
rect 4295 4644 4988 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4672 5687 4675
rect 5675 4644 6500 4672
rect 5675 4641 5687 4644
rect 5629 4635 5687 4641
rect 3976 4607 4034 4613
rect 3976 4604 3988 4607
rect 3620 4576 3988 4604
rect 3513 4567 3571 4573
rect 3976 4573 3988 4576
rect 4022 4573 4034 4607
rect 3976 4567 4034 4573
rect 4062 4564 4068 4616
rect 4120 4604 4126 4616
rect 4120 4576 5764 4604
rect 4120 4564 4126 4576
rect 5626 4496 5632 4548
rect 5684 4496 5690 4548
rect 1544 4440 2774 4468
rect 1544 4428 1550 4440
rect 3234 4428 3240 4480
rect 3292 4428 3298 4480
rect 3418 4428 3424 4480
rect 3476 4468 3482 4480
rect 5644 4468 5672 4496
rect 3476 4440 5672 4468
rect 5736 4468 5764 4576
rect 5810 4564 5816 4616
rect 5868 4604 5874 4616
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 5868 4576 6009 4604
rect 5868 4564 5874 4576
rect 5997 4573 6009 4576
rect 6043 4573 6055 4607
rect 5997 4567 6055 4573
rect 6178 4564 6184 4616
rect 6236 4604 6242 4616
rect 6472 4615 6500 4644
rect 7190 4632 7196 4684
rect 7248 4672 7254 4684
rect 8588 4681 8616 4712
rect 8573 4675 8631 4681
rect 8573 4672 8585 4675
rect 7248 4644 8585 4672
rect 7248 4632 7254 4644
rect 8573 4641 8585 4644
rect 8619 4641 8631 4675
rect 8573 4635 8631 4641
rect 9490 4632 9496 4684
rect 9548 4672 9554 4684
rect 11072 4672 11100 4712
rect 11238 4700 11244 4752
rect 11296 4740 11302 4752
rect 11532 4740 11560 4768
rect 11296 4712 11468 4740
rect 11532 4712 11750 4740
rect 11296 4700 11302 4712
rect 9548 4644 11100 4672
rect 11149 4675 11207 4681
rect 9548 4632 9554 4644
rect 11149 4641 11161 4675
rect 11195 4672 11207 4675
rect 11330 4672 11336 4684
rect 11195 4644 11336 4672
rect 11195 4641 11207 4644
rect 11149 4635 11207 4641
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 11440 4681 11468 4712
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4641 11483 4675
rect 11425 4635 11483 4641
rect 6324 4607 6382 4613
rect 6324 4604 6336 4607
rect 6236 4576 6336 4604
rect 6236 4564 6242 4576
rect 6324 4573 6336 4576
rect 6370 4573 6382 4607
rect 6324 4567 6382 4573
rect 6460 4609 6518 4615
rect 6460 4575 6472 4609
rect 6506 4575 6518 4609
rect 6460 4569 6518 4575
rect 6733 4607 6791 4613
rect 6733 4573 6745 4607
rect 6779 4604 6791 4607
rect 8294 4604 8300 4616
rect 6779 4576 8300 4604
rect 6779 4573 6791 4576
rect 6733 4567 6791 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4604 8723 4607
rect 8846 4604 8852 4616
rect 8711 4576 8852 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 8846 4564 8852 4576
rect 8904 4564 8910 4616
rect 9030 4613 9036 4616
rect 8992 4607 9036 4613
rect 8992 4573 9004 4607
rect 8992 4567 9036 4573
rect 9030 4564 9036 4567
rect 9088 4564 9094 4616
rect 9128 4609 9186 4615
rect 9128 4575 9140 4609
rect 9174 4604 9186 4609
rect 9214 4604 9220 4616
rect 9174 4576 9220 4604
rect 9174 4575 9186 4576
rect 9128 4569 9186 4575
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4604 9459 4607
rect 11440 4604 11468 4635
rect 11606 4632 11612 4684
rect 11664 4632 11670 4684
rect 11722 4672 11750 4712
rect 13722 4700 13728 4752
rect 13780 4700 13786 4752
rect 18325 4743 18383 4749
rect 18325 4709 18337 4743
rect 18371 4740 18383 4743
rect 18966 4740 18972 4752
rect 18371 4712 18972 4740
rect 18371 4709 18383 4712
rect 18325 4703 18383 4709
rect 18966 4700 18972 4712
rect 19024 4700 19030 4752
rect 24136 4740 24164 4780
rect 24213 4777 24225 4811
rect 24259 4808 24271 4811
rect 24486 4808 24492 4820
rect 24259 4780 24492 4808
rect 24259 4777 24271 4780
rect 24213 4771 24271 4777
rect 24486 4768 24492 4780
rect 24544 4768 24550 4820
rect 24581 4811 24639 4817
rect 24581 4777 24593 4811
rect 24627 4808 24639 4811
rect 26234 4808 26240 4820
rect 24627 4780 26240 4808
rect 24627 4777 24639 4780
rect 24581 4771 24639 4777
rect 26234 4768 26240 4780
rect 26292 4768 26298 4820
rect 29178 4808 29184 4820
rect 26344 4780 29184 4808
rect 26344 4740 26372 4780
rect 29178 4768 29184 4780
rect 29236 4768 29242 4820
rect 21744 4712 22324 4740
rect 24136 4712 26372 4740
rect 12345 4675 12403 4681
rect 11722 4644 12020 4672
rect 11992 4622 12020 4644
rect 12345 4641 12357 4675
rect 12391 4672 12403 4675
rect 13538 4672 13544 4684
rect 12391 4644 13544 4672
rect 12391 4641 12403 4644
rect 12345 4635 12403 4641
rect 13538 4632 13544 4644
rect 13596 4632 13602 4684
rect 13740 4672 13768 4700
rect 14553 4675 14611 4681
rect 14553 4672 14565 4675
rect 13740 4644 14565 4672
rect 14553 4641 14565 4644
rect 14599 4641 14611 4675
rect 14553 4635 14611 4641
rect 15933 4675 15991 4681
rect 15933 4641 15945 4675
rect 15979 4672 15991 4675
rect 16945 4675 17003 4681
rect 15979 4644 16715 4672
rect 15979 4641 15991 4644
rect 15933 4635 15991 4641
rect 12072 4625 12130 4631
rect 12072 4622 12084 4625
rect 11882 4604 11888 4616
rect 9447 4576 11284 4604
rect 11440 4576 11888 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 8389 4539 8447 4545
rect 8389 4505 8401 4539
rect 8435 4536 8447 4539
rect 8478 4536 8484 4548
rect 8435 4508 8484 4536
rect 8435 4505 8447 4508
rect 8389 4499 8447 4505
rect 8478 4496 8484 4508
rect 8536 4496 8542 4548
rect 11256 4545 11284 4576
rect 11882 4564 11888 4576
rect 11940 4564 11946 4616
rect 11992 4594 12084 4622
rect 12072 4591 12084 4594
rect 12118 4591 12130 4625
rect 12072 4585 12130 4591
rect 13817 4607 13875 4613
rect 13817 4573 13829 4607
rect 13863 4604 13875 4607
rect 13998 4604 14004 4616
rect 13863 4576 14004 4604
rect 13863 4573 13875 4576
rect 13817 4567 13875 4573
rect 13998 4564 14004 4576
rect 14056 4564 14062 4616
rect 14274 4564 14280 4616
rect 14332 4604 14338 4616
rect 14332 4576 14377 4604
rect 14332 4564 14338 4576
rect 16206 4564 16212 4616
rect 16264 4564 16270 4616
rect 16687 4615 16715 4644
rect 16945 4641 16957 4675
rect 16991 4672 17003 4675
rect 17218 4672 17224 4684
rect 16991 4644 17224 4672
rect 16991 4641 17003 4644
rect 16945 4635 17003 4641
rect 17218 4632 17224 4644
rect 17276 4632 17282 4684
rect 18046 4632 18052 4684
rect 18104 4632 18110 4684
rect 18414 4632 18420 4684
rect 18472 4672 18478 4684
rect 19058 4672 19064 4684
rect 18472 4644 19064 4672
rect 18472 4632 18478 4644
rect 19058 4632 19064 4644
rect 19116 4632 19122 4684
rect 20438 4672 20444 4684
rect 19490 4644 20444 4672
rect 16672 4609 16730 4615
rect 16672 4575 16684 4609
rect 16718 4575 16730 4609
rect 16672 4569 16730 4575
rect 11241 4539 11299 4545
rect 11241 4505 11253 4539
rect 11287 4505 11299 4539
rect 18064 4536 18092 4632
rect 18693 4607 18751 4613
rect 18693 4573 18705 4607
rect 18739 4604 18751 4607
rect 18782 4604 18788 4616
rect 18739 4576 18788 4604
rect 18739 4573 18751 4576
rect 18693 4567 18751 4573
rect 18782 4564 18788 4576
rect 18840 4564 18846 4616
rect 19490 4613 19518 4644
rect 20438 4632 20444 4644
rect 20496 4632 20502 4684
rect 20530 4632 20536 4684
rect 20588 4672 20594 4684
rect 21744 4681 21772 4712
rect 21453 4675 21511 4681
rect 21453 4672 21465 4675
rect 20588 4644 21465 4672
rect 20588 4632 20594 4644
rect 21453 4641 21465 4644
rect 21499 4672 21511 4675
rect 21729 4675 21787 4681
rect 21729 4672 21741 4675
rect 21499 4644 21741 4672
rect 21499 4641 21511 4644
rect 21453 4635 21511 4641
rect 21729 4641 21741 4644
rect 21775 4641 21787 4675
rect 21729 4635 21787 4641
rect 21910 4632 21916 4684
rect 21968 4672 21974 4684
rect 22005 4675 22063 4681
rect 22005 4672 22017 4675
rect 21968 4644 22017 4672
rect 21968 4632 21974 4644
rect 22005 4641 22017 4644
rect 22051 4641 22063 4675
rect 22005 4635 22063 4641
rect 22189 4675 22247 4681
rect 22189 4641 22201 4675
rect 22235 4641 22247 4675
rect 22296 4672 22324 4712
rect 27522 4700 27528 4752
rect 27580 4740 27586 4752
rect 27580 4712 28028 4740
rect 27580 4700 27586 4712
rect 28000 4684 28028 4712
rect 22296 4644 22876 4672
rect 22189 4635 22247 4641
rect 18969 4607 19027 4613
rect 18969 4573 18981 4607
rect 19015 4573 19027 4607
rect 18969 4567 19027 4573
rect 19475 4607 19533 4613
rect 19475 4573 19487 4607
rect 19521 4573 19533 4607
rect 19475 4567 19533 4573
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4604 19763 4607
rect 20162 4604 20168 4616
rect 19751 4576 20168 4604
rect 19751 4573 19763 4576
rect 19705 4567 19763 4573
rect 18874 4536 18880 4548
rect 18064 4508 18880 4536
rect 11241 4499 11299 4505
rect 18874 4496 18880 4508
rect 18932 4536 18938 4548
rect 18984 4536 19012 4567
rect 20162 4564 20168 4576
rect 20220 4564 20226 4616
rect 22204 4548 22232 4635
rect 22554 4613 22560 4616
rect 22516 4607 22560 4613
rect 22516 4573 22528 4607
rect 22516 4567 22560 4573
rect 22554 4564 22560 4567
rect 22612 4564 22618 4616
rect 22652 4609 22710 4615
rect 22652 4575 22664 4609
rect 22698 4604 22710 4609
rect 22738 4604 22744 4616
rect 22698 4576 22744 4604
rect 22698 4575 22710 4576
rect 22652 4569 22710 4575
rect 22738 4564 22744 4576
rect 22796 4564 22802 4616
rect 22848 4604 22876 4644
rect 22922 4632 22928 4684
rect 22980 4632 22986 4684
rect 23566 4632 23572 4684
rect 23624 4672 23630 4684
rect 24765 4675 24823 4681
rect 24765 4672 24777 4675
rect 23624 4644 24777 4672
rect 23624 4632 23630 4644
rect 24765 4641 24777 4644
rect 24811 4672 24823 4675
rect 27065 4675 27123 4681
rect 27065 4672 27077 4675
rect 24811 4644 27077 4672
rect 24811 4641 24823 4644
rect 24765 4635 24823 4641
rect 27065 4641 27077 4644
rect 27111 4672 27123 4675
rect 27890 4672 27896 4684
rect 27111 4644 27896 4672
rect 27111 4641 27123 4644
rect 27065 4635 27123 4641
rect 27890 4632 27896 4644
rect 27948 4632 27954 4684
rect 27982 4632 27988 4684
rect 28040 4632 28046 4684
rect 28721 4675 28779 4681
rect 28721 4641 28733 4675
rect 28767 4672 28779 4675
rect 30098 4672 30104 4684
rect 28767 4644 30104 4672
rect 28767 4641 28779 4644
rect 28721 4635 28779 4641
rect 30098 4632 30104 4644
rect 30156 4632 30162 4684
rect 25222 4604 25228 4616
rect 22848 4576 25228 4604
rect 25222 4564 25228 4576
rect 25280 4564 25286 4616
rect 28350 4613 28356 4616
rect 28312 4607 28356 4613
rect 28312 4573 28324 4607
rect 28312 4567 28356 4573
rect 28350 4564 28356 4567
rect 28408 4564 28414 4616
rect 28534 4613 28540 4616
rect 28491 4607 28540 4613
rect 28491 4573 28503 4607
rect 28537 4573 28540 4607
rect 28491 4567 28540 4573
rect 28534 4564 28540 4567
rect 28592 4564 28598 4616
rect 18932 4508 19012 4536
rect 20364 4508 22048 4536
rect 18932 4496 18938 4508
rect 9858 4468 9864 4480
rect 5736 4440 9864 4468
rect 3476 4428 3482 4440
rect 9858 4428 9864 4440
rect 9916 4428 9922 4480
rect 10689 4471 10747 4477
rect 10689 4437 10701 4471
rect 10735 4468 10747 4471
rect 12158 4468 12164 4480
rect 10735 4440 12164 4468
rect 10735 4437 10747 4440
rect 10689 4431 10747 4437
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 17402 4468 17408 4480
rect 13872 4440 17408 4468
rect 13872 4428 13878 4440
rect 17402 4428 17408 4440
rect 17460 4468 17466 4480
rect 20364 4468 20392 4508
rect 22020 4480 22048 4508
rect 22186 4496 22192 4548
rect 22244 4496 22250 4548
rect 25774 4496 25780 4548
rect 25832 4536 25838 4548
rect 29825 4539 29883 4545
rect 25832 4508 27016 4536
rect 25832 4496 25838 4508
rect 17460 4440 20392 4468
rect 17460 4428 17466 4440
rect 20990 4428 20996 4480
rect 21048 4428 21054 4480
rect 21266 4428 21272 4480
rect 21324 4428 21330 4480
rect 21542 4428 21548 4480
rect 21600 4428 21606 4480
rect 21818 4428 21824 4480
rect 21876 4428 21882 4480
rect 22002 4428 22008 4480
rect 22060 4428 22066 4480
rect 23658 4428 23664 4480
rect 23716 4468 23722 4480
rect 24762 4468 24768 4480
rect 23716 4440 24768 4468
rect 23716 4428 23722 4440
rect 24762 4428 24768 4440
rect 24820 4428 24826 4480
rect 25038 4428 25044 4480
rect 25096 4428 25102 4480
rect 25958 4428 25964 4480
rect 26016 4468 26022 4480
rect 26786 4468 26792 4480
rect 26016 4440 26792 4468
rect 26016 4428 26022 4440
rect 26786 4428 26792 4440
rect 26844 4428 26850 4480
rect 26878 4428 26884 4480
rect 26936 4428 26942 4480
rect 26988 4468 27016 4508
rect 29825 4505 29837 4539
rect 29871 4505 29883 4539
rect 29825 4499 29883 4505
rect 29840 4468 29868 4499
rect 26988 4440 29868 4468
rect 552 4378 30912 4400
rect 552 4326 4193 4378
rect 4245 4326 4257 4378
rect 4309 4326 4321 4378
rect 4373 4326 4385 4378
rect 4437 4326 4449 4378
rect 4501 4326 11783 4378
rect 11835 4326 11847 4378
rect 11899 4326 11911 4378
rect 11963 4326 11975 4378
rect 12027 4326 12039 4378
rect 12091 4326 19373 4378
rect 19425 4326 19437 4378
rect 19489 4326 19501 4378
rect 19553 4326 19565 4378
rect 19617 4326 19629 4378
rect 19681 4326 26963 4378
rect 27015 4326 27027 4378
rect 27079 4326 27091 4378
rect 27143 4326 27155 4378
rect 27207 4326 27219 4378
rect 27271 4326 30912 4378
rect 552 4304 30912 4326
rect 1394 4224 1400 4276
rect 1452 4264 1458 4276
rect 1854 4264 1860 4276
rect 1452 4236 1860 4264
rect 1452 4224 1458 4236
rect 1854 4224 1860 4236
rect 1912 4264 1918 4276
rect 1912 4236 2774 4264
rect 1912 4224 1918 4236
rect 934 4088 940 4140
rect 992 4088 998 4140
rect 2746 4128 2774 4236
rect 3234 4224 3240 4276
rect 3292 4264 3298 4276
rect 6546 4264 6552 4276
rect 3292 4236 6552 4264
rect 3292 4224 3298 4236
rect 6546 4224 6552 4236
rect 6604 4224 6610 4276
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8941 4267 8999 4273
rect 8941 4264 8953 4267
rect 8352 4236 8953 4264
rect 8352 4224 8358 4236
rect 8941 4233 8953 4236
rect 8987 4233 8999 4267
rect 8941 4227 8999 4233
rect 9766 4224 9772 4276
rect 9824 4264 9830 4276
rect 9824 4236 11560 4264
rect 9824 4224 9830 4236
rect 8386 4156 8392 4208
rect 8444 4196 8450 4208
rect 8444 4168 9812 4196
rect 8444 4156 8450 4168
rect 3513 4131 3571 4137
rect 3513 4128 3525 4131
rect 1458 4119 2176 4128
rect 1433 4113 2176 4119
rect 1433 4079 1445 4113
rect 1479 4100 2176 4113
rect 2746 4100 3525 4128
rect 1479 4079 1491 4100
rect 1433 4073 1491 4079
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4060 1731 4063
rect 1762 4060 1768 4072
rect 1719 4032 1768 4060
rect 1719 4029 1731 4032
rect 1673 4023 1731 4029
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 2148 4060 2176 4100
rect 3513 4097 3525 4100
rect 3559 4128 3571 4131
rect 3602 4128 3608 4140
rect 3559 4100 3608 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 4338 4135 4344 4140
rect 4295 4129 4344 4135
rect 4295 4095 4307 4129
rect 4341 4095 4344 4129
rect 4295 4089 4344 4095
rect 4338 4088 4344 4089
rect 4396 4088 4402 4140
rect 4522 4088 4528 4140
rect 4580 4088 4586 4140
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 6460 4131 6518 4137
rect 6460 4128 6472 4131
rect 5592 4100 6472 4128
rect 5592 4088 5598 4100
rect 6460 4097 6472 4100
rect 6506 4097 6518 4131
rect 6460 4091 6518 4097
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4128 8171 4131
rect 8570 4128 8576 4140
rect 8159 4100 8576 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 8662 4088 8668 4140
rect 8720 4088 8726 4140
rect 2774 4060 2780 4072
rect 2148 4032 2780 4060
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 3237 4063 3295 4069
rect 3237 4029 3249 4063
rect 3283 4060 3295 4063
rect 3283 4032 3372 4060
rect 3283 4029 3295 4032
rect 3237 4023 3295 4029
rect 3344 3936 3372 4032
rect 3786 4020 3792 4072
rect 3844 4020 3850 4072
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 5997 4063 6055 4069
rect 5997 4060 6009 4063
rect 5868 4032 6009 4060
rect 5868 4020 5874 4032
rect 5997 4029 6009 4032
rect 6043 4029 6055 4063
rect 5997 4023 6055 4029
rect 6730 4020 6736 4072
rect 6788 4020 6794 4072
rect 7466 4020 7472 4072
rect 7524 4020 7530 4072
rect 8389 4063 8447 4069
rect 8389 4029 8401 4063
rect 8435 4029 8447 4063
rect 8389 4023 8447 4029
rect 5902 3952 5908 4004
rect 5960 3952 5966 4004
rect 1403 3927 1461 3933
rect 1403 3893 1415 3927
rect 1449 3924 1461 3927
rect 1670 3924 1676 3936
rect 1449 3896 1676 3924
rect 1449 3893 1461 3896
rect 1403 3887 1461 3893
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 2774 3884 2780 3936
rect 2832 3884 2838 3936
rect 3326 3884 3332 3936
rect 3384 3884 3390 3936
rect 4255 3927 4313 3933
rect 4255 3893 4267 3927
rect 4301 3924 4313 3927
rect 4522 3924 4528 3936
rect 4301 3896 4528 3924
rect 4301 3893 4313 3896
rect 4255 3887 4313 3893
rect 4522 3884 4528 3896
rect 4580 3884 4586 3936
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 6463 3927 6521 3933
rect 6463 3924 6475 3927
rect 6328 3896 6475 3924
rect 6328 3884 6334 3896
rect 6463 3893 6475 3896
rect 6509 3893 6521 3927
rect 7484 3924 7512 4020
rect 8404 3992 8432 4023
rect 8938 4020 8944 4072
rect 8996 4020 9002 4072
rect 9122 4020 9128 4072
rect 9180 4020 9186 4072
rect 9784 4069 9812 4168
rect 9858 4156 9864 4208
rect 9916 4156 9922 4208
rect 10042 4156 10048 4208
rect 10100 4156 10106 4208
rect 11532 4196 11560 4236
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 11977 4267 12035 4273
rect 11977 4264 11989 4267
rect 11756 4236 11989 4264
rect 11756 4224 11762 4236
rect 11977 4233 11989 4236
rect 12023 4233 12035 4267
rect 17678 4264 17684 4276
rect 11977 4227 12035 4233
rect 12406 4236 17684 4264
rect 12406 4196 12434 4236
rect 17678 4224 17684 4236
rect 17736 4224 17742 4276
rect 17770 4224 17776 4276
rect 17828 4264 17834 4276
rect 20530 4264 20536 4276
rect 17828 4236 20536 4264
rect 17828 4224 17834 4236
rect 20530 4224 20536 4236
rect 20588 4224 20594 4276
rect 21266 4264 21272 4276
rect 20691 4236 21272 4264
rect 11532 4168 12434 4196
rect 10060 4128 10088 4156
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 10060 4100 10149 4128
rect 10137 4097 10149 4100
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 10600 4131 10658 4137
rect 10600 4128 10612 4131
rect 10376 4100 10612 4128
rect 10376 4088 10382 4100
rect 10600 4097 10612 4100
rect 10646 4097 10658 4131
rect 10600 4091 10658 4097
rect 10778 4088 10784 4140
rect 10836 4128 10842 4140
rect 10873 4131 10931 4137
rect 10873 4128 10885 4131
rect 10836 4100 10885 4128
rect 10836 4088 10842 4100
rect 10873 4097 10885 4100
rect 10919 4097 10931 4131
rect 10873 4091 10931 4097
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 11606 4128 11612 4140
rect 11296 4100 11612 4128
rect 11296 4088 11302 4100
rect 11606 4088 11612 4100
rect 11664 4128 11670 4140
rect 12066 4128 12072 4140
rect 11664 4100 12072 4128
rect 11664 4088 11670 4100
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12250 4088 12256 4140
rect 12308 4128 12314 4140
rect 12529 4131 12587 4137
rect 12529 4128 12541 4131
rect 12308 4100 12541 4128
rect 12308 4088 12314 4100
rect 12529 4097 12541 4100
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 16117 4131 16175 4137
rect 14516 4100 14561 4128
rect 14516 4088 14522 4100
rect 16117 4097 16129 4131
rect 16163 4128 16175 4131
rect 16672 4131 16730 4137
rect 16672 4128 16684 4131
rect 16163 4100 16684 4128
rect 16163 4097 16175 4100
rect 16117 4091 16175 4097
rect 16672 4097 16684 4100
rect 16718 4097 16730 4131
rect 16672 4091 16730 4097
rect 18325 4131 18383 4137
rect 18325 4097 18337 4131
rect 18371 4128 18383 4131
rect 19156 4131 19214 4137
rect 19156 4128 19168 4131
rect 18371 4100 19168 4128
rect 18371 4097 18383 4100
rect 18325 4091 18383 4097
rect 19156 4097 19168 4100
rect 19202 4097 19214 4131
rect 19156 4091 19214 4097
rect 19429 4131 19487 4137
rect 19429 4097 19441 4131
rect 19475 4128 19487 4131
rect 20691 4128 20719 4236
rect 21266 4224 21272 4236
rect 21324 4224 21330 4276
rect 22296 4168 25176 4196
rect 19475 4100 20719 4128
rect 20809 4131 20867 4137
rect 19475 4097 19487 4100
rect 19429 4091 19487 4097
rect 20809 4097 20821 4131
rect 20855 4128 20867 4131
rect 21364 4131 21422 4137
rect 21364 4128 21376 4131
rect 20855 4100 21376 4128
rect 20855 4097 20867 4100
rect 20809 4091 20867 4097
rect 21364 4097 21376 4100
rect 21410 4097 21422 4131
rect 21364 4091 21422 4097
rect 21450 4088 21456 4140
rect 21508 4088 21514 4140
rect 21542 4088 21548 4140
rect 21600 4128 21606 4140
rect 21637 4131 21695 4137
rect 21637 4128 21649 4131
rect 21600 4100 21649 4128
rect 21600 4088 21606 4100
rect 21637 4097 21649 4100
rect 21683 4097 21695 4131
rect 21637 4091 21695 4097
rect 22002 4088 22008 4140
rect 22060 4128 22066 4140
rect 22296 4128 22324 4168
rect 25148 4137 25176 4168
rect 25133 4131 25191 4137
rect 22060 4100 22324 4128
rect 23768 4100 24348 4128
rect 22060 4088 22066 4100
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4060 9551 4063
rect 9769 4063 9827 4069
rect 9539 4032 9720 4060
rect 9539 4029 9551 4032
rect 9493 4023 9551 4029
rect 8956 3992 8984 4020
rect 8404 3964 8984 3992
rect 9140 3924 9168 4020
rect 7484 3896 9168 3924
rect 6463 3887 6521 3893
rect 9306 3884 9312 3936
rect 9364 3884 9370 3936
rect 9398 3884 9404 3936
rect 9456 3924 9462 3936
rect 9585 3927 9643 3933
rect 9585 3924 9597 3927
rect 9456 3896 9597 3924
rect 9456 3884 9462 3896
rect 9585 3893 9597 3896
rect 9631 3893 9643 3927
rect 9692 3924 9720 4032
rect 9769 4029 9781 4063
rect 9815 4029 9827 4063
rect 9769 4023 9827 4029
rect 10045 4063 10103 4069
rect 10045 4029 10057 4063
rect 10091 4060 10103 4063
rect 10410 4060 10416 4072
rect 10091 4032 10416 4060
rect 10091 4029 10103 4032
rect 10045 4023 10103 4029
rect 9784 3992 9812 4023
rect 10134 3992 10140 4004
rect 9784 3964 10140 3992
rect 10134 3952 10140 3964
rect 10192 3952 10198 4004
rect 10244 3924 10272 4032
rect 10410 4020 10416 4032
rect 10468 4060 10474 4072
rect 10468 4032 11560 4060
rect 10468 4020 10474 4032
rect 11532 3992 11560 4032
rect 11882 4020 11888 4072
rect 11940 4060 11946 4072
rect 12345 4063 12403 4069
rect 12345 4060 12357 4063
rect 11940 4032 12357 4060
rect 11940 4020 11946 4032
rect 12345 4029 12357 4032
rect 12391 4060 12403 4063
rect 12710 4060 12716 4072
rect 12391 4032 12716 4060
rect 12391 4029 12403 4032
rect 12345 4023 12403 4029
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 13906 4020 13912 4072
rect 13964 4020 13970 4072
rect 13998 4020 14004 4072
rect 14056 4020 14062 4072
rect 14734 4020 14740 4072
rect 14792 4020 14798 4072
rect 16206 4020 16212 4072
rect 16264 4020 16270 4072
rect 16945 4063 17003 4069
rect 16945 4060 16957 4063
rect 16316 4032 16957 4060
rect 12434 3992 12440 4004
rect 11532 3964 12440 3992
rect 12434 3952 12440 3964
rect 12492 3952 12498 4004
rect 12989 3995 13047 4001
rect 12989 3961 13001 3995
rect 13035 3992 13047 3995
rect 14016 3992 14044 4020
rect 13035 3964 14044 3992
rect 13035 3961 13047 3964
rect 12989 3955 13047 3961
rect 15470 3952 15476 4004
rect 15528 3992 15534 4004
rect 16316 3992 16344 4032
rect 16945 4029 16957 4032
rect 16991 4029 17003 4063
rect 16945 4023 17003 4029
rect 18690 4020 18696 4072
rect 18748 4060 18754 4072
rect 18966 4060 18972 4072
rect 18748 4032 18972 4060
rect 18748 4020 18754 4032
rect 18966 4020 18972 4032
rect 19024 4020 19030 4072
rect 20898 4020 20904 4072
rect 20956 4020 20962 4072
rect 21228 4063 21286 4069
rect 21228 4029 21240 4063
rect 21274 4060 21286 4063
rect 21468 4060 21496 4088
rect 23768 4072 23796 4100
rect 21274 4032 21496 4060
rect 23109 4063 23167 4069
rect 21274 4029 21286 4032
rect 21228 4023 21286 4029
rect 23109 4029 23121 4063
rect 23155 4060 23167 4063
rect 23566 4060 23572 4072
rect 23155 4032 23572 4060
rect 23155 4029 23167 4032
rect 23109 4023 23167 4029
rect 23566 4020 23572 4032
rect 23624 4020 23630 4072
rect 23750 4020 23756 4072
rect 23808 4020 23814 4072
rect 24029 4063 24087 4069
rect 24029 4029 24041 4063
rect 24075 4060 24087 4063
rect 24210 4060 24216 4072
rect 24075 4032 24216 4060
rect 24075 4029 24087 4032
rect 24029 4023 24087 4029
rect 24210 4020 24216 4032
rect 24268 4020 24274 4072
rect 24320 4069 24348 4100
rect 25133 4097 25145 4131
rect 25179 4097 25191 4131
rect 25133 4091 25191 4097
rect 26142 4088 26148 4140
rect 26200 4128 26206 4140
rect 26424 4131 26482 4137
rect 26424 4128 26436 4131
rect 26200 4100 26436 4128
rect 26200 4088 26206 4100
rect 26424 4097 26436 4100
rect 26470 4097 26482 4131
rect 26424 4091 26482 4097
rect 26510 4088 26516 4140
rect 26568 4088 26574 4140
rect 26602 4088 26608 4140
rect 26660 4128 26666 4140
rect 26697 4131 26755 4137
rect 26697 4128 26709 4131
rect 26660 4100 26709 4128
rect 26660 4088 26666 4100
rect 26697 4097 26709 4100
rect 26743 4097 26755 4131
rect 29546 4128 29552 4140
rect 26697 4091 26755 4097
rect 29012 4100 29552 4128
rect 24305 4063 24363 4069
rect 24305 4029 24317 4063
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 24578 4020 24584 4072
rect 24636 4020 24642 4072
rect 24854 4020 24860 4072
rect 24912 4020 24918 4072
rect 25958 4020 25964 4072
rect 26016 4020 26022 4072
rect 26528 4060 26556 4088
rect 27430 4060 27436 4072
rect 26528 4032 27436 4060
rect 27430 4020 27436 4032
rect 27488 4020 27494 4072
rect 28166 4020 28172 4072
rect 28224 4020 28230 4072
rect 29012 4069 29040 4100
rect 29546 4088 29552 4100
rect 29604 4088 29610 4140
rect 28997 4063 29055 4069
rect 28997 4029 29009 4063
rect 29043 4029 29055 4063
rect 28997 4023 29055 4029
rect 15528 3964 16344 3992
rect 15528 3952 15534 3964
rect 22554 3952 22560 4004
rect 22612 3992 22618 4004
rect 23385 3995 23443 4001
rect 23385 3992 23397 3995
rect 22612 3964 23397 3992
rect 22612 3952 22618 3964
rect 23385 3961 23397 3964
rect 23431 3992 23443 3995
rect 23431 3964 24072 3992
rect 23431 3961 23443 3964
rect 23385 3955 23443 3961
rect 24044 3936 24072 3964
rect 27356 3964 29224 3992
rect 9692 3896 10272 3924
rect 9585 3887 9643 3893
rect 10594 3884 10600 3936
rect 10652 3933 10658 3936
rect 10652 3924 10661 3933
rect 10652 3896 10697 3924
rect 10652 3887 10661 3896
rect 10652 3884 10658 3887
rect 12066 3884 12072 3936
rect 12124 3924 12130 3936
rect 13081 3927 13139 3933
rect 13081 3924 13093 3927
rect 12124 3896 13093 3924
rect 12124 3884 12130 3896
rect 13081 3893 13093 3896
rect 13127 3893 13139 3927
rect 13081 3887 13139 3893
rect 13722 3884 13728 3936
rect 13780 3884 13786 3936
rect 14274 3884 14280 3936
rect 14332 3924 14338 3936
rect 14467 3927 14525 3933
rect 14467 3924 14479 3927
rect 14332 3896 14479 3924
rect 14332 3884 14338 3896
rect 14467 3893 14479 3896
rect 14513 3893 14525 3927
rect 14467 3887 14525 3893
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 16675 3927 16733 3933
rect 16675 3924 16687 3927
rect 16632 3896 16687 3924
rect 16632 3884 16638 3896
rect 16675 3893 16687 3896
rect 16721 3893 16733 3927
rect 16675 3887 16733 3893
rect 18782 3884 18788 3936
rect 18840 3924 18846 3936
rect 19159 3927 19217 3933
rect 19159 3924 19171 3927
rect 18840 3896 19171 3924
rect 18840 3884 18846 3896
rect 19159 3893 19171 3896
rect 19205 3893 19217 3927
rect 19159 3887 19217 3893
rect 22738 3884 22744 3936
rect 22796 3884 22802 3936
rect 22922 3884 22928 3936
rect 22980 3924 22986 3936
rect 23845 3927 23903 3933
rect 23845 3924 23857 3927
rect 22980 3896 23857 3924
rect 22980 3884 22986 3896
rect 23845 3893 23857 3896
rect 23891 3893 23903 3927
rect 23845 3887 23903 3893
rect 24026 3884 24032 3936
rect 24084 3884 24090 3936
rect 24118 3884 24124 3936
rect 24176 3884 24182 3936
rect 24394 3884 24400 3936
rect 24452 3884 24458 3936
rect 24670 3884 24676 3936
rect 24728 3884 24734 3936
rect 25498 3884 25504 3936
rect 25556 3884 25562 3936
rect 26418 3884 26424 3936
rect 26476 3933 26482 3936
rect 26476 3924 26485 3933
rect 26476 3896 26521 3924
rect 26476 3887 26485 3896
rect 26476 3884 26482 3887
rect 26602 3884 26608 3936
rect 26660 3924 26666 3936
rect 27356 3924 27384 3964
rect 26660 3896 27384 3924
rect 26660 3884 26666 3896
rect 27522 3884 27528 3936
rect 27580 3924 27586 3936
rect 27801 3927 27859 3933
rect 27801 3924 27813 3927
rect 27580 3896 27813 3924
rect 27580 3884 27586 3896
rect 27801 3893 27813 3896
rect 27847 3893 27859 3927
rect 27801 3887 27859 3893
rect 28350 3884 28356 3936
rect 28408 3884 28414 3936
rect 29196 3933 29224 3964
rect 29181 3927 29239 3933
rect 29181 3893 29193 3927
rect 29227 3893 29239 3927
rect 29181 3887 29239 3893
rect 552 3834 31072 3856
rect 552 3782 7988 3834
rect 8040 3782 8052 3834
rect 8104 3782 8116 3834
rect 8168 3782 8180 3834
rect 8232 3782 8244 3834
rect 8296 3782 15578 3834
rect 15630 3782 15642 3834
rect 15694 3782 15706 3834
rect 15758 3782 15770 3834
rect 15822 3782 15834 3834
rect 15886 3782 23168 3834
rect 23220 3782 23232 3834
rect 23284 3782 23296 3834
rect 23348 3782 23360 3834
rect 23412 3782 23424 3834
rect 23476 3782 30758 3834
rect 30810 3782 30822 3834
rect 30874 3782 30886 3834
rect 30938 3782 30950 3834
rect 31002 3782 31014 3834
rect 31066 3782 31072 3834
rect 552 3760 31072 3782
rect 1029 3723 1087 3729
rect 1029 3689 1041 3723
rect 1075 3720 1087 3723
rect 6730 3720 6736 3732
rect 1075 3692 6736 3720
rect 1075 3689 1087 3692
rect 1029 3683 1087 3689
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 6923 3723 6981 3729
rect 6923 3720 6935 3723
rect 6880 3692 6935 3720
rect 6880 3680 6886 3692
rect 6923 3689 6935 3692
rect 6969 3720 6981 3723
rect 8662 3720 8668 3732
rect 6969 3692 8668 3720
rect 6969 3689 6981 3692
rect 6923 3683 6981 3689
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 10594 3720 10600 3732
rect 9088 3692 10600 3720
rect 9088 3680 9094 3692
rect 10594 3680 10600 3692
rect 10652 3720 10658 3732
rect 11517 3723 11575 3729
rect 10652 3692 11284 3720
rect 10652 3680 10658 3692
rect 2774 3652 2780 3664
rect 2746 3612 2780 3652
rect 2832 3612 2838 3664
rect 3421 3655 3479 3661
rect 3421 3621 3433 3655
rect 3467 3652 3479 3655
rect 3602 3652 3608 3664
rect 3467 3624 3608 3652
rect 3467 3621 3479 3624
rect 3421 3615 3479 3621
rect 3602 3612 3608 3624
rect 3660 3612 3666 3664
rect 5000 3624 6592 3652
rect 1213 3587 1271 3593
rect 1213 3584 1225 3587
rect 1044 3556 1225 3584
rect 1044 3528 1072 3556
rect 1213 3553 1225 3556
rect 1259 3553 1271 3587
rect 2746 3584 2774 3612
rect 1213 3547 1271 3553
rect 1964 3556 2774 3584
rect 1801 3537 1859 3543
rect 1801 3534 1813 3537
rect 1026 3476 1032 3528
rect 1084 3476 1090 3528
rect 1670 3525 1676 3528
rect 1305 3519 1363 3525
rect 1305 3485 1317 3519
rect 1351 3485 1363 3519
rect 1305 3479 1363 3485
rect 1632 3519 1676 3525
rect 1632 3485 1644 3519
rect 1632 3479 1676 3485
rect 1320 3380 1348 3479
rect 1670 3476 1676 3479
rect 1728 3476 1734 3528
rect 1780 3503 1813 3534
rect 1847 3516 1859 3537
rect 1964 3516 1992 3556
rect 4062 3544 4068 3596
rect 4120 3584 4126 3596
rect 5000 3584 5028 3624
rect 4120 3556 5028 3584
rect 4120 3544 4126 3556
rect 5350 3544 5356 3596
rect 5408 3544 5414 3596
rect 5997 3587 6055 3593
rect 5997 3553 6009 3587
rect 6043 3584 6055 3587
rect 6454 3584 6460 3596
rect 6043 3556 6460 3584
rect 6043 3553 6055 3556
rect 5997 3547 6055 3553
rect 6454 3544 6460 3556
rect 6512 3544 6518 3596
rect 6564 3584 6592 3624
rect 10134 3612 10140 3664
rect 10192 3652 10198 3664
rect 11256 3661 11284 3692
rect 11517 3689 11529 3723
rect 11563 3720 11575 3723
rect 14093 3723 14151 3729
rect 11563 3692 12204 3720
rect 11563 3689 11575 3692
rect 11517 3683 11575 3689
rect 11241 3655 11299 3661
rect 10192 3624 11100 3652
rect 10192 3612 10198 3624
rect 7193 3587 7251 3593
rect 6564 3556 7144 3584
rect 3976 3537 4034 3543
rect 1847 3503 1992 3516
rect 1780 3488 1992 3503
rect 2038 3476 2044 3528
rect 2096 3476 2102 3528
rect 3234 3476 3240 3528
rect 3292 3516 3298 3528
rect 3513 3519 3571 3525
rect 3513 3516 3525 3519
rect 3292 3488 3525 3516
rect 3292 3476 3298 3488
rect 3513 3485 3525 3488
rect 3559 3485 3571 3519
rect 3513 3479 3571 3485
rect 3694 3476 3700 3528
rect 3752 3518 3758 3528
rect 3840 3519 3898 3525
rect 3840 3518 3852 3519
rect 3752 3490 3852 3518
rect 3752 3476 3758 3490
rect 3840 3485 3852 3490
rect 3886 3485 3898 3519
rect 3976 3503 3988 3537
rect 4022 3516 4034 3537
rect 4154 3516 4160 3528
rect 4022 3503 4160 3516
rect 3976 3497 4160 3503
rect 3991 3488 4160 3497
rect 3840 3479 3898 3485
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 5368 3516 5396 3544
rect 4295 3488 5396 3516
rect 5629 3519 5687 3525
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 5629 3485 5641 3519
rect 5675 3516 5687 3519
rect 6270 3516 6276 3528
rect 5675 3488 6276 3516
rect 5675 3485 5687 3488
rect 5629 3479 5687 3485
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 7006 3525 7012 3528
rect 6963 3519 7012 3525
rect 6963 3485 6975 3519
rect 7009 3485 7012 3519
rect 6963 3479 7012 3485
rect 7006 3476 7012 3479
rect 7064 3476 7070 3528
rect 7116 3516 7144 3556
rect 7193 3553 7205 3587
rect 7239 3584 7251 3587
rect 7558 3584 7564 3596
rect 7239 3556 7564 3584
rect 7239 3553 7251 3556
rect 7193 3547 7251 3553
rect 7558 3544 7564 3556
rect 7616 3544 7622 3596
rect 8573 3587 8631 3593
rect 8573 3553 8585 3587
rect 8619 3584 8631 3587
rect 8619 3556 9171 3584
rect 8619 3553 8631 3556
rect 8573 3547 8631 3553
rect 8294 3516 8300 3528
rect 7116 3488 8300 3516
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 8665 3519 8723 3525
rect 8665 3485 8677 3519
rect 8711 3516 8723 3519
rect 8846 3516 8852 3528
rect 8711 3488 8852 3516
rect 8711 3485 8723 3488
rect 8665 3479 8723 3485
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 9030 3525 9036 3528
rect 8992 3519 9036 3525
rect 8992 3485 9004 3519
rect 8992 3479 9036 3485
rect 9030 3476 9036 3479
rect 9088 3476 9094 3528
rect 9143 3527 9171 3556
rect 9398 3544 9404 3596
rect 9456 3544 9462 3596
rect 9674 3544 9680 3596
rect 9732 3584 9738 3596
rect 10226 3584 10232 3596
rect 9732 3556 10232 3584
rect 9732 3544 9738 3556
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 10965 3587 11023 3593
rect 10965 3553 10977 3587
rect 11011 3553 11023 3587
rect 11072 3584 11100 3624
rect 11241 3621 11253 3655
rect 11287 3621 11299 3655
rect 11241 3615 11299 3621
rect 11701 3587 11759 3593
rect 11701 3584 11713 3587
rect 11072 3556 11713 3584
rect 10965 3547 11023 3553
rect 11701 3553 11713 3556
rect 11747 3584 11759 3587
rect 11977 3587 12035 3593
rect 11977 3584 11989 3587
rect 11747 3556 11989 3584
rect 11747 3553 11759 3556
rect 11701 3547 11759 3553
rect 11977 3553 11989 3556
rect 12023 3553 12035 3587
rect 11977 3547 12035 3553
rect 9128 3521 9186 3527
rect 9128 3487 9140 3521
rect 9174 3487 9186 3521
rect 9128 3481 9186 3487
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 9582 3516 9588 3528
rect 9364 3488 9588 3516
rect 9364 3476 9370 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10980 3516 11008 3547
rect 11882 3516 11888 3528
rect 10980 3488 11888 3516
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 5810 3408 5816 3460
rect 5868 3448 5874 3460
rect 6181 3451 6239 3457
rect 6181 3448 6193 3451
rect 5868 3420 6193 3448
rect 5868 3408 5874 3420
rect 6181 3417 6193 3420
rect 6227 3417 6239 3451
rect 6181 3411 6239 3417
rect 10505 3451 10563 3457
rect 10505 3417 10517 3451
rect 10551 3448 10563 3451
rect 11992 3448 12020 3547
rect 12066 3544 12072 3596
rect 12124 3544 12130 3596
rect 12176 3584 12204 3692
rect 14093 3689 14105 3723
rect 14139 3720 14151 3723
rect 14458 3720 14464 3732
rect 14139 3692 14464 3720
rect 14139 3689 14151 3692
rect 14093 3683 14151 3689
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 15841 3723 15899 3729
rect 15841 3720 15853 3723
rect 15028 3692 15853 3720
rect 15028 3661 15056 3692
rect 15841 3689 15853 3692
rect 15887 3720 15899 3723
rect 16206 3720 16212 3732
rect 15887 3692 16212 3720
rect 15887 3689 15899 3692
rect 15841 3683 15899 3689
rect 16206 3680 16212 3692
rect 16264 3680 16270 3732
rect 27065 3723 27123 3729
rect 27065 3720 27077 3723
rect 16408 3692 19012 3720
rect 15013 3655 15071 3661
rect 15013 3621 15025 3655
rect 15059 3621 15071 3655
rect 15013 3615 15071 3621
rect 15565 3655 15623 3661
rect 15565 3621 15577 3655
rect 15611 3652 15623 3655
rect 16408 3652 16436 3692
rect 18984 3664 19012 3692
rect 19076 3692 27077 3720
rect 15611 3624 16436 3652
rect 16485 3655 16543 3661
rect 15611 3621 15623 3624
rect 15565 3615 15623 3621
rect 16485 3621 16497 3655
rect 16531 3652 16543 3655
rect 16574 3652 16580 3664
rect 16531 3624 16580 3652
rect 16531 3621 16543 3624
rect 16485 3615 16543 3621
rect 16574 3612 16580 3624
rect 16632 3612 16638 3664
rect 18966 3612 18972 3664
rect 19024 3612 19030 3664
rect 12805 3587 12863 3593
rect 12805 3584 12817 3587
rect 12176 3556 12817 3584
rect 12805 3553 12817 3556
rect 12851 3553 12863 3587
rect 12805 3547 12863 3553
rect 13262 3544 13268 3596
rect 13320 3584 13326 3596
rect 14461 3587 14519 3593
rect 14461 3584 14473 3587
rect 13320 3556 14473 3584
rect 13320 3544 13326 3556
rect 14461 3553 14473 3556
rect 14507 3553 14519 3587
rect 14461 3547 14519 3553
rect 16209 3587 16267 3593
rect 16209 3553 16221 3587
rect 16255 3584 16267 3587
rect 17497 3587 17555 3593
rect 16255 3556 17448 3584
rect 16255 3553 16267 3556
rect 16209 3547 16267 3553
rect 12250 3476 12256 3528
rect 12308 3516 12314 3528
rect 12396 3519 12454 3525
rect 12396 3516 12408 3519
rect 12308 3488 12408 3516
rect 12308 3476 12314 3488
rect 12396 3485 12408 3488
rect 12442 3485 12454 3519
rect 12396 3479 12454 3485
rect 12526 3476 12532 3528
rect 12584 3476 12590 3528
rect 15286 3476 15292 3528
rect 15344 3516 15350 3528
rect 16758 3516 16764 3528
rect 15344 3488 16764 3516
rect 15344 3476 15350 3488
rect 16758 3476 16764 3488
rect 16816 3476 16822 3528
rect 17126 3525 17132 3528
rect 17088 3519 17132 3525
rect 17088 3485 17100 3519
rect 17088 3479 17132 3485
rect 17126 3476 17132 3479
rect 17184 3476 17190 3528
rect 17218 3476 17224 3528
rect 17276 3525 17282 3528
rect 17276 3519 17325 3525
rect 17276 3485 17279 3519
rect 17313 3485 17325 3519
rect 17420 3516 17448 3556
rect 17497 3553 17509 3587
rect 17543 3584 17555 3587
rect 19076 3584 19104 3692
rect 27065 3689 27077 3692
rect 27111 3689 27123 3723
rect 28166 3720 28172 3732
rect 27065 3683 27123 3689
rect 27172 3692 28172 3720
rect 20898 3612 20904 3664
rect 20956 3652 20962 3664
rect 21361 3655 21419 3661
rect 21361 3652 21373 3655
rect 20956 3624 21373 3652
rect 20956 3612 20962 3624
rect 21361 3621 21373 3624
rect 21407 3621 21419 3655
rect 21361 3615 21419 3621
rect 21634 3612 21640 3664
rect 21692 3612 21698 3664
rect 25222 3612 25228 3664
rect 25280 3652 25286 3664
rect 25280 3624 25360 3652
rect 25280 3612 25286 3624
rect 19334 3593 19340 3596
rect 17543 3556 19104 3584
rect 19296 3587 19340 3593
rect 17543 3553 17555 3556
rect 17497 3547 17555 3553
rect 19296 3553 19308 3587
rect 19296 3547 19340 3553
rect 19334 3544 19340 3547
rect 19392 3544 19398 3596
rect 21085 3587 21143 3593
rect 19628 3556 20852 3584
rect 18414 3516 18420 3528
rect 17420 3488 18420 3516
rect 17276 3479 17325 3485
rect 17276 3476 17282 3479
rect 18414 3476 18420 3488
rect 18472 3476 18478 3528
rect 18598 3476 18604 3528
rect 18656 3516 18662 3528
rect 18874 3516 18880 3528
rect 18656 3488 18880 3516
rect 18656 3476 18662 3488
rect 18874 3476 18880 3488
rect 18932 3516 18938 3528
rect 18969 3519 19027 3525
rect 18969 3516 18981 3519
rect 18932 3488 18981 3516
rect 18932 3476 18938 3488
rect 18969 3485 18981 3488
rect 19015 3485 19027 3519
rect 18969 3479 19027 3485
rect 19475 3519 19533 3525
rect 19475 3485 19487 3519
rect 19521 3516 19533 3519
rect 19628 3516 19656 3556
rect 19521 3488 19656 3516
rect 19705 3519 19763 3525
rect 19521 3485 19533 3488
rect 19475 3479 19533 3485
rect 19705 3485 19717 3519
rect 19751 3516 19763 3519
rect 20622 3516 20628 3528
rect 19751 3488 20628 3516
rect 19751 3485 19763 3488
rect 19705 3479 19763 3485
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 12066 3448 12072 3460
rect 10551 3420 11928 3448
rect 11992 3420 12072 3448
rect 10551 3417 10563 3420
rect 10505 3411 10563 3417
rect 1578 3380 1584 3392
rect 1320 3352 1584 3380
rect 1578 3340 1584 3352
rect 1636 3340 1642 3392
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 3694 3380 3700 3392
rect 1728 3352 3700 3380
rect 1728 3340 1734 3352
rect 3694 3340 3700 3352
rect 3752 3340 3758 3392
rect 4338 3340 4344 3392
rect 4396 3380 4402 3392
rect 4614 3380 4620 3392
rect 4396 3352 4620 3380
rect 4396 3340 4402 3352
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 6362 3340 6368 3392
rect 6420 3380 6426 3392
rect 8938 3380 8944 3392
rect 6420 3352 8944 3380
rect 6420 3340 6426 3352
rect 8938 3340 8944 3352
rect 8996 3380 9002 3392
rect 11606 3380 11612 3392
rect 8996 3352 11612 3380
rect 8996 3340 9002 3352
rect 11606 3340 11612 3352
rect 11664 3340 11670 3392
rect 11698 3340 11704 3392
rect 11756 3380 11762 3392
rect 11793 3383 11851 3389
rect 11793 3380 11805 3383
rect 11756 3352 11805 3380
rect 11756 3340 11762 3352
rect 11793 3349 11805 3352
rect 11839 3349 11851 3383
rect 11900 3380 11928 3420
rect 12066 3408 12072 3420
rect 12124 3408 12130 3460
rect 14090 3408 14096 3460
rect 14148 3448 14154 3460
rect 15197 3451 15255 3457
rect 15197 3448 15209 3451
rect 14148 3420 15209 3448
rect 14148 3408 14154 3420
rect 15197 3417 15209 3420
rect 15243 3417 15255 3451
rect 20824 3448 20852 3556
rect 21085 3553 21097 3587
rect 21131 3584 21143 3587
rect 21652 3584 21680 3612
rect 25332 3608 25360 3624
rect 25516 3624 26740 3652
rect 25409 3611 25467 3617
rect 25409 3608 25421 3611
rect 22554 3593 22560 3596
rect 22005 3587 22063 3593
rect 22005 3584 22017 3587
rect 21131 3556 21680 3584
rect 21928 3556 22017 3584
rect 21131 3553 21143 3556
rect 21085 3547 21143 3553
rect 21928 3528 21956 3556
rect 22005 3553 22017 3556
rect 22051 3553 22063 3587
rect 22005 3547 22063 3553
rect 22516 3587 22560 3593
rect 22516 3553 22528 3587
rect 22516 3547 22560 3553
rect 22554 3544 22560 3547
rect 22612 3544 22618 3596
rect 22922 3544 22928 3596
rect 22980 3544 22986 3596
rect 24673 3587 24731 3593
rect 24581 3571 24639 3577
rect 24581 3537 24593 3571
rect 24627 3537 24639 3571
rect 24673 3553 24685 3587
rect 24719 3584 24731 3587
rect 24762 3584 24768 3596
rect 24719 3556 24768 3584
rect 24719 3553 24731 3556
rect 24673 3547 24731 3553
rect 24762 3544 24768 3556
rect 24820 3544 24826 3596
rect 25332 3580 25421 3608
rect 25409 3577 25421 3580
rect 25455 3608 25467 3611
rect 25516 3608 25544 3624
rect 25455 3580 25544 3608
rect 25455 3577 25467 3580
rect 25409 3571 25467 3577
rect 25590 3544 25596 3596
rect 25648 3584 25654 3596
rect 25685 3587 25743 3593
rect 25685 3584 25697 3587
rect 25648 3556 25697 3584
rect 25648 3544 25654 3556
rect 25685 3553 25697 3556
rect 25731 3553 25743 3587
rect 25685 3547 25743 3553
rect 25866 3544 25872 3596
rect 25924 3584 25930 3596
rect 26712 3593 26740 3624
rect 25961 3587 26019 3593
rect 25961 3584 25973 3587
rect 25924 3556 25973 3584
rect 25924 3544 25930 3556
rect 25961 3553 25973 3556
rect 26007 3553 26019 3587
rect 25961 3547 26019 3553
rect 26697 3587 26755 3593
rect 26697 3553 26709 3587
rect 26743 3584 26755 3587
rect 27172 3584 27200 3692
rect 28166 3680 28172 3692
rect 28224 3680 28230 3732
rect 28994 3680 29000 3732
rect 29052 3720 29058 3732
rect 29733 3723 29791 3729
rect 29733 3720 29745 3723
rect 29052 3692 29745 3720
rect 29052 3680 29058 3692
rect 29733 3689 29745 3692
rect 29779 3689 29791 3723
rect 29733 3683 29791 3689
rect 27264 3624 27844 3652
rect 27264 3593 27292 3624
rect 26743 3556 27200 3584
rect 27249 3587 27307 3593
rect 26743 3553 26755 3556
rect 26697 3547 26755 3553
rect 27249 3553 27261 3587
rect 27295 3553 27307 3587
rect 27249 3547 27307 3553
rect 27341 3587 27399 3593
rect 27341 3553 27353 3587
rect 27387 3584 27399 3587
rect 27430 3584 27436 3596
rect 27387 3556 27436 3584
rect 27387 3553 27399 3556
rect 27341 3547 27399 3553
rect 27430 3544 27436 3556
rect 27488 3544 27494 3596
rect 24581 3531 24639 3537
rect 21910 3476 21916 3528
rect 21968 3476 21974 3528
rect 22186 3476 22192 3528
rect 22244 3476 22250 3528
rect 22652 3521 22710 3527
rect 22652 3487 22664 3521
rect 22698 3516 22710 3521
rect 22738 3516 22744 3528
rect 22698 3488 22744 3516
rect 22698 3487 22710 3488
rect 22652 3481 22710 3487
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 20824 3420 22094 3448
rect 15197 3411 15255 3417
rect 22066 3392 22094 3420
rect 12526 3380 12532 3392
rect 11900 3352 12532 3380
rect 11793 3343 11851 3349
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 13630 3340 13636 3392
rect 13688 3380 13694 3392
rect 14553 3383 14611 3389
rect 14553 3380 14565 3383
rect 13688 3352 14565 3380
rect 13688 3340 13694 3352
rect 14553 3349 14565 3352
rect 14599 3349 14611 3383
rect 14553 3343 14611 3349
rect 14642 3340 14648 3392
rect 14700 3380 14706 3392
rect 18601 3383 18659 3389
rect 18601 3380 18613 3383
rect 14700 3352 18613 3380
rect 14700 3340 14706 3352
rect 18601 3349 18613 3352
rect 18647 3349 18659 3383
rect 18601 3343 18659 3349
rect 18966 3340 18972 3392
rect 19024 3380 19030 3392
rect 21453 3383 21511 3389
rect 21453 3380 21465 3383
rect 19024 3352 21465 3380
rect 19024 3340 19030 3352
rect 21453 3349 21465 3352
rect 21499 3349 21511 3383
rect 21453 3343 21511 3349
rect 21542 3340 21548 3392
rect 21600 3380 21606 3392
rect 21821 3383 21879 3389
rect 21821 3380 21833 3383
rect 21600 3352 21833 3380
rect 21600 3340 21606 3352
rect 21821 3349 21833 3352
rect 21867 3349 21879 3383
rect 22066 3352 22100 3392
rect 21821 3343 21879 3349
rect 22094 3340 22100 3352
rect 22152 3340 22158 3392
rect 22204 3380 22232 3476
rect 23842 3380 23848 3392
rect 22204 3352 23848 3380
rect 23842 3340 23848 3352
rect 23900 3340 23906 3392
rect 24210 3340 24216 3392
rect 24268 3340 24274 3392
rect 24397 3383 24455 3389
rect 24397 3349 24409 3383
rect 24443 3380 24455 3383
rect 24486 3380 24492 3392
rect 24443 3352 24492 3380
rect 24443 3349 24455 3352
rect 24397 3343 24455 3349
rect 24486 3340 24492 3352
rect 24544 3340 24550 3392
rect 24596 3380 24624 3531
rect 24946 3476 24952 3528
rect 25004 3476 25010 3528
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 27525 3519 27583 3525
rect 27525 3516 27537 3519
rect 26568 3488 27537 3516
rect 26568 3476 26574 3488
rect 27525 3485 27537 3488
rect 27571 3485 27583 3519
rect 27525 3479 27583 3485
rect 25590 3448 25596 3460
rect 25148 3420 25596 3448
rect 25148 3380 25176 3420
rect 25590 3408 25596 3420
rect 25648 3408 25654 3460
rect 25774 3408 25780 3460
rect 25832 3408 25838 3460
rect 24596 3352 25176 3380
rect 25222 3340 25228 3392
rect 25280 3340 25286 3392
rect 25498 3340 25504 3392
rect 25556 3340 25562 3392
rect 25866 3340 25872 3392
rect 25924 3380 25930 3392
rect 26513 3383 26571 3389
rect 26513 3380 26525 3383
rect 25924 3352 26525 3380
rect 25924 3340 25930 3352
rect 26513 3349 26525 3352
rect 26559 3349 26571 3383
rect 27816 3380 27844 3624
rect 27893 3587 27951 3593
rect 27893 3553 27905 3587
rect 27939 3584 27951 3587
rect 27982 3584 27988 3596
rect 27939 3556 27988 3584
rect 27939 3553 27951 3556
rect 27893 3547 27951 3553
rect 27982 3544 27988 3556
rect 28040 3544 28046 3596
rect 28220 3587 28278 3593
rect 28220 3553 28232 3587
rect 28266 3584 28278 3587
rect 28266 3556 28488 3584
rect 28266 3553 28278 3556
rect 28220 3547 28278 3553
rect 28460 3528 28488 3556
rect 28626 3544 28632 3596
rect 28684 3544 28690 3596
rect 28350 3476 28356 3528
rect 28408 3476 28414 3528
rect 28442 3476 28448 3528
rect 28500 3476 28506 3528
rect 29546 3408 29552 3460
rect 29604 3408 29610 3460
rect 29564 3380 29592 3408
rect 27816 3352 29592 3380
rect 26513 3343 26571 3349
rect 552 3290 30912 3312
rect 552 3238 4193 3290
rect 4245 3238 4257 3290
rect 4309 3238 4321 3290
rect 4373 3238 4385 3290
rect 4437 3238 4449 3290
rect 4501 3238 11783 3290
rect 11835 3238 11847 3290
rect 11899 3238 11911 3290
rect 11963 3238 11975 3290
rect 12027 3238 12039 3290
rect 12091 3238 19373 3290
rect 19425 3238 19437 3290
rect 19489 3238 19501 3290
rect 19553 3238 19565 3290
rect 19617 3238 19629 3290
rect 19681 3238 26963 3290
rect 27015 3238 27027 3290
rect 27079 3238 27091 3290
rect 27143 3238 27155 3290
rect 27207 3238 27219 3290
rect 27271 3238 30912 3290
rect 552 3216 30912 3238
rect 1578 3136 1584 3188
rect 1636 3176 1642 3188
rect 2961 3179 3019 3185
rect 1636 3148 2360 3176
rect 1636 3136 1642 3148
rect 2332 3108 2360 3148
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 3050 3176 3056 3188
rect 3007 3148 3056 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 3234 3136 3240 3188
rect 3292 3136 3298 3188
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 6362 3176 6368 3188
rect 3384 3148 6368 3176
rect 3384 3136 3390 3148
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 9674 3176 9680 3188
rect 8128 3148 9680 3176
rect 3252 3108 3280 3136
rect 2332 3080 3280 3108
rect 934 3000 940 3052
rect 992 3000 998 3052
rect 2958 3040 2964 3052
rect 1458 3031 2964 3040
rect 1433 3025 2964 3031
rect 1433 2991 1445 3025
rect 1479 3012 2964 3025
rect 1479 2991 1491 3012
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 1433 2985 1491 2991
rect 1670 2932 1676 2984
rect 1728 2932 1734 2984
rect 3344 2981 3372 3136
rect 3602 3068 3608 3120
rect 3660 3068 3666 3120
rect 3620 3040 3648 3068
rect 4344 3043 4402 3049
rect 4344 3040 4356 3043
rect 3620 3012 4356 3040
rect 4344 3009 4356 3012
rect 4390 3009 4402 3043
rect 4344 3003 4402 3009
rect 4617 3043 4675 3049
rect 4617 3009 4629 3043
rect 4663 3040 4675 3043
rect 5258 3040 5264 3052
rect 4663 3012 5264 3040
rect 4663 3009 4675 3012
rect 4617 3003 4675 3009
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 5810 3000 5816 3052
rect 5868 3000 5874 3052
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3040 6055 3043
rect 6552 3043 6610 3049
rect 6552 3040 6564 3043
rect 6043 3012 6564 3040
rect 6043 3009 6055 3012
rect 5997 3003 6055 3009
rect 6552 3009 6564 3012
rect 6598 3009 6610 3043
rect 6552 3003 6610 3009
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3040 6883 3043
rect 8128 3040 8156 3148
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 9916 3148 11008 3176
rect 9916 3136 9922 3148
rect 6871 3012 8156 3040
rect 8205 3043 8263 3049
rect 6871 3009 6883 3012
rect 6825 3003 6883 3009
rect 8205 3009 8217 3043
rect 8251 3040 8263 3043
rect 9496 3043 9554 3049
rect 9496 3040 9508 3043
rect 8251 3012 9508 3040
rect 8251 3009 8263 3012
rect 8205 3003 8263 3009
rect 9496 3009 9508 3012
rect 9542 3009 9554 3043
rect 9496 3003 9554 3009
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 9640 3012 9812 3040
rect 9640 3000 9646 3012
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2972 3663 2975
rect 3694 2972 3700 2984
rect 3651 2944 3700 2972
rect 3651 2941 3663 2944
rect 3605 2935 3663 2941
rect 3694 2932 3700 2944
rect 3752 2932 3758 2984
rect 3881 2975 3939 2981
rect 3881 2941 3893 2975
rect 3927 2972 3939 2975
rect 5828 2972 5856 3000
rect 3927 2944 5856 2972
rect 6089 2975 6147 2981
rect 3927 2941 3939 2944
rect 3881 2935 3939 2941
rect 6089 2941 6101 2975
rect 6135 2972 6147 2975
rect 6454 2972 6460 2984
rect 6135 2944 6460 2972
rect 6135 2941 6147 2944
rect 6089 2935 6147 2941
rect 1403 2839 1461 2845
rect 1403 2805 1415 2839
rect 1449 2836 1461 2839
rect 1762 2836 1768 2848
rect 1449 2808 1768 2836
rect 1449 2805 1461 2808
rect 1403 2799 1461 2805
rect 1762 2796 1768 2808
rect 1820 2796 1826 2848
rect 1946 2796 1952 2848
rect 2004 2836 2010 2848
rect 3896 2836 3924 2935
rect 6454 2932 6460 2944
rect 6512 2972 6518 2984
rect 8573 2975 8631 2981
rect 6512 2944 7512 2972
rect 6512 2932 6518 2944
rect 6178 2864 6184 2916
rect 6236 2864 6242 2916
rect 2004 2808 3924 2836
rect 2004 2796 2010 2808
rect 4154 2796 4160 2848
rect 4212 2836 4218 2848
rect 4347 2839 4405 2845
rect 4347 2836 4359 2839
rect 4212 2808 4359 2836
rect 4212 2796 4218 2808
rect 4347 2805 4359 2808
rect 4393 2836 4405 2839
rect 6196 2836 6224 2864
rect 4393 2808 6224 2836
rect 6555 2839 6613 2845
rect 4393 2805 4405 2808
rect 4347 2799 4405 2805
rect 6555 2805 6567 2839
rect 6601 2836 6613 2839
rect 6914 2836 6920 2848
rect 6601 2808 6920 2836
rect 6601 2805 6613 2808
rect 6555 2799 6613 2805
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7484 2836 7512 2944
rect 8573 2941 8585 2975
rect 8619 2972 8631 2975
rect 8846 2972 8852 2984
rect 8619 2944 8852 2972
rect 8619 2941 8631 2944
rect 8573 2935 8631 2941
rect 8846 2932 8852 2944
rect 8904 2972 8910 2984
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 8904 2944 9045 2972
rect 8904 2932 8910 2944
rect 9033 2941 9045 2944
rect 9079 2972 9091 2975
rect 9306 2972 9312 2984
rect 9079 2944 9312 2972
rect 9079 2941 9091 2944
rect 9033 2935 9091 2941
rect 9306 2932 9312 2944
rect 9364 2932 9370 2984
rect 9784 2981 9812 3012
rect 9769 2975 9827 2981
rect 9769 2941 9781 2975
rect 9815 2941 9827 2975
rect 9769 2935 9827 2941
rect 10980 2904 11008 3148
rect 11698 3136 11704 3188
rect 11756 3176 11762 3188
rect 14734 3176 14740 3188
rect 11756 3148 14740 3176
rect 11756 3136 11762 3148
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 16574 3136 16580 3188
rect 16632 3176 16638 3188
rect 17126 3176 17132 3188
rect 16632 3148 17132 3176
rect 16632 3136 16638 3148
rect 17126 3136 17132 3148
rect 17184 3136 17190 3188
rect 21542 3176 21548 3188
rect 20640 3148 21548 3176
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 11704 3043 11762 3049
rect 11704 3040 11716 3043
rect 11195 3012 11716 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 11704 3009 11716 3012
rect 11750 3009 11762 3043
rect 11704 3003 11762 3009
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 13357 3043 13415 3049
rect 11848 3012 12434 3040
rect 11848 3000 11854 3012
rect 11238 2932 11244 2984
rect 11296 2932 11302 2984
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11348 2944 11989 2972
rect 11348 2904 11376 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 12406 2972 12434 3012
rect 13357 3009 13369 3043
rect 13403 3040 13415 3043
rect 14556 3043 14614 3049
rect 14556 3040 14568 3043
rect 13403 3012 14568 3040
rect 13403 3009 13415 3012
rect 13357 3003 13415 3009
rect 14556 3009 14568 3012
rect 14602 3009 14614 3043
rect 14556 3003 14614 3009
rect 16209 3043 16267 3049
rect 16209 3009 16221 3043
rect 16255 3040 16267 3043
rect 16764 3043 16822 3049
rect 16764 3040 16776 3043
rect 16255 3012 16776 3040
rect 16255 3009 16267 3012
rect 16209 3003 16267 3009
rect 16764 3009 16776 3012
rect 16810 3009 16822 3043
rect 16764 3003 16822 3009
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3040 18475 3043
rect 19156 3043 19214 3049
rect 19156 3040 19168 3043
rect 18463 3012 19168 3040
rect 18463 3009 18475 3012
rect 18417 3003 18475 3009
rect 19156 3009 19168 3012
rect 19202 3009 19214 3043
rect 19156 3003 19214 3009
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3040 19487 3043
rect 20640 3040 20668 3148
rect 21542 3136 21548 3148
rect 21600 3136 21606 3188
rect 22094 3136 22100 3188
rect 22152 3176 22158 3188
rect 22152 3148 28212 3176
rect 22152 3136 22158 3148
rect 28184 3120 28212 3148
rect 28166 3068 28172 3120
rect 28224 3068 28230 3120
rect 19475 3012 20668 3040
rect 20809 3043 20867 3049
rect 19475 3009 19487 3012
rect 19429 3003 19487 3009
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 21364 3043 21422 3049
rect 21364 3040 21376 3043
rect 20855 3012 21376 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 21364 3009 21376 3012
rect 21410 3009 21422 3043
rect 21364 3003 21422 3009
rect 21450 3000 21456 3052
rect 21508 3000 21514 3052
rect 21637 3043 21695 3049
rect 21637 3009 21649 3043
rect 21683 3040 21695 3043
rect 21818 3040 21824 3052
rect 21683 3012 21824 3040
rect 21683 3009 21695 3012
rect 21637 3003 21695 3009
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 23017 3043 23075 3049
rect 23017 3009 23029 3043
rect 23063 3040 23075 3043
rect 24308 3043 24366 3049
rect 24308 3040 24320 3043
rect 23063 3012 24320 3040
rect 23063 3009 23075 3012
rect 23017 3003 23075 3009
rect 24308 3009 24320 3012
rect 24354 3009 24366 3043
rect 24308 3003 24366 3009
rect 24486 3000 24492 3052
rect 24544 3040 24550 3052
rect 24581 3043 24639 3049
rect 24581 3040 24593 3043
rect 24544 3012 24593 3040
rect 24544 3000 24550 3012
rect 24581 3009 24593 3012
rect 24627 3009 24639 3043
rect 25958 3040 25964 3052
rect 24581 3003 24639 3009
rect 25792 3012 25964 3040
rect 13541 2975 13599 2981
rect 13541 2972 13553 2975
rect 12406 2944 13553 2972
rect 11977 2935 12035 2941
rect 13541 2941 13553 2944
rect 13587 2972 13599 2975
rect 13630 2972 13636 2984
rect 13587 2944 13636 2972
rect 13587 2941 13599 2944
rect 13541 2935 13599 2941
rect 13630 2932 13636 2944
rect 13688 2932 13694 2984
rect 14090 2932 14096 2984
rect 14148 2932 14154 2984
rect 14182 2932 14188 2984
rect 14240 2972 14246 2984
rect 14420 2975 14478 2981
rect 14420 2972 14432 2975
rect 14240 2944 14432 2972
rect 14240 2932 14246 2944
rect 14420 2941 14432 2944
rect 14466 2941 14478 2975
rect 14420 2935 14478 2941
rect 14826 2932 14832 2984
rect 14884 2932 14890 2984
rect 16666 2981 16672 2984
rect 16301 2975 16359 2981
rect 16301 2972 16313 2975
rect 16224 2944 16313 2972
rect 10980 2876 11376 2904
rect 13817 2907 13875 2913
rect 13817 2873 13829 2907
rect 13863 2904 13875 2907
rect 14200 2904 14228 2932
rect 16224 2916 16252 2944
rect 16301 2941 16313 2944
rect 16347 2941 16359 2975
rect 16301 2935 16359 2941
rect 16628 2975 16672 2981
rect 16628 2941 16640 2975
rect 16628 2935 16672 2941
rect 16666 2932 16672 2935
rect 16724 2932 16730 2984
rect 17034 2932 17040 2984
rect 17092 2932 17098 2984
rect 18506 2932 18512 2984
rect 18564 2972 18570 2984
rect 18690 2972 18696 2984
rect 18564 2944 18696 2972
rect 18564 2932 18570 2944
rect 18690 2932 18696 2944
rect 18748 2972 18754 2984
rect 18966 2972 18972 2984
rect 18748 2944 18972 2972
rect 18748 2932 18754 2944
rect 18966 2932 18972 2944
rect 19024 2932 19030 2984
rect 20898 2932 20904 2984
rect 20956 2932 20962 2984
rect 21228 2975 21286 2981
rect 21228 2941 21240 2975
rect 21274 2972 21286 2975
rect 21468 2972 21496 3000
rect 25792 2984 25820 3012
rect 25958 3000 25964 3012
rect 26016 3040 26022 3052
rect 26418 3049 26424 3052
rect 26053 3043 26111 3049
rect 26053 3040 26065 3043
rect 26016 3012 26065 3040
rect 26016 3000 26022 3012
rect 26053 3009 26065 3012
rect 26099 3009 26111 3043
rect 26053 3003 26111 3009
rect 26380 3043 26424 3049
rect 26380 3009 26392 3043
rect 26380 3003 26424 3009
rect 26418 3000 26424 3003
rect 26476 3000 26482 3052
rect 26516 3043 26574 3049
rect 26516 3009 26528 3043
rect 26562 3009 26574 3043
rect 26516 3003 26574 3009
rect 22002 2972 22008 2984
rect 21274 2944 22008 2972
rect 21274 2941 21286 2944
rect 21228 2935 21286 2941
rect 22002 2932 22008 2944
rect 22060 2932 22066 2984
rect 23201 2975 23259 2981
rect 23201 2941 23213 2975
rect 23247 2972 23259 2975
rect 23842 2972 23848 2984
rect 23247 2944 23848 2972
rect 23247 2941 23259 2944
rect 23201 2935 23259 2941
rect 23842 2932 23848 2944
rect 23900 2932 23906 2984
rect 25774 2932 25780 2984
rect 25832 2932 25838 2984
rect 26531 2972 26559 3003
rect 26694 3000 26700 3052
rect 26752 3040 26758 3052
rect 26789 3043 26847 3049
rect 26789 3040 26801 3043
rect 26752 3012 26801 3040
rect 26752 3000 26758 3012
rect 26789 3009 26801 3012
rect 26835 3009 26847 3043
rect 26789 3003 26847 3009
rect 26970 3000 26976 3052
rect 27028 3000 27034 3052
rect 28997 3043 29055 3049
rect 28997 3009 29009 3043
rect 29043 3040 29055 3043
rect 29086 3040 29092 3052
rect 29043 3012 29092 3040
rect 29043 3009 29055 3012
rect 28997 3003 29055 3009
rect 29086 3000 29092 3012
rect 29144 3000 29150 3052
rect 26988 2972 27016 3000
rect 26531 2944 27016 2972
rect 29270 2932 29276 2984
rect 29328 2932 29334 2984
rect 13863 2876 14228 2904
rect 13863 2873 13875 2876
rect 13817 2867 13875 2873
rect 16206 2864 16212 2916
rect 16264 2864 16270 2916
rect 8386 2836 8392 2848
rect 7484 2808 8392 2836
rect 8386 2796 8392 2808
rect 8444 2836 8450 2848
rect 8665 2839 8723 2845
rect 8665 2836 8677 2839
rect 8444 2808 8677 2836
rect 8444 2796 8450 2808
rect 8665 2805 8677 2808
rect 8711 2805 8723 2839
rect 8665 2799 8723 2805
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9499 2839 9557 2845
rect 9499 2836 9511 2839
rect 9088 2808 9511 2836
rect 9088 2796 9094 2808
rect 9499 2805 9511 2808
rect 9545 2805 9557 2839
rect 9499 2799 9557 2805
rect 11707 2839 11765 2845
rect 11707 2805 11719 2839
rect 11753 2836 11765 2839
rect 11974 2836 11980 2848
rect 11753 2808 11980 2836
rect 11753 2805 11765 2808
rect 11707 2799 11765 2805
rect 11974 2796 11980 2808
rect 12032 2836 12038 2848
rect 12250 2836 12256 2848
rect 12032 2808 12256 2836
rect 12032 2796 12038 2808
rect 12250 2796 12256 2808
rect 12308 2796 12314 2848
rect 18782 2796 18788 2848
rect 18840 2836 18846 2848
rect 19159 2839 19217 2845
rect 19159 2836 19171 2839
rect 18840 2808 19171 2836
rect 18840 2796 18846 2808
rect 19159 2805 19171 2808
rect 19205 2805 19217 2839
rect 20916 2836 20944 2932
rect 22664 2876 22876 2904
rect 22664 2836 22692 2876
rect 20916 2808 22692 2836
rect 22848 2836 22876 2876
rect 25958 2864 25964 2916
rect 26016 2864 26022 2916
rect 23293 2839 23351 2845
rect 23293 2836 23305 2839
rect 22848 2808 23305 2836
rect 19159 2799 19217 2805
rect 23293 2805 23305 2808
rect 23339 2805 23351 2839
rect 23293 2799 23351 2805
rect 24118 2796 24124 2848
rect 24176 2836 24182 2848
rect 24311 2839 24369 2845
rect 24311 2836 24323 2839
rect 24176 2808 24323 2836
rect 24176 2796 24182 2808
rect 24311 2805 24323 2808
rect 24357 2805 24369 2839
rect 24311 2799 24369 2805
rect 26786 2796 26792 2848
rect 26844 2836 26850 2848
rect 27893 2839 27951 2845
rect 27893 2836 27905 2839
rect 26844 2808 27905 2836
rect 26844 2796 26850 2808
rect 27893 2805 27905 2808
rect 27939 2805 27951 2839
rect 27893 2799 27951 2805
rect 552 2746 31072 2768
rect 552 2694 7988 2746
rect 8040 2694 8052 2746
rect 8104 2694 8116 2746
rect 8168 2694 8180 2746
rect 8232 2694 8244 2746
rect 8296 2694 15578 2746
rect 15630 2694 15642 2746
rect 15694 2694 15706 2746
rect 15758 2694 15770 2746
rect 15822 2694 15834 2746
rect 15886 2694 23168 2746
rect 23220 2694 23232 2746
rect 23284 2694 23296 2746
rect 23348 2694 23360 2746
rect 23412 2694 23424 2746
rect 23476 2694 30758 2746
rect 30810 2694 30822 2746
rect 30874 2694 30886 2746
rect 30938 2694 30950 2746
rect 31002 2694 31014 2746
rect 31066 2694 31072 2746
rect 552 2672 31072 2694
rect 1495 2635 1553 2641
rect 1495 2601 1507 2635
rect 1541 2632 1553 2635
rect 2038 2632 2044 2644
rect 1541 2604 2044 2632
rect 1541 2601 1553 2604
rect 1495 2595 1553 2601
rect 2038 2592 2044 2604
rect 2096 2592 2102 2644
rect 3053 2635 3111 2641
rect 2746 2604 3004 2632
rect 1029 2499 1087 2505
rect 1029 2465 1041 2499
rect 1075 2496 1087 2499
rect 1854 2496 1860 2508
rect 1075 2468 1860 2496
rect 1075 2465 1087 2468
rect 1029 2459 1087 2465
rect 1854 2456 1860 2468
rect 1912 2456 1918 2508
rect 1535 2431 1593 2437
rect 1535 2397 1547 2431
rect 1581 2428 1593 2431
rect 1670 2428 1676 2440
rect 1581 2400 1676 2428
rect 1581 2397 1593 2400
rect 1535 2391 1593 2397
rect 1670 2388 1676 2400
rect 1728 2388 1734 2440
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 2746 2428 2774 2604
rect 2976 2496 3004 2604
rect 3053 2601 3065 2635
rect 3099 2632 3111 2635
rect 4062 2632 4068 2644
rect 3099 2604 4068 2632
rect 3099 2601 3111 2604
rect 3053 2595 3111 2601
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 4614 2592 4620 2644
rect 4672 2632 4678 2644
rect 5077 2635 5135 2641
rect 5077 2632 5089 2635
rect 4672 2604 5089 2632
rect 4672 2592 4678 2604
rect 5077 2601 5089 2604
rect 5123 2601 5135 2635
rect 5077 2595 5135 2601
rect 6178 2592 6184 2644
rect 6236 2632 6242 2644
rect 6279 2635 6337 2641
rect 6279 2632 6291 2635
rect 6236 2604 6291 2632
rect 6236 2592 6242 2604
rect 6279 2601 6291 2604
rect 6325 2632 6337 2635
rect 6638 2632 6644 2644
rect 6325 2604 6644 2632
rect 6325 2601 6337 2604
rect 6279 2595 6337 2601
rect 6638 2592 6644 2604
rect 6696 2592 6702 2644
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 7653 2635 7711 2641
rect 7653 2632 7665 2635
rect 7064 2604 7665 2632
rect 7064 2592 7070 2604
rect 7653 2601 7665 2604
rect 7699 2601 7711 2635
rect 7653 2595 7711 2601
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 9131 2635 9189 2641
rect 9131 2632 9143 2635
rect 9088 2604 9143 2632
rect 9088 2592 9094 2604
rect 9131 2601 9143 2604
rect 9177 2601 9189 2635
rect 9131 2595 9189 2601
rect 9306 2592 9312 2644
rect 9364 2632 9370 2644
rect 10042 2632 10048 2644
rect 9364 2604 10048 2632
rect 9364 2592 9370 2604
rect 10042 2592 10048 2604
rect 10100 2632 10106 2644
rect 11149 2635 11207 2641
rect 11149 2632 11161 2635
rect 10100 2604 11161 2632
rect 10100 2592 10106 2604
rect 11149 2601 11161 2604
rect 11195 2601 11207 2635
rect 11149 2595 11207 2601
rect 11514 2592 11520 2644
rect 11572 2632 11578 2644
rect 15286 2632 15292 2644
rect 11572 2604 15292 2632
rect 11572 2592 11578 2604
rect 15286 2592 15292 2604
rect 15344 2592 15350 2644
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 16675 2635 16733 2641
rect 16675 2632 16687 2635
rect 16632 2604 16687 2632
rect 16632 2592 16638 2604
rect 16675 2601 16687 2604
rect 16721 2601 16733 2635
rect 16675 2595 16733 2601
rect 17218 2592 17224 2644
rect 17276 2632 17282 2644
rect 21634 2632 21640 2644
rect 17276 2604 21640 2632
rect 17276 2592 17282 2604
rect 21634 2592 21640 2604
rect 21692 2592 21698 2644
rect 21735 2635 21793 2641
rect 21735 2601 21747 2635
rect 21781 2632 21793 2635
rect 22002 2632 22008 2644
rect 21781 2604 22008 2632
rect 21781 2601 21793 2604
rect 21735 2595 21793 2601
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 23842 2592 23848 2644
rect 23900 2592 23906 2644
rect 24210 2592 24216 2644
rect 24268 2592 24274 2644
rect 25774 2592 25780 2644
rect 25832 2632 25838 2644
rect 27617 2635 27675 2641
rect 27617 2632 27629 2635
rect 25832 2604 27629 2632
rect 25832 2592 25838 2604
rect 27617 2601 27629 2604
rect 27663 2601 27675 2635
rect 27617 2595 27675 2601
rect 28442 2592 28448 2644
rect 28500 2641 28506 2644
rect 28500 2595 28509 2641
rect 28500 2592 28506 2595
rect 29362 2592 29368 2644
rect 29420 2632 29426 2644
rect 29825 2635 29883 2641
rect 29825 2632 29837 2635
rect 29420 2604 29837 2632
rect 29420 2592 29426 2604
rect 29825 2601 29837 2604
rect 29871 2601 29883 2635
rect 29825 2595 29883 2601
rect 8297 2567 8355 2573
rect 8297 2533 8309 2567
rect 8343 2564 8355 2567
rect 8662 2564 8668 2576
rect 8343 2536 8668 2564
rect 8343 2533 8355 2536
rect 8297 2527 8355 2533
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 10781 2567 10839 2573
rect 10781 2533 10793 2567
rect 10827 2564 10839 2567
rect 10827 2536 11750 2564
rect 10827 2533 10839 2536
rect 10781 2527 10839 2533
rect 3564 2499 3622 2505
rect 2976 2468 3464 2496
rect 3436 2440 3464 2468
rect 3564 2465 3576 2499
rect 3610 2496 3622 2499
rect 5629 2499 5687 2505
rect 3610 2468 4108 2496
rect 3610 2465 3622 2468
rect 3564 2459 3622 2465
rect 4080 2440 4108 2468
rect 5629 2465 5641 2499
rect 5675 2496 5687 2499
rect 7650 2496 7656 2508
rect 5675 2468 7656 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 8021 2499 8079 2505
rect 8021 2465 8033 2499
rect 8067 2496 8079 2499
rect 8754 2496 8760 2508
rect 8067 2468 8760 2496
rect 8067 2465 8079 2468
rect 8021 2459 8079 2465
rect 8754 2456 8760 2468
rect 8812 2456 8818 2508
rect 9306 2496 9312 2508
rect 9054 2468 9312 2496
rect 1811 2400 2774 2428
rect 3237 2431 3295 2437
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 3237 2397 3249 2431
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 3252 2292 3280 2391
rect 3418 2388 3424 2440
rect 3476 2388 3482 2440
rect 3786 2437 3792 2440
rect 3743 2431 3792 2437
rect 3743 2397 3755 2431
rect 3789 2397 3792 2431
rect 3743 2391 3792 2397
rect 3786 2388 3792 2391
rect 3844 2388 3850 2440
rect 3970 2388 3976 2440
rect 4028 2388 4034 2440
rect 4062 2388 4068 2440
rect 4120 2388 4126 2440
rect 5810 2388 5816 2440
rect 5868 2388 5874 2440
rect 6270 2388 6276 2440
rect 6328 2428 6334 2440
rect 6328 2400 6373 2428
rect 6328 2388 6334 2400
rect 6546 2388 6552 2440
rect 6604 2388 6610 2440
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2428 8723 2431
rect 9054 2428 9082 2468
rect 9306 2456 9312 2468
rect 9364 2456 9370 2508
rect 9398 2456 9404 2508
rect 9456 2456 9462 2508
rect 11057 2499 11115 2505
rect 11057 2465 11069 2499
rect 11103 2496 11115 2499
rect 11238 2496 11244 2508
rect 11103 2468 11244 2496
rect 11103 2465 11115 2468
rect 11057 2459 11115 2465
rect 11238 2456 11244 2468
rect 11296 2496 11302 2508
rect 11609 2499 11667 2505
rect 11609 2496 11621 2499
rect 11296 2468 11621 2496
rect 11296 2456 11302 2468
rect 11609 2465 11621 2468
rect 11655 2465 11667 2499
rect 11722 2496 11750 2536
rect 20530 2524 20536 2576
rect 20588 2524 20594 2576
rect 11992 2496 12115 2500
rect 11722 2472 12115 2496
rect 11722 2468 12020 2472
rect 11609 2459 11667 2465
rect 8711 2400 9082 2428
rect 8711 2397 8723 2400
rect 8665 2391 8723 2397
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 11974 2437 11980 2440
rect 11936 2431 11980 2437
rect 11936 2428 11948 2431
rect 11848 2400 11948 2428
rect 11848 2388 11854 2400
rect 11936 2397 11948 2400
rect 11936 2391 11980 2397
rect 11974 2388 11980 2391
rect 12032 2388 12038 2440
rect 12087 2439 12115 2472
rect 13725 2499 13783 2505
rect 13725 2465 13737 2499
rect 13771 2496 13783 2499
rect 13771 2468 14320 2496
rect 13771 2465 13783 2468
rect 13725 2459 13783 2465
rect 12072 2433 12130 2439
rect 12072 2399 12084 2433
rect 12118 2399 12130 2433
rect 12072 2393 12130 2399
rect 12158 2388 12164 2440
rect 12216 2428 12222 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12216 2400 12357 2428
rect 12216 2388 12222 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 13817 2431 13875 2437
rect 13817 2397 13829 2431
rect 13863 2428 13875 2431
rect 13998 2428 14004 2440
rect 13863 2400 14004 2428
rect 13863 2397 13875 2400
rect 13817 2391 13875 2397
rect 13998 2388 14004 2400
rect 14056 2388 14062 2440
rect 14182 2437 14188 2440
rect 14144 2431 14188 2437
rect 14144 2397 14156 2431
rect 14144 2391 14188 2397
rect 14182 2388 14188 2391
rect 14240 2388 14246 2440
rect 14292 2437 14320 2468
rect 16114 2456 16120 2508
rect 16172 2496 16178 2508
rect 16209 2499 16267 2505
rect 16209 2496 16221 2499
rect 16172 2468 16221 2496
rect 16172 2456 16178 2468
rect 16209 2465 16221 2468
rect 16255 2465 16267 2499
rect 16209 2459 16267 2465
rect 18414 2456 18420 2508
rect 18472 2456 18478 2508
rect 18782 2505 18788 2508
rect 18744 2499 18788 2505
rect 18744 2465 18756 2499
rect 18744 2459 18788 2465
rect 18782 2456 18788 2459
rect 18840 2456 18846 2508
rect 19242 2456 19248 2508
rect 19300 2496 19306 2508
rect 20625 2499 20683 2505
rect 20625 2496 20637 2499
rect 19300 2468 20637 2496
rect 19300 2456 19306 2468
rect 20625 2465 20637 2468
rect 20671 2465 20683 2499
rect 20625 2459 20683 2465
rect 18880 2449 18938 2455
rect 14280 2431 14338 2437
rect 14280 2397 14292 2431
rect 14326 2397 14338 2431
rect 14280 2391 14338 2397
rect 14550 2388 14556 2440
rect 14608 2388 14614 2440
rect 15933 2431 15991 2437
rect 15933 2397 15945 2431
rect 15979 2428 15991 2431
rect 16672 2431 16730 2437
rect 16672 2428 16684 2431
rect 15979 2400 16684 2428
rect 15979 2397 15991 2400
rect 15933 2391 15991 2397
rect 16672 2397 16684 2400
rect 16718 2397 16730 2431
rect 16672 2391 16730 2397
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2428 17003 2431
rect 18325 2431 18383 2437
rect 16991 2400 18276 2428
rect 16991 2397 17003 2400
rect 16945 2391 17003 2397
rect 11072 2332 11652 2360
rect 3510 2292 3516 2304
rect 3252 2264 3516 2292
rect 3510 2252 3516 2264
rect 3568 2292 3574 2304
rect 5350 2292 5356 2304
rect 3568 2264 5356 2292
rect 3568 2252 3574 2264
rect 5350 2252 5356 2264
rect 5408 2252 5414 2304
rect 5445 2295 5503 2301
rect 5445 2261 5457 2295
rect 5491 2292 5503 2295
rect 11072 2292 11100 2332
rect 5491 2264 11100 2292
rect 11624 2292 11652 2332
rect 12158 2292 12164 2304
rect 11624 2264 12164 2292
rect 5491 2261 5503 2264
rect 5445 2255 5503 2261
rect 12158 2252 12164 2264
rect 12216 2252 12222 2304
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 16482 2292 16488 2304
rect 13596 2264 16488 2292
rect 13596 2252 13602 2264
rect 16482 2252 16488 2264
rect 16540 2252 16546 2304
rect 18248 2292 18276 2400
rect 18325 2397 18337 2431
rect 18371 2428 18383 2431
rect 18880 2428 18892 2449
rect 18371 2415 18892 2428
rect 18926 2415 18938 2449
rect 18371 2409 18938 2415
rect 18371 2400 18920 2409
rect 18371 2397 18383 2400
rect 18325 2391 18383 2397
rect 19150 2388 19156 2440
rect 19208 2388 19214 2440
rect 20640 2360 20668 2459
rect 20898 2456 20904 2508
rect 20956 2496 20962 2508
rect 21269 2499 21327 2505
rect 21269 2496 21281 2499
rect 20956 2468 21281 2496
rect 20956 2456 20962 2468
rect 21269 2465 21281 2468
rect 21315 2465 21327 2499
rect 21269 2459 21327 2465
rect 22738 2456 22744 2508
rect 22796 2496 22802 2508
rect 23569 2499 23627 2505
rect 23569 2496 23581 2499
rect 22796 2468 23581 2496
rect 22796 2456 22802 2468
rect 23569 2465 23581 2468
rect 23615 2496 23627 2499
rect 24026 2496 24032 2508
rect 23615 2468 24032 2496
rect 23615 2465 23627 2468
rect 23569 2459 23627 2465
rect 24026 2456 24032 2468
rect 24084 2496 24090 2508
rect 24121 2499 24179 2505
rect 24121 2496 24133 2499
rect 24084 2468 24133 2496
rect 24084 2456 24090 2468
rect 24121 2465 24133 2468
rect 24167 2465 24179 2499
rect 24228 2496 24256 2592
rect 27430 2564 27436 2576
rect 26252 2536 27436 2564
rect 26252 2508 26280 2536
rect 24857 2499 24915 2505
rect 24228 2468 24660 2496
rect 24121 2459 24179 2465
rect 20809 2431 20867 2437
rect 20809 2397 20821 2431
rect 20855 2428 20867 2431
rect 21450 2428 21456 2440
rect 20855 2400 21456 2428
rect 20855 2397 20867 2400
rect 20809 2391 20867 2397
rect 21450 2388 21456 2400
rect 21508 2388 21514 2440
rect 21732 2433 21790 2439
rect 21732 2399 21744 2433
rect 21778 2428 21790 2433
rect 21818 2428 21824 2440
rect 21778 2400 21824 2428
rect 21778 2399 21790 2400
rect 21732 2393 21790 2399
rect 21818 2388 21824 2400
rect 21876 2388 21882 2440
rect 22005 2431 22063 2437
rect 22005 2397 22017 2431
rect 22051 2428 22063 2431
rect 22830 2428 22836 2440
rect 22051 2400 22836 2428
rect 22051 2397 22063 2400
rect 22005 2391 22063 2397
rect 22830 2388 22836 2400
rect 22888 2388 22894 2440
rect 22922 2388 22928 2440
rect 22980 2428 22986 2440
rect 24394 2428 24400 2440
rect 22980 2400 24400 2428
rect 22980 2388 22986 2400
rect 24394 2388 24400 2400
rect 24452 2437 24458 2440
rect 24632 2439 24660 2468
rect 24857 2465 24869 2499
rect 24903 2496 24915 2499
rect 25222 2496 25228 2508
rect 24903 2468 25228 2496
rect 24903 2465 24915 2468
rect 24857 2459 24915 2465
rect 25222 2456 25228 2468
rect 25280 2456 25286 2508
rect 26234 2456 26240 2508
rect 26292 2456 26298 2508
rect 26712 2505 26740 2536
rect 27430 2524 27436 2536
rect 27488 2524 27494 2576
rect 27540 2536 28120 2564
rect 26605 2499 26663 2505
rect 26605 2465 26617 2499
rect 26651 2465 26663 2499
rect 26605 2459 26663 2465
rect 26697 2499 26755 2505
rect 26697 2465 26709 2499
rect 26743 2465 26755 2499
rect 26697 2459 26755 2465
rect 24452 2431 24506 2437
rect 24452 2397 24460 2431
rect 24494 2397 24506 2431
rect 24452 2391 24506 2397
rect 24617 2433 24675 2439
rect 24617 2399 24629 2433
rect 24663 2399 24675 2433
rect 24617 2393 24675 2399
rect 24452 2388 24458 2391
rect 24946 2388 24952 2440
rect 25004 2428 25010 2440
rect 26050 2428 26056 2440
rect 25004 2400 26056 2428
rect 25004 2388 25010 2400
rect 26050 2388 26056 2400
rect 26108 2388 26114 2440
rect 26326 2388 26332 2440
rect 26384 2428 26390 2440
rect 26620 2428 26648 2459
rect 27246 2456 27252 2508
rect 27304 2496 27310 2508
rect 27341 2499 27399 2505
rect 27341 2496 27353 2499
rect 27304 2468 27353 2496
rect 27304 2456 27310 2468
rect 27341 2465 27353 2468
rect 27387 2496 27399 2499
rect 27387 2468 27476 2496
rect 27387 2465 27399 2468
rect 27341 2459 27399 2465
rect 27448 2440 27476 2468
rect 26384 2400 26648 2428
rect 26384 2388 26390 2400
rect 21082 2360 21088 2372
rect 20640 2332 21088 2360
rect 21082 2320 21088 2332
rect 21140 2320 21146 2372
rect 23658 2360 23664 2372
rect 22664 2332 23664 2360
rect 20622 2292 20628 2304
rect 18248 2264 20628 2292
rect 20622 2252 20628 2264
rect 20680 2252 20686 2304
rect 20806 2252 20812 2304
rect 20864 2292 20870 2304
rect 22664 2292 22692 2332
rect 23658 2320 23664 2332
rect 23716 2320 23722 2372
rect 26421 2363 26479 2369
rect 26421 2360 26433 2363
rect 25516 2332 26433 2360
rect 20864 2264 22692 2292
rect 23293 2295 23351 2301
rect 20864 2252 20870 2264
rect 23293 2261 23305 2295
rect 23339 2292 23351 2295
rect 23934 2292 23940 2304
rect 23339 2264 23940 2292
rect 23339 2261 23351 2264
rect 23293 2255 23351 2261
rect 23934 2252 23940 2264
rect 23992 2252 23998 2304
rect 24578 2252 24584 2304
rect 24636 2292 24642 2304
rect 25516 2292 25544 2332
rect 26421 2329 26433 2332
rect 26467 2329 26479 2363
rect 26620 2360 26648 2400
rect 26786 2388 26792 2440
rect 26844 2428 26850 2440
rect 26881 2431 26939 2437
rect 26881 2428 26893 2431
rect 26844 2400 26893 2428
rect 26844 2388 26850 2400
rect 26881 2397 26893 2400
rect 26927 2397 26939 2431
rect 26881 2391 26939 2397
rect 27430 2388 27436 2440
rect 27488 2388 27494 2440
rect 27540 2360 27568 2536
rect 27982 2456 27988 2508
rect 28040 2456 28046 2508
rect 28092 2496 28120 2536
rect 28092 2468 28580 2496
rect 27614 2388 27620 2440
rect 27672 2428 27678 2440
rect 28448 2431 28506 2437
rect 28448 2428 28460 2431
rect 27672 2400 28460 2428
rect 27672 2388 27678 2400
rect 28448 2397 28460 2400
rect 28494 2397 28506 2431
rect 28552 2428 28580 2468
rect 28718 2456 28724 2508
rect 28776 2456 28782 2508
rect 29086 2428 29092 2440
rect 28552 2400 29092 2428
rect 28448 2391 28506 2397
rect 29086 2388 29092 2400
rect 29144 2428 29150 2440
rect 29454 2428 29460 2440
rect 29144 2400 29460 2428
rect 29144 2388 29150 2400
rect 29454 2388 29460 2400
rect 29512 2388 29518 2440
rect 26620 2332 27568 2360
rect 26421 2323 26479 2329
rect 24636 2264 25544 2292
rect 24636 2252 24642 2264
rect 25590 2252 25596 2304
rect 25648 2292 25654 2304
rect 25961 2295 26019 2301
rect 25961 2292 25973 2295
rect 25648 2264 25973 2292
rect 25648 2252 25654 2264
rect 25961 2261 25973 2264
rect 26007 2261 26019 2295
rect 25961 2255 26019 2261
rect 26050 2252 26056 2304
rect 26108 2292 26114 2304
rect 29362 2292 29368 2304
rect 26108 2264 29368 2292
rect 26108 2252 26114 2264
rect 29362 2252 29368 2264
rect 29420 2252 29426 2304
rect 552 2202 30912 2224
rect 552 2150 4193 2202
rect 4245 2150 4257 2202
rect 4309 2150 4321 2202
rect 4373 2150 4385 2202
rect 4437 2150 4449 2202
rect 4501 2150 11783 2202
rect 11835 2150 11847 2202
rect 11899 2150 11911 2202
rect 11963 2150 11975 2202
rect 12027 2150 12039 2202
rect 12091 2150 19373 2202
rect 19425 2150 19437 2202
rect 19489 2150 19501 2202
rect 19553 2150 19565 2202
rect 19617 2150 19629 2202
rect 19681 2150 26963 2202
rect 27015 2150 27027 2202
rect 27079 2150 27091 2202
rect 27143 2150 27155 2202
rect 27207 2150 27219 2202
rect 27271 2150 30912 2202
rect 552 2128 30912 2150
rect 1670 2048 1676 2100
rect 1728 2088 1734 2100
rect 3237 2091 3295 2097
rect 1728 2060 2774 2088
rect 1728 2048 1734 2060
rect 1443 1955 1501 1961
rect 1443 1921 1455 1955
rect 1489 1952 1501 1955
rect 2314 1952 2320 1964
rect 1489 1924 2320 1952
rect 1489 1921 1501 1924
rect 1443 1915 1501 1921
rect 2314 1912 2320 1924
rect 2372 1912 2378 1964
rect 2746 1952 2774 2060
rect 3237 2057 3249 2091
rect 3283 2088 3295 2091
rect 3878 2088 3884 2100
rect 3283 2060 3884 2088
rect 3283 2057 3295 2060
rect 3237 2051 3295 2057
rect 3878 2048 3884 2060
rect 3936 2048 3942 2100
rect 3970 2048 3976 2100
rect 4028 2088 4034 2100
rect 9858 2088 9864 2100
rect 4028 2060 9864 2088
rect 4028 2048 4034 2060
rect 9858 2048 9864 2060
rect 9916 2048 9922 2100
rect 11974 2048 11980 2100
rect 12032 2088 12038 2100
rect 13538 2088 13544 2100
rect 12032 2060 13544 2088
rect 12032 2048 12038 2060
rect 13538 2048 13544 2060
rect 13596 2048 13602 2100
rect 13633 2091 13691 2097
rect 13633 2057 13645 2091
rect 13679 2088 13691 2091
rect 14826 2088 14832 2100
rect 13679 2060 14832 2088
rect 13679 2057 13691 2060
rect 13633 2051 13691 2057
rect 14826 2048 14832 2060
rect 14884 2048 14890 2100
rect 17034 2048 17040 2100
rect 17092 2088 17098 2100
rect 18325 2091 18383 2097
rect 18325 2088 18337 2091
rect 17092 2060 18337 2088
rect 17092 2048 17098 2060
rect 18325 2057 18337 2060
rect 18371 2057 18383 2091
rect 18325 2051 18383 2057
rect 19150 2048 19156 2100
rect 19208 2088 19214 2100
rect 23109 2091 23167 2097
rect 23109 2088 23121 2091
rect 19208 2060 23121 2088
rect 19208 2048 19214 2060
rect 23109 2057 23121 2060
rect 23155 2057 23167 2091
rect 25869 2091 25927 2097
rect 25869 2088 25881 2091
rect 23109 2051 23167 2057
rect 23216 2060 25881 2088
rect 11238 2020 11244 2032
rect 10428 1992 11244 2020
rect 3878 1961 3884 1964
rect 3840 1955 3884 1961
rect 2746 1924 3648 1952
rect 934 1844 940 1896
rect 992 1884 998 1896
rect 1578 1884 1584 1896
rect 992 1856 1584 1884
rect 992 1844 998 1856
rect 1578 1844 1584 1856
rect 1636 1844 1642 1896
rect 1673 1887 1731 1893
rect 1673 1853 1685 1887
rect 1719 1884 1731 1887
rect 2590 1884 2596 1896
rect 1719 1856 2596 1884
rect 1719 1853 1731 1856
rect 1673 1847 1731 1853
rect 2590 1844 2596 1856
rect 2648 1844 2654 1896
rect 3421 1887 3479 1893
rect 3421 1853 3433 1887
rect 3467 1853 3479 1887
rect 3421 1847 3479 1853
rect 3050 1776 3056 1828
rect 3108 1776 3114 1828
rect 1394 1708 1400 1760
rect 1452 1757 1458 1760
rect 1452 1748 1461 1757
rect 1452 1720 1497 1748
rect 1452 1711 1461 1720
rect 1452 1708 1458 1711
rect 2038 1708 2044 1760
rect 2096 1748 2102 1760
rect 3436 1748 3464 1847
rect 3510 1844 3516 1896
rect 3568 1844 3574 1896
rect 3620 1884 3648 1924
rect 3840 1921 3852 1955
rect 3840 1915 3884 1921
rect 3878 1912 3884 1915
rect 3936 1912 3942 1964
rect 3976 1953 4034 1959
rect 3976 1919 3988 1953
rect 4022 1952 4034 1953
rect 4062 1952 4068 1964
rect 4022 1924 4068 1952
rect 4022 1919 4034 1924
rect 3976 1913 4034 1919
rect 4062 1912 4068 1924
rect 4120 1912 4126 1964
rect 4249 1955 4307 1961
rect 4249 1921 4261 1955
rect 4295 1952 4307 1955
rect 5442 1952 5448 1964
rect 4295 1924 5448 1952
rect 4295 1921 4307 1924
rect 4249 1915 4307 1921
rect 5442 1912 5448 1924
rect 5500 1912 5506 1964
rect 6089 1955 6147 1961
rect 6089 1921 6101 1955
rect 6135 1952 6147 1955
rect 6454 1952 6460 1964
rect 6135 1924 6460 1952
rect 6135 1921 6147 1924
rect 6089 1915 6147 1921
rect 6454 1912 6460 1924
rect 6512 1912 6518 1964
rect 6552 1955 6610 1961
rect 6552 1921 6564 1955
rect 6598 1921 6610 1955
rect 6552 1915 6610 1921
rect 3620 1856 5396 1884
rect 4982 1776 4988 1828
rect 5040 1776 5046 1828
rect 5000 1748 5028 1776
rect 5368 1757 5396 1856
rect 5994 1844 6000 1896
rect 6052 1884 6058 1896
rect 6567 1884 6595 1915
rect 6638 1912 6644 1964
rect 6696 1912 6702 1964
rect 6822 1912 6828 1964
rect 6880 1912 6886 1964
rect 8205 1955 8263 1961
rect 8205 1921 8217 1955
rect 8251 1952 8263 1955
rect 9496 1955 9554 1961
rect 9496 1952 9508 1955
rect 8251 1924 9508 1952
rect 8251 1921 8263 1924
rect 8205 1915 8263 1921
rect 9496 1921 9508 1924
rect 9542 1921 9554 1955
rect 9496 1915 9554 1921
rect 9674 1912 9680 1964
rect 9732 1952 9738 1964
rect 9769 1955 9827 1961
rect 9769 1952 9781 1955
rect 9732 1924 9781 1952
rect 9732 1912 9738 1924
rect 9769 1921 9781 1924
rect 9815 1921 9827 1955
rect 9769 1915 9827 1921
rect 9858 1912 9864 1964
rect 9916 1952 9922 1964
rect 10428 1952 10456 1992
rect 11238 1980 11244 1992
rect 11296 1980 11302 2032
rect 23014 1980 23020 2032
rect 23072 2020 23078 2032
rect 23216 2020 23244 2060
rect 25869 2057 25881 2060
rect 25915 2057 25927 2091
rect 25869 2051 25927 2057
rect 28166 2048 28172 2100
rect 28224 2048 28230 2100
rect 29178 2048 29184 2100
rect 29236 2048 29242 2100
rect 29457 2091 29515 2097
rect 29457 2057 29469 2091
rect 29503 2088 29515 2091
rect 29638 2088 29644 2100
rect 29503 2060 29644 2088
rect 29503 2057 29515 2060
rect 29457 2051 29515 2057
rect 29638 2048 29644 2060
rect 29696 2048 29702 2100
rect 23750 2020 23756 2032
rect 23072 1992 23244 2020
rect 23308 1992 23756 2020
rect 23072 1980 23078 1992
rect 9916 1924 10456 1952
rect 11149 1955 11207 1961
rect 9916 1912 9922 1924
rect 11149 1921 11161 1955
rect 11195 1952 11207 1955
rect 11704 1955 11762 1961
rect 11704 1952 11716 1955
rect 11195 1924 11716 1952
rect 11195 1921 11207 1924
rect 11149 1915 11207 1921
rect 11704 1921 11716 1924
rect 11750 1921 11762 1955
rect 11704 1915 11762 1921
rect 13357 1955 13415 1961
rect 13357 1921 13369 1955
rect 13403 1952 13415 1955
rect 14372 1955 14430 1961
rect 14372 1952 14384 1955
rect 13403 1924 14384 1952
rect 13403 1921 13415 1924
rect 13357 1915 13415 1921
rect 14372 1921 14384 1924
rect 14418 1921 14430 1955
rect 14372 1915 14430 1921
rect 16114 1912 16120 1964
rect 16172 1912 16178 1964
rect 18233 1955 18291 1961
rect 16224 1943 16620 1952
rect 16224 1937 16638 1943
rect 16224 1924 16592 1937
rect 6052 1856 6595 1884
rect 6656 1884 6684 1912
rect 8389 1887 8447 1893
rect 6656 1856 7512 1884
rect 6052 1844 6058 1856
rect 7484 1816 7512 1856
rect 8389 1853 8401 1887
rect 8435 1884 8447 1887
rect 8754 1884 8760 1896
rect 8435 1856 8760 1884
rect 8435 1853 8447 1856
rect 8389 1847 8447 1853
rect 8754 1844 8760 1856
rect 8812 1844 8818 1896
rect 8846 1844 8852 1896
rect 8904 1884 8910 1896
rect 9033 1887 9091 1893
rect 9033 1884 9045 1887
rect 8904 1856 9045 1884
rect 8904 1844 8910 1856
rect 9033 1853 9045 1856
rect 9079 1884 9091 1887
rect 9306 1884 9312 1896
rect 9079 1856 9312 1884
rect 9079 1853 9091 1856
rect 9033 1847 9091 1853
rect 9306 1844 9312 1856
rect 9364 1844 9370 1896
rect 11241 1887 11299 1893
rect 11241 1853 11253 1887
rect 11287 1884 11299 1887
rect 11330 1884 11336 1896
rect 11287 1856 11336 1884
rect 11287 1853 11299 1856
rect 11241 1847 11299 1853
rect 11330 1844 11336 1856
rect 11388 1884 11394 1896
rect 11606 1884 11612 1896
rect 11388 1856 11612 1884
rect 11388 1844 11394 1856
rect 11606 1844 11612 1856
rect 11664 1844 11670 1896
rect 11974 1844 11980 1896
rect 12032 1844 12038 1896
rect 12434 1844 12440 1896
rect 12492 1884 12498 1896
rect 13817 1887 13875 1893
rect 13817 1884 13829 1887
rect 12492 1856 13829 1884
rect 12492 1844 12498 1856
rect 13817 1853 13829 1856
rect 13863 1853 13875 1887
rect 13817 1847 13875 1853
rect 13906 1844 13912 1896
rect 13964 1844 13970 1896
rect 14645 1887 14703 1893
rect 14645 1884 14657 1887
rect 14016 1856 14657 1884
rect 8665 1819 8723 1825
rect 8665 1816 8677 1819
rect 7484 1788 8677 1816
rect 8665 1785 8677 1788
rect 8711 1785 8723 1819
rect 8665 1779 8723 1785
rect 13538 1776 13544 1828
rect 13596 1816 13602 1828
rect 14016 1816 14044 1856
rect 14645 1853 14657 1856
rect 14691 1853 14703 1887
rect 14645 1847 14703 1853
rect 16025 1887 16083 1893
rect 16025 1853 16037 1887
rect 16071 1884 16083 1887
rect 16224 1884 16252 1924
rect 16580 1903 16592 1924
rect 16626 1903 16638 1937
rect 18233 1921 18245 1955
rect 18279 1952 18291 1955
rect 19156 1955 19214 1961
rect 19156 1952 19168 1955
rect 18279 1924 19168 1952
rect 18279 1921 18291 1924
rect 18233 1915 18291 1921
rect 19156 1921 19168 1924
rect 19202 1921 19214 1955
rect 19156 1915 19214 1921
rect 19242 1912 19248 1964
rect 19300 1952 19306 1964
rect 20714 1952 20720 1964
rect 19300 1924 20720 1952
rect 19300 1912 19306 1924
rect 20714 1912 20720 1924
rect 20772 1912 20778 1964
rect 20809 1955 20867 1961
rect 20809 1921 20821 1955
rect 20855 1952 20867 1955
rect 21364 1955 21422 1961
rect 21364 1952 21376 1955
rect 20855 1924 21376 1952
rect 20855 1921 20867 1924
rect 20809 1915 20867 1921
rect 21364 1921 21376 1924
rect 21410 1921 21422 1955
rect 21364 1915 21422 1921
rect 21450 1912 21456 1964
rect 21508 1912 21514 1964
rect 21637 1955 21695 1961
rect 21637 1921 21649 1955
rect 21683 1952 21695 1955
rect 23106 1952 23112 1964
rect 21683 1924 23112 1952
rect 21683 1921 21695 1924
rect 21637 1915 21695 1921
rect 23106 1912 23112 1924
rect 23164 1912 23170 1964
rect 23308 1952 23336 1992
rect 23750 1980 23756 1992
rect 23808 1980 23814 2032
rect 23658 1952 23664 1964
rect 23216 1924 23336 1952
rect 23400 1924 23664 1952
rect 16580 1897 16638 1903
rect 16071 1856 16252 1884
rect 16071 1853 16083 1856
rect 16025 1847 16083 1853
rect 16850 1844 16856 1896
rect 16908 1844 16914 1896
rect 18509 1887 18567 1893
rect 18509 1853 18521 1887
rect 18555 1853 18567 1887
rect 18509 1847 18567 1853
rect 13596 1788 14044 1816
rect 13596 1776 13602 1788
rect 2096 1720 5028 1748
rect 5353 1751 5411 1757
rect 2096 1708 2102 1720
rect 5353 1717 5365 1751
rect 5399 1717 5411 1751
rect 5353 1711 5411 1717
rect 5994 1708 6000 1760
rect 6052 1708 6058 1760
rect 6555 1751 6613 1757
rect 6555 1717 6567 1751
rect 6601 1748 6613 1751
rect 6914 1748 6920 1760
rect 6601 1720 6920 1748
rect 6601 1717 6613 1720
rect 6555 1711 6613 1717
rect 6914 1708 6920 1720
rect 6972 1708 6978 1760
rect 9030 1708 9036 1760
rect 9088 1748 9094 1760
rect 9499 1751 9557 1757
rect 9499 1748 9511 1751
rect 9088 1720 9511 1748
rect 9088 1708 9094 1720
rect 9499 1717 9511 1720
rect 9545 1717 9557 1751
rect 9499 1711 9557 1717
rect 9674 1708 9680 1760
rect 9732 1748 9738 1760
rect 10410 1748 10416 1760
rect 9732 1720 10416 1748
rect 9732 1708 9738 1720
rect 10410 1708 10416 1720
rect 10468 1708 10474 1760
rect 11698 1708 11704 1760
rect 11756 1757 11762 1760
rect 11756 1748 11765 1757
rect 11756 1720 11801 1748
rect 11756 1711 11765 1720
rect 11756 1708 11762 1711
rect 14182 1708 14188 1760
rect 14240 1748 14246 1760
rect 14375 1751 14433 1757
rect 14375 1748 14387 1751
rect 14240 1720 14387 1748
rect 14240 1708 14246 1720
rect 14375 1717 14387 1720
rect 14421 1717 14433 1751
rect 14375 1711 14433 1717
rect 16574 1708 16580 1760
rect 16632 1757 16638 1760
rect 16632 1748 16641 1757
rect 18524 1748 18552 1847
rect 18690 1844 18696 1896
rect 18748 1844 18754 1896
rect 18782 1844 18788 1896
rect 18840 1884 18846 1896
rect 19020 1887 19078 1893
rect 19020 1884 19032 1887
rect 18840 1856 19032 1884
rect 18840 1844 18846 1856
rect 19020 1853 19032 1856
rect 19066 1853 19078 1887
rect 19020 1847 19078 1853
rect 19426 1844 19432 1896
rect 19484 1844 19490 1896
rect 20898 1844 20904 1896
rect 20956 1844 20962 1896
rect 21228 1887 21286 1893
rect 21228 1853 21240 1887
rect 21274 1884 21286 1887
rect 21468 1884 21496 1912
rect 23216 1884 23244 1924
rect 21274 1856 21496 1884
rect 22664 1856 23244 1884
rect 23293 1887 23351 1893
rect 21274 1853 21286 1856
rect 21228 1847 21286 1853
rect 22664 1828 22692 1856
rect 23293 1853 23305 1887
rect 23339 1884 23351 1887
rect 23400 1884 23428 1924
rect 23658 1912 23664 1924
rect 23716 1912 23722 1964
rect 23339 1856 23428 1884
rect 23569 1887 23627 1893
rect 23339 1853 23351 1856
rect 23293 1847 23351 1853
rect 23569 1853 23581 1887
rect 23615 1884 23627 1887
rect 23768 1884 23796 1980
rect 23952 1943 24348 1952
rect 23952 1937 24366 1943
rect 23952 1924 24320 1937
rect 23615 1856 23796 1884
rect 23615 1853 23627 1856
rect 23569 1847 23627 1853
rect 23842 1844 23848 1896
rect 23900 1844 23906 1896
rect 22646 1776 22652 1828
rect 22704 1776 22710 1828
rect 23017 1819 23075 1825
rect 23017 1785 23029 1819
rect 23063 1816 23075 1819
rect 23952 1816 23980 1924
rect 24308 1903 24320 1924
rect 24354 1903 24366 1937
rect 24486 1912 24492 1964
rect 24544 1952 24550 1964
rect 24581 1955 24639 1961
rect 24581 1952 24593 1955
rect 24544 1924 24593 1952
rect 24544 1912 24550 1924
rect 24581 1921 24593 1924
rect 24627 1921 24639 1955
rect 26329 1955 26387 1961
rect 24581 1915 24639 1921
rect 25792 1950 26096 1952
rect 26329 1950 26341 1955
rect 25792 1924 26341 1950
rect 24308 1897 24366 1903
rect 25792 1896 25820 1924
rect 26068 1922 26341 1924
rect 26329 1921 26341 1922
rect 26375 1921 26387 1955
rect 26329 1915 26387 1921
rect 26835 1955 26893 1961
rect 26835 1921 26847 1955
rect 26881 1952 26893 1955
rect 27706 1952 27712 1964
rect 26881 1924 27712 1952
rect 26881 1921 26893 1924
rect 26835 1915 26893 1921
rect 27706 1912 27712 1924
rect 27764 1912 27770 1964
rect 28810 1912 28816 1964
rect 28868 1952 28874 1964
rect 28868 1924 29316 1952
rect 28868 1912 28874 1924
rect 25774 1844 25780 1896
rect 25832 1844 25838 1896
rect 26229 1887 26287 1893
rect 26229 1884 26241 1887
rect 25884 1856 26241 1884
rect 23063 1788 23980 1816
rect 23063 1785 23075 1788
rect 23017 1779 23075 1785
rect 21910 1748 21916 1760
rect 16632 1720 16677 1748
rect 18524 1720 21916 1748
rect 16632 1711 16641 1720
rect 16632 1708 16638 1711
rect 21910 1708 21916 1720
rect 21968 1708 21974 1760
rect 23106 1708 23112 1760
rect 23164 1748 23170 1760
rect 23385 1751 23443 1757
rect 23385 1748 23397 1751
rect 23164 1720 23397 1748
rect 23164 1708 23170 1720
rect 23385 1717 23397 1720
rect 23431 1717 23443 1751
rect 23385 1711 23443 1717
rect 24118 1708 24124 1760
rect 24176 1748 24182 1760
rect 24311 1751 24369 1757
rect 24311 1748 24323 1751
rect 24176 1720 24323 1748
rect 24176 1708 24182 1720
rect 24311 1717 24323 1720
rect 24357 1717 24369 1751
rect 24311 1711 24369 1717
rect 24486 1708 24492 1760
rect 24544 1748 24550 1760
rect 25884 1748 25912 1856
rect 26229 1853 26241 1856
rect 26275 1853 26287 1887
rect 26229 1847 26287 1853
rect 26252 1816 26280 1847
rect 26418 1844 26424 1896
rect 26476 1884 26482 1896
rect 26656 1887 26714 1893
rect 26656 1884 26668 1887
rect 26476 1856 26668 1884
rect 26476 1844 26482 1856
rect 26656 1853 26668 1856
rect 26702 1853 26714 1887
rect 26656 1847 26714 1853
rect 26970 1844 26976 1896
rect 27028 1884 27034 1896
rect 27065 1887 27123 1893
rect 27065 1884 27077 1887
rect 27028 1856 27077 1884
rect 27028 1844 27034 1856
rect 27065 1853 27077 1856
rect 27111 1853 27123 1887
rect 28537 1887 28595 1893
rect 28537 1884 28549 1887
rect 27065 1847 27123 1853
rect 27724 1856 28549 1884
rect 26326 1816 26332 1828
rect 26252 1788 26332 1816
rect 26326 1776 26332 1788
rect 26384 1776 26390 1828
rect 24544 1720 25912 1748
rect 24544 1708 24550 1720
rect 26050 1708 26056 1760
rect 26108 1708 26114 1760
rect 26418 1708 26424 1760
rect 26476 1748 26482 1760
rect 27724 1748 27752 1856
rect 28537 1853 28549 1856
rect 28583 1884 28595 1887
rect 28828 1884 28856 1912
rect 28583 1856 28856 1884
rect 28583 1853 28595 1856
rect 28537 1847 28595 1853
rect 28994 1844 29000 1896
rect 29052 1893 29058 1896
rect 29288 1893 29316 1924
rect 29052 1884 29064 1893
rect 29273 1887 29331 1893
rect 29052 1856 29097 1884
rect 29052 1847 29064 1856
rect 29273 1853 29285 1887
rect 29319 1853 29331 1887
rect 29273 1847 29331 1853
rect 29052 1844 29058 1847
rect 26476 1720 27752 1748
rect 26476 1708 26482 1720
rect 28718 1708 28724 1760
rect 28776 1708 28782 1760
rect 552 1658 31072 1680
rect 552 1606 7988 1658
rect 8040 1606 8052 1658
rect 8104 1606 8116 1658
rect 8168 1606 8180 1658
rect 8232 1606 8244 1658
rect 8296 1606 15578 1658
rect 15630 1606 15642 1658
rect 15694 1606 15706 1658
rect 15758 1606 15770 1658
rect 15822 1606 15834 1658
rect 15886 1606 23168 1658
rect 23220 1606 23232 1658
rect 23284 1606 23296 1658
rect 23348 1606 23360 1658
rect 23412 1606 23424 1658
rect 23476 1606 30758 1658
rect 30810 1606 30822 1658
rect 30874 1606 30886 1658
rect 30938 1606 30950 1658
rect 31002 1606 31014 1658
rect 31066 1606 31072 1658
rect 552 1584 31072 1606
rect 845 1547 903 1553
rect 845 1513 857 1547
rect 891 1544 903 1547
rect 1118 1544 1124 1556
rect 891 1516 1124 1544
rect 891 1513 903 1516
rect 845 1507 903 1513
rect 1118 1504 1124 1516
rect 1176 1504 1182 1556
rect 1210 1504 1216 1556
rect 1268 1544 1274 1556
rect 1268 1516 2452 1544
rect 1268 1504 1274 1516
rect 2314 1476 2320 1488
rect 952 1448 2320 1476
rect 952 1272 980 1448
rect 2314 1436 2320 1448
rect 2372 1436 2378 1488
rect 2424 1476 2452 1516
rect 2590 1504 2596 1556
rect 2648 1544 2654 1556
rect 2648 1516 3096 1544
rect 2648 1504 2654 1516
rect 3068 1476 3096 1516
rect 3142 1504 3148 1556
rect 3200 1504 3206 1556
rect 4706 1544 4712 1556
rect 3252 1516 4712 1544
rect 3252 1476 3280 1516
rect 4706 1504 4712 1516
rect 4764 1504 4770 1556
rect 5350 1504 5356 1556
rect 5408 1544 5414 1556
rect 5408 1516 6592 1544
rect 5408 1504 5414 1516
rect 2424 1448 2912 1476
rect 3068 1448 3280 1476
rect 1026 1368 1032 1420
rect 1084 1368 1090 1420
rect 1305 1411 1363 1417
rect 1305 1377 1317 1411
rect 1351 1408 1363 1411
rect 2038 1408 2044 1420
rect 1351 1380 2044 1408
rect 1351 1377 1363 1380
rect 1305 1371 1363 1377
rect 2038 1368 2044 1380
rect 2096 1368 2102 1420
rect 2884 1417 2912 1448
rect 3326 1436 3332 1488
rect 3384 1436 3390 1488
rect 5810 1436 5816 1488
rect 5868 1476 5874 1488
rect 5905 1479 5963 1485
rect 5905 1476 5917 1479
rect 5868 1448 5917 1476
rect 5868 1436 5874 1448
rect 5905 1445 5917 1448
rect 5951 1445 5963 1479
rect 6270 1476 6276 1488
rect 5905 1439 5963 1445
rect 6012 1448 6276 1476
rect 2593 1411 2651 1417
rect 2593 1408 2605 1411
rect 2240 1380 2605 1408
rect 1044 1340 1072 1368
rect 2240 1340 2268 1380
rect 2593 1377 2605 1380
rect 2639 1377 2651 1411
rect 2593 1371 2651 1377
rect 2869 1411 2927 1417
rect 2869 1377 2881 1411
rect 2915 1377 2927 1411
rect 2869 1371 2927 1377
rect 3053 1411 3111 1417
rect 3053 1377 3065 1411
rect 3099 1408 3111 1411
rect 3344 1408 3372 1436
rect 5629 1411 5687 1417
rect 3099 1380 5120 1408
rect 3099 1377 3111 1380
rect 3053 1371 3111 1377
rect 1044 1312 2268 1340
rect 2317 1343 2375 1349
rect 2317 1309 2329 1343
rect 2363 1340 2375 1343
rect 2363 1312 3464 1340
rect 2363 1309 2375 1312
rect 2317 1303 2375 1309
rect 1121 1275 1179 1281
rect 1121 1272 1133 1275
rect 952 1244 1133 1272
rect 1121 1241 1133 1244
rect 1167 1241 1179 1275
rect 1121 1235 1179 1241
rect 1949 1275 2007 1281
rect 1949 1241 1961 1275
rect 1995 1272 2007 1275
rect 3234 1272 3240 1284
rect 1995 1244 3240 1272
rect 1995 1241 2007 1244
rect 1949 1235 2007 1241
rect 3234 1232 3240 1244
rect 3292 1232 3298 1284
rect 2222 1164 2228 1216
rect 2280 1204 2286 1216
rect 2409 1207 2467 1213
rect 2409 1204 2421 1207
rect 2280 1176 2421 1204
rect 2280 1164 2286 1176
rect 2409 1173 2421 1176
rect 2455 1173 2467 1207
rect 2409 1167 2467 1173
rect 2682 1164 2688 1216
rect 2740 1164 2746 1216
rect 3436 1204 3464 1312
rect 3510 1300 3516 1352
rect 3568 1300 3574 1352
rect 3878 1349 3884 1352
rect 3840 1343 3884 1349
rect 3840 1309 3852 1343
rect 3840 1303 3884 1309
rect 3878 1300 3884 1303
rect 3936 1300 3942 1352
rect 3970 1300 3976 1352
rect 4028 1340 4034 1352
rect 4028 1312 4073 1340
rect 4028 1300 4034 1312
rect 4246 1300 4252 1352
rect 4304 1300 4310 1352
rect 5092 1340 5120 1380
rect 5629 1377 5641 1411
rect 5675 1408 5687 1411
rect 6012 1408 6040 1448
rect 6270 1436 6276 1448
rect 6328 1436 6334 1488
rect 5675 1380 6040 1408
rect 5675 1377 5687 1380
rect 5629 1371 5687 1377
rect 6454 1368 6460 1420
rect 6512 1368 6518 1420
rect 6564 1408 6592 1516
rect 6914 1504 6920 1556
rect 6972 1553 6978 1556
rect 6972 1544 6981 1553
rect 8481 1547 8539 1553
rect 6972 1516 8248 1544
rect 6972 1507 6981 1516
rect 6972 1504 6978 1507
rect 8220 1488 8248 1516
rect 8481 1513 8493 1547
rect 8527 1544 8539 1547
rect 9122 1544 9128 1556
rect 8527 1516 9128 1544
rect 8527 1513 8539 1516
rect 8481 1507 8539 1513
rect 9122 1504 9128 1516
rect 9180 1504 9186 1556
rect 11514 1544 11520 1556
rect 10336 1516 11520 1544
rect 8202 1436 8208 1488
rect 8260 1436 8266 1488
rect 10336 1408 10364 1516
rect 11514 1504 11520 1516
rect 11572 1504 11578 1556
rect 11698 1504 11704 1556
rect 11756 1544 11762 1556
rect 12075 1547 12133 1553
rect 12075 1544 12087 1547
rect 11756 1516 12087 1544
rect 11756 1504 11762 1516
rect 12075 1513 12087 1516
rect 12121 1513 12133 1547
rect 12075 1507 12133 1513
rect 12250 1504 12256 1556
rect 12308 1544 12314 1556
rect 14366 1544 14372 1556
rect 12308 1516 14372 1544
rect 12308 1504 12314 1516
rect 14366 1504 14372 1516
rect 14424 1504 14430 1556
rect 16574 1504 16580 1556
rect 16632 1544 16638 1556
rect 16675 1547 16733 1553
rect 16675 1544 16687 1547
rect 16632 1516 16687 1544
rect 16632 1504 16638 1516
rect 16675 1513 16687 1516
rect 16721 1513 16733 1547
rect 16675 1507 16733 1513
rect 18782 1504 18788 1556
rect 18840 1544 18846 1556
rect 18883 1547 18941 1553
rect 18883 1544 18895 1547
rect 18840 1516 18895 1544
rect 18840 1504 18846 1516
rect 18883 1513 18895 1516
rect 18929 1513 18941 1547
rect 18883 1507 18941 1513
rect 19426 1504 19432 1556
rect 19484 1544 19490 1556
rect 20901 1547 20959 1553
rect 20901 1544 20913 1547
rect 19484 1516 20913 1544
rect 19484 1504 19490 1516
rect 20901 1513 20913 1516
rect 20947 1513 20959 1547
rect 20901 1507 20959 1513
rect 21542 1504 21548 1556
rect 21600 1544 21606 1556
rect 21735 1547 21793 1553
rect 21735 1544 21747 1547
rect 21600 1516 21747 1544
rect 21600 1504 21606 1516
rect 21735 1513 21747 1516
rect 21781 1513 21793 1547
rect 21735 1507 21793 1513
rect 26878 1504 26884 1556
rect 26936 1544 26942 1556
rect 27430 1544 27436 1556
rect 26936 1516 27436 1544
rect 26936 1504 26942 1516
rect 27430 1504 27436 1516
rect 27488 1544 27494 1556
rect 27488 1516 27844 1544
rect 27488 1504 27494 1516
rect 10410 1436 10416 1488
rect 10468 1436 10474 1488
rect 10781 1479 10839 1485
rect 10781 1445 10793 1479
rect 10827 1476 10839 1479
rect 20533 1479 20591 1485
rect 10827 1448 11750 1476
rect 10827 1445 10839 1448
rect 10781 1439 10839 1445
rect 6564 1380 10364 1408
rect 10428 1408 10456 1436
rect 11149 1411 11207 1417
rect 11149 1408 11161 1411
rect 10428 1380 11161 1408
rect 11149 1377 11161 1380
rect 11195 1408 11207 1411
rect 11517 1411 11575 1417
rect 11517 1408 11529 1411
rect 11195 1380 11529 1408
rect 11195 1377 11207 1380
rect 11149 1371 11207 1377
rect 11517 1377 11529 1380
rect 11563 1377 11575 1411
rect 11517 1371 11575 1377
rect 11606 1368 11612 1420
rect 11664 1368 11670 1420
rect 6181 1343 6239 1349
rect 6181 1340 6193 1343
rect 5092 1312 6193 1340
rect 6181 1309 6193 1312
rect 6227 1309 6239 1343
rect 6181 1303 6239 1309
rect 6914 1300 6920 1352
rect 6972 1300 6978 1352
rect 7193 1343 7251 1349
rect 7193 1309 7205 1343
rect 7239 1340 7251 1343
rect 8570 1340 8576 1352
rect 7239 1312 8576 1340
rect 7239 1309 7251 1312
rect 7193 1303 7251 1309
rect 8570 1300 8576 1312
rect 8628 1300 8634 1352
rect 8665 1343 8723 1349
rect 8665 1309 8677 1343
rect 8711 1340 8723 1343
rect 8846 1340 8852 1352
rect 8711 1312 8852 1340
rect 8711 1309 8723 1312
rect 8665 1303 8723 1309
rect 8846 1300 8852 1312
rect 8904 1300 8910 1352
rect 9030 1349 9036 1352
rect 8992 1343 9036 1349
rect 8992 1309 9004 1343
rect 8992 1303 9036 1309
rect 9030 1300 9036 1303
rect 9088 1300 9094 1352
rect 9171 1343 9229 1349
rect 9171 1309 9183 1343
rect 9217 1340 9229 1343
rect 9306 1340 9312 1352
rect 9217 1312 9312 1340
rect 9217 1309 9229 1312
rect 9171 1303 9229 1309
rect 9306 1300 9312 1312
rect 9364 1300 9370 1352
rect 9401 1343 9459 1349
rect 9401 1309 9413 1343
rect 9447 1340 9459 1343
rect 11722 1340 11750 1448
rect 20533 1445 20545 1479
rect 20579 1476 20591 1479
rect 23566 1476 23572 1488
rect 20579 1448 21404 1476
rect 20579 1445 20591 1448
rect 20533 1439 20591 1445
rect 11882 1368 11888 1420
rect 11940 1408 11946 1420
rect 13725 1411 13783 1417
rect 11940 1380 12388 1408
rect 11940 1368 11946 1380
rect 12360 1349 12388 1380
rect 13725 1377 13737 1411
rect 13771 1408 13783 1411
rect 13771 1380 14320 1408
rect 13771 1377 13783 1380
rect 13725 1371 13783 1377
rect 12072 1343 12130 1349
rect 12072 1340 12084 1343
rect 9447 1312 11008 1340
rect 11722 1312 12084 1340
rect 9447 1309 9459 1312
rect 9401 1303 9459 1309
rect 10980 1281 11008 1312
rect 12072 1309 12084 1312
rect 12118 1309 12130 1343
rect 12072 1303 12130 1309
rect 12345 1343 12403 1349
rect 12345 1309 12357 1343
rect 12391 1309 12403 1343
rect 12345 1303 12403 1309
rect 13814 1300 13820 1352
rect 13872 1300 13878 1352
rect 14182 1349 14188 1352
rect 14144 1343 14188 1349
rect 14144 1309 14156 1343
rect 14144 1303 14188 1309
rect 14182 1300 14188 1303
rect 14240 1300 14246 1352
rect 14292 1349 14320 1380
rect 16114 1368 16120 1420
rect 16172 1408 16178 1420
rect 16209 1411 16267 1417
rect 16209 1408 16221 1411
rect 16172 1380 16221 1408
rect 16172 1368 16178 1380
rect 16209 1377 16221 1380
rect 16255 1377 16267 1411
rect 16209 1371 16267 1377
rect 18325 1411 18383 1417
rect 18325 1377 18337 1411
rect 18371 1408 18383 1411
rect 18371 1380 18920 1408
rect 18371 1377 18383 1380
rect 18325 1371 18383 1377
rect 14280 1343 14338 1349
rect 14280 1309 14292 1343
rect 14326 1309 14338 1343
rect 14280 1303 14338 1309
rect 14366 1300 14372 1352
rect 14424 1340 14430 1352
rect 14553 1343 14611 1349
rect 14553 1340 14565 1343
rect 14424 1312 14565 1340
rect 14424 1300 14430 1312
rect 14553 1309 14565 1312
rect 14599 1309 14611 1343
rect 14553 1303 14611 1309
rect 15933 1343 15991 1349
rect 15933 1309 15945 1343
rect 15979 1340 15991 1343
rect 16672 1343 16730 1349
rect 16672 1340 16684 1343
rect 15979 1312 16684 1340
rect 15979 1309 15991 1312
rect 15933 1303 15991 1309
rect 16672 1309 16684 1312
rect 16718 1309 16730 1343
rect 16672 1303 16730 1309
rect 16942 1300 16948 1352
rect 17000 1300 17006 1352
rect 17034 1300 17040 1352
rect 17092 1340 17098 1352
rect 18417 1343 18475 1349
rect 17092 1312 18368 1340
rect 17092 1300 17098 1312
rect 10965 1275 11023 1281
rect 4908 1244 6132 1272
rect 3970 1204 3976 1216
rect 3436 1176 3976 1204
rect 3970 1164 3976 1176
rect 4028 1164 4034 1216
rect 4062 1164 4068 1216
rect 4120 1204 4126 1216
rect 4908 1204 4936 1244
rect 4120 1176 4936 1204
rect 6104 1204 6132 1244
rect 10965 1241 10977 1275
rect 11011 1241 11023 1275
rect 10965 1235 11023 1241
rect 7650 1204 7656 1216
rect 6104 1176 7656 1204
rect 4120 1164 4126 1176
rect 7650 1164 7656 1176
rect 7708 1164 7714 1216
rect 11333 1207 11391 1213
rect 11333 1173 11345 1207
rect 11379 1204 11391 1207
rect 12066 1204 12072 1216
rect 11379 1176 12072 1204
rect 11379 1173 11391 1176
rect 11333 1167 11391 1173
rect 12066 1164 12072 1176
rect 12124 1164 12130 1216
rect 12158 1164 12164 1216
rect 12216 1204 12222 1216
rect 14550 1204 14556 1216
rect 12216 1176 14556 1204
rect 12216 1164 12222 1176
rect 14550 1164 14556 1176
rect 14608 1164 14614 1216
rect 18340 1204 18368 1312
rect 18417 1309 18429 1343
rect 18463 1340 18475 1343
rect 18598 1340 18604 1352
rect 18463 1312 18604 1340
rect 18463 1309 18475 1312
rect 18417 1303 18475 1309
rect 18598 1300 18604 1312
rect 18656 1300 18662 1352
rect 18892 1349 18920 1380
rect 20806 1368 20812 1420
rect 20864 1368 20870 1420
rect 21082 1368 21088 1420
rect 21140 1368 21146 1420
rect 18880 1343 18938 1349
rect 18880 1309 18892 1343
rect 18926 1309 18938 1343
rect 18880 1303 18938 1309
rect 19153 1343 19211 1349
rect 19153 1309 19165 1343
rect 19199 1340 19211 1343
rect 19199 1312 20852 1340
rect 19199 1309 19211 1312
rect 19153 1303 19211 1309
rect 20824 1272 20852 1312
rect 20990 1300 20996 1352
rect 21048 1340 21054 1352
rect 21269 1343 21327 1349
rect 21269 1340 21281 1343
rect 21048 1312 21281 1340
rect 21048 1300 21054 1312
rect 21269 1309 21281 1312
rect 21315 1309 21327 1343
rect 21376 1340 21404 1448
rect 23400 1448 23572 1476
rect 23400 1417 23428 1448
rect 23566 1436 23572 1448
rect 23624 1436 23630 1488
rect 24946 1436 24952 1488
rect 25004 1476 25010 1488
rect 25774 1476 25780 1488
rect 25004 1448 25780 1476
rect 25004 1436 25010 1448
rect 25774 1436 25780 1448
rect 25832 1436 25838 1488
rect 26510 1476 26516 1488
rect 25884 1448 26516 1476
rect 23385 1411 23443 1417
rect 23385 1377 23397 1411
rect 23431 1377 23443 1411
rect 23385 1371 23443 1377
rect 23804 1411 23862 1417
rect 23804 1377 23816 1411
rect 23850 1408 23862 1411
rect 23850 1380 24164 1408
rect 23850 1377 23862 1380
rect 23804 1371 23862 1377
rect 21732 1361 21790 1367
rect 21732 1340 21744 1361
rect 21376 1327 21744 1340
rect 21778 1327 21790 1361
rect 24136 1352 24164 1380
rect 24854 1368 24860 1420
rect 24912 1408 24918 1420
rect 25884 1408 25912 1448
rect 26510 1436 26516 1448
rect 26568 1436 26574 1488
rect 24912 1380 25912 1408
rect 24912 1368 24918 1380
rect 25958 1368 25964 1420
rect 26016 1408 26022 1420
rect 26807 1408 26927 1412
rect 26016 1384 26927 1408
rect 26016 1380 26835 1384
rect 26016 1368 26022 1380
rect 21376 1321 21790 1327
rect 22005 1343 22063 1349
rect 21376 1312 21772 1321
rect 21269 1303 21327 1309
rect 22005 1309 22017 1343
rect 22051 1340 22063 1343
rect 23477 1343 23535 1349
rect 22051 1312 23428 1340
rect 22051 1309 22063 1312
rect 22005 1303 22063 1309
rect 20898 1272 20904 1284
rect 20548 1244 20760 1272
rect 20824 1244 20904 1272
rect 20548 1204 20576 1244
rect 18340 1176 20576 1204
rect 20622 1164 20628 1216
rect 20680 1164 20686 1216
rect 20732 1204 20760 1244
rect 20898 1232 20904 1244
rect 20956 1232 20962 1284
rect 23400 1216 23428 1312
rect 23477 1309 23489 1343
rect 23523 1342 23535 1343
rect 23523 1340 23612 1342
rect 23658 1340 23664 1352
rect 23523 1314 23664 1340
rect 23523 1309 23535 1314
rect 23584 1312 23664 1314
rect 23477 1303 23535 1309
rect 23658 1300 23664 1312
rect 23716 1300 23722 1352
rect 23934 1300 23940 1352
rect 23992 1340 23998 1352
rect 23992 1312 24037 1340
rect 23992 1300 23998 1312
rect 24118 1300 24124 1352
rect 24176 1300 24182 1352
rect 24213 1343 24271 1349
rect 24213 1309 24225 1343
rect 24259 1340 24271 1343
rect 25406 1340 25412 1352
rect 24259 1312 25412 1340
rect 24259 1309 24271 1312
rect 24213 1303 24271 1309
rect 25406 1300 25412 1312
rect 25464 1300 25470 1352
rect 26421 1343 26479 1349
rect 26421 1309 26433 1343
rect 26467 1309 26479 1343
rect 26421 1303 26479 1309
rect 25682 1272 25688 1284
rect 24872 1244 25688 1272
rect 23014 1204 23020 1216
rect 20732 1176 23020 1204
rect 23014 1164 23020 1176
rect 23072 1164 23078 1216
rect 23382 1164 23388 1216
rect 23440 1164 23446 1216
rect 24026 1164 24032 1216
rect 24084 1204 24090 1216
rect 24872 1204 24900 1244
rect 25682 1232 25688 1244
rect 25740 1272 25746 1284
rect 25961 1275 26019 1281
rect 25961 1272 25973 1275
rect 25740 1244 25973 1272
rect 25740 1232 25746 1244
rect 25961 1241 25973 1244
rect 26007 1272 26019 1275
rect 26436 1272 26464 1303
rect 26602 1300 26608 1352
rect 26660 1340 26666 1352
rect 26899 1351 26927 1384
rect 26748 1343 26806 1349
rect 26748 1340 26760 1343
rect 26660 1312 26760 1340
rect 26660 1300 26666 1312
rect 26748 1309 26760 1312
rect 26794 1309 26806 1343
rect 26748 1303 26806 1309
rect 26884 1345 26942 1351
rect 26884 1311 26896 1345
rect 26930 1311 26942 1345
rect 26884 1305 26942 1311
rect 26970 1300 26976 1352
rect 27028 1340 27034 1352
rect 27157 1343 27215 1349
rect 27157 1340 27169 1343
rect 27028 1312 27169 1340
rect 27028 1300 27034 1312
rect 27157 1309 27169 1312
rect 27203 1309 27215 1343
rect 27157 1303 27215 1309
rect 26007 1244 26464 1272
rect 27816 1272 27844 1516
rect 27982 1504 27988 1556
rect 28040 1544 28046 1556
rect 28261 1547 28319 1553
rect 28261 1544 28273 1547
rect 28040 1516 28273 1544
rect 28040 1504 28046 1516
rect 28261 1513 28273 1516
rect 28307 1513 28319 1547
rect 28261 1507 28319 1513
rect 28350 1504 28356 1556
rect 28408 1544 28414 1556
rect 29089 1547 29147 1553
rect 29089 1544 29101 1547
rect 28408 1516 28948 1544
rect 28408 1504 28414 1516
rect 28920 1476 28948 1516
rect 29012 1516 29101 1544
rect 29012 1476 29040 1516
rect 29089 1513 29101 1516
rect 29135 1513 29147 1547
rect 29089 1507 29147 1513
rect 29362 1504 29368 1556
rect 29420 1544 29426 1556
rect 29641 1547 29699 1553
rect 29641 1544 29653 1547
rect 29420 1516 29653 1544
rect 29420 1504 29426 1516
rect 29641 1513 29653 1516
rect 29687 1513 29699 1547
rect 29641 1507 29699 1513
rect 28920 1448 29040 1476
rect 28626 1368 28632 1420
rect 28684 1412 28690 1420
rect 28684 1401 28856 1412
rect 28905 1411 28963 1417
rect 28684 1395 28871 1401
rect 28684 1384 28825 1395
rect 28684 1368 28690 1384
rect 28813 1361 28825 1384
rect 28859 1361 28871 1395
rect 28905 1377 28917 1411
rect 28951 1408 28963 1411
rect 28994 1408 29000 1420
rect 28951 1380 29000 1408
rect 28951 1377 28963 1380
rect 28905 1371 28963 1377
rect 28994 1368 29000 1380
rect 29052 1368 29058 1420
rect 29181 1412 29239 1417
rect 29181 1411 29316 1412
rect 29181 1377 29193 1411
rect 29227 1408 29316 1411
rect 29362 1408 29368 1420
rect 29227 1384 29368 1408
rect 29227 1377 29239 1384
rect 29288 1380 29368 1384
rect 29181 1371 29239 1377
rect 29362 1368 29368 1380
rect 29420 1368 29426 1420
rect 29457 1411 29515 1417
rect 29457 1377 29469 1411
rect 29503 1377 29515 1411
rect 29457 1371 29515 1377
rect 28813 1355 28871 1361
rect 29012 1340 29040 1368
rect 29472 1340 29500 1371
rect 29012 1312 29500 1340
rect 29917 1275 29975 1281
rect 29917 1272 29929 1275
rect 27816 1244 28856 1272
rect 26007 1241 26019 1244
rect 25961 1235 26019 1241
rect 24084 1176 24900 1204
rect 24084 1164 24090 1176
rect 25314 1164 25320 1216
rect 25372 1164 25378 1216
rect 26142 1164 26148 1216
rect 26200 1204 26206 1216
rect 26970 1204 26976 1216
rect 26200 1176 26976 1204
rect 26200 1164 26206 1176
rect 26970 1164 26976 1176
rect 27028 1164 27034 1216
rect 28626 1164 28632 1216
rect 28684 1164 28690 1216
rect 28828 1204 28856 1244
rect 28966 1244 29929 1272
rect 28966 1204 28994 1244
rect 29917 1241 29929 1244
rect 29963 1241 29975 1275
rect 29917 1235 29975 1241
rect 28828 1176 28994 1204
rect 29362 1164 29368 1216
rect 29420 1164 29426 1216
rect 552 1114 30912 1136
rect 552 1062 4193 1114
rect 4245 1062 4257 1114
rect 4309 1062 4321 1114
rect 4373 1062 4385 1114
rect 4437 1062 4449 1114
rect 4501 1062 11783 1114
rect 11835 1062 11847 1114
rect 11899 1062 11911 1114
rect 11963 1062 11975 1114
rect 12027 1062 12039 1114
rect 12091 1062 19373 1114
rect 19425 1062 19437 1114
rect 19489 1062 19501 1114
rect 19553 1062 19565 1114
rect 19617 1062 19629 1114
rect 19681 1062 26963 1114
rect 27015 1062 27027 1114
rect 27079 1062 27091 1114
rect 27143 1062 27155 1114
rect 27207 1062 27219 1114
rect 27271 1062 30912 1114
rect 552 1040 30912 1062
rect 2961 1003 3019 1009
rect 2961 969 2973 1003
rect 3007 1000 3019 1003
rect 6914 1000 6920 1012
rect 3007 972 6920 1000
rect 3007 969 3019 972
rect 2961 963 3019 969
rect 6914 960 6920 972
rect 6972 960 6978 1012
rect 7650 960 7656 1012
rect 7708 960 7714 1012
rect 9306 960 9312 1012
rect 9364 1000 9370 1012
rect 10229 1003 10287 1009
rect 10229 1000 10241 1003
rect 9364 972 10241 1000
rect 9364 960 9370 972
rect 10229 969 10241 972
rect 10275 969 10287 1003
rect 10229 963 10287 969
rect 10594 960 10600 1012
rect 10652 960 10658 1012
rect 10965 1003 11023 1009
rect 10965 969 10977 1003
rect 11011 1000 11023 1003
rect 12158 1000 12164 1012
rect 11011 972 12164 1000
rect 11011 969 11023 972
rect 10965 963 11023 969
rect 12158 960 12164 972
rect 12216 960 12222 1012
rect 12342 960 12348 1012
rect 12400 1000 12406 1012
rect 13265 1003 13323 1009
rect 12400 972 13216 1000
rect 12400 960 12406 972
rect 5166 932 5172 944
rect 2976 904 5172 932
rect 934 824 940 876
rect 992 824 998 876
rect 1448 855 1624 864
rect 1433 849 1624 855
rect 1433 815 1445 849
rect 1479 836 1624 849
rect 1479 815 1491 836
rect 1433 809 1491 815
rect 1596 796 1624 836
rect 1670 824 1676 876
rect 1728 824 1734 876
rect 2976 796 3004 904
rect 5166 892 5172 904
rect 5224 892 5230 944
rect 13188 932 13216 972
rect 13265 969 13277 1003
rect 13311 1000 13323 1003
rect 13354 1000 13360 1012
rect 13311 972 13360 1000
rect 13311 969 13323 972
rect 13265 963 13323 969
rect 13354 960 13360 972
rect 13412 960 13418 1012
rect 13538 960 13544 1012
rect 13596 960 13602 1012
rect 16117 1003 16175 1009
rect 13648 972 16068 1000
rect 13648 932 13676 972
rect 13188 904 13676 932
rect 16040 932 16068 972
rect 16117 969 16129 1003
rect 16163 1000 16175 1003
rect 16850 1000 16856 1012
rect 16163 972 16856 1000
rect 16163 969 16175 972
rect 16117 963 16175 969
rect 16850 960 16856 972
rect 16908 960 16914 1012
rect 16942 960 16948 1012
rect 17000 1000 17006 1012
rect 18693 1003 18751 1009
rect 18693 1000 18705 1003
rect 17000 972 18705 1000
rect 17000 960 17006 972
rect 18693 969 18705 972
rect 18739 969 18751 1003
rect 20438 1000 20444 1012
rect 18693 963 18751 969
rect 18892 972 20444 1000
rect 16206 932 16212 944
rect 16040 904 16212 932
rect 16206 892 16212 904
rect 16264 892 16270 944
rect 17954 892 17960 944
rect 18012 932 18018 944
rect 18892 932 18920 972
rect 20438 960 20444 972
rect 20496 960 20502 1012
rect 25314 1000 25320 1012
rect 20640 972 25320 1000
rect 18012 904 18920 932
rect 18012 892 18018 904
rect 6270 824 6276 876
rect 6328 824 6334 876
rect 6638 824 6644 876
rect 6696 864 6702 876
rect 6696 836 8340 864
rect 6696 824 6702 836
rect 1596 768 3004 796
rect 3602 756 3608 808
rect 3660 796 3666 808
rect 3881 799 3939 805
rect 3881 796 3893 799
rect 3660 768 3893 796
rect 3660 756 3666 768
rect 3881 765 3893 768
rect 3927 796 3939 799
rect 4982 796 4988 808
rect 3927 768 4988 796
rect 3927 765 3939 768
rect 3881 759 3939 765
rect 4982 756 4988 768
rect 5040 756 5046 808
rect 5626 756 5632 808
rect 5684 756 5690 808
rect 5810 756 5816 808
rect 5868 756 5874 808
rect 6549 799 6607 805
rect 6549 765 6561 799
rect 6595 796 6607 799
rect 7834 796 7840 808
rect 6595 768 7840 796
rect 6595 765 6607 768
rect 6549 759 6607 765
rect 7834 756 7840 768
rect 7892 756 7898 808
rect 8312 796 8340 836
rect 8386 824 8392 876
rect 8444 824 8450 876
rect 8852 867 8910 873
rect 8852 864 8864 867
rect 8496 836 8864 864
rect 8496 796 8524 836
rect 8852 833 8864 836
rect 8898 833 8910 867
rect 8852 827 8910 833
rect 10502 824 10508 876
rect 10560 864 10566 876
rect 11606 864 11612 876
rect 10560 836 11612 864
rect 10560 824 10566 836
rect 8312 768 8524 796
rect 9030 756 9036 808
rect 9088 796 9094 808
rect 10796 805 10824 836
rect 11606 824 11612 836
rect 11664 824 11670 876
rect 11747 867 11805 873
rect 11747 833 11759 867
rect 11793 864 11805 867
rect 12066 864 12072 876
rect 11793 836 12072 864
rect 11793 833 11805 836
rect 11747 827 11805 833
rect 12066 824 12072 836
rect 12124 824 12130 876
rect 14366 871 14372 876
rect 14323 865 14372 871
rect 13556 836 13860 864
rect 9125 799 9183 805
rect 9125 796 9137 799
rect 9088 768 9137 796
rect 9088 756 9094 768
rect 9125 765 9137 768
rect 9171 765 9183 799
rect 9125 759 9183 765
rect 10781 799 10839 805
rect 10781 765 10793 799
rect 10827 765 10839 799
rect 10781 759 10839 765
rect 11146 756 11152 808
rect 11204 756 11210 808
rect 11241 799 11299 805
rect 11241 765 11253 799
rect 11287 796 11299 799
rect 11882 796 11888 808
rect 11287 768 11888 796
rect 11287 765 11299 768
rect 11241 759 11299 765
rect 11256 728 11284 759
rect 11882 756 11888 768
rect 11940 756 11946 808
rect 11977 799 12035 805
rect 11977 765 11989 799
rect 12023 796 12035 799
rect 12250 796 12256 808
rect 12023 768 12256 796
rect 12023 765 12035 768
rect 11977 759 12035 765
rect 12250 756 12256 768
rect 12308 756 12314 808
rect 11164 700 11284 728
rect 1394 620 1400 672
rect 1452 669 1458 672
rect 1452 660 1461 669
rect 1452 632 1497 660
rect 1452 623 1461 632
rect 1452 620 1458 623
rect 1670 620 1676 672
rect 1728 660 1734 672
rect 3513 663 3571 669
rect 3513 660 3525 663
rect 1728 632 3525 660
rect 1728 620 1734 632
rect 3513 629 3525 632
rect 3559 660 3571 663
rect 5350 660 5356 672
rect 3559 632 5356 660
rect 3559 629 3571 632
rect 3513 623 3571 629
rect 5350 620 5356 632
rect 5408 620 5414 672
rect 5442 620 5448 672
rect 5500 620 5506 672
rect 6279 663 6337 669
rect 6279 629 6291 663
rect 6325 660 6337 663
rect 7558 660 7564 672
rect 6325 632 7564 660
rect 6325 629 6337 632
rect 6279 623 6337 629
rect 7558 620 7564 632
rect 7616 620 7622 672
rect 8294 620 8300 672
rect 8352 660 8358 672
rect 8855 663 8913 669
rect 8855 660 8867 663
rect 8352 632 8867 660
rect 8352 620 8358 632
rect 8855 629 8867 632
rect 8901 629 8913 663
rect 8855 623 8913 629
rect 9122 620 9128 672
rect 9180 660 9186 672
rect 11164 660 11192 700
rect 9180 632 11192 660
rect 9180 620 9186 632
rect 11330 620 11336 672
rect 11388 660 11394 672
rect 11707 663 11765 669
rect 11707 660 11719 663
rect 11388 632 11719 660
rect 11388 620 11394 632
rect 11707 629 11719 632
rect 11753 660 11765 663
rect 12066 660 12072 672
rect 11753 632 12072 660
rect 11753 629 11765 632
rect 11707 623 11765 629
rect 12066 620 12072 632
rect 12124 620 12130 672
rect 12250 620 12256 672
rect 12308 660 12314 672
rect 13556 660 13584 836
rect 13832 808 13860 836
rect 14323 831 14335 865
rect 14369 831 14372 865
rect 14323 825 14372 831
rect 14366 824 14372 825
rect 14424 824 14430 876
rect 16899 867 16957 873
rect 16899 833 16911 867
rect 16945 864 16957 867
rect 17034 864 17040 876
rect 16945 836 17040 864
rect 16945 833 16957 836
rect 16899 827 16957 833
rect 17034 824 17040 836
rect 17092 824 17098 876
rect 17129 867 17187 873
rect 17129 833 17141 867
rect 17175 864 17187 867
rect 18782 864 18788 876
rect 17175 836 18788 864
rect 17175 833 17187 836
rect 17129 827 17187 833
rect 18782 824 18788 836
rect 18840 824 18846 876
rect 13722 805 13728 808
rect 13717 796 13728 805
rect 13683 768 13728 796
rect 13717 759 13728 768
rect 13722 756 13728 759
rect 13780 756 13786 808
rect 13814 756 13820 808
rect 13872 756 13878 808
rect 14144 799 14202 805
rect 14144 765 14156 799
rect 14190 796 14202 799
rect 14458 796 14464 808
rect 14190 768 14464 796
rect 14190 765 14202 768
rect 14144 759 14202 765
rect 14458 756 14464 768
rect 14516 756 14522 808
rect 14553 799 14611 805
rect 14553 765 14565 799
rect 14599 796 14611 799
rect 15010 796 15016 808
rect 14599 768 15016 796
rect 14599 765 14611 768
rect 14553 759 14611 765
rect 15010 756 15016 768
rect 15068 756 15074 808
rect 16298 756 16304 808
rect 16356 756 16362 808
rect 16390 756 16396 808
rect 16448 756 16454 808
rect 18892 805 18920 904
rect 19475 867 19533 873
rect 19475 833 19487 867
rect 19521 864 19533 867
rect 20640 864 20668 972
rect 25314 960 25320 972
rect 25372 960 25378 1012
rect 25406 960 25412 1012
rect 25464 1000 25470 1012
rect 26421 1003 26479 1009
rect 26421 1000 26433 1003
rect 25464 972 26433 1000
rect 25464 960 25470 972
rect 26421 969 26433 972
rect 26467 969 26479 1003
rect 26421 963 26479 969
rect 28534 960 28540 1012
rect 28592 960 28598 1012
rect 20898 892 20904 944
rect 20956 932 20962 944
rect 21269 935 21327 941
rect 21269 932 21281 935
rect 20956 904 21281 932
rect 20956 892 20962 904
rect 21269 901 21281 904
rect 21315 901 21327 935
rect 21269 895 21327 901
rect 25498 892 25504 944
rect 25556 932 25562 944
rect 26142 932 26148 944
rect 25556 904 26148 932
rect 25556 892 25562 904
rect 26142 892 26148 904
rect 26200 892 26206 944
rect 19521 836 20668 864
rect 19521 833 19533 836
rect 19475 827 19533 833
rect 20806 824 20812 876
rect 20864 864 20870 876
rect 21542 864 21548 876
rect 20864 836 21548 864
rect 20864 824 20870 836
rect 21542 824 21548 836
rect 21600 824 21606 876
rect 22051 867 22109 873
rect 22051 833 22063 867
rect 22097 864 22109 867
rect 22097 836 23520 864
rect 22097 833 22109 836
rect 22051 827 22109 833
rect 18877 799 18935 805
rect 18877 765 18889 799
rect 18923 765 18935 799
rect 18877 759 18935 765
rect 18969 799 19027 805
rect 18969 765 18981 799
rect 19015 765 19027 799
rect 18969 759 19027 765
rect 19705 799 19763 805
rect 19705 765 19717 799
rect 19751 796 19763 799
rect 21266 796 21272 808
rect 19751 768 21272 796
rect 19751 765 19763 768
rect 19705 759 19763 765
rect 15933 731 15991 737
rect 15933 697 15945 731
rect 15979 728 15991 731
rect 16482 728 16488 740
rect 15979 700 16488 728
rect 15979 697 15991 700
rect 15933 691 15991 697
rect 16482 688 16488 700
rect 16540 688 16546 740
rect 18156 700 18368 728
rect 12308 632 13584 660
rect 12308 620 12314 632
rect 13630 620 13636 672
rect 13688 660 13694 672
rect 16859 663 16917 669
rect 16859 660 16871 663
rect 13688 632 16871 660
rect 13688 620 13694 632
rect 16859 629 16871 632
rect 16905 660 16917 663
rect 18156 660 18184 700
rect 16905 632 18184 660
rect 16905 629 16917 632
rect 16859 623 16917 629
rect 18230 620 18236 672
rect 18288 620 18294 672
rect 18340 660 18368 700
rect 18414 688 18420 740
rect 18472 728 18478 740
rect 18984 728 19012 759
rect 21266 756 21272 768
rect 21324 756 21330 808
rect 21453 799 21511 805
rect 21453 765 21465 799
rect 21499 765 21511 799
rect 21453 759 21511 765
rect 18472 700 19012 728
rect 18472 688 18478 700
rect 20438 688 20444 740
rect 20496 728 20502 740
rect 21468 728 21496 759
rect 21634 756 21640 808
rect 21692 796 21698 808
rect 21872 799 21930 805
rect 21872 796 21884 799
rect 21692 768 21884 796
rect 21692 756 21698 768
rect 21872 765 21884 768
rect 21918 765 21930 799
rect 21872 759 21930 765
rect 22281 799 22339 805
rect 22281 765 22293 799
rect 22327 796 22339 799
rect 23014 796 23020 808
rect 22327 768 23020 796
rect 22327 765 22339 768
rect 22281 759 22339 765
rect 23014 756 23020 768
rect 23072 756 23078 808
rect 20496 700 21496 728
rect 23492 728 23520 836
rect 23566 824 23572 876
rect 23624 864 23630 876
rect 24308 867 24366 873
rect 24308 864 24320 867
rect 23624 836 24320 864
rect 23624 824 23630 836
rect 24308 833 24320 836
rect 24354 833 24366 867
rect 24308 827 24366 833
rect 24578 824 24584 876
rect 24636 824 24642 876
rect 25222 824 25228 876
rect 25280 824 25286 876
rect 26418 824 26424 876
rect 26476 824 26482 876
rect 26697 867 26755 873
rect 26697 833 26709 867
rect 26743 864 26755 867
rect 26878 864 26884 876
rect 26743 836 26884 864
rect 26743 833 26755 836
rect 26697 827 26755 833
rect 26878 824 26884 836
rect 26936 824 26942 876
rect 27203 867 27261 873
rect 27203 833 27215 867
rect 27249 833 27261 867
rect 27203 827 27261 833
rect 23658 756 23664 808
rect 23716 756 23722 808
rect 23842 756 23848 808
rect 23900 756 23906 808
rect 24486 796 24492 808
rect 23958 768 24492 796
rect 23750 728 23756 740
rect 23492 700 23756 728
rect 20496 688 20502 700
rect 19435 663 19493 669
rect 19435 660 19447 663
rect 18340 632 19447 660
rect 19435 629 19447 632
rect 19481 660 19493 663
rect 20530 660 20536 672
rect 19481 632 20536 660
rect 19481 629 19493 632
rect 19435 623 19493 629
rect 20530 620 20536 632
rect 20588 620 20594 672
rect 20806 620 20812 672
rect 20864 620 20870 672
rect 21468 660 21496 700
rect 23750 688 23756 700
rect 23808 688 23814 740
rect 23958 660 23986 768
rect 24486 756 24492 768
rect 24544 756 24550 808
rect 25240 728 25268 824
rect 26237 799 26295 805
rect 26237 765 26249 799
rect 26283 796 26295 799
rect 26436 796 26464 824
rect 26283 768 26464 796
rect 26283 765 26295 768
rect 26237 759 26295 765
rect 26602 756 26608 808
rect 26660 756 26666 808
rect 26786 756 26792 808
rect 26844 796 26850 808
rect 27024 799 27082 805
rect 27024 796 27036 799
rect 26844 768 27036 796
rect 26844 756 26850 768
rect 27024 765 27036 768
rect 27070 765 27082 799
rect 27218 796 27246 827
rect 27338 824 27344 876
rect 27396 864 27402 876
rect 27433 867 27491 873
rect 27433 864 27445 867
rect 27396 836 27445 864
rect 27396 824 27402 836
rect 27433 833 27445 836
rect 27479 833 27491 867
rect 27433 827 27491 833
rect 27522 796 27528 808
rect 27218 768 27528 796
rect 27024 759 27082 765
rect 27522 756 27528 768
rect 27580 756 27586 808
rect 28997 799 29055 805
rect 28997 765 29009 799
rect 29043 796 29055 799
rect 29454 796 29460 808
rect 29043 768 29460 796
rect 29043 765 29055 768
rect 28997 759 29055 765
rect 29454 756 29460 768
rect 29512 756 29518 808
rect 25240 700 26832 728
rect 21468 632 23986 660
rect 24118 620 24124 672
rect 24176 660 24182 672
rect 24311 663 24369 669
rect 24311 660 24323 663
rect 24176 632 24323 660
rect 24176 620 24182 632
rect 24311 629 24323 632
rect 24357 629 24369 663
rect 24311 623 24369 629
rect 25682 620 25688 672
rect 25740 620 25746 672
rect 26050 620 26056 672
rect 26108 620 26114 672
rect 26804 660 26832 700
rect 29181 663 29239 669
rect 29181 660 29193 663
rect 26804 632 29193 660
rect 29181 629 29193 632
rect 29227 629 29239 663
rect 29181 623 29239 629
rect 552 570 31072 592
rect 552 518 7988 570
rect 8040 518 8052 570
rect 8104 518 8116 570
rect 8168 518 8180 570
rect 8232 518 8244 570
rect 8296 518 15578 570
rect 15630 518 15642 570
rect 15694 518 15706 570
rect 15758 518 15770 570
rect 15822 518 15834 570
rect 15886 518 23168 570
rect 23220 518 23232 570
rect 23284 518 23296 570
rect 23348 518 23360 570
rect 23412 518 23424 570
rect 23476 518 30758 570
rect 30810 518 30822 570
rect 30874 518 30886 570
rect 30938 518 30950 570
rect 31002 518 31014 570
rect 31066 518 31072 570
rect 552 496 31072 518
rect 3970 416 3976 468
rect 4028 456 4034 468
rect 6914 456 6920 468
rect 4028 428 6920 456
rect 4028 416 4034 428
rect 6914 416 6920 428
rect 6972 416 6978 468
rect 7558 416 7564 468
rect 7616 416 7622 468
rect 7834 416 7840 468
rect 7892 456 7898 468
rect 20714 456 20720 468
rect 7892 428 20720 456
rect 7892 416 7898 428
rect 20714 416 20720 428
rect 20772 416 20778 468
rect 23750 416 23756 468
rect 23808 456 23814 468
rect 25590 456 25596 468
rect 23808 428 25596 456
rect 23808 416 23814 428
rect 25590 416 25596 428
rect 25648 416 25654 468
rect 7576 388 7604 416
rect 13630 388 13636 400
rect 7576 360 13636 388
rect 13630 348 13636 360
rect 13688 348 13694 400
rect 14458 348 14464 400
rect 14516 388 14522 400
rect 18598 388 18604 400
rect 14516 360 18604 388
rect 14516 348 14522 360
rect 18598 348 18604 360
rect 18656 348 18662 400
rect 23014 348 23020 400
rect 23072 388 23078 400
rect 25866 388 25872 400
rect 23072 360 25872 388
rect 23072 348 23078 360
rect 25866 348 25872 360
rect 25924 348 25930 400
rect 5442 280 5448 332
rect 5500 320 5506 332
rect 11514 320 11520 332
rect 5500 292 11520 320
rect 5500 280 5506 292
rect 11514 280 11520 292
rect 11572 280 11578 332
rect 11606 280 11612 332
rect 11664 320 11670 332
rect 13722 320 13728 332
rect 11664 292 13728 320
rect 11664 280 11670 292
rect 13722 280 13728 292
rect 13780 280 13786 332
rect 13814 280 13820 332
rect 13872 320 13878 332
rect 18506 320 18512 332
rect 13872 292 18512 320
rect 13872 280 13878 292
rect 18506 280 18512 292
rect 18564 280 18570 332
rect 22830 280 22836 332
rect 22888 320 22894 332
rect 26050 320 26056 332
rect 22888 292 26056 320
rect 22888 280 22894 292
rect 26050 280 26056 292
rect 26108 280 26114 332
rect 5994 212 6000 264
rect 6052 252 6058 264
rect 9030 252 9036 264
rect 6052 224 9036 252
rect 6052 212 6058 224
rect 9030 212 9036 224
rect 9088 252 9094 264
rect 12342 252 12348 264
rect 9088 224 12348 252
rect 9088 212 9094 224
rect 12342 212 12348 224
rect 12400 212 12406 264
rect 21266 212 21272 264
rect 21324 252 21330 264
rect 28626 252 28632 264
rect 21324 224 28632 252
rect 21324 212 21330 224
rect 28626 212 28632 224
rect 28684 212 28690 264
rect 5074 144 5080 196
rect 5132 144 5138 196
rect 5350 144 5356 196
rect 5408 184 5414 196
rect 15378 184 15384 196
rect 5408 156 15384 184
rect 5408 144 5414 156
rect 15378 144 15384 156
rect 15436 144 15442 196
rect 18782 144 18788 196
rect 18840 184 18846 196
rect 28350 184 28356 196
rect 18840 156 28356 184
rect 18840 144 18846 156
rect 28350 144 28356 156
rect 28408 144 28414 196
rect 5092 116 5120 144
rect 9122 116 9128 128
rect 5092 88 9128 116
rect 9122 76 9128 88
rect 9180 76 9186 128
rect 22738 116 22744 128
rect 18432 88 22744 116
rect 18432 60 18460 88
rect 22738 76 22744 88
rect 22796 76 22802 128
rect 5810 8 5816 60
rect 5868 48 5874 60
rect 16390 48 16396 60
rect 5868 20 16396 48
rect 5868 8 5874 20
rect 16390 8 16396 20
rect 16448 48 16454 60
rect 18414 48 18420 60
rect 16448 20 18420 48
rect 16448 8 16454 20
rect 18414 8 18420 20
rect 18472 8 18478 60
rect 18598 8 18604 60
rect 18656 48 18662 60
rect 19702 48 19708 60
rect 18656 20 19708 48
rect 18656 8 18662 20
rect 19702 8 19708 20
rect 19760 48 19766 60
rect 26786 48 26792 60
rect 19760 20 26792 48
rect 19760 8 19766 20
rect 26786 8 26792 20
rect 26844 8 26850 60
<< via1 >>
rect 1952 22244 2004 22296
rect 8852 22244 8904 22296
rect 4068 22176 4120 22228
rect 9680 22244 9732 22296
rect 18788 22244 18840 22296
rect 23572 22244 23624 22296
rect 9128 22176 9180 22228
rect 9772 22176 9824 22228
rect 3056 22108 3108 22160
rect 12900 22176 12952 22228
rect 12808 22108 12860 22160
rect 5264 22040 5316 22092
rect 9588 22040 9640 22092
rect 12440 22040 12492 22092
rect 18512 22176 18564 22228
rect 22376 22176 22428 22228
rect 22468 22176 22520 22228
rect 25964 22244 26016 22296
rect 23756 22176 23808 22228
rect 28724 22176 28776 22228
rect 18604 22108 18656 22160
rect 28080 22108 28132 22160
rect 28172 22040 28224 22092
rect 12624 21972 12676 22024
rect 2136 21836 2188 21888
rect 2504 21836 2556 21888
rect 3792 21836 3844 21888
rect 7196 21904 7248 21956
rect 16120 21904 16172 21956
rect 8760 21836 8812 21888
rect 8852 21836 8904 21888
rect 12532 21836 12584 21888
rect 13728 21836 13780 21888
rect 18420 21904 18472 21956
rect 19248 21904 19300 21956
rect 28356 21972 28408 22024
rect 23296 21904 23348 21956
rect 16672 21836 16724 21888
rect 21364 21836 21416 21888
rect 22284 21836 22336 21888
rect 26608 21836 26660 21888
rect 30472 21836 30524 21888
rect 4193 21734 4245 21786
rect 4257 21734 4309 21786
rect 4321 21734 4373 21786
rect 4385 21734 4437 21786
rect 4449 21734 4501 21786
rect 11783 21734 11835 21786
rect 11847 21734 11899 21786
rect 11911 21734 11963 21786
rect 11975 21734 12027 21786
rect 12039 21734 12091 21786
rect 19373 21734 19425 21786
rect 19437 21734 19489 21786
rect 19501 21734 19553 21786
rect 19565 21734 19617 21786
rect 19629 21734 19681 21786
rect 26963 21734 27015 21786
rect 27027 21734 27079 21786
rect 27091 21734 27143 21786
rect 27155 21734 27207 21786
rect 27219 21734 27271 21786
rect 2780 21632 2832 21684
rect 8208 21632 8260 21684
rect 5540 21564 5592 21616
rect 3424 21496 3476 21548
rect 1676 21471 1728 21480
rect 1676 21437 1685 21471
rect 1685 21437 1719 21471
rect 1719 21437 1728 21471
rect 1676 21428 1728 21437
rect 3240 21471 3292 21480
rect 3240 21437 3249 21471
rect 3249 21437 3283 21471
rect 3283 21437 3292 21471
rect 3240 21428 3292 21437
rect 8944 21496 8996 21548
rect 9128 21539 9180 21548
rect 9128 21505 9137 21539
rect 9137 21505 9171 21539
rect 9171 21505 9180 21539
rect 9128 21496 9180 21505
rect 9496 21496 9548 21548
rect 3976 21471 4028 21480
rect 3976 21437 3985 21471
rect 3985 21437 4019 21471
rect 4019 21437 4028 21471
rect 3976 21428 4028 21437
rect 4804 21428 4856 21480
rect 5540 21428 5592 21480
rect 5908 21428 5960 21480
rect 8208 21471 8260 21480
rect 8208 21437 8217 21471
rect 8217 21437 8251 21471
rect 8251 21437 8260 21471
rect 8208 21428 8260 21437
rect 8392 21471 8444 21480
rect 8392 21437 8401 21471
rect 8401 21437 8435 21471
rect 8435 21437 8444 21471
rect 8392 21428 8444 21437
rect 1400 21335 1452 21344
rect 1400 21301 1415 21335
rect 1415 21301 1449 21335
rect 1449 21301 1452 21335
rect 1400 21292 1452 21301
rect 3516 21292 3568 21344
rect 5448 21335 5500 21344
rect 5448 21301 5457 21335
rect 5457 21301 5491 21335
rect 5491 21301 5500 21335
rect 5448 21292 5500 21301
rect 7564 21360 7616 21412
rect 8668 21428 8720 21480
rect 9404 21428 9456 21480
rect 10692 21428 10744 21480
rect 10876 21428 10928 21480
rect 10968 21471 11020 21480
rect 10968 21437 10977 21471
rect 10977 21437 11011 21471
rect 11011 21437 11020 21471
rect 10968 21428 11020 21437
rect 11060 21428 11112 21480
rect 11612 21428 11664 21480
rect 12532 21632 12584 21684
rect 12808 21675 12860 21684
rect 12808 21641 12817 21675
rect 12817 21641 12851 21675
rect 12851 21641 12860 21675
rect 12808 21632 12860 21641
rect 16120 21632 16172 21684
rect 13912 21564 13964 21616
rect 12624 21496 12676 21548
rect 13268 21496 13320 21548
rect 13728 21496 13780 21548
rect 14096 21428 14148 21480
rect 14372 21428 14424 21480
rect 14648 21428 14700 21480
rect 6184 21292 6236 21344
rect 6276 21335 6328 21344
rect 6276 21301 6291 21335
rect 6291 21301 6325 21335
rect 6325 21301 6328 21335
rect 6276 21292 6328 21301
rect 6644 21292 6696 21344
rect 7840 21292 7892 21344
rect 8484 21292 8536 21344
rect 10048 21292 10100 21344
rect 10600 21335 10652 21344
rect 10600 21301 10609 21335
rect 10609 21301 10643 21335
rect 10643 21301 10652 21335
rect 10600 21292 10652 21301
rect 11336 21292 11388 21344
rect 13176 21335 13228 21344
rect 13176 21301 13185 21335
rect 13185 21301 13219 21335
rect 13219 21301 13228 21335
rect 13176 21292 13228 21301
rect 13360 21292 13412 21344
rect 15936 21403 15988 21412
rect 15936 21369 15945 21403
rect 15945 21369 15979 21403
rect 15979 21369 15988 21403
rect 15936 21360 15988 21369
rect 16672 21564 16724 21616
rect 18512 21632 18564 21684
rect 18788 21564 18840 21616
rect 19892 21632 19944 21684
rect 21088 21632 21140 21684
rect 21640 21564 21692 21616
rect 22008 21564 22060 21616
rect 18604 21428 18656 21480
rect 19340 21471 19392 21480
rect 19340 21437 19349 21471
rect 19349 21437 19383 21471
rect 19383 21437 19392 21471
rect 19340 21428 19392 21437
rect 19432 21471 19484 21480
rect 19432 21437 19441 21471
rect 19441 21437 19475 21471
rect 19475 21437 19484 21471
rect 19432 21428 19484 21437
rect 21548 21496 21600 21548
rect 25964 21564 26016 21616
rect 19800 21428 19852 21480
rect 21272 21471 21324 21480
rect 21272 21437 21281 21471
rect 21281 21437 21315 21471
rect 21315 21437 21324 21471
rect 21272 21428 21324 21437
rect 21456 21471 21508 21480
rect 21456 21437 21465 21471
rect 21465 21437 21499 21471
rect 21499 21437 21508 21471
rect 21456 21428 21508 21437
rect 22192 21471 22244 21480
rect 22192 21437 22201 21471
rect 22201 21437 22235 21471
rect 22235 21437 22244 21471
rect 22192 21428 22244 21437
rect 23756 21496 23808 21548
rect 23940 21496 23992 21548
rect 24032 21539 24084 21548
rect 24032 21505 24041 21539
rect 24041 21505 24075 21539
rect 24075 21505 24084 21539
rect 24032 21496 24084 21505
rect 24492 21539 24544 21548
rect 24492 21505 24501 21539
rect 24501 21505 24535 21539
rect 24535 21505 24544 21539
rect 24492 21496 24544 21505
rect 24584 21496 24636 21548
rect 25412 21496 25464 21548
rect 27528 21496 27580 21548
rect 23296 21360 23348 21412
rect 23572 21471 23624 21480
rect 23572 21437 23581 21471
rect 23581 21437 23615 21471
rect 23615 21437 23624 21471
rect 23572 21428 23624 21437
rect 23664 21471 23716 21480
rect 23664 21437 23673 21471
rect 23673 21437 23707 21471
rect 23707 21437 23716 21471
rect 23664 21428 23716 21437
rect 24860 21428 24912 21480
rect 25044 21471 25096 21480
rect 25044 21437 25053 21471
rect 25053 21437 25087 21471
rect 25087 21437 25096 21471
rect 25044 21428 25096 21437
rect 23848 21360 23900 21412
rect 19156 21335 19208 21344
rect 19156 21301 19165 21335
rect 19165 21301 19199 21335
rect 19199 21301 19208 21335
rect 19156 21292 19208 21301
rect 20996 21335 21048 21344
rect 20996 21301 21005 21335
rect 21005 21301 21039 21335
rect 21039 21301 21048 21335
rect 20996 21292 21048 21301
rect 22008 21292 22060 21344
rect 26240 21428 26292 21480
rect 26608 21471 26660 21480
rect 26608 21437 26617 21471
rect 26617 21437 26651 21471
rect 26651 21437 26660 21471
rect 26608 21428 26660 21437
rect 26792 21428 26844 21480
rect 27896 21428 27948 21480
rect 26148 21360 26200 21412
rect 24032 21292 24084 21344
rect 25320 21292 25372 21344
rect 25688 21335 25740 21344
rect 25688 21301 25697 21335
rect 25697 21301 25731 21335
rect 25731 21301 25740 21335
rect 25688 21292 25740 21301
rect 25872 21292 25924 21344
rect 26424 21335 26476 21344
rect 26424 21301 26433 21335
rect 26433 21301 26467 21335
rect 26467 21301 26476 21335
rect 26424 21292 26476 21301
rect 28540 21335 28592 21344
rect 28540 21301 28549 21335
rect 28549 21301 28583 21335
rect 28583 21301 28592 21335
rect 28540 21292 28592 21301
rect 30012 21292 30064 21344
rect 30288 21335 30340 21344
rect 30288 21301 30297 21335
rect 30297 21301 30331 21335
rect 30331 21301 30340 21335
rect 30288 21292 30340 21301
rect 31300 21292 31352 21344
rect 7988 21190 8040 21242
rect 8052 21190 8104 21242
rect 8116 21190 8168 21242
rect 8180 21190 8232 21242
rect 8244 21190 8296 21242
rect 15578 21190 15630 21242
rect 15642 21190 15694 21242
rect 15706 21190 15758 21242
rect 15770 21190 15822 21242
rect 15834 21190 15886 21242
rect 23168 21190 23220 21242
rect 23232 21190 23284 21242
rect 23296 21190 23348 21242
rect 23360 21190 23412 21242
rect 23424 21190 23476 21242
rect 30758 21190 30810 21242
rect 30822 21190 30874 21242
rect 30886 21190 30938 21242
rect 30950 21190 31002 21242
rect 31014 21190 31066 21242
rect 7932 21088 7984 21140
rect 1952 21063 2004 21072
rect 1952 21029 1961 21063
rect 1961 21029 1995 21063
rect 1995 21029 2004 21063
rect 1952 21020 2004 21029
rect 2136 21063 2188 21072
rect 2136 21029 2145 21063
rect 2145 21029 2179 21063
rect 2179 21029 2188 21063
rect 2136 21020 2188 21029
rect 5264 21063 5316 21072
rect 5264 21029 5273 21063
rect 5273 21029 5307 21063
rect 5307 21029 5316 21063
rect 5264 21020 5316 21029
rect 5816 21020 5868 21072
rect 1124 20952 1176 21004
rect 1400 20952 1452 21004
rect 2964 20995 3016 21004
rect 2964 20961 2966 20995
rect 2966 20961 3016 20995
rect 2964 20952 3016 20961
rect 3792 20952 3844 21004
rect 4988 20952 5040 21004
rect 6000 20995 6052 21004
rect 6000 20961 6009 20995
rect 6009 20961 6043 20995
rect 6043 20961 6052 20995
rect 6000 20952 6052 20961
rect 6092 20952 6144 21004
rect 7196 21020 7248 21072
rect 8576 21088 8628 21140
rect 8760 21088 8812 21140
rect 10600 21088 10652 21140
rect 11520 21088 11572 21140
rect 12348 21088 12400 21140
rect 12440 21088 12492 21140
rect 15200 21088 15252 21140
rect 17960 21088 18012 21140
rect 19432 21088 19484 21140
rect 19984 21088 20036 21140
rect 21272 21088 21324 21140
rect 22192 21088 22244 21140
rect 8024 20952 8076 21004
rect 10968 21020 11020 21072
rect 11060 21020 11112 21072
rect 2780 20884 2832 20936
rect 3056 20911 3101 20936
rect 3101 20911 3108 20936
rect 3056 20884 3108 20911
rect 3700 20884 3752 20936
rect 7656 20884 7708 20936
rect 8300 20927 8352 20936
rect 8300 20893 8309 20927
rect 8309 20893 8343 20927
rect 8343 20893 8352 20927
rect 8300 20884 8352 20893
rect 8668 20927 8720 20936
rect 8668 20893 8670 20927
rect 8670 20893 8720 20927
rect 8668 20884 8720 20893
rect 9680 20952 9732 21004
rect 8852 20884 8904 20936
rect 10784 20952 10836 21004
rect 14648 21020 14700 21072
rect 11520 20952 11572 21004
rect 10508 20884 10560 20936
rect 11796 20884 11848 20936
rect 4068 20748 4120 20800
rect 4528 20748 4580 20800
rect 5264 20748 5316 20800
rect 5816 20791 5868 20800
rect 5816 20757 5825 20791
rect 5825 20757 5859 20791
rect 5859 20757 5868 20791
rect 5816 20748 5868 20757
rect 7472 20748 7524 20800
rect 7748 20748 7800 20800
rect 11244 20816 11296 20868
rect 10968 20791 11020 20800
rect 10968 20757 10977 20791
rect 10977 20757 11011 20791
rect 11011 20757 11020 20791
rect 10968 20748 11020 20757
rect 11152 20748 11204 20800
rect 13544 20995 13596 21004
rect 13544 20961 13553 20995
rect 13553 20961 13587 20995
rect 13587 20961 13596 20995
rect 13544 20952 13596 20961
rect 14280 20952 14332 21004
rect 14832 20952 14884 21004
rect 18144 20952 18196 21004
rect 18420 20995 18472 21004
rect 18420 20961 18429 20995
rect 18429 20961 18463 20995
rect 18463 20961 18472 20995
rect 18420 20952 18472 20961
rect 19248 21020 19300 21072
rect 22836 21020 22888 21072
rect 25320 21131 25372 21140
rect 25320 21097 25329 21131
rect 25329 21097 25363 21131
rect 25363 21097 25372 21131
rect 25320 21088 25372 21097
rect 30288 21088 30340 21140
rect 30472 21131 30524 21140
rect 30472 21097 30481 21131
rect 30481 21097 30515 21131
rect 30515 21097 30524 21131
rect 30472 21088 30524 21097
rect 16396 20927 16448 20936
rect 16396 20893 16405 20927
rect 16405 20893 16439 20927
rect 16439 20893 16448 20927
rect 20720 20952 20772 21004
rect 16396 20884 16448 20893
rect 15108 20748 15160 20800
rect 15292 20748 15344 20800
rect 16488 20748 16540 20800
rect 19708 20884 19760 20936
rect 23112 20952 23164 21004
rect 21272 20927 21324 20936
rect 21272 20893 21281 20927
rect 21281 20893 21315 20927
rect 21315 20893 21324 20927
rect 21272 20884 21324 20893
rect 25136 20952 25188 21004
rect 28080 21063 28132 21072
rect 28080 21029 28089 21063
rect 28089 21029 28123 21063
rect 28123 21029 28132 21063
rect 28080 21020 28132 21029
rect 28540 21020 28592 21072
rect 20536 20748 20588 20800
rect 20996 20748 21048 20800
rect 21916 20748 21968 20800
rect 22192 20748 22244 20800
rect 28356 20995 28408 21004
rect 28356 20961 28365 20995
rect 28365 20961 28399 20995
rect 28399 20961 28408 20995
rect 28356 20952 28408 20961
rect 24768 20816 24820 20868
rect 26056 20884 26108 20936
rect 26332 20884 26384 20936
rect 28264 20884 28316 20936
rect 28448 20927 28500 20936
rect 28448 20893 28457 20927
rect 28457 20893 28491 20927
rect 28491 20893 28500 20927
rect 28448 20884 28500 20893
rect 28816 20927 28868 20936
rect 28816 20893 28818 20927
rect 28818 20893 28868 20927
rect 28816 20884 28868 20893
rect 29000 20884 29052 20936
rect 29552 20884 29604 20936
rect 25688 20816 25740 20868
rect 28172 20859 28224 20868
rect 28172 20825 28181 20859
rect 28181 20825 28215 20859
rect 28215 20825 28224 20859
rect 28172 20816 28224 20825
rect 24308 20748 24360 20800
rect 25872 20748 25924 20800
rect 29644 20748 29696 20800
rect 4193 20646 4245 20698
rect 4257 20646 4309 20698
rect 4321 20646 4373 20698
rect 4385 20646 4437 20698
rect 4449 20646 4501 20698
rect 11783 20646 11835 20698
rect 11847 20646 11899 20698
rect 11911 20646 11963 20698
rect 11975 20646 12027 20698
rect 12039 20646 12091 20698
rect 19373 20646 19425 20698
rect 19437 20646 19489 20698
rect 19501 20646 19553 20698
rect 19565 20646 19617 20698
rect 19629 20646 19681 20698
rect 26963 20646 27015 20698
rect 27027 20646 27079 20698
rect 27091 20646 27143 20698
rect 27155 20646 27207 20698
rect 27219 20646 27271 20698
rect 2780 20408 2832 20460
rect 4528 20408 4580 20460
rect 4620 20451 4672 20460
rect 4620 20417 4629 20451
rect 4629 20417 4663 20451
rect 4663 20417 4672 20451
rect 4620 20408 4672 20417
rect 7288 20544 7340 20596
rect 7932 20587 7984 20596
rect 7932 20553 7941 20587
rect 7941 20553 7975 20587
rect 7975 20553 7984 20587
rect 7932 20544 7984 20553
rect 1216 20340 1268 20392
rect 1584 20383 1636 20392
rect 1584 20349 1593 20383
rect 1593 20349 1627 20383
rect 1627 20349 1636 20383
rect 1584 20340 1636 20349
rect 4712 20340 4764 20392
rect 6184 20340 6236 20392
rect 6644 20408 6696 20460
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 6828 20408 6880 20417
rect 10324 20544 10376 20596
rect 10508 20587 10560 20596
rect 10508 20553 10517 20587
rect 10517 20553 10551 20587
rect 10551 20553 10560 20587
rect 10508 20544 10560 20553
rect 8852 20408 8904 20460
rect 10232 20408 10284 20460
rect 1308 20247 1360 20256
rect 1308 20213 1323 20247
rect 1323 20213 1357 20247
rect 1357 20213 1360 20247
rect 1308 20204 1360 20213
rect 3608 20204 3660 20256
rect 8392 20272 8444 20324
rect 9128 20340 9180 20392
rect 12532 20544 12584 20596
rect 13176 20544 13228 20596
rect 13820 20476 13872 20528
rect 10968 20408 11020 20460
rect 11060 20408 11112 20460
rect 14280 20476 14332 20528
rect 19248 20544 19300 20596
rect 23020 20544 23072 20596
rect 14648 20408 14700 20460
rect 15200 20408 15252 20460
rect 23572 20476 23624 20528
rect 25320 20476 25372 20528
rect 26332 20519 26384 20528
rect 26332 20485 26341 20519
rect 26341 20485 26375 20519
rect 26375 20485 26384 20519
rect 26332 20476 26384 20485
rect 15936 20408 15988 20460
rect 18788 20408 18840 20460
rect 19708 20408 19760 20460
rect 11704 20340 11756 20392
rect 4252 20204 4304 20256
rect 6184 20204 6236 20256
rect 7564 20204 7616 20256
rect 9312 20204 9364 20256
rect 10600 20204 10652 20256
rect 11428 20204 11480 20256
rect 11796 20204 11848 20256
rect 12992 20315 13044 20324
rect 12992 20281 13001 20315
rect 13001 20281 13035 20315
rect 13035 20281 13044 20315
rect 12992 20272 13044 20281
rect 14280 20383 14332 20392
rect 14280 20349 14289 20383
rect 14289 20349 14323 20383
rect 14323 20349 14332 20383
rect 14280 20340 14332 20349
rect 12164 20204 12216 20256
rect 14832 20272 14884 20324
rect 15292 20272 15344 20324
rect 15936 20204 15988 20256
rect 16856 20204 16908 20256
rect 17500 20247 17552 20256
rect 17500 20213 17509 20247
rect 17509 20213 17543 20247
rect 17543 20213 17552 20247
rect 17500 20204 17552 20213
rect 17960 20315 18012 20324
rect 17960 20281 17969 20315
rect 17969 20281 18003 20315
rect 18003 20281 18012 20315
rect 17960 20272 18012 20281
rect 20720 20340 20772 20392
rect 19524 20272 19576 20324
rect 21272 20340 21324 20392
rect 25136 20340 25188 20392
rect 25412 20340 25464 20392
rect 28540 20408 28592 20460
rect 29184 20408 29236 20460
rect 25964 20340 26016 20392
rect 27344 20340 27396 20392
rect 29276 20340 29328 20392
rect 29460 20383 29512 20392
rect 29460 20349 29469 20383
rect 29469 20349 29503 20383
rect 29503 20349 29512 20383
rect 29460 20340 29512 20349
rect 29736 20408 29788 20460
rect 21548 20204 21600 20256
rect 23112 20272 23164 20324
rect 24124 20272 24176 20324
rect 22468 20204 22520 20256
rect 24860 20204 24912 20256
rect 28172 20204 28224 20256
rect 28816 20204 28868 20256
rect 30012 20272 30064 20324
rect 31392 20272 31444 20324
rect 29644 20204 29696 20256
rect 29828 20204 29880 20256
rect 7988 20102 8040 20154
rect 8052 20102 8104 20154
rect 8116 20102 8168 20154
rect 8180 20102 8232 20154
rect 8244 20102 8296 20154
rect 15578 20102 15630 20154
rect 15642 20102 15694 20154
rect 15706 20102 15758 20154
rect 15770 20102 15822 20154
rect 15834 20102 15886 20154
rect 23168 20102 23220 20154
rect 23232 20102 23284 20154
rect 23296 20102 23348 20154
rect 23360 20102 23412 20154
rect 23424 20102 23476 20154
rect 30758 20102 30810 20154
rect 30822 20102 30874 20154
rect 30886 20102 30938 20154
rect 30950 20102 31002 20154
rect 31014 20102 31066 20154
rect 1400 20000 1452 20052
rect 3424 20000 3476 20052
rect 4252 20000 4304 20052
rect 6000 19932 6052 19984
rect 848 19839 900 19848
rect 848 19805 857 19839
rect 857 19805 891 19839
rect 891 19805 900 19839
rect 848 19796 900 19805
rect 1584 19839 1636 19848
rect 1584 19805 1593 19839
rect 1593 19805 1627 19839
rect 1627 19805 1636 19839
rect 1584 19796 1636 19805
rect 5632 19907 5684 19916
rect 5632 19873 5641 19907
rect 5641 19873 5675 19907
rect 5675 19873 5684 19907
rect 5632 19864 5684 19873
rect 2964 19796 3016 19848
rect 3240 19796 3292 19848
rect 3608 19796 3660 19848
rect 3700 19796 3752 19848
rect 5264 19796 5316 19848
rect 5356 19796 5408 19848
rect 5908 19839 5960 19848
rect 5908 19805 5917 19839
rect 5917 19805 5951 19839
rect 5951 19805 5960 19839
rect 5908 19796 5960 19805
rect 6092 19796 6144 19848
rect 6276 19839 6328 19848
rect 6276 19805 6278 19839
rect 6278 19805 6328 19839
rect 6276 19796 6328 19805
rect 6644 19839 6696 19848
rect 6644 19805 6653 19839
rect 6653 19805 6687 19839
rect 6687 19805 6696 19839
rect 6644 19796 6696 19805
rect 8944 20043 8996 20052
rect 8944 20009 8959 20043
rect 8959 20009 8993 20043
rect 8993 20009 8996 20043
rect 8944 20000 8996 20009
rect 9220 20000 9272 20052
rect 11152 20000 11204 20052
rect 12256 20000 12308 20052
rect 12440 20000 12492 20052
rect 13544 20000 13596 20052
rect 15200 20000 15252 20052
rect 15292 20000 15344 20052
rect 8300 19864 8352 19916
rect 8392 19864 8444 19916
rect 11704 19932 11756 19984
rect 13728 19932 13780 19984
rect 16120 20000 16172 20052
rect 19800 20000 19852 20052
rect 20536 20043 20588 20052
rect 20536 20009 20545 20043
rect 20545 20009 20579 20043
rect 20579 20009 20588 20043
rect 20536 20000 20588 20009
rect 21088 20043 21140 20052
rect 21088 20009 21097 20043
rect 21097 20009 21131 20043
rect 21131 20009 21140 20043
rect 21088 20000 21140 20009
rect 11796 19864 11848 19916
rect 2872 19660 2924 19712
rect 5080 19703 5132 19712
rect 5080 19669 5089 19703
rect 5089 19669 5123 19703
rect 5123 19669 5132 19703
rect 5080 19660 5132 19669
rect 6828 19660 6880 19712
rect 8300 19703 8352 19712
rect 8300 19669 8309 19703
rect 8309 19669 8343 19703
rect 8343 19669 8352 19703
rect 8300 19660 8352 19669
rect 9220 19839 9272 19848
rect 9220 19805 9229 19839
rect 9229 19805 9263 19839
rect 9263 19805 9272 19839
rect 9220 19796 9272 19805
rect 10784 19660 10836 19712
rect 11980 19796 12032 19848
rect 12624 19839 12676 19848
rect 12624 19805 12636 19839
rect 12636 19805 12670 19839
rect 12670 19805 12676 19839
rect 12624 19796 12676 19805
rect 12808 19796 12860 19848
rect 14556 19864 14608 19916
rect 14832 19864 14884 19916
rect 14372 19839 14424 19848
rect 14372 19805 14381 19839
rect 14381 19805 14415 19839
rect 14415 19805 14424 19839
rect 14372 19796 14424 19805
rect 15568 19864 15620 19916
rect 16212 19932 16264 19984
rect 16396 19932 16448 19984
rect 21456 20000 21508 20052
rect 21548 20000 21600 20052
rect 23940 20000 23992 20052
rect 24124 20000 24176 20052
rect 25136 20000 25188 20052
rect 28816 20043 28868 20052
rect 28816 20009 28831 20043
rect 28831 20009 28865 20043
rect 28865 20009 28868 20043
rect 28816 20000 28868 20009
rect 17960 19864 18012 19916
rect 20628 19907 20680 19916
rect 20628 19873 20637 19907
rect 20637 19873 20671 19907
rect 20671 19873 20680 19907
rect 20628 19864 20680 19873
rect 20904 19907 20956 19916
rect 20904 19873 20913 19907
rect 20913 19873 20947 19907
rect 20947 19873 20956 19907
rect 20904 19864 20956 19873
rect 21548 19907 21600 19916
rect 21548 19873 21557 19907
rect 21557 19873 21591 19907
rect 21591 19873 21600 19907
rect 21548 19864 21600 19873
rect 16120 19796 16172 19848
rect 16856 19796 16908 19848
rect 17224 19839 17276 19848
rect 17224 19805 17233 19839
rect 17233 19805 17267 19839
rect 17267 19805 17276 19839
rect 17224 19796 17276 19805
rect 18696 19839 18748 19848
rect 18696 19805 18705 19839
rect 18705 19805 18739 19839
rect 18739 19805 18748 19839
rect 18696 19796 18748 19805
rect 20720 19796 20772 19848
rect 12808 19660 12860 19712
rect 13084 19660 13136 19712
rect 15292 19660 15344 19712
rect 16304 19728 16356 19780
rect 19892 19728 19944 19780
rect 22192 19907 22244 19916
rect 22192 19873 22201 19907
rect 22201 19873 22235 19907
rect 22235 19873 22244 19907
rect 22192 19864 22244 19873
rect 22468 19839 22520 19848
rect 22468 19805 22477 19839
rect 22477 19805 22511 19839
rect 22511 19805 22520 19839
rect 27344 19864 27396 19916
rect 28448 19864 28500 19916
rect 22468 19796 22520 19805
rect 24400 19839 24452 19848
rect 24400 19805 24409 19839
rect 24409 19805 24443 19839
rect 24443 19805 24452 19839
rect 24400 19796 24452 19805
rect 24676 19839 24728 19848
rect 24676 19805 24685 19839
rect 24685 19805 24719 19839
rect 24719 19805 24728 19839
rect 24676 19796 24728 19805
rect 26884 19796 26936 19848
rect 27528 19796 27580 19848
rect 28908 19796 28960 19848
rect 29092 19839 29144 19848
rect 29092 19805 29101 19839
rect 29101 19805 29135 19839
rect 29135 19805 29144 19839
rect 29092 19796 29144 19805
rect 21364 19703 21416 19712
rect 21364 19669 21373 19703
rect 21373 19669 21407 19703
rect 21407 19669 21416 19703
rect 21364 19660 21416 19669
rect 27988 19703 28040 19712
rect 27988 19669 27997 19703
rect 27997 19669 28031 19703
rect 28031 19669 28040 19703
rect 27988 19660 28040 19669
rect 28080 19660 28132 19712
rect 30472 19660 30524 19712
rect 4193 19558 4245 19610
rect 4257 19558 4309 19610
rect 4321 19558 4373 19610
rect 4385 19558 4437 19610
rect 4449 19558 4501 19610
rect 11783 19558 11835 19610
rect 11847 19558 11899 19610
rect 11911 19558 11963 19610
rect 11975 19558 12027 19610
rect 12039 19558 12091 19610
rect 19373 19558 19425 19610
rect 19437 19558 19489 19610
rect 19501 19558 19553 19610
rect 19565 19558 19617 19610
rect 19629 19558 19681 19610
rect 26963 19558 27015 19610
rect 27027 19558 27079 19610
rect 27091 19558 27143 19610
rect 27155 19558 27207 19610
rect 27219 19558 27271 19610
rect 5080 19456 5132 19508
rect 6092 19456 6144 19508
rect 848 19320 900 19372
rect 2044 19320 2096 19372
rect 2964 19320 3016 19372
rect 3240 19363 3292 19372
rect 3240 19329 3249 19363
rect 3249 19329 3283 19363
rect 3283 19329 3292 19363
rect 3240 19320 3292 19329
rect 8300 19456 8352 19508
rect 1952 19252 2004 19304
rect 3148 19252 3200 19304
rect 3884 19252 3936 19304
rect 3976 19295 4028 19304
rect 3976 19261 3985 19295
rect 3985 19261 4019 19295
rect 4019 19261 4028 19295
rect 3976 19252 4028 19261
rect 4252 19252 4304 19304
rect 5356 19295 5408 19304
rect 5356 19261 5365 19295
rect 5365 19261 5399 19295
rect 5399 19261 5408 19295
rect 5356 19252 5408 19261
rect 6092 19320 6144 19372
rect 7656 19320 7708 19372
rect 4712 19184 4764 19236
rect 6644 19252 6696 19304
rect 7380 19252 7432 19304
rect 8392 19295 8444 19304
rect 8392 19261 8401 19295
rect 8401 19261 8435 19295
rect 8435 19261 8444 19295
rect 8392 19252 8444 19261
rect 8576 19320 8628 19372
rect 8944 19320 8996 19372
rect 9496 19320 9548 19372
rect 9588 19252 9640 19304
rect 10232 19499 10284 19508
rect 10232 19465 10241 19499
rect 10241 19465 10275 19499
rect 10275 19465 10284 19499
rect 10232 19456 10284 19465
rect 11244 19456 11296 19508
rect 11980 19456 12032 19508
rect 12348 19456 12400 19508
rect 12992 19456 13044 19508
rect 14464 19456 14516 19508
rect 18052 19499 18104 19508
rect 18052 19465 18061 19499
rect 18061 19465 18095 19499
rect 18095 19465 18104 19499
rect 18052 19456 18104 19465
rect 22468 19456 22520 19508
rect 23020 19456 23072 19508
rect 12164 19320 12216 19372
rect 14372 19320 14424 19372
rect 11060 19252 11112 19304
rect 1400 19159 1452 19168
rect 1400 19125 1415 19159
rect 1415 19125 1449 19159
rect 1449 19125 1452 19159
rect 1400 19116 1452 19125
rect 5172 19116 5224 19168
rect 6276 19116 6328 19168
rect 8484 19184 8536 19236
rect 10232 19184 10284 19236
rect 10876 19184 10928 19236
rect 11888 19252 11940 19304
rect 13084 19252 13136 19304
rect 13176 19252 13228 19304
rect 13544 19295 13596 19304
rect 13544 19261 13553 19295
rect 13553 19261 13587 19295
rect 13587 19261 13596 19295
rect 13544 19252 13596 19261
rect 14280 19295 14332 19304
rect 14280 19261 14289 19295
rect 14289 19261 14323 19295
rect 14323 19261 14332 19295
rect 14280 19252 14332 19261
rect 15936 19363 15988 19372
rect 15936 19329 15945 19363
rect 15945 19329 15979 19363
rect 15979 19329 15988 19363
rect 15936 19320 15988 19329
rect 22008 19320 22060 19372
rect 26424 19456 26476 19508
rect 16028 19252 16080 19304
rect 16212 19295 16264 19304
rect 16212 19261 16221 19295
rect 16221 19261 16255 19295
rect 16255 19261 16264 19295
rect 16212 19252 16264 19261
rect 16856 19252 16908 19304
rect 15108 19184 15160 19236
rect 8760 19116 8812 19168
rect 8852 19159 8904 19168
rect 8852 19125 8867 19159
rect 8867 19125 8901 19159
rect 8901 19125 8904 19159
rect 8852 19116 8904 19125
rect 9036 19116 9088 19168
rect 12348 19116 12400 19168
rect 12440 19116 12492 19168
rect 14188 19116 14240 19168
rect 17776 19227 17828 19236
rect 17776 19193 17785 19227
rect 17785 19193 17819 19227
rect 17819 19193 17828 19227
rect 17776 19184 17828 19193
rect 18236 19295 18288 19304
rect 18236 19261 18245 19295
rect 18245 19261 18279 19295
rect 18279 19261 18288 19295
rect 18236 19252 18288 19261
rect 18328 19252 18380 19304
rect 21180 19252 21232 19304
rect 21824 19252 21876 19304
rect 21364 19184 21416 19236
rect 18328 19159 18380 19168
rect 18328 19125 18337 19159
rect 18337 19125 18371 19159
rect 18371 19125 18380 19159
rect 18328 19116 18380 19125
rect 20076 19159 20128 19168
rect 20076 19125 20085 19159
rect 20085 19125 20119 19159
rect 20119 19125 20128 19159
rect 20076 19116 20128 19125
rect 20812 19159 20864 19168
rect 20812 19125 20821 19159
rect 20821 19125 20855 19159
rect 20855 19125 20864 19159
rect 20812 19116 20864 19125
rect 21088 19159 21140 19168
rect 21088 19125 21097 19159
rect 21097 19125 21131 19159
rect 21131 19125 21140 19159
rect 21088 19116 21140 19125
rect 22192 19116 22244 19168
rect 23572 19159 23624 19168
rect 23572 19125 23581 19159
rect 23581 19125 23615 19159
rect 23615 19125 23624 19159
rect 23572 19116 23624 19125
rect 23756 19252 23808 19304
rect 23848 19252 23900 19304
rect 24308 19295 24360 19304
rect 24308 19261 24317 19295
rect 24317 19261 24351 19295
rect 24351 19261 24360 19295
rect 24308 19252 24360 19261
rect 24584 19252 24636 19304
rect 23756 19116 23808 19168
rect 24124 19184 24176 19236
rect 25688 19252 25740 19304
rect 26056 19252 26108 19304
rect 26884 19295 26936 19304
rect 26884 19261 26893 19295
rect 26893 19261 26927 19295
rect 26927 19261 26936 19295
rect 26884 19252 26936 19261
rect 26240 19184 26292 19236
rect 28724 19295 28776 19304
rect 28724 19261 28733 19295
rect 28733 19261 28767 19295
rect 28767 19261 28776 19295
rect 28724 19252 28776 19261
rect 29184 19252 29236 19304
rect 30564 19295 30616 19304
rect 30564 19261 30573 19295
rect 30573 19261 30607 19295
rect 30607 19261 30616 19295
rect 30564 19252 30616 19261
rect 29460 19184 29512 19236
rect 29644 19184 29696 19236
rect 25136 19159 25188 19168
rect 25136 19125 25151 19159
rect 25151 19125 25185 19159
rect 25185 19125 25188 19159
rect 25136 19116 25188 19125
rect 26516 19159 26568 19168
rect 26516 19125 26525 19159
rect 26525 19125 26559 19159
rect 26559 19125 26568 19159
rect 26516 19116 26568 19125
rect 26700 19116 26752 19168
rect 28632 19116 28684 19168
rect 30104 19159 30156 19168
rect 30104 19125 30113 19159
rect 30113 19125 30147 19159
rect 30147 19125 30156 19159
rect 30104 19116 30156 19125
rect 30196 19116 30248 19168
rect 30380 19159 30432 19168
rect 30380 19125 30389 19159
rect 30389 19125 30423 19159
rect 30423 19125 30432 19159
rect 30380 19116 30432 19125
rect 7988 19014 8040 19066
rect 8052 19014 8104 19066
rect 8116 19014 8168 19066
rect 8180 19014 8232 19066
rect 8244 19014 8296 19066
rect 15578 19014 15630 19066
rect 15642 19014 15694 19066
rect 15706 19014 15758 19066
rect 15770 19014 15822 19066
rect 15834 19014 15886 19066
rect 23168 19014 23220 19066
rect 23232 19014 23284 19066
rect 23296 19014 23348 19066
rect 23360 19014 23412 19066
rect 23424 19014 23476 19066
rect 30758 19014 30810 19066
rect 30822 19014 30874 19066
rect 30886 19014 30938 19066
rect 30950 19014 31002 19066
rect 31014 19014 31066 19066
rect 1216 18844 1268 18896
rect 1308 18844 1360 18896
rect 4252 18955 4304 18964
rect 4252 18921 4261 18955
rect 4261 18921 4295 18955
rect 4295 18921 4304 18955
rect 4252 18912 4304 18921
rect 1032 18819 1084 18828
rect 1032 18785 1041 18819
rect 1041 18785 1075 18819
rect 1075 18785 1084 18819
rect 1032 18776 1084 18785
rect 1124 18819 1176 18828
rect 1124 18785 1133 18819
rect 1133 18785 1167 18819
rect 1167 18785 1176 18819
rect 1124 18776 1176 18785
rect 4620 18844 4672 18896
rect 4712 18887 4764 18896
rect 4712 18853 4721 18887
rect 4721 18853 4755 18887
rect 4755 18853 4764 18887
rect 4712 18844 4764 18853
rect 6276 18912 6328 18964
rect 9312 18912 9364 18964
rect 7656 18844 7708 18896
rect 1584 18708 1636 18760
rect 3516 18776 3568 18828
rect 3792 18776 3844 18828
rect 5356 18776 5408 18828
rect 2412 18751 2464 18760
rect 2412 18717 2421 18751
rect 2421 18717 2455 18751
rect 2455 18717 2464 18751
rect 2412 18708 2464 18717
rect 2964 18708 3016 18760
rect 5540 18708 5592 18760
rect 848 18640 900 18692
rect 6276 18751 6328 18760
rect 6276 18717 6278 18751
rect 6278 18717 6328 18751
rect 3884 18572 3936 18624
rect 4068 18572 4120 18624
rect 6276 18708 6328 18717
rect 6368 18751 6420 18760
rect 6368 18717 6380 18751
rect 6380 18717 6414 18751
rect 6414 18717 6420 18751
rect 6368 18708 6420 18717
rect 7748 18776 7800 18828
rect 8760 18844 8812 18896
rect 13176 18912 13228 18964
rect 13452 18912 13504 18964
rect 14188 18912 14240 18964
rect 15292 18912 15344 18964
rect 16212 18912 16264 18964
rect 18052 18912 18104 18964
rect 8300 18776 8352 18828
rect 8944 18776 8996 18828
rect 8392 18708 8444 18760
rect 8484 18708 8536 18760
rect 9036 18708 9088 18760
rect 10508 18776 10560 18828
rect 10876 18708 10928 18760
rect 11152 18819 11204 18828
rect 11152 18785 11161 18819
rect 11161 18785 11195 18819
rect 11195 18785 11204 18819
rect 11152 18776 11204 18785
rect 11244 18776 11296 18828
rect 11428 18708 11480 18760
rect 11704 18708 11756 18760
rect 12164 18751 12216 18760
rect 12164 18717 12166 18751
rect 12166 18717 12216 18751
rect 12164 18708 12216 18717
rect 14188 18819 14240 18828
rect 14188 18785 14197 18819
rect 14197 18785 14231 18819
rect 14231 18785 14240 18819
rect 14188 18776 14240 18785
rect 14648 18776 14700 18828
rect 16028 18776 16080 18828
rect 19984 18844 20036 18896
rect 22192 18912 22244 18964
rect 23480 18912 23532 18964
rect 23848 18912 23900 18964
rect 24400 18912 24452 18964
rect 24492 18912 24544 18964
rect 25688 18912 25740 18964
rect 26792 18912 26844 18964
rect 30380 18912 30432 18964
rect 30472 18955 30524 18964
rect 30472 18921 30481 18955
rect 30481 18921 30515 18955
rect 30515 18921 30524 18955
rect 30472 18912 30524 18921
rect 12532 18751 12584 18760
rect 12532 18717 12541 18751
rect 12541 18717 12575 18751
rect 12575 18717 12584 18751
rect 12532 18708 12584 18717
rect 14464 18708 14516 18760
rect 16212 18751 16264 18760
rect 16212 18717 16221 18751
rect 16221 18717 16255 18751
rect 16255 18717 16264 18751
rect 16212 18708 16264 18717
rect 16304 18708 16356 18760
rect 16856 18708 16908 18760
rect 17500 18776 17552 18828
rect 18144 18708 18196 18760
rect 18696 18751 18748 18760
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 7564 18640 7616 18692
rect 6092 18572 6144 18624
rect 8208 18572 8260 18624
rect 10784 18640 10836 18692
rect 15384 18640 15436 18692
rect 21824 18776 21876 18828
rect 22468 18708 22520 18760
rect 22652 18751 22704 18760
rect 22652 18717 22661 18751
rect 22661 18717 22695 18751
rect 22695 18717 22704 18751
rect 22652 18708 22704 18717
rect 24400 18776 24452 18828
rect 24676 18708 24728 18760
rect 26332 18708 26384 18760
rect 27068 18708 27120 18760
rect 9772 18572 9824 18624
rect 11060 18572 11112 18624
rect 12992 18572 13044 18624
rect 14556 18572 14608 18624
rect 19800 18572 19852 18624
rect 20260 18572 20312 18624
rect 21732 18572 21784 18624
rect 26148 18640 26200 18692
rect 22284 18572 22336 18624
rect 23480 18572 23532 18624
rect 24400 18572 24452 18624
rect 24492 18572 24544 18624
rect 27068 18572 27120 18624
rect 27620 18572 27672 18624
rect 27804 18572 27856 18624
rect 28816 18776 28868 18828
rect 29184 18776 29236 18828
rect 28632 18640 28684 18692
rect 30196 18683 30248 18692
rect 30196 18649 30205 18683
rect 30205 18649 30239 18683
rect 30239 18649 30248 18683
rect 30196 18640 30248 18649
rect 30380 18572 30432 18624
rect 4193 18470 4245 18522
rect 4257 18470 4309 18522
rect 4321 18470 4373 18522
rect 4385 18470 4437 18522
rect 4449 18470 4501 18522
rect 11783 18470 11835 18522
rect 11847 18470 11899 18522
rect 11911 18470 11963 18522
rect 11975 18470 12027 18522
rect 12039 18470 12091 18522
rect 19373 18470 19425 18522
rect 19437 18470 19489 18522
rect 19501 18470 19553 18522
rect 19565 18470 19617 18522
rect 19629 18470 19681 18522
rect 26963 18470 27015 18522
rect 27027 18470 27079 18522
rect 27091 18470 27143 18522
rect 27155 18470 27207 18522
rect 27219 18470 27271 18522
rect 2412 18368 2464 18420
rect 2964 18411 3016 18420
rect 2964 18377 2973 18411
rect 2973 18377 3007 18411
rect 3007 18377 3016 18411
rect 2964 18368 3016 18377
rect 3332 18368 3384 18420
rect 3516 18368 3568 18420
rect 5724 18368 5776 18420
rect 6368 18368 6420 18420
rect 6460 18368 6512 18420
rect 10692 18368 10744 18420
rect 12624 18411 12676 18420
rect 12624 18377 12633 18411
rect 12633 18377 12667 18411
rect 12667 18377 12676 18411
rect 12624 18368 12676 18377
rect 12256 18300 12308 18352
rect 17224 18411 17276 18420
rect 17224 18377 17233 18411
rect 17233 18377 17267 18411
rect 17267 18377 17276 18411
rect 17224 18368 17276 18377
rect 17500 18368 17552 18420
rect 22744 18368 22796 18420
rect 23480 18368 23532 18420
rect 23756 18368 23808 18420
rect 18236 18300 18288 18352
rect 848 18232 900 18284
rect 3148 18232 3200 18284
rect 2412 18164 2464 18216
rect 3240 18164 3292 18216
rect 4068 18232 4120 18284
rect 4252 18275 4304 18284
rect 4252 18241 4254 18275
rect 4254 18241 4304 18275
rect 4252 18232 4304 18241
rect 4344 18275 4396 18284
rect 4344 18241 4356 18275
rect 4356 18241 4390 18275
rect 4390 18241 4396 18275
rect 4344 18232 4396 18241
rect 5356 18232 5408 18284
rect 5632 18232 5684 18284
rect 8392 18232 8444 18284
rect 8576 18275 8628 18284
rect 8576 18241 8585 18275
rect 8585 18241 8619 18275
rect 8619 18241 8628 18275
rect 8576 18232 8628 18241
rect 8760 18232 8812 18284
rect 9128 18232 9180 18284
rect 3884 18207 3936 18216
rect 3884 18173 3893 18207
rect 3893 18173 3927 18207
rect 3927 18173 3936 18207
rect 3884 18164 3936 18173
rect 6092 18207 6144 18216
rect 6092 18173 6101 18207
rect 6101 18173 6135 18207
rect 6135 18173 6144 18207
rect 6092 18164 6144 18173
rect 6736 18164 6788 18216
rect 8484 18096 8536 18148
rect 1400 18071 1452 18080
rect 1400 18037 1415 18071
rect 1415 18037 1449 18071
rect 1449 18037 1452 18071
rect 1400 18028 1452 18037
rect 3332 18028 3384 18080
rect 6184 18028 6236 18080
rect 6460 18028 6512 18080
rect 6828 18028 6880 18080
rect 8392 18028 8444 18080
rect 11336 18232 11388 18284
rect 10784 18207 10836 18216
rect 10784 18173 10793 18207
rect 10793 18173 10827 18207
rect 10827 18173 10836 18207
rect 10784 18164 10836 18173
rect 13728 18232 13780 18284
rect 14004 18257 14056 18284
rect 14004 18232 14049 18257
rect 14049 18232 14056 18257
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 16028 18232 16080 18284
rect 16488 18232 16540 18284
rect 10232 18096 10284 18148
rect 13544 18207 13596 18216
rect 13544 18173 13553 18207
rect 13553 18173 13587 18207
rect 13587 18173 13596 18207
rect 13544 18164 13596 18173
rect 14648 18164 14700 18216
rect 16396 18164 16448 18216
rect 18052 18207 18104 18216
rect 18052 18173 18061 18207
rect 18061 18173 18095 18207
rect 18095 18173 18104 18207
rect 18052 18164 18104 18173
rect 18144 18164 18196 18216
rect 19892 18300 19944 18352
rect 20628 18232 20680 18284
rect 22836 18232 22888 18284
rect 24216 18232 24268 18284
rect 20260 18164 20312 18216
rect 8852 18028 8904 18080
rect 11428 18028 11480 18080
rect 13820 18028 13872 18080
rect 15108 18028 15160 18080
rect 15568 18071 15620 18080
rect 15568 18037 15577 18071
rect 15577 18037 15611 18071
rect 15611 18037 15620 18071
rect 15568 18028 15620 18037
rect 16212 18028 16264 18080
rect 19156 18096 19208 18148
rect 19892 18096 19944 18148
rect 20076 18096 20128 18148
rect 20996 18164 21048 18216
rect 22928 18164 22980 18216
rect 23664 18207 23716 18216
rect 23664 18173 23673 18207
rect 23673 18173 23707 18207
rect 23707 18173 23716 18207
rect 23664 18164 23716 18173
rect 24584 18300 24636 18352
rect 28264 18411 28316 18420
rect 28264 18377 28273 18411
rect 28273 18377 28307 18411
rect 28307 18377 28316 18411
rect 28264 18368 28316 18377
rect 24860 18232 24912 18284
rect 26884 18275 26936 18284
rect 26884 18241 26893 18275
rect 26893 18241 26927 18275
rect 26927 18241 26936 18275
rect 26884 18232 26936 18241
rect 27896 18232 27948 18284
rect 23940 18139 23992 18148
rect 23940 18105 23949 18139
rect 23949 18105 23983 18139
rect 23983 18105 23992 18139
rect 23940 18096 23992 18105
rect 25412 18207 25464 18216
rect 25412 18173 25421 18207
rect 25421 18173 25455 18207
rect 25455 18173 25464 18207
rect 25412 18164 25464 18173
rect 26608 18164 26660 18216
rect 28724 18164 28776 18216
rect 28632 18096 28684 18148
rect 29184 18164 29236 18216
rect 29368 18164 29420 18216
rect 30196 18164 30248 18216
rect 20352 18028 20404 18080
rect 21548 18028 21600 18080
rect 21732 18028 21784 18080
rect 23388 18028 23440 18080
rect 24308 18028 24360 18080
rect 24952 18028 25004 18080
rect 25136 18071 25188 18080
rect 25136 18037 25151 18071
rect 25151 18037 25185 18071
rect 25185 18037 25188 18071
rect 25136 18028 25188 18037
rect 26424 18028 26476 18080
rect 29644 18028 29696 18080
rect 29920 18028 29972 18080
rect 30288 18071 30340 18080
rect 30288 18037 30297 18071
rect 30297 18037 30331 18071
rect 30331 18037 30340 18071
rect 30288 18028 30340 18037
rect 7988 17926 8040 17978
rect 8052 17926 8104 17978
rect 8116 17926 8168 17978
rect 8180 17926 8232 17978
rect 8244 17926 8296 17978
rect 15578 17926 15630 17978
rect 15642 17926 15694 17978
rect 15706 17926 15758 17978
rect 15770 17926 15822 17978
rect 15834 17926 15886 17978
rect 23168 17926 23220 17978
rect 23232 17926 23284 17978
rect 23296 17926 23348 17978
rect 23360 17926 23412 17978
rect 23424 17926 23476 17978
rect 30758 17926 30810 17978
rect 30822 17926 30874 17978
rect 30886 17926 30938 17978
rect 30950 17926 31002 17978
rect 31014 17926 31066 17978
rect 1400 17867 1452 17876
rect 1400 17833 1415 17867
rect 1415 17833 1449 17867
rect 1449 17833 1452 17867
rect 1400 17824 1452 17833
rect 2780 17867 2832 17876
rect 2780 17833 2789 17867
rect 2789 17833 2823 17867
rect 2823 17833 2832 17867
rect 2780 17824 2832 17833
rect 3516 17824 3568 17876
rect 4252 17824 4304 17876
rect 4528 17824 4580 17876
rect 8392 17824 8444 17876
rect 5632 17799 5684 17808
rect 5632 17765 5641 17799
rect 5641 17765 5675 17799
rect 5675 17765 5684 17799
rect 5632 17756 5684 17765
rect 848 17688 900 17740
rect 2964 17688 3016 17740
rect 3608 17688 3660 17740
rect 4344 17688 4396 17740
rect 4896 17688 4948 17740
rect 3424 17620 3476 17672
rect 3884 17620 3936 17672
rect 4068 17620 4120 17672
rect 5172 17620 5224 17672
rect 3792 17484 3844 17536
rect 6276 17688 6328 17740
rect 6368 17731 6420 17740
rect 6368 17697 6377 17731
rect 6377 17697 6411 17731
rect 6411 17697 6420 17731
rect 6368 17688 6420 17697
rect 8760 17756 8812 17808
rect 12348 17824 12400 17876
rect 16028 17824 16080 17876
rect 16764 17824 16816 17876
rect 18328 17824 18380 17876
rect 8484 17688 8536 17740
rect 6184 17620 6236 17672
rect 6828 17663 6880 17672
rect 6828 17629 6830 17663
rect 6830 17629 6880 17663
rect 6828 17620 6880 17629
rect 7012 17620 7064 17672
rect 7196 17663 7248 17672
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 8576 17620 8628 17672
rect 8852 17620 8904 17672
rect 9036 17663 9088 17672
rect 9036 17629 9038 17663
rect 9038 17629 9088 17663
rect 9036 17620 9088 17629
rect 10140 17688 10192 17740
rect 10968 17688 11020 17740
rect 11152 17731 11204 17740
rect 11152 17697 11161 17731
rect 11161 17697 11195 17731
rect 11195 17697 11204 17731
rect 11152 17688 11204 17697
rect 16856 17756 16908 17808
rect 9220 17620 9272 17672
rect 13912 17688 13964 17740
rect 11520 17620 11572 17672
rect 11704 17620 11756 17672
rect 12164 17663 12216 17672
rect 12164 17629 12166 17663
rect 12166 17629 12216 17663
rect 12164 17620 12216 17629
rect 14832 17688 14884 17740
rect 16396 17688 16448 17740
rect 14280 17663 14332 17672
rect 9220 17484 9272 17536
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 14924 17620 14976 17672
rect 16488 17620 16540 17672
rect 17316 17663 17368 17672
rect 17316 17629 17318 17663
rect 17318 17629 17368 17663
rect 17316 17620 17368 17629
rect 17500 17620 17552 17672
rect 16764 17552 16816 17604
rect 13452 17484 13504 17536
rect 13636 17527 13688 17536
rect 13636 17493 13645 17527
rect 13645 17493 13679 17527
rect 13679 17493 13688 17527
rect 13636 17484 13688 17493
rect 13912 17484 13964 17536
rect 14464 17484 14516 17536
rect 16304 17484 16356 17536
rect 24124 17756 24176 17808
rect 18696 17688 18748 17740
rect 19892 17688 19944 17740
rect 20352 17688 20404 17740
rect 21088 17731 21140 17740
rect 21088 17697 21097 17731
rect 21097 17697 21131 17731
rect 21131 17697 21140 17731
rect 21088 17688 21140 17697
rect 21640 17731 21692 17740
rect 21640 17697 21642 17731
rect 21642 17697 21692 17731
rect 21640 17688 21692 17697
rect 22100 17688 22152 17740
rect 23756 17731 23808 17740
rect 23756 17697 23765 17731
rect 23765 17697 23799 17731
rect 23799 17697 23808 17731
rect 23756 17688 23808 17697
rect 24032 17731 24084 17740
rect 24032 17697 24041 17731
rect 24041 17697 24075 17731
rect 24075 17697 24084 17731
rect 24032 17688 24084 17697
rect 24400 17824 24452 17876
rect 25136 17824 25188 17876
rect 26516 17824 26568 17876
rect 27160 17824 27212 17876
rect 28724 17824 28776 17876
rect 30656 17824 30708 17876
rect 28632 17756 28684 17808
rect 28816 17756 28868 17808
rect 29368 17756 29420 17808
rect 26792 17731 26844 17740
rect 26792 17697 26794 17731
rect 26794 17697 26844 17731
rect 21732 17663 21784 17672
rect 21732 17629 21744 17663
rect 21744 17629 21778 17663
rect 21778 17629 21784 17663
rect 21732 17620 21784 17629
rect 18788 17527 18840 17536
rect 18788 17493 18797 17527
rect 18797 17493 18831 17527
rect 18831 17493 18840 17527
rect 18788 17484 18840 17493
rect 18972 17484 19024 17536
rect 20628 17484 20680 17536
rect 20720 17527 20772 17536
rect 20720 17493 20729 17527
rect 20729 17493 20763 17527
rect 20763 17493 20772 17527
rect 20720 17484 20772 17493
rect 20996 17484 21048 17536
rect 21088 17484 21140 17536
rect 23020 17552 23072 17604
rect 23112 17527 23164 17536
rect 23112 17493 23121 17527
rect 23121 17493 23155 17527
rect 23155 17493 23164 17527
rect 23112 17484 23164 17493
rect 24032 17552 24084 17604
rect 24492 17620 24544 17672
rect 24768 17620 24820 17672
rect 25964 17620 26016 17672
rect 26332 17620 26384 17672
rect 26792 17688 26844 17697
rect 27160 17731 27212 17740
rect 27160 17697 27169 17731
rect 27169 17697 27203 17731
rect 27203 17697 27212 17731
rect 27160 17688 27212 17697
rect 26884 17665 26936 17672
rect 26884 17631 26896 17665
rect 26896 17631 26930 17665
rect 26930 17631 26936 17665
rect 26884 17620 26936 17631
rect 29644 17620 29696 17672
rect 26332 17484 26384 17536
rect 28356 17484 28408 17536
rect 29920 17484 29972 17536
rect 30012 17484 30064 17536
rect 4193 17382 4245 17434
rect 4257 17382 4309 17434
rect 4321 17382 4373 17434
rect 4385 17382 4437 17434
rect 4449 17382 4501 17434
rect 11783 17382 11835 17434
rect 11847 17382 11899 17434
rect 11911 17382 11963 17434
rect 11975 17382 12027 17434
rect 12039 17382 12091 17434
rect 19373 17382 19425 17434
rect 19437 17382 19489 17434
rect 19501 17382 19553 17434
rect 19565 17382 19617 17434
rect 19629 17382 19681 17434
rect 26963 17382 27015 17434
rect 27027 17382 27079 17434
rect 27091 17382 27143 17434
rect 27155 17382 27207 17434
rect 27219 17382 27271 17434
rect 2872 17280 2924 17332
rect 3792 17280 3844 17332
rect 3884 17280 3936 17332
rect 3332 17144 3384 17196
rect 5448 17144 5500 17196
rect 1308 17076 1360 17128
rect 2136 17076 2188 17128
rect 3700 17076 3752 17128
rect 7196 17280 7248 17332
rect 8392 17255 8444 17264
rect 8392 17221 8401 17255
rect 8401 17221 8435 17255
rect 8435 17221 8444 17255
rect 8392 17212 8444 17221
rect 8576 17212 8628 17264
rect 10508 17323 10560 17332
rect 10508 17289 10517 17323
rect 10517 17289 10551 17323
rect 10551 17289 10560 17323
rect 10508 17280 10560 17289
rect 10876 17323 10928 17332
rect 10876 17289 10885 17323
rect 10885 17289 10919 17323
rect 10919 17289 10928 17323
rect 10876 17280 10928 17289
rect 6184 17076 6236 17128
rect 6460 17119 6512 17128
rect 6460 17085 6462 17119
rect 6462 17085 6512 17119
rect 6460 17076 6512 17085
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 8484 17076 8536 17128
rect 1400 16983 1452 16992
rect 1400 16949 1415 16983
rect 1415 16949 1449 16983
rect 1449 16949 1452 16983
rect 1400 16940 1452 16949
rect 5632 17008 5684 17060
rect 5816 17008 5868 17060
rect 9404 17187 9456 17196
rect 9404 17153 9413 17187
rect 9413 17153 9447 17187
rect 9447 17153 9456 17187
rect 9404 17144 9456 17153
rect 11520 17144 11572 17196
rect 13452 17144 13504 17196
rect 13912 17280 13964 17332
rect 14188 17212 14240 17264
rect 9680 17076 9732 17128
rect 10600 17076 10652 17128
rect 10876 17008 10928 17060
rect 14004 17076 14056 17128
rect 18972 17323 19024 17332
rect 18972 17289 18981 17323
rect 18981 17289 19015 17323
rect 19015 17289 19024 17323
rect 18972 17280 19024 17289
rect 21916 17280 21968 17332
rect 22008 17280 22060 17332
rect 19064 17212 19116 17264
rect 19524 17255 19576 17264
rect 19524 17221 19533 17255
rect 19533 17221 19567 17255
rect 19567 17221 19576 17255
rect 19524 17212 19576 17221
rect 19708 17212 19760 17264
rect 17868 17144 17920 17196
rect 18696 17187 18748 17196
rect 18696 17153 18705 17187
rect 18705 17153 18739 17187
rect 18739 17153 18748 17187
rect 18696 17144 18748 17153
rect 14832 17076 14884 17128
rect 15936 17076 15988 17128
rect 16488 17076 16540 17128
rect 16764 17119 16816 17128
rect 16764 17085 16766 17119
rect 16766 17085 16816 17119
rect 16764 17076 16816 17085
rect 17040 17076 17092 17128
rect 18144 17076 18196 17128
rect 13176 17008 13228 17060
rect 13912 17008 13964 17060
rect 19340 17076 19392 17128
rect 23020 17212 23072 17264
rect 23204 17280 23256 17332
rect 23572 17144 23624 17196
rect 4528 16940 4580 16992
rect 6184 16940 6236 16992
rect 9036 16940 9088 16992
rect 12072 16940 12124 16992
rect 13084 16983 13136 16992
rect 13084 16949 13093 16983
rect 13093 16949 13127 16983
rect 13127 16949 13136 16983
rect 13084 16940 13136 16949
rect 14188 16940 14240 16992
rect 14832 16940 14884 16992
rect 16672 16940 16724 16992
rect 17040 16940 17092 16992
rect 18236 16983 18288 16992
rect 18236 16949 18245 16983
rect 18245 16949 18279 16983
rect 18279 16949 18288 16983
rect 18236 16940 18288 16949
rect 20260 17076 20312 17128
rect 20352 17119 20404 17128
rect 20352 17085 20361 17119
rect 20361 17085 20395 17119
rect 20395 17085 20404 17119
rect 20352 17076 20404 17085
rect 19892 17008 19944 17060
rect 19984 17008 20036 17060
rect 20628 17076 20680 17128
rect 20996 17076 21048 17128
rect 23112 17076 23164 17128
rect 22652 17051 22704 17060
rect 22652 17017 22661 17051
rect 22661 17017 22695 17051
rect 22695 17017 22704 17051
rect 22652 17008 22704 17017
rect 23020 17008 23072 17060
rect 23848 17119 23900 17128
rect 23848 17085 23857 17119
rect 23857 17085 23891 17119
rect 23891 17085 23900 17119
rect 23848 17076 23900 17085
rect 24216 17076 24268 17128
rect 25412 17280 25464 17332
rect 26240 17280 26292 17332
rect 27252 17280 27304 17332
rect 28724 17280 28776 17332
rect 29368 17280 29420 17332
rect 30564 17280 30616 17332
rect 27528 17144 27580 17196
rect 28632 17212 28684 17264
rect 25780 17119 25832 17128
rect 25780 17085 25789 17119
rect 25789 17085 25823 17119
rect 25823 17085 25832 17119
rect 25780 17076 25832 17085
rect 25964 17076 26016 17128
rect 27344 17076 27396 17128
rect 30288 17144 30340 17196
rect 28724 17076 28776 17128
rect 29644 17119 29696 17128
rect 29644 17085 29653 17119
rect 29653 17085 29687 17119
rect 29687 17085 29696 17119
rect 29644 17076 29696 17085
rect 22192 16983 22244 16992
rect 22192 16949 22201 16983
rect 22201 16949 22235 16983
rect 22235 16949 22244 16983
rect 22192 16940 22244 16949
rect 23848 16940 23900 16992
rect 25136 17008 25188 17060
rect 28264 17008 28316 17060
rect 28632 17008 28684 17060
rect 30104 17051 30156 17060
rect 26148 16940 26200 16992
rect 26700 16940 26752 16992
rect 27252 16940 27304 16992
rect 27712 16983 27764 16992
rect 27712 16949 27721 16983
rect 27721 16949 27755 16983
rect 27755 16949 27764 16983
rect 27712 16940 27764 16949
rect 28724 16983 28776 16992
rect 28724 16949 28733 16983
rect 28733 16949 28767 16983
rect 28767 16949 28776 16983
rect 28724 16940 28776 16949
rect 29368 16940 29420 16992
rect 30104 17017 30113 17051
rect 30113 17017 30147 17051
rect 30147 17017 30156 17051
rect 30104 17008 30156 17017
rect 29920 16983 29972 16992
rect 29920 16949 29929 16983
rect 29929 16949 29963 16983
rect 29963 16949 29972 16983
rect 29920 16940 29972 16949
rect 7988 16838 8040 16890
rect 8052 16838 8104 16890
rect 8116 16838 8168 16890
rect 8180 16838 8232 16890
rect 8244 16838 8296 16890
rect 15578 16838 15630 16890
rect 15642 16838 15694 16890
rect 15706 16838 15758 16890
rect 15770 16838 15822 16890
rect 15834 16838 15886 16890
rect 23168 16838 23220 16890
rect 23232 16838 23284 16890
rect 23296 16838 23348 16890
rect 23360 16838 23412 16890
rect 23424 16838 23476 16890
rect 30758 16838 30810 16890
rect 30822 16838 30874 16890
rect 30886 16838 30938 16890
rect 30950 16838 31002 16890
rect 31014 16838 31066 16890
rect 2872 16736 2924 16788
rect 940 16643 992 16652
rect 940 16609 949 16643
rect 949 16609 983 16643
rect 983 16609 992 16643
rect 940 16600 992 16609
rect 4160 16736 4212 16788
rect 4712 16736 4764 16788
rect 4896 16736 4948 16788
rect 6920 16736 6972 16788
rect 7012 16736 7064 16788
rect 8576 16736 8628 16788
rect 10968 16736 11020 16788
rect 12348 16736 12400 16788
rect 12808 16736 12860 16788
rect 10048 16668 10100 16720
rect 1676 16575 1728 16584
rect 1676 16541 1685 16575
rect 1685 16541 1719 16575
rect 1719 16541 1728 16575
rect 1676 16532 1728 16541
rect 2780 16532 2832 16584
rect 3240 16532 3292 16584
rect 3516 16575 3568 16584
rect 3516 16541 3525 16575
rect 3525 16541 3559 16575
rect 3559 16541 3568 16575
rect 3516 16532 3568 16541
rect 3884 16575 3936 16584
rect 3884 16541 3886 16575
rect 3886 16541 3936 16575
rect 3884 16532 3936 16541
rect 5724 16600 5776 16652
rect 8668 16600 8720 16652
rect 9312 16643 9364 16652
rect 9312 16609 9321 16643
rect 9321 16609 9355 16643
rect 9355 16609 9364 16643
rect 9312 16600 9364 16609
rect 11428 16668 11480 16720
rect 5816 16575 5868 16584
rect 5816 16541 5825 16575
rect 5825 16541 5859 16575
rect 5859 16541 5868 16575
rect 5816 16532 5868 16541
rect 6184 16575 6236 16584
rect 6184 16541 6186 16575
rect 6186 16541 6236 16575
rect 6184 16532 6236 16541
rect 6276 16577 6328 16584
rect 6276 16543 6288 16577
rect 6288 16543 6322 16577
rect 6322 16543 6328 16577
rect 6276 16532 6328 16543
rect 6644 16532 6696 16584
rect 8944 16575 8996 16584
rect 2412 16464 2464 16516
rect 2320 16396 2372 16448
rect 7288 16396 7340 16448
rect 8944 16541 8946 16575
rect 8946 16541 8996 16575
rect 8944 16532 8996 16541
rect 9772 16532 9824 16584
rect 11152 16532 11204 16584
rect 11520 16600 11572 16652
rect 16396 16779 16448 16788
rect 16396 16745 16405 16779
rect 16405 16745 16439 16779
rect 16439 16745 16448 16779
rect 16396 16736 16448 16745
rect 16580 16736 16632 16788
rect 11980 16575 12032 16584
rect 11980 16541 11982 16575
rect 11982 16541 12032 16575
rect 11980 16532 12032 16541
rect 14464 16600 14516 16652
rect 12348 16575 12400 16584
rect 12348 16541 12357 16575
rect 12357 16541 12391 16575
rect 12391 16541 12400 16575
rect 12348 16532 12400 16541
rect 14004 16532 14056 16584
rect 14188 16575 14240 16584
rect 14188 16541 14190 16575
rect 14190 16541 14240 16575
rect 14188 16532 14240 16541
rect 16304 16643 16356 16652
rect 16304 16609 16313 16643
rect 16313 16609 16347 16643
rect 16347 16609 16356 16643
rect 16304 16600 16356 16609
rect 17316 16736 17368 16788
rect 18144 16736 18196 16788
rect 16856 16643 16908 16652
rect 16856 16609 16865 16643
rect 16865 16609 16899 16643
rect 16899 16609 16908 16643
rect 16856 16600 16908 16609
rect 19064 16711 19116 16720
rect 19064 16677 19073 16711
rect 19073 16677 19107 16711
rect 19107 16677 19116 16711
rect 19064 16668 19116 16677
rect 24124 16736 24176 16788
rect 10048 16464 10100 16516
rect 11428 16464 11480 16516
rect 9036 16396 9088 16448
rect 9496 16396 9548 16448
rect 13820 16396 13872 16448
rect 14464 16396 14516 16448
rect 16120 16439 16172 16448
rect 16120 16405 16129 16439
rect 16129 16405 16163 16439
rect 16163 16405 16172 16439
rect 16120 16396 16172 16405
rect 17224 16532 17276 16584
rect 20628 16668 20680 16720
rect 26424 16736 26476 16788
rect 19340 16643 19392 16652
rect 19340 16609 19349 16643
rect 19349 16609 19383 16643
rect 19383 16609 19392 16643
rect 19340 16600 19392 16609
rect 19800 16600 19852 16652
rect 21088 16600 21140 16652
rect 17132 16396 17184 16448
rect 20352 16532 20404 16584
rect 21640 16575 21692 16584
rect 21640 16541 21642 16575
rect 21642 16541 21692 16575
rect 21640 16532 21692 16541
rect 21916 16532 21968 16584
rect 22652 16532 22704 16584
rect 23940 16643 23992 16652
rect 23940 16609 23949 16643
rect 23949 16609 23983 16643
rect 23983 16609 23992 16643
rect 23940 16600 23992 16609
rect 24032 16600 24084 16652
rect 19708 16396 19760 16448
rect 20076 16396 20128 16448
rect 20996 16439 21048 16448
rect 20996 16405 21005 16439
rect 21005 16405 21039 16439
rect 21039 16405 21048 16439
rect 20996 16396 21048 16405
rect 21272 16396 21324 16448
rect 24308 16532 24360 16584
rect 24584 16577 24636 16584
rect 24584 16543 24596 16577
rect 24596 16543 24630 16577
rect 24630 16543 24636 16577
rect 24952 16600 25004 16652
rect 25872 16600 25924 16652
rect 28816 16668 28868 16720
rect 29184 16779 29236 16788
rect 29184 16745 29193 16779
rect 29193 16745 29227 16779
rect 29227 16745 29236 16779
rect 29184 16736 29236 16745
rect 29920 16736 29972 16788
rect 30380 16779 30432 16788
rect 30380 16745 30389 16779
rect 30389 16745 30423 16779
rect 30423 16745 30432 16779
rect 30380 16736 30432 16745
rect 29644 16668 29696 16720
rect 27436 16600 27488 16652
rect 24584 16532 24636 16543
rect 27896 16532 27948 16584
rect 28080 16643 28132 16652
rect 28080 16609 28089 16643
rect 28089 16609 28123 16643
rect 28123 16609 28132 16643
rect 28080 16600 28132 16609
rect 28172 16600 28224 16652
rect 30288 16600 30340 16652
rect 30380 16600 30432 16652
rect 31116 16600 31168 16652
rect 22836 16464 22888 16516
rect 22744 16396 22796 16448
rect 23572 16396 23624 16448
rect 23756 16464 23808 16516
rect 23940 16464 23992 16516
rect 26056 16396 26108 16448
rect 26332 16396 26384 16448
rect 26792 16439 26844 16448
rect 26792 16405 26801 16439
rect 26801 16405 26835 16439
rect 26835 16405 26844 16439
rect 26792 16396 26844 16405
rect 27160 16439 27212 16448
rect 27160 16405 27169 16439
rect 27169 16405 27203 16439
rect 27203 16405 27212 16439
rect 27160 16396 27212 16405
rect 4193 16294 4245 16346
rect 4257 16294 4309 16346
rect 4321 16294 4373 16346
rect 4385 16294 4437 16346
rect 4449 16294 4501 16346
rect 11783 16294 11835 16346
rect 11847 16294 11899 16346
rect 11911 16294 11963 16346
rect 11975 16294 12027 16346
rect 12039 16294 12091 16346
rect 19373 16294 19425 16346
rect 19437 16294 19489 16346
rect 19501 16294 19553 16346
rect 19565 16294 19617 16346
rect 19629 16294 19681 16346
rect 26963 16294 27015 16346
rect 27027 16294 27079 16346
rect 27091 16294 27143 16346
rect 27155 16294 27207 16346
rect 27219 16294 27271 16346
rect 2044 16192 2096 16244
rect 4252 16192 4304 16244
rect 4620 16192 4672 16244
rect 4712 16192 4764 16244
rect 1308 15988 1360 16040
rect 2504 15988 2556 16040
rect 3332 16031 3384 16040
rect 3332 15997 3341 16031
rect 3341 15997 3375 16031
rect 3375 15997 3384 16031
rect 3332 15988 3384 15997
rect 6460 16056 6512 16108
rect 4436 15988 4488 16040
rect 4528 16031 4580 16040
rect 4528 15997 4537 16031
rect 4537 15997 4571 16031
rect 4571 15997 4580 16031
rect 4528 15988 4580 15997
rect 6092 16031 6144 16040
rect 6092 15997 6101 16031
rect 6101 15997 6135 16031
rect 6135 15997 6144 16031
rect 6092 15988 6144 15997
rect 9772 16192 9824 16244
rect 13084 16192 13136 16244
rect 14372 16192 14424 16244
rect 14832 16192 14884 16244
rect 10968 16167 11020 16176
rect 10968 16133 10977 16167
rect 10977 16133 11011 16167
rect 11011 16133 11020 16167
rect 10968 16124 11020 16133
rect 11060 16124 11112 16176
rect 5264 15920 5316 15972
rect 8668 16031 8720 16040
rect 8668 15997 8677 16031
rect 8677 15997 8711 16031
rect 8711 15997 8720 16031
rect 8668 15988 8720 15997
rect 8944 15988 8996 16040
rect 9864 15988 9916 16040
rect 11520 16056 11572 16108
rect 11704 16097 11756 16108
rect 11704 16063 11716 16097
rect 11716 16063 11750 16097
rect 11750 16063 11756 16097
rect 11704 16056 11756 16063
rect 1400 15895 1452 15904
rect 1400 15861 1415 15895
rect 1415 15861 1449 15895
rect 1449 15861 1452 15895
rect 1400 15852 1452 15861
rect 3608 15895 3660 15904
rect 3608 15861 3617 15895
rect 3617 15861 3651 15895
rect 3651 15861 3660 15895
rect 3608 15852 3660 15861
rect 3884 15852 3936 15904
rect 6460 15852 6512 15904
rect 8392 15895 8444 15904
rect 8392 15861 8401 15895
rect 8401 15861 8435 15895
rect 8435 15861 8444 15895
rect 8392 15852 8444 15861
rect 9036 15852 9088 15904
rect 10508 15895 10560 15904
rect 10508 15861 10517 15895
rect 10517 15861 10551 15895
rect 10551 15861 10560 15895
rect 10508 15852 10560 15861
rect 12716 15988 12768 16040
rect 14556 16056 14608 16108
rect 18236 16192 18288 16244
rect 16120 16056 16172 16108
rect 16488 15988 16540 16040
rect 17868 16056 17920 16108
rect 19800 16192 19852 16244
rect 20352 16192 20404 16244
rect 26608 16192 26660 16244
rect 26792 16192 26844 16244
rect 27712 16192 27764 16244
rect 17224 15988 17276 16040
rect 19984 16099 20036 16108
rect 19984 16065 19986 16099
rect 19986 16065 20036 16099
rect 19984 16056 20036 16065
rect 19432 16031 19484 16040
rect 19432 15997 19441 16031
rect 19441 15997 19475 16031
rect 19475 15997 19484 16031
rect 19432 15988 19484 15997
rect 20260 15988 20312 16040
rect 20996 16056 21048 16108
rect 22284 16056 22336 16108
rect 23756 16056 23808 16108
rect 24216 16056 24268 16108
rect 24400 16056 24452 16108
rect 11152 15852 11204 15904
rect 11888 15852 11940 15904
rect 12072 15852 12124 15904
rect 13084 15895 13136 15904
rect 13084 15861 13093 15895
rect 13093 15861 13127 15895
rect 13127 15861 13136 15895
rect 13084 15852 13136 15861
rect 14004 15852 14056 15904
rect 14188 15852 14240 15904
rect 14464 15852 14516 15904
rect 14924 15852 14976 15904
rect 15292 15852 15344 15904
rect 16764 15852 16816 15904
rect 17040 15852 17092 15904
rect 17132 15852 17184 15904
rect 19248 15895 19300 15904
rect 19248 15861 19257 15895
rect 19257 15861 19291 15895
rect 19291 15861 19300 15895
rect 19248 15852 19300 15861
rect 20352 15852 20404 15904
rect 22744 15988 22796 16040
rect 23480 15988 23532 16040
rect 23664 15988 23716 16040
rect 23848 16031 23900 16040
rect 23848 15997 23857 16031
rect 23857 15997 23891 16031
rect 23891 15997 23900 16031
rect 23848 15988 23900 15997
rect 28264 16056 28316 16108
rect 24584 16031 24636 16040
rect 24584 15997 24593 16031
rect 24593 15997 24627 16031
rect 24627 15997 24636 16031
rect 24584 15988 24636 15997
rect 25964 15988 26016 16040
rect 23848 15852 23900 15904
rect 24308 15895 24360 15904
rect 24308 15861 24323 15895
rect 24323 15861 24357 15895
rect 24357 15861 24360 15895
rect 26700 15988 26752 16040
rect 26792 16031 26844 16040
rect 26792 15997 26801 16031
rect 26801 15997 26835 16031
rect 26835 15997 26844 16031
rect 26792 15988 26844 15997
rect 27252 15988 27304 16040
rect 27436 15988 27488 16040
rect 27804 15920 27856 15972
rect 24308 15852 24360 15861
rect 26332 15852 26384 15904
rect 26700 15852 26752 15904
rect 28816 15852 28868 15904
rect 30380 16192 30432 16244
rect 30472 16192 30524 16244
rect 30104 16099 30156 16108
rect 30104 16065 30113 16099
rect 30113 16065 30147 16099
rect 30147 16065 30156 16099
rect 30104 16056 30156 16065
rect 29184 15988 29236 16040
rect 29736 15988 29788 16040
rect 30196 15988 30248 16040
rect 30196 15852 30248 15904
rect 30472 15895 30524 15904
rect 30472 15861 30481 15895
rect 30481 15861 30515 15895
rect 30515 15861 30524 15895
rect 30472 15852 30524 15861
rect 7988 15750 8040 15802
rect 8052 15750 8104 15802
rect 8116 15750 8168 15802
rect 8180 15750 8232 15802
rect 8244 15750 8296 15802
rect 15578 15750 15630 15802
rect 15642 15750 15694 15802
rect 15706 15750 15758 15802
rect 15770 15750 15822 15802
rect 15834 15750 15886 15802
rect 23168 15750 23220 15802
rect 23232 15750 23284 15802
rect 23296 15750 23348 15802
rect 23360 15750 23412 15802
rect 23424 15750 23476 15802
rect 30758 15750 30810 15802
rect 30822 15750 30874 15802
rect 30886 15750 30938 15802
rect 30950 15750 31002 15802
rect 31014 15750 31066 15802
rect 1400 15648 1452 15700
rect 3148 15691 3200 15700
rect 3148 15657 3157 15691
rect 3157 15657 3191 15691
rect 3191 15657 3200 15691
rect 3148 15648 3200 15657
rect 5632 15623 5684 15632
rect 5632 15589 5641 15623
rect 5641 15589 5675 15623
rect 5675 15589 5684 15623
rect 5632 15580 5684 15589
rect 6460 15580 6512 15632
rect 7932 15580 7984 15632
rect 1676 15444 1728 15496
rect 2412 15444 2464 15496
rect 940 15351 992 15360
rect 940 15317 949 15351
rect 949 15317 983 15351
rect 983 15317 992 15351
rect 940 15308 992 15317
rect 1308 15308 1360 15360
rect 3608 15512 3660 15564
rect 4252 15555 4304 15564
rect 4252 15521 4261 15555
rect 4261 15521 4295 15555
rect 4295 15521 4304 15555
rect 4252 15512 4304 15521
rect 4344 15512 4396 15564
rect 13084 15648 13136 15700
rect 13452 15648 13504 15700
rect 15936 15648 15988 15700
rect 16396 15648 16448 15700
rect 18788 15648 18840 15700
rect 20352 15648 20404 15700
rect 11336 15580 11388 15632
rect 3884 15487 3936 15496
rect 3884 15453 3886 15487
rect 3886 15453 3936 15487
rect 3884 15444 3936 15453
rect 6000 15444 6052 15496
rect 8392 15512 8444 15564
rect 6092 15376 6144 15428
rect 7196 15487 7248 15496
rect 7196 15453 7205 15487
rect 7205 15453 7239 15487
rect 7239 15453 7248 15487
rect 7196 15444 7248 15453
rect 9036 15487 9088 15496
rect 9036 15453 9038 15487
rect 9038 15453 9088 15487
rect 9036 15444 9088 15453
rect 9220 15444 9272 15496
rect 9496 15444 9548 15496
rect 10968 15444 11020 15496
rect 11520 15580 11572 15632
rect 11888 15555 11940 15564
rect 11888 15521 11890 15555
rect 11890 15521 11940 15555
rect 11888 15512 11940 15521
rect 12256 15487 12308 15496
rect 12256 15453 12265 15487
rect 12265 15453 12299 15487
rect 12299 15453 12308 15487
rect 12256 15444 12308 15453
rect 3792 15308 3844 15360
rect 4344 15308 4396 15360
rect 4712 15308 4764 15360
rect 4896 15308 4948 15360
rect 8300 15351 8352 15360
rect 8300 15317 8309 15351
rect 8309 15317 8343 15351
rect 8343 15317 8352 15351
rect 8300 15308 8352 15317
rect 8668 15308 8720 15360
rect 14004 15444 14056 15496
rect 14464 15512 14516 15564
rect 14556 15555 14608 15564
rect 14556 15521 14565 15555
rect 14565 15521 14599 15555
rect 14599 15521 14608 15555
rect 14556 15512 14608 15521
rect 14832 15512 14884 15564
rect 16580 15555 16632 15564
rect 16580 15521 16589 15555
rect 16589 15521 16623 15555
rect 16623 15521 16632 15555
rect 16580 15512 16632 15521
rect 16396 15444 16448 15496
rect 13728 15376 13780 15428
rect 10140 15308 10192 15360
rect 11060 15308 11112 15360
rect 12164 15308 12216 15360
rect 13360 15351 13412 15360
rect 13360 15317 13369 15351
rect 13369 15317 13403 15351
rect 13403 15317 13412 15351
rect 13360 15308 13412 15317
rect 13636 15308 13688 15360
rect 16120 15419 16172 15428
rect 16120 15385 16129 15419
rect 16129 15385 16163 15419
rect 16163 15385 16172 15419
rect 16120 15376 16172 15385
rect 17040 15580 17092 15632
rect 17224 15444 17276 15496
rect 20720 15512 20772 15564
rect 18972 15444 19024 15496
rect 19616 15444 19668 15496
rect 16856 15376 16908 15428
rect 17408 15308 17460 15360
rect 18880 15351 18932 15360
rect 18880 15317 18889 15351
rect 18889 15317 18923 15351
rect 18923 15317 18932 15351
rect 18880 15308 18932 15317
rect 23020 15580 23072 15632
rect 24584 15648 24636 15700
rect 26792 15648 26844 15700
rect 27344 15648 27396 15700
rect 27804 15648 27856 15700
rect 23480 15580 23532 15632
rect 21272 15487 21324 15496
rect 21272 15453 21281 15487
rect 21281 15453 21315 15487
rect 21315 15453 21324 15487
rect 21272 15444 21324 15453
rect 21456 15444 21508 15496
rect 21640 15487 21692 15496
rect 21640 15453 21642 15487
rect 21642 15453 21692 15487
rect 21640 15444 21692 15453
rect 23572 15512 23624 15564
rect 24308 15512 24360 15564
rect 26240 15580 26292 15632
rect 26608 15580 26660 15632
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22008 15444 22060 15453
rect 23664 15444 23716 15496
rect 23848 15487 23900 15496
rect 23848 15453 23850 15487
rect 23850 15453 23900 15487
rect 23848 15444 23900 15453
rect 24676 15444 24728 15496
rect 26056 15512 26108 15564
rect 26240 15444 26292 15496
rect 21916 15308 21968 15360
rect 25964 15308 26016 15360
rect 26792 15376 26844 15428
rect 28356 15555 28408 15564
rect 28356 15521 28358 15555
rect 28358 15521 28408 15555
rect 28356 15512 28408 15521
rect 29368 15512 29420 15564
rect 28632 15444 28684 15496
rect 29828 15444 29880 15496
rect 29552 15376 29604 15428
rect 29736 15376 29788 15428
rect 28356 15308 28408 15360
rect 28540 15308 28592 15360
rect 4193 15206 4245 15258
rect 4257 15206 4309 15258
rect 4321 15206 4373 15258
rect 4385 15206 4437 15258
rect 4449 15206 4501 15258
rect 11783 15206 11835 15258
rect 11847 15206 11899 15258
rect 11911 15206 11963 15258
rect 11975 15206 12027 15258
rect 12039 15206 12091 15258
rect 19373 15206 19425 15258
rect 19437 15206 19489 15258
rect 19501 15206 19553 15258
rect 19565 15206 19617 15258
rect 19629 15206 19681 15258
rect 26963 15206 27015 15258
rect 27027 15206 27079 15258
rect 27091 15206 27143 15258
rect 27155 15206 27207 15258
rect 27219 15206 27271 15258
rect 1676 15104 1728 15156
rect 2964 15147 3016 15156
rect 2964 15113 2973 15147
rect 2973 15113 3007 15147
rect 3007 15113 3016 15147
rect 2964 15104 3016 15113
rect 4252 15104 4304 15156
rect 1308 14968 1360 15020
rect 3516 14968 3568 15020
rect 3792 14968 3844 15020
rect 8300 15104 8352 15156
rect 7932 15036 7984 15088
rect 10876 15104 10928 15156
rect 11796 15104 11848 15156
rect 15384 15104 15436 15156
rect 16212 15104 16264 15156
rect 17132 15104 17184 15156
rect 20260 15104 20312 15156
rect 20352 15104 20404 15156
rect 23388 15104 23440 15156
rect 23480 15104 23532 15156
rect 26516 15104 26568 15156
rect 6276 14968 6328 15020
rect 9036 15011 9088 15020
rect 2688 14900 2740 14952
rect 3700 14900 3752 14952
rect 4160 14900 4212 14952
rect 6092 14943 6144 14952
rect 6092 14909 6101 14943
rect 6101 14909 6135 14943
rect 6135 14909 6144 14943
rect 6092 14900 6144 14909
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 7288 14900 7340 14952
rect 8484 14900 8536 14952
rect 1400 14807 1452 14816
rect 1400 14773 1415 14807
rect 1415 14773 1449 14807
rect 1449 14773 1452 14807
rect 1400 14764 1452 14773
rect 3884 14764 3936 14816
rect 6460 14764 6512 14816
rect 6920 14764 6972 14816
rect 8668 14943 8720 14952
rect 8668 14909 8677 14943
rect 8677 14909 8711 14943
rect 8711 14909 8720 14943
rect 8668 14900 8720 14909
rect 9036 14977 9038 15011
rect 9038 14977 9088 15011
rect 9036 14968 9088 14977
rect 9220 14968 9272 15020
rect 9404 14943 9456 14952
rect 9404 14909 9413 14943
rect 9413 14909 9447 14943
rect 9447 14909 9456 14943
rect 9404 14900 9456 14909
rect 10324 14900 10376 14952
rect 10876 14900 10928 14952
rect 11060 14900 11112 14952
rect 11336 14900 11388 14952
rect 11796 14968 11848 15020
rect 13912 15079 13964 15088
rect 13912 15045 13921 15079
rect 13921 15045 13955 15079
rect 13955 15045 13964 15079
rect 13912 15036 13964 15045
rect 14096 15036 14148 15088
rect 13636 14968 13688 15020
rect 12440 14900 12492 14952
rect 12624 14900 12676 14952
rect 13452 14832 13504 14884
rect 13728 14832 13780 14884
rect 11336 14764 11388 14816
rect 11704 14807 11756 14816
rect 11704 14773 11719 14807
rect 11719 14773 11753 14807
rect 11753 14773 11756 14807
rect 14280 14900 14332 14952
rect 14464 14900 14516 14952
rect 14004 14832 14056 14884
rect 15200 14900 15252 14952
rect 15292 14943 15344 14952
rect 15292 14909 15301 14943
rect 15301 14909 15335 14943
rect 15335 14909 15344 14943
rect 15292 14900 15344 14909
rect 11704 14764 11756 14773
rect 14096 14764 14148 14816
rect 14372 14764 14424 14816
rect 14924 14764 14976 14816
rect 16396 14807 16448 14816
rect 16396 14773 16405 14807
rect 16405 14773 16439 14807
rect 16439 14773 16448 14807
rect 16396 14764 16448 14773
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 19432 15036 19484 15088
rect 23848 15036 23900 15088
rect 26424 15036 26476 15088
rect 27344 15104 27396 15156
rect 28356 15104 28408 15156
rect 28540 15104 28592 15156
rect 29000 15104 29052 15156
rect 29460 15104 29512 15156
rect 30656 15104 30708 15156
rect 29368 15036 29420 15088
rect 29920 15079 29972 15088
rect 29920 15045 29929 15079
rect 29929 15045 29963 15079
rect 29963 15045 29972 15079
rect 29920 15036 29972 15045
rect 19984 14968 20036 15020
rect 17592 14900 17644 14952
rect 18788 14900 18840 14952
rect 17960 14832 18012 14884
rect 19708 14900 19760 14952
rect 20352 14943 20404 14952
rect 20352 14909 20361 14943
rect 20361 14909 20395 14943
rect 20395 14909 20404 14943
rect 20352 14900 20404 14909
rect 22928 14968 22980 15020
rect 23664 14968 23716 15020
rect 24768 14968 24820 15020
rect 24952 14968 25004 15020
rect 23572 14900 23624 14952
rect 22100 14832 22152 14884
rect 24676 14900 24728 14952
rect 27068 14968 27120 15020
rect 18788 14764 18840 14816
rect 19156 14764 19208 14816
rect 20628 14764 20680 14816
rect 21180 14764 21232 14816
rect 21548 14764 21600 14816
rect 22744 14764 22796 14816
rect 22928 14764 22980 14816
rect 26148 14764 26200 14816
rect 26608 14900 26660 14952
rect 26792 14900 26844 14952
rect 27252 14968 27304 15020
rect 27344 14900 27396 14952
rect 29000 14900 29052 14952
rect 29184 14900 29236 14952
rect 30012 14900 30064 14952
rect 30196 14900 30248 14952
rect 30472 14900 30524 14952
rect 27436 14764 27488 14816
rect 27712 14764 27764 14816
rect 7988 14662 8040 14714
rect 8052 14662 8104 14714
rect 8116 14662 8168 14714
rect 8180 14662 8232 14714
rect 8244 14662 8296 14714
rect 15578 14662 15630 14714
rect 15642 14662 15694 14714
rect 15706 14662 15758 14714
rect 15770 14662 15822 14714
rect 15834 14662 15886 14714
rect 23168 14662 23220 14714
rect 23232 14662 23284 14714
rect 23296 14662 23348 14714
rect 23360 14662 23412 14714
rect 23424 14662 23476 14714
rect 30758 14662 30810 14714
rect 30822 14662 30874 14714
rect 30886 14662 30938 14714
rect 30950 14662 31002 14714
rect 31014 14662 31066 14714
rect 1124 14467 1176 14476
rect 1124 14433 1133 14467
rect 1133 14433 1167 14467
rect 1167 14433 1176 14467
rect 1124 14424 1176 14433
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 4068 14603 4120 14612
rect 4068 14569 4077 14603
rect 4077 14569 4111 14603
rect 4111 14569 4120 14603
rect 4068 14560 4120 14569
rect 4528 14560 4580 14612
rect 5080 14560 5132 14612
rect 4620 14492 4672 14544
rect 1492 14399 1544 14408
rect 1492 14365 1501 14399
rect 1501 14365 1535 14399
rect 1535 14365 1544 14399
rect 1492 14356 1544 14365
rect 1768 14356 1820 14408
rect 2044 14356 2096 14408
rect 2228 14399 2280 14408
rect 2228 14365 2237 14399
rect 2237 14365 2271 14399
rect 2271 14365 2280 14399
rect 2228 14356 2280 14365
rect 3240 14356 3292 14408
rect 4252 14467 4304 14476
rect 4252 14433 4261 14467
rect 4261 14433 4295 14467
rect 4295 14433 4304 14467
rect 4252 14424 4304 14433
rect 4436 14424 4488 14476
rect 6828 14560 6880 14612
rect 9036 14560 9088 14612
rect 9864 14560 9916 14612
rect 5816 14492 5868 14544
rect 5172 14424 5224 14476
rect 5264 14424 5316 14476
rect 5448 14424 5500 14476
rect 6184 14424 6236 14476
rect 6276 14356 6328 14408
rect 6644 14424 6696 14476
rect 8484 14424 8536 14476
rect 8760 14424 8812 14476
rect 10324 14492 10376 14544
rect 10784 14560 10836 14612
rect 12164 14560 12216 14612
rect 13360 14560 13412 14612
rect 9772 14467 9824 14476
rect 9772 14433 9781 14467
rect 9781 14433 9815 14467
rect 9815 14433 9824 14467
rect 9772 14424 9824 14433
rect 6828 14399 6880 14408
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 7196 14399 7248 14408
rect 7196 14365 7198 14399
rect 7198 14365 7248 14399
rect 7196 14356 7248 14365
rect 7288 14399 7340 14408
rect 7288 14365 7300 14399
rect 7300 14365 7334 14399
rect 7334 14365 7340 14399
rect 7288 14356 7340 14365
rect 7564 14399 7616 14408
rect 7564 14365 7573 14399
rect 7573 14365 7607 14399
rect 7607 14365 7616 14399
rect 7564 14356 7616 14365
rect 8576 14356 8628 14408
rect 10600 14424 10652 14476
rect 10692 14424 10744 14476
rect 10876 14424 10928 14476
rect 11428 14424 11480 14476
rect 12624 14424 12676 14476
rect 13176 14424 13228 14476
rect 11336 14356 11388 14408
rect 11796 14356 11848 14408
rect 16396 14560 16448 14612
rect 16488 14603 16540 14612
rect 16488 14569 16497 14603
rect 16497 14569 16531 14603
rect 16531 14569 16540 14603
rect 16488 14560 16540 14569
rect 16672 14603 16724 14612
rect 16672 14569 16681 14603
rect 16681 14569 16715 14603
rect 16715 14569 16724 14603
rect 16672 14560 16724 14569
rect 17040 14560 17092 14612
rect 17960 14560 18012 14612
rect 18788 14603 18840 14612
rect 18788 14569 18797 14603
rect 18797 14569 18831 14603
rect 18831 14569 18840 14603
rect 18788 14560 18840 14569
rect 21548 14560 21600 14612
rect 21640 14560 21692 14612
rect 22100 14560 22152 14612
rect 25412 14560 25464 14612
rect 26976 14560 27028 14612
rect 27620 14560 27672 14612
rect 28356 14560 28408 14612
rect 29184 14560 29236 14612
rect 29276 14560 29328 14612
rect 15384 14492 15436 14544
rect 13912 14424 13964 14476
rect 15016 14424 15068 14476
rect 6368 14288 6420 14340
rect 3516 14263 3568 14272
rect 3516 14229 3525 14263
rect 3525 14229 3559 14263
rect 3559 14229 3568 14263
rect 3516 14220 3568 14229
rect 3792 14220 3844 14272
rect 4068 14220 4120 14272
rect 5724 14220 5776 14272
rect 5816 14263 5868 14272
rect 5816 14229 5825 14263
rect 5825 14229 5859 14263
rect 5859 14229 5868 14263
rect 5816 14220 5868 14229
rect 5908 14220 5960 14272
rect 6736 14288 6788 14340
rect 9680 14288 9732 14340
rect 8760 14220 8812 14272
rect 10692 14220 10744 14272
rect 12256 14220 12308 14272
rect 12348 14220 12400 14272
rect 14004 14356 14056 14408
rect 14372 14356 14424 14408
rect 14464 14356 14516 14408
rect 16304 14356 16356 14408
rect 18328 14424 18380 14476
rect 14188 14220 14240 14272
rect 15016 14220 15068 14272
rect 16028 14220 16080 14272
rect 16488 14220 16540 14272
rect 17408 14356 17460 14408
rect 19432 14467 19484 14476
rect 19432 14433 19441 14467
rect 19441 14433 19475 14467
rect 19475 14433 19484 14467
rect 19432 14424 19484 14433
rect 21272 14467 21324 14476
rect 21272 14433 21281 14467
rect 21281 14433 21315 14467
rect 21315 14433 21324 14467
rect 21272 14424 21324 14433
rect 23848 14467 23900 14476
rect 23848 14433 23850 14467
rect 23850 14433 23900 14467
rect 23848 14424 23900 14433
rect 24124 14424 24176 14476
rect 24492 14424 24544 14476
rect 25964 14424 26016 14476
rect 26424 14467 26476 14476
rect 26424 14433 26433 14467
rect 26433 14433 26467 14467
rect 26467 14433 26476 14467
rect 26424 14424 26476 14433
rect 21180 14356 21232 14408
rect 21916 14356 21968 14408
rect 22008 14399 22060 14408
rect 22008 14365 22017 14399
rect 22017 14365 22051 14399
rect 22051 14365 22060 14399
rect 22008 14356 22060 14365
rect 23664 14356 23716 14408
rect 24860 14356 24912 14408
rect 26700 14424 26752 14476
rect 28172 14492 28224 14544
rect 27988 14424 28040 14476
rect 29184 14424 29236 14476
rect 31300 14492 31352 14544
rect 30012 14424 30064 14476
rect 30196 14424 30248 14476
rect 27068 14356 27120 14408
rect 27528 14356 27580 14408
rect 20536 14288 20588 14340
rect 18144 14220 18196 14272
rect 21272 14220 21324 14272
rect 24032 14220 24084 14272
rect 26792 14220 26844 14272
rect 26976 14220 27028 14272
rect 28632 14220 28684 14272
rect 4193 14118 4245 14170
rect 4257 14118 4309 14170
rect 4321 14118 4373 14170
rect 4385 14118 4437 14170
rect 4449 14118 4501 14170
rect 11783 14118 11835 14170
rect 11847 14118 11899 14170
rect 11911 14118 11963 14170
rect 11975 14118 12027 14170
rect 12039 14118 12091 14170
rect 19373 14118 19425 14170
rect 19437 14118 19489 14170
rect 19501 14118 19553 14170
rect 19565 14118 19617 14170
rect 19629 14118 19681 14170
rect 26963 14118 27015 14170
rect 27027 14118 27079 14170
rect 27091 14118 27143 14170
rect 27155 14118 27207 14170
rect 27219 14118 27271 14170
rect 1124 14016 1176 14068
rect 2044 13880 2096 13932
rect 2780 14059 2832 14068
rect 2780 14025 2789 14059
rect 2789 14025 2823 14059
rect 2823 14025 2832 14059
rect 2780 14016 2832 14025
rect 3424 14016 3476 14068
rect 5724 14016 5776 14068
rect 5816 14016 5868 14068
rect 3608 13948 3660 14000
rect 1216 13812 1268 13864
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 2504 13812 2556 13864
rect 4528 13880 4580 13932
rect 6920 14016 6972 14068
rect 7012 14016 7064 14068
rect 7748 14016 7800 14068
rect 8944 14016 8996 14068
rect 9220 14059 9272 14068
rect 9220 14025 9229 14059
rect 9229 14025 9263 14059
rect 9263 14025 9272 14059
rect 9220 14016 9272 14025
rect 9312 14016 9364 14068
rect 8852 13948 8904 14000
rect 12348 14016 12400 14068
rect 12440 14059 12492 14068
rect 12440 14025 12449 14059
rect 12449 14025 12483 14059
rect 12483 14025 12492 14059
rect 12440 14016 12492 14025
rect 12532 14016 12584 14068
rect 11704 13948 11756 14000
rect 6460 13923 6512 13932
rect 3884 13855 3936 13864
rect 3884 13821 3893 13855
rect 3893 13821 3927 13855
rect 3927 13821 3936 13855
rect 3884 13812 3936 13821
rect 4252 13812 4304 13864
rect 5080 13812 5132 13864
rect 6092 13855 6144 13864
rect 6092 13821 6101 13855
rect 6101 13821 6135 13855
rect 6135 13821 6144 13855
rect 6092 13812 6144 13821
rect 6460 13889 6462 13923
rect 6462 13889 6512 13923
rect 6460 13880 6512 13889
rect 8944 13855 8996 13864
rect 8944 13821 8953 13855
rect 8953 13821 8987 13855
rect 8987 13821 8996 13855
rect 8944 13812 8996 13821
rect 9404 13812 9456 13864
rect 9680 13855 9732 13864
rect 9680 13821 9689 13855
rect 9689 13821 9723 13855
rect 9723 13821 9732 13855
rect 9680 13812 9732 13821
rect 9956 13812 10008 13864
rect 10140 13923 10192 13932
rect 10140 13889 10152 13923
rect 10152 13889 10186 13923
rect 10186 13889 10192 13923
rect 10140 13880 10192 13889
rect 12072 13880 12124 13932
rect 10416 13855 10468 13864
rect 10416 13821 10425 13855
rect 10425 13821 10459 13855
rect 10459 13821 10468 13855
rect 10416 13812 10468 13821
rect 11520 13812 11572 13864
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 12716 13991 12768 14000
rect 12716 13957 12725 13991
rect 12725 13957 12759 13991
rect 12759 13957 12768 13991
rect 12716 13948 12768 13957
rect 12624 13855 12676 13864
rect 12624 13821 12633 13855
rect 12633 13821 12667 13855
rect 12667 13821 12676 13855
rect 12624 13812 12676 13821
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 13912 14059 13964 14068
rect 13912 14025 13921 14059
rect 13921 14025 13955 14059
rect 13955 14025 13964 14059
rect 13912 14016 13964 14025
rect 14096 13948 14148 14000
rect 1400 13719 1452 13728
rect 1400 13685 1415 13719
rect 1415 13685 1449 13719
rect 1449 13685 1452 13719
rect 1400 13676 1452 13685
rect 3976 13676 4028 13728
rect 9588 13676 9640 13728
rect 10692 13676 10744 13728
rect 11520 13676 11572 13728
rect 12716 13744 12768 13796
rect 13728 13744 13780 13796
rect 14096 13855 14148 13864
rect 14096 13821 14105 13855
rect 14105 13821 14139 13855
rect 14139 13821 14148 13855
rect 14096 13812 14148 13821
rect 14188 13855 14240 13864
rect 14188 13821 14197 13855
rect 14197 13821 14231 13855
rect 14231 13821 14240 13855
rect 14188 13812 14240 13821
rect 18880 14016 18932 14068
rect 18972 14059 19024 14068
rect 18972 14025 18981 14059
rect 18981 14025 19015 14059
rect 19015 14025 19024 14059
rect 18972 14016 19024 14025
rect 20352 14016 20404 14068
rect 22928 14016 22980 14068
rect 23020 14059 23072 14068
rect 23020 14025 23029 14059
rect 23029 14025 23063 14059
rect 23063 14025 23072 14059
rect 23020 14016 23072 14025
rect 16948 13880 17000 13932
rect 23572 13948 23624 14000
rect 15200 13812 15252 13864
rect 16488 13812 16540 13864
rect 17040 13812 17092 13864
rect 17960 13812 18012 13864
rect 18880 13855 18932 13864
rect 18880 13821 18889 13855
rect 18889 13821 18923 13855
rect 18923 13821 18932 13855
rect 18880 13812 18932 13821
rect 19156 13855 19208 13864
rect 19156 13821 19165 13855
rect 19165 13821 19199 13855
rect 19199 13821 19208 13855
rect 19156 13812 19208 13821
rect 13912 13744 13964 13796
rect 19892 13855 19944 13864
rect 19892 13821 19901 13855
rect 19901 13821 19935 13855
rect 19935 13821 19944 13855
rect 19892 13812 19944 13821
rect 20168 13812 20220 13864
rect 20260 13812 20312 13864
rect 20628 13855 20680 13864
rect 20628 13821 20637 13855
rect 20637 13821 20671 13855
rect 20671 13821 20680 13855
rect 20628 13812 20680 13821
rect 22284 13812 22336 13864
rect 23756 13880 23808 13932
rect 24860 13923 24912 13932
rect 23020 13744 23072 13796
rect 24400 13855 24452 13864
rect 24400 13821 24409 13855
rect 24409 13821 24443 13855
rect 24443 13821 24452 13855
rect 24400 13812 24452 13821
rect 24860 13889 24862 13923
rect 24862 13889 24912 13923
rect 24860 13880 24912 13889
rect 26884 14016 26936 14068
rect 28080 14016 28132 14068
rect 29092 14016 29144 14068
rect 29736 14016 29788 14068
rect 30564 14016 30616 14068
rect 14556 13676 14608 13728
rect 14924 13676 14976 13728
rect 17132 13676 17184 13728
rect 18236 13719 18288 13728
rect 18236 13685 18245 13719
rect 18245 13685 18279 13719
rect 18279 13685 18288 13719
rect 18236 13676 18288 13685
rect 18696 13719 18748 13728
rect 18696 13685 18705 13719
rect 18705 13685 18739 13719
rect 18739 13685 18748 13719
rect 18696 13676 18748 13685
rect 19248 13676 19300 13728
rect 19800 13676 19852 13728
rect 20260 13676 20312 13728
rect 20904 13676 20956 13728
rect 22836 13676 22888 13728
rect 24308 13744 24360 13796
rect 25688 13812 25740 13864
rect 26148 13812 26200 13864
rect 26424 13812 26476 13864
rect 26884 13880 26936 13932
rect 27620 13880 27672 13932
rect 24584 13744 24636 13796
rect 25320 13676 25372 13728
rect 25596 13676 25648 13728
rect 26056 13676 26108 13728
rect 27068 13676 27120 13728
rect 28172 13812 28224 13864
rect 29644 13948 29696 14000
rect 29920 13880 29972 13932
rect 30472 13880 30524 13932
rect 29552 13744 29604 13796
rect 30104 13744 30156 13796
rect 28172 13676 28224 13728
rect 28816 13676 28868 13728
rect 7988 13574 8040 13626
rect 8052 13574 8104 13626
rect 8116 13574 8168 13626
rect 8180 13574 8232 13626
rect 8244 13574 8296 13626
rect 15578 13574 15630 13626
rect 15642 13574 15694 13626
rect 15706 13574 15758 13626
rect 15770 13574 15822 13626
rect 15834 13574 15886 13626
rect 23168 13574 23220 13626
rect 23232 13574 23284 13626
rect 23296 13574 23348 13626
rect 23360 13574 23412 13626
rect 23424 13574 23476 13626
rect 30758 13574 30810 13626
rect 30822 13574 30874 13626
rect 30886 13574 30938 13626
rect 30950 13574 31002 13626
rect 31014 13574 31066 13626
rect 1768 13515 1820 13524
rect 1768 13481 1783 13515
rect 1783 13481 1817 13515
rect 1817 13481 1820 13515
rect 1768 13472 1820 13481
rect 3976 13515 4028 13524
rect 3976 13481 3991 13515
rect 3991 13481 4025 13515
rect 4025 13481 4028 13515
rect 3976 13472 4028 13481
rect 6552 13515 6604 13524
rect 6552 13481 6561 13515
rect 6561 13481 6595 13515
rect 6595 13481 6604 13515
rect 6552 13472 6604 13481
rect 8760 13472 8812 13524
rect 9404 13472 9456 13524
rect 9864 13472 9916 13524
rect 1124 13268 1176 13320
rect 1308 13311 1360 13320
rect 1308 13277 1317 13311
rect 1317 13277 1351 13311
rect 1351 13277 1360 13311
rect 1308 13268 1360 13277
rect 1492 13268 1544 13320
rect 3148 13336 3200 13388
rect 3332 13268 3384 13320
rect 5632 13447 5684 13456
rect 5632 13413 5641 13447
rect 5641 13413 5675 13447
rect 5675 13413 5684 13447
rect 5632 13404 5684 13413
rect 6276 13404 6328 13456
rect 5080 13268 5132 13320
rect 5356 13268 5408 13320
rect 6828 13379 6880 13388
rect 6828 13345 6837 13379
rect 6837 13345 6871 13379
rect 6871 13345 6880 13379
rect 6828 13336 6880 13345
rect 9312 13447 9364 13456
rect 9312 13413 9321 13447
rect 9321 13413 9355 13447
rect 9355 13413 9364 13447
rect 9312 13404 9364 13413
rect 6644 13268 6696 13320
rect 6368 13200 6420 13252
rect 7196 13311 7248 13320
rect 7196 13277 7198 13311
rect 7198 13277 7248 13311
rect 7196 13268 7248 13277
rect 7288 13311 7340 13320
rect 7288 13277 7300 13311
rect 7300 13277 7334 13311
rect 7334 13277 7340 13311
rect 7288 13268 7340 13277
rect 1032 13175 1084 13184
rect 1032 13141 1041 13175
rect 1041 13141 1075 13175
rect 1075 13141 1084 13175
rect 1032 13132 1084 13141
rect 3332 13132 3384 13184
rect 3884 13132 3936 13184
rect 4252 13132 4304 13184
rect 5908 13132 5960 13184
rect 6276 13175 6328 13184
rect 6276 13141 6285 13175
rect 6285 13141 6319 13175
rect 6319 13141 6328 13175
rect 6276 13132 6328 13141
rect 7472 13132 7524 13184
rect 8852 13175 8904 13184
rect 8852 13141 8861 13175
rect 8861 13141 8895 13175
rect 8895 13141 8904 13175
rect 8852 13132 8904 13141
rect 9864 13379 9916 13388
rect 9864 13345 9873 13379
rect 9873 13345 9907 13379
rect 9907 13345 9916 13379
rect 9864 13336 9916 13345
rect 10876 13472 10928 13524
rect 10968 13472 11020 13524
rect 11612 13472 11664 13524
rect 11704 13472 11756 13524
rect 12716 13472 12768 13524
rect 13268 13472 13320 13524
rect 14280 13472 14332 13524
rect 16396 13472 16448 13524
rect 16580 13472 16632 13524
rect 17132 13472 17184 13524
rect 17684 13472 17736 13524
rect 9772 13268 9824 13320
rect 11152 13336 11204 13388
rect 11520 13404 11572 13456
rect 11888 13404 11940 13456
rect 11980 13379 12032 13388
rect 11980 13345 11989 13379
rect 11989 13345 12023 13379
rect 12023 13345 12032 13379
rect 11980 13336 12032 13345
rect 12532 13404 12584 13456
rect 13912 13404 13964 13456
rect 10784 13268 10836 13320
rect 12440 13311 12492 13320
rect 12440 13277 12449 13311
rect 12449 13277 12483 13311
rect 12483 13277 12492 13311
rect 12440 13268 12492 13277
rect 15476 13336 15528 13388
rect 15752 13336 15804 13388
rect 12992 13268 13044 13320
rect 13268 13268 13320 13320
rect 13912 13268 13964 13320
rect 14924 13268 14976 13320
rect 10416 13200 10468 13252
rect 10692 13200 10744 13252
rect 11060 13200 11112 13252
rect 9312 13132 9364 13184
rect 9496 13132 9548 13184
rect 10232 13132 10284 13184
rect 10508 13132 10560 13184
rect 11520 13243 11572 13252
rect 11520 13209 11529 13243
rect 11529 13209 11563 13243
rect 11563 13209 11572 13243
rect 11520 13200 11572 13209
rect 11888 13132 11940 13184
rect 12256 13132 12308 13184
rect 16028 13336 16080 13388
rect 16120 13379 16172 13388
rect 16120 13345 16129 13379
rect 16129 13345 16163 13379
rect 16163 13345 16172 13379
rect 16120 13336 16172 13345
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 17040 13379 17092 13388
rect 17040 13345 17049 13379
rect 17049 13345 17083 13379
rect 17083 13345 17092 13379
rect 17040 13336 17092 13345
rect 18512 13404 18564 13456
rect 25320 13472 25372 13524
rect 26332 13472 26384 13524
rect 26424 13472 26476 13524
rect 26884 13515 26936 13524
rect 26884 13481 26899 13515
rect 26899 13481 26933 13515
rect 26933 13481 26936 13515
rect 26884 13472 26936 13481
rect 27068 13472 27120 13524
rect 17408 13336 17460 13388
rect 18696 13336 18748 13388
rect 19984 13336 20036 13388
rect 20260 13336 20312 13388
rect 20536 13336 20588 13388
rect 21272 13268 21324 13320
rect 21732 13336 21784 13388
rect 24032 13447 24084 13456
rect 24032 13413 24041 13447
rect 24041 13413 24075 13447
rect 24075 13413 24084 13447
rect 24032 13404 24084 13413
rect 24216 13404 24268 13456
rect 23572 13336 23624 13388
rect 21640 13268 21692 13320
rect 22192 13268 22244 13320
rect 22284 13268 22336 13320
rect 24124 13311 24176 13320
rect 24124 13277 24133 13311
rect 24133 13277 24167 13311
rect 24167 13277 24176 13311
rect 24124 13268 24176 13277
rect 24400 13268 24452 13320
rect 24492 13268 24544 13320
rect 24676 13268 24728 13320
rect 26516 13336 26568 13388
rect 27620 13336 27672 13388
rect 28264 13515 28316 13524
rect 28264 13481 28273 13515
rect 28273 13481 28307 13515
rect 28307 13481 28316 13515
rect 28264 13472 28316 13481
rect 28172 13404 28224 13456
rect 28632 13404 28684 13456
rect 16396 13200 16448 13252
rect 14280 13175 14332 13184
rect 14280 13141 14289 13175
rect 14289 13141 14323 13175
rect 14323 13141 14332 13175
rect 14280 13132 14332 13141
rect 15752 13175 15804 13184
rect 15752 13141 15761 13175
rect 15761 13141 15795 13175
rect 15795 13141 15804 13175
rect 15752 13132 15804 13141
rect 15844 13132 15896 13184
rect 16672 13132 16724 13184
rect 20076 13200 20128 13252
rect 19340 13132 19392 13184
rect 19984 13132 20036 13184
rect 20352 13132 20404 13184
rect 21824 13132 21876 13184
rect 21916 13132 21968 13184
rect 23756 13132 23808 13184
rect 27528 13132 27580 13184
rect 28816 13132 28868 13184
rect 4193 13030 4245 13082
rect 4257 13030 4309 13082
rect 4321 13030 4373 13082
rect 4385 13030 4437 13082
rect 4449 13030 4501 13082
rect 11783 13030 11835 13082
rect 11847 13030 11899 13082
rect 11911 13030 11963 13082
rect 11975 13030 12027 13082
rect 12039 13030 12091 13082
rect 19373 13030 19425 13082
rect 19437 13030 19489 13082
rect 19501 13030 19553 13082
rect 19565 13030 19617 13082
rect 19629 13030 19681 13082
rect 26963 13030 27015 13082
rect 27027 13030 27079 13082
rect 27091 13030 27143 13082
rect 27155 13030 27207 13082
rect 27219 13030 27271 13082
rect 1676 12928 1728 12980
rect 3148 12928 3200 12980
rect 3516 12928 3568 12980
rect 3884 12928 3936 12980
rect 7288 12928 7340 12980
rect 7656 12928 7708 12980
rect 9312 12928 9364 12980
rect 10048 12928 10100 12980
rect 12348 12928 12400 12980
rect 1308 12792 1360 12844
rect 2136 12724 2188 12776
rect 3056 12835 3108 12844
rect 3056 12801 3065 12835
rect 3065 12801 3099 12835
rect 3099 12801 3108 12835
rect 3056 12792 3108 12801
rect 3332 12792 3384 12844
rect 3424 12792 3476 12844
rect 4252 12792 4304 12844
rect 5356 12792 5408 12844
rect 11244 12860 11296 12912
rect 12072 12860 12124 12912
rect 12716 12928 12768 12980
rect 12808 12928 12860 12980
rect 12992 12928 13044 12980
rect 13176 12928 13228 12980
rect 13636 12928 13688 12980
rect 14096 12928 14148 12980
rect 10048 12792 10100 12844
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 10508 12792 10560 12844
rect 12256 12792 12308 12844
rect 14372 12860 14424 12912
rect 16764 12971 16816 12980
rect 16764 12937 16773 12971
rect 16773 12937 16807 12971
rect 16807 12937 16816 12971
rect 16764 12928 16816 12937
rect 16856 12928 16908 12980
rect 3516 12767 3568 12776
rect 3516 12733 3525 12767
rect 3525 12733 3559 12767
rect 3559 12733 3568 12767
rect 3516 12724 3568 12733
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 5632 12724 5684 12776
rect 6184 12724 6236 12776
rect 7196 12724 7248 12776
rect 8760 12724 8812 12776
rect 9128 12724 9180 12776
rect 1676 12588 1728 12640
rect 2596 12588 2648 12640
rect 8484 12699 8536 12708
rect 8484 12665 8493 12699
rect 8493 12665 8527 12699
rect 8527 12665 8536 12699
rect 8484 12656 8536 12665
rect 9312 12767 9364 12776
rect 9312 12733 9321 12767
rect 9321 12733 9355 12767
rect 9355 12733 9364 12767
rect 9312 12724 9364 12733
rect 9680 12767 9732 12776
rect 9680 12733 9689 12767
rect 9689 12733 9723 12767
rect 9723 12733 9732 12767
rect 9680 12724 9732 12733
rect 11612 12724 11664 12776
rect 11980 12724 12032 12776
rect 12348 12767 12400 12776
rect 12348 12733 12365 12767
rect 12365 12733 12399 12767
rect 12399 12733 12400 12767
rect 12348 12724 12400 12733
rect 11152 12656 11204 12708
rect 13176 12724 13228 12776
rect 13636 12792 13688 12844
rect 13912 12792 13964 12844
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 14924 12835 14976 12844
rect 14924 12801 14926 12835
rect 14926 12801 14976 12835
rect 14924 12792 14976 12801
rect 13820 12724 13872 12776
rect 15752 12792 15804 12844
rect 18236 12792 18288 12844
rect 16304 12724 16356 12776
rect 20628 12928 20680 12980
rect 23572 12928 23624 12980
rect 24492 12928 24544 12980
rect 25688 12971 25740 12980
rect 25688 12937 25697 12971
rect 25697 12937 25731 12971
rect 25731 12937 25740 12971
rect 25688 12928 25740 12937
rect 26608 12928 26660 12980
rect 22928 12860 22980 12912
rect 23756 12860 23808 12912
rect 19892 12792 19944 12844
rect 20812 12835 20864 12844
rect 20812 12801 20824 12835
rect 20824 12801 20858 12835
rect 20858 12801 20864 12835
rect 20812 12792 20864 12801
rect 3976 12588 4028 12640
rect 4896 12588 4948 12640
rect 7472 12588 7524 12640
rect 8576 12631 8628 12640
rect 8576 12597 8585 12631
rect 8585 12597 8619 12631
rect 8619 12597 8628 12631
rect 8576 12588 8628 12597
rect 9036 12588 9088 12640
rect 9588 12588 9640 12640
rect 12256 12588 12308 12640
rect 12348 12588 12400 12640
rect 13176 12631 13228 12640
rect 13176 12597 13185 12631
rect 13185 12597 13219 12631
rect 13219 12597 13228 12631
rect 13176 12588 13228 12597
rect 14004 12656 14056 12708
rect 18052 12656 18104 12708
rect 18328 12699 18380 12708
rect 18328 12665 18337 12699
rect 18337 12665 18371 12699
rect 18371 12665 18380 12699
rect 18328 12656 18380 12665
rect 19800 12724 19852 12776
rect 20260 12767 20312 12776
rect 20260 12733 20269 12767
rect 20269 12733 20303 12767
rect 20303 12733 20312 12767
rect 20260 12724 20312 12733
rect 20352 12767 20404 12776
rect 20352 12733 20361 12767
rect 20361 12733 20395 12767
rect 20395 12733 20404 12767
rect 20352 12724 20404 12733
rect 20904 12724 20956 12776
rect 22008 12792 22060 12844
rect 22192 12792 22244 12844
rect 23848 12835 23900 12844
rect 23848 12801 23857 12835
rect 23857 12801 23891 12835
rect 23891 12801 23900 12835
rect 23848 12792 23900 12801
rect 24124 12792 24176 12844
rect 21088 12767 21140 12776
rect 21088 12733 21097 12767
rect 21097 12733 21131 12767
rect 21131 12733 21140 12767
rect 21088 12724 21140 12733
rect 14556 12588 14608 12640
rect 14832 12588 14884 12640
rect 16948 12588 17000 12640
rect 18696 12631 18748 12640
rect 18696 12597 18705 12631
rect 18705 12597 18739 12631
rect 18739 12597 18748 12631
rect 18696 12588 18748 12597
rect 19708 12588 19760 12640
rect 21180 12588 21232 12640
rect 21456 12588 21508 12640
rect 22836 12724 22888 12776
rect 23112 12724 23164 12776
rect 23756 12724 23808 12776
rect 24492 12792 24544 12844
rect 28908 12928 28960 12980
rect 29828 12971 29880 12980
rect 29828 12937 29837 12971
rect 29837 12937 29871 12971
rect 29871 12937 29880 12971
rect 29828 12928 29880 12937
rect 24400 12724 24452 12776
rect 26424 12724 26476 12776
rect 27804 12792 27856 12844
rect 29552 12792 29604 12844
rect 29368 12656 29420 12708
rect 24124 12588 24176 12640
rect 24216 12588 24268 12640
rect 26148 12588 26200 12640
rect 26516 12588 26568 12640
rect 27436 12588 27488 12640
rect 28080 12588 28132 12640
rect 28632 12588 28684 12640
rect 30012 12767 30064 12776
rect 30012 12733 30013 12767
rect 30013 12733 30047 12767
rect 30047 12733 30064 12767
rect 30012 12724 30064 12733
rect 7988 12486 8040 12538
rect 8052 12486 8104 12538
rect 8116 12486 8168 12538
rect 8180 12486 8232 12538
rect 8244 12486 8296 12538
rect 15578 12486 15630 12538
rect 15642 12486 15694 12538
rect 15706 12486 15758 12538
rect 15770 12486 15822 12538
rect 15834 12486 15886 12538
rect 23168 12486 23220 12538
rect 23232 12486 23284 12538
rect 23296 12486 23348 12538
rect 23360 12486 23412 12538
rect 23424 12486 23476 12538
rect 30758 12486 30810 12538
rect 30822 12486 30874 12538
rect 30886 12486 30938 12538
rect 30950 12486 31002 12538
rect 31014 12486 31066 12538
rect 1032 12384 1084 12436
rect 1952 12384 2004 12436
rect 3976 12427 4028 12436
rect 3976 12393 3991 12427
rect 3991 12393 4025 12427
rect 4025 12393 4028 12427
rect 3976 12384 4028 12393
rect 5264 12384 5316 12436
rect 5724 12384 5776 12436
rect 6092 12384 6144 12436
rect 2872 12248 2924 12300
rect 1308 12223 1360 12232
rect 1308 12189 1317 12223
rect 1317 12189 1351 12223
rect 1351 12189 1360 12223
rect 1308 12180 1360 12189
rect 1676 12223 1728 12232
rect 1676 12189 1678 12223
rect 1678 12189 1728 12223
rect 1676 12180 1728 12189
rect 1860 12180 1912 12232
rect 1952 12180 2004 12232
rect 3332 12180 3384 12232
rect 4160 12248 4212 12300
rect 5080 12180 5132 12232
rect 1584 12044 1636 12096
rect 1768 12044 1820 12096
rect 6000 12044 6052 12096
rect 6092 12087 6144 12096
rect 6092 12053 6101 12087
rect 6101 12053 6135 12087
rect 6135 12053 6144 12087
rect 6092 12044 6144 12053
rect 6368 12248 6420 12300
rect 6828 12384 6880 12436
rect 7196 12384 7248 12436
rect 7472 12384 7524 12436
rect 7932 12384 7984 12436
rect 8576 12384 8628 12436
rect 8760 12384 8812 12436
rect 10048 12384 10100 12436
rect 10784 12384 10836 12436
rect 11336 12384 11388 12436
rect 6828 12223 6880 12232
rect 6828 12189 6830 12223
rect 6830 12189 6880 12223
rect 6828 12180 6880 12189
rect 6920 12223 6972 12232
rect 6920 12189 6932 12223
rect 6932 12189 6966 12223
rect 6966 12189 6972 12223
rect 6920 12180 6972 12189
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 9036 12223 9088 12232
rect 9036 12189 9038 12223
rect 9038 12189 9088 12223
rect 9036 12180 9088 12189
rect 10876 12248 10928 12300
rect 6736 12044 6788 12096
rect 8208 12044 8260 12096
rect 10416 12180 10468 12232
rect 11612 12316 11664 12368
rect 11980 12384 12032 12436
rect 12808 12384 12860 12436
rect 13636 12384 13688 12436
rect 14924 12384 14976 12436
rect 15292 12427 15344 12436
rect 15292 12393 15301 12427
rect 15301 12393 15335 12427
rect 15335 12393 15344 12427
rect 15292 12384 15344 12393
rect 15384 12384 15436 12436
rect 11796 12316 11848 12368
rect 17040 12384 17092 12436
rect 19156 12384 19208 12436
rect 20168 12384 20220 12436
rect 21088 12384 21140 12436
rect 21180 12384 21232 12436
rect 21548 12384 21600 12436
rect 22008 12384 22060 12436
rect 23388 12384 23440 12436
rect 24216 12384 24268 12436
rect 25780 12384 25832 12436
rect 26148 12384 26200 12436
rect 27436 12384 27488 12436
rect 27896 12384 27948 12436
rect 29000 12384 29052 12436
rect 12072 12248 12124 12300
rect 12532 12291 12584 12300
rect 12532 12257 12541 12291
rect 12541 12257 12575 12291
rect 12575 12257 12584 12291
rect 12532 12248 12584 12257
rect 13176 12248 13228 12300
rect 13728 12248 13780 12300
rect 13912 12248 13964 12300
rect 15108 12248 15160 12300
rect 15200 12291 15252 12300
rect 15200 12257 15209 12291
rect 15209 12257 15243 12291
rect 15243 12257 15252 12291
rect 15200 12248 15252 12257
rect 11520 12087 11572 12096
rect 11520 12053 11529 12087
rect 11529 12053 11563 12087
rect 11563 12053 11572 12087
rect 11520 12044 11572 12053
rect 16028 12248 16080 12300
rect 16396 12248 16448 12300
rect 17224 12291 17276 12300
rect 17224 12257 17233 12291
rect 17233 12257 17267 12291
rect 17267 12257 17276 12291
rect 17224 12248 17276 12257
rect 17592 12248 17644 12300
rect 12900 12044 12952 12096
rect 13084 12044 13136 12096
rect 13912 12044 13964 12096
rect 14372 12087 14424 12096
rect 14372 12053 14381 12087
rect 14381 12053 14415 12087
rect 14415 12053 14424 12087
rect 14372 12044 14424 12053
rect 14740 12087 14792 12096
rect 14740 12053 14749 12087
rect 14749 12053 14783 12087
rect 14783 12053 14792 12087
rect 14740 12044 14792 12053
rect 15016 12087 15068 12096
rect 15016 12053 15025 12087
rect 15025 12053 15059 12087
rect 15059 12053 15068 12087
rect 15016 12044 15068 12053
rect 15568 12112 15620 12164
rect 16396 12112 16448 12164
rect 18052 12223 18104 12232
rect 18052 12189 18061 12223
rect 18061 12189 18095 12223
rect 18095 12189 18104 12223
rect 18052 12180 18104 12189
rect 18512 12223 18564 12232
rect 18512 12189 18524 12223
rect 18524 12189 18558 12223
rect 18558 12189 18564 12223
rect 18512 12180 18564 12189
rect 18696 12248 18748 12300
rect 19248 12248 19300 12300
rect 21364 12248 21416 12300
rect 21548 12248 21600 12300
rect 23848 12248 23900 12300
rect 24124 12248 24176 12300
rect 25412 12248 25464 12300
rect 25964 12248 26016 12300
rect 26148 12248 26200 12300
rect 26424 12291 26476 12300
rect 26424 12257 26433 12291
rect 26433 12257 26467 12291
rect 26467 12257 26476 12291
rect 26424 12248 26476 12257
rect 28540 12248 28592 12300
rect 16580 12044 16632 12096
rect 17040 12087 17092 12096
rect 17040 12053 17049 12087
rect 17049 12053 17083 12087
rect 17083 12053 17092 12087
rect 17040 12044 17092 12053
rect 18880 12044 18932 12096
rect 19800 12180 19852 12232
rect 20352 12180 20404 12232
rect 21180 12044 21232 12096
rect 21732 12223 21784 12232
rect 21732 12189 21744 12223
rect 21744 12189 21778 12223
rect 21778 12189 21784 12223
rect 21732 12180 21784 12189
rect 21824 12180 21876 12232
rect 23020 12180 23072 12232
rect 23940 12223 23992 12232
rect 23940 12189 23952 12223
rect 23952 12189 23986 12223
rect 23986 12189 23992 12223
rect 23940 12180 23992 12189
rect 30472 12248 30524 12300
rect 26884 12223 26936 12232
rect 26884 12189 26896 12223
rect 26896 12189 26930 12223
rect 26930 12189 26936 12223
rect 26884 12180 26936 12189
rect 28080 12180 28132 12232
rect 21916 12044 21968 12096
rect 22652 12044 22704 12096
rect 29368 12180 29420 12232
rect 28816 12044 28868 12096
rect 4193 11942 4245 11994
rect 4257 11942 4309 11994
rect 4321 11942 4373 11994
rect 4385 11942 4437 11994
rect 4449 11942 4501 11994
rect 11783 11942 11835 11994
rect 11847 11942 11899 11994
rect 11911 11942 11963 11994
rect 11975 11942 12027 11994
rect 12039 11942 12091 11994
rect 19373 11942 19425 11994
rect 19437 11942 19489 11994
rect 19501 11942 19553 11994
rect 19565 11942 19617 11994
rect 19629 11942 19681 11994
rect 26963 11942 27015 11994
rect 27027 11942 27079 11994
rect 27091 11942 27143 11994
rect 27155 11942 27207 11994
rect 27219 11942 27271 11994
rect 4436 11840 4488 11892
rect 4988 11840 5040 11892
rect 5356 11883 5408 11892
rect 5356 11849 5365 11883
rect 5365 11849 5399 11883
rect 5399 11849 5408 11883
rect 5356 11840 5408 11849
rect 3240 11772 3292 11824
rect 1492 11704 1544 11756
rect 3700 11704 3752 11756
rect 3884 11704 3936 11756
rect 6092 11840 6144 11892
rect 7564 11840 7616 11892
rect 7380 11772 7432 11824
rect 5908 11704 5960 11756
rect 6092 11704 6144 11756
rect 1216 11636 1268 11688
rect 1768 11636 1820 11688
rect 3332 11679 3384 11688
rect 3332 11645 3341 11679
rect 3341 11645 3375 11679
rect 3375 11645 3384 11679
rect 3332 11636 3384 11645
rect 4804 11636 4856 11688
rect 5632 11636 5684 11688
rect 5816 11636 5868 11688
rect 7932 11679 7984 11688
rect 7932 11645 7941 11679
rect 7941 11645 7975 11679
rect 7975 11645 7984 11679
rect 7932 11636 7984 11645
rect 8208 11679 8260 11688
rect 8208 11645 8217 11679
rect 8217 11645 8251 11679
rect 8251 11645 8260 11679
rect 8208 11636 8260 11645
rect 3424 11568 3476 11620
rect 8576 11679 8628 11688
rect 8576 11645 8585 11679
rect 8585 11645 8619 11679
rect 8619 11645 8628 11679
rect 8576 11636 8628 11645
rect 8852 11704 8904 11756
rect 11520 11840 11572 11892
rect 11612 11840 11664 11892
rect 12716 11840 12768 11892
rect 16028 11840 16080 11892
rect 18512 11840 18564 11892
rect 13084 11772 13136 11824
rect 11520 11704 11572 11756
rect 12348 11704 12400 11756
rect 12440 11704 12492 11756
rect 13544 11772 13596 11824
rect 15108 11772 15160 11824
rect 16304 11772 16356 11824
rect 21732 11840 21784 11892
rect 21916 11840 21968 11892
rect 8760 11636 8812 11688
rect 11244 11679 11296 11688
rect 11244 11645 11253 11679
rect 11253 11645 11287 11679
rect 11287 11645 11296 11679
rect 11244 11636 11296 11645
rect 11612 11636 11664 11688
rect 11796 11636 11848 11688
rect 11888 11636 11940 11688
rect 14280 11747 14332 11756
rect 14280 11713 14289 11747
rect 14289 11713 14323 11747
rect 14323 11713 14332 11747
rect 14280 11704 14332 11713
rect 13544 11679 13596 11688
rect 13544 11645 13553 11679
rect 13553 11645 13587 11679
rect 13587 11645 13596 11679
rect 13544 11636 13596 11645
rect 13636 11636 13688 11688
rect 14556 11636 14608 11688
rect 15108 11636 15160 11688
rect 16764 11704 16816 11756
rect 16948 11704 17000 11756
rect 17040 11704 17092 11756
rect 20996 11772 21048 11824
rect 16672 11636 16724 11688
rect 18328 11636 18380 11688
rect 18880 11704 18932 11756
rect 19432 11747 19484 11756
rect 19432 11713 19441 11747
rect 19441 11713 19475 11747
rect 19475 11713 19484 11747
rect 19432 11704 19484 11713
rect 21916 11704 21968 11756
rect 18972 11636 19024 11688
rect 22284 11679 22336 11688
rect 22284 11645 22293 11679
rect 22293 11645 22327 11679
rect 22327 11645 22336 11679
rect 22284 11636 22336 11645
rect 22744 11636 22796 11688
rect 13360 11611 13412 11620
rect 13360 11577 13369 11611
rect 13369 11577 13403 11611
rect 13403 11577 13412 11611
rect 13360 11568 13412 11577
rect 1400 11543 1452 11552
rect 1400 11509 1415 11543
rect 1415 11509 1449 11543
rect 1449 11509 1452 11543
rect 1400 11500 1452 11509
rect 1768 11500 1820 11552
rect 3976 11500 4028 11552
rect 4896 11500 4948 11552
rect 5816 11500 5868 11552
rect 6000 11543 6052 11552
rect 6000 11509 6015 11543
rect 6015 11509 6049 11543
rect 6049 11509 6052 11543
rect 6000 11500 6052 11509
rect 7012 11500 7064 11552
rect 7748 11543 7800 11552
rect 7748 11509 7757 11543
rect 7757 11509 7791 11543
rect 7791 11509 7800 11543
rect 7748 11500 7800 11509
rect 8392 11543 8444 11552
rect 8392 11509 8401 11543
rect 8401 11509 8435 11543
rect 8435 11509 8444 11543
rect 8392 11500 8444 11509
rect 8852 11543 8904 11552
rect 8852 11509 8861 11543
rect 8861 11509 8895 11543
rect 8895 11509 8904 11543
rect 8852 11500 8904 11509
rect 9036 11500 9088 11552
rect 9404 11500 9456 11552
rect 12256 11500 12308 11552
rect 23940 11840 23992 11892
rect 24676 11840 24728 11892
rect 26516 11840 26568 11892
rect 26792 11840 26844 11892
rect 27528 11840 27580 11892
rect 28632 11883 28684 11892
rect 28632 11849 28641 11883
rect 28641 11849 28675 11883
rect 28675 11849 28684 11883
rect 28632 11840 28684 11849
rect 24124 11704 24176 11756
rect 24676 11679 24728 11688
rect 24676 11645 24685 11679
rect 24685 11645 24719 11679
rect 24719 11645 24728 11679
rect 24676 11636 24728 11645
rect 26056 11704 26108 11756
rect 28172 11704 28224 11756
rect 25688 11636 25740 11688
rect 24400 11568 24452 11620
rect 24768 11568 24820 11620
rect 15016 11500 15068 11552
rect 16120 11543 16172 11552
rect 16120 11509 16129 11543
rect 16129 11509 16163 11543
rect 16163 11509 16172 11543
rect 16120 11500 16172 11509
rect 17132 11500 17184 11552
rect 19156 11543 19208 11552
rect 19156 11509 19171 11543
rect 19171 11509 19205 11543
rect 19205 11509 19208 11543
rect 19156 11500 19208 11509
rect 22008 11543 22060 11552
rect 22008 11509 22023 11543
rect 22023 11509 22057 11543
rect 22057 11509 22060 11543
rect 22008 11500 22060 11509
rect 27528 11636 27580 11688
rect 27620 11636 27672 11688
rect 29644 11772 29696 11824
rect 26608 11500 26660 11552
rect 28264 11543 28316 11552
rect 28264 11509 28273 11543
rect 28273 11509 28307 11543
rect 28307 11509 28316 11543
rect 28264 11500 28316 11509
rect 28540 11500 28592 11552
rect 7988 11398 8040 11450
rect 8052 11398 8104 11450
rect 8116 11398 8168 11450
rect 8180 11398 8232 11450
rect 8244 11398 8296 11450
rect 15578 11398 15630 11450
rect 15642 11398 15694 11450
rect 15706 11398 15758 11450
rect 15770 11398 15822 11450
rect 15834 11398 15886 11450
rect 23168 11398 23220 11450
rect 23232 11398 23284 11450
rect 23296 11398 23348 11450
rect 23360 11398 23412 11450
rect 23424 11398 23476 11450
rect 30758 11398 30810 11450
rect 30822 11398 30874 11450
rect 30886 11398 30938 11450
rect 30950 11398 31002 11450
rect 31014 11398 31066 11450
rect 940 11296 992 11348
rect 2136 11296 2188 11348
rect 4528 11296 4580 11348
rect 4804 11339 4856 11348
rect 4804 11305 4813 11339
rect 4813 11305 4847 11339
rect 4847 11305 4856 11339
rect 4804 11296 4856 11305
rect 1400 11092 1452 11144
rect 1676 11092 1728 11144
rect 2136 11160 2188 11212
rect 3884 11228 3936 11280
rect 4436 11228 4488 11280
rect 4620 11228 4672 11280
rect 5080 11228 5132 11280
rect 5724 11296 5776 11348
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 5356 11160 5408 11212
rect 6368 11160 6420 11212
rect 6460 11160 6512 11212
rect 6736 11203 6788 11212
rect 6736 11169 6745 11203
rect 6745 11169 6779 11203
rect 6779 11169 6788 11203
rect 6736 11160 6788 11169
rect 8208 11296 8260 11348
rect 8668 11296 8720 11348
rect 9588 11296 9640 11348
rect 6000 11092 6052 11144
rect 6920 11092 6972 11144
rect 7748 11160 7800 11212
rect 8576 11160 8628 11212
rect 8944 11203 8996 11212
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 9496 11160 9548 11212
rect 11060 11228 11112 11280
rect 10508 11160 10560 11212
rect 10784 11160 10836 11212
rect 12072 11339 12124 11348
rect 12072 11305 12081 11339
rect 12081 11305 12115 11339
rect 12115 11305 12124 11339
rect 12072 11296 12124 11305
rect 12256 11296 12308 11348
rect 14740 11296 14792 11348
rect 9864 11092 9916 11144
rect 12348 11228 12400 11280
rect 3240 11024 3292 11076
rect 6368 11067 6420 11076
rect 6368 11033 6377 11067
rect 6377 11033 6411 11067
rect 6411 11033 6420 11067
rect 6368 11024 6420 11033
rect 12164 11092 12216 11144
rect 1860 10956 1912 11008
rect 3148 10956 3200 11008
rect 3792 10956 3844 11008
rect 4068 10956 4120 11008
rect 4620 10956 4672 11008
rect 4804 10956 4856 11008
rect 10140 11024 10192 11076
rect 10508 11067 10560 11076
rect 10508 11033 10517 11067
rect 10517 11033 10551 11067
rect 10551 11033 10560 11067
rect 10508 11024 10560 11033
rect 10968 11067 11020 11076
rect 10968 11033 10977 11067
rect 10977 11033 11011 11067
rect 11011 11033 11020 11067
rect 10968 11024 11020 11033
rect 11060 11024 11112 11076
rect 12440 11135 12492 11144
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 15108 11296 15160 11348
rect 16120 11296 16172 11348
rect 16304 11296 16356 11348
rect 17132 11296 17184 11348
rect 15384 11228 15436 11280
rect 15476 11203 15528 11212
rect 15476 11169 15485 11203
rect 15485 11169 15519 11203
rect 15519 11169 15528 11203
rect 15476 11160 15528 11169
rect 12440 11092 12492 11101
rect 13544 11092 13596 11144
rect 16028 11160 16080 11212
rect 18972 11296 19024 11348
rect 22284 11296 22336 11348
rect 22468 11296 22520 11348
rect 18972 11160 19024 11212
rect 19524 11160 19576 11212
rect 19800 11203 19852 11212
rect 19800 11169 19809 11203
rect 19809 11169 19843 11203
rect 19843 11169 19852 11203
rect 19800 11160 19852 11169
rect 21088 11228 21140 11280
rect 25688 11296 25740 11348
rect 26700 11296 26752 11348
rect 27436 11296 27488 11348
rect 20904 11160 20956 11212
rect 21824 11203 21876 11212
rect 21824 11169 21833 11203
rect 21833 11169 21867 11203
rect 21867 11169 21876 11203
rect 21824 11160 21876 11169
rect 22008 11160 22060 11212
rect 16672 11092 16724 11144
rect 12348 11024 12400 11076
rect 14188 11024 14240 11076
rect 14464 11024 14516 11076
rect 9128 10999 9180 11008
rect 9128 10965 9137 10999
rect 9137 10965 9171 10999
rect 9171 10965 9180 10999
rect 9128 10956 9180 10965
rect 9496 10956 9548 11008
rect 11244 10956 11296 11008
rect 11428 10999 11480 11008
rect 11428 10965 11437 10999
rect 11437 10965 11471 10999
rect 11471 10965 11480 10999
rect 11428 10956 11480 10965
rect 11520 10956 11572 11008
rect 14648 10999 14700 11008
rect 14648 10965 14657 10999
rect 14657 10965 14691 10999
rect 14691 10965 14700 10999
rect 14648 10956 14700 10965
rect 14924 11067 14976 11076
rect 14924 11033 14933 11067
rect 14933 11033 14967 11067
rect 14967 11033 14976 11067
rect 14924 11024 14976 11033
rect 20812 11092 20864 11144
rect 20996 11092 21048 11144
rect 22560 11092 22612 11144
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 24400 11092 24452 11144
rect 24768 11160 24820 11212
rect 24860 11135 24912 11144
rect 24860 11101 24869 11135
rect 24869 11101 24903 11135
rect 24903 11101 24912 11135
rect 24860 11092 24912 11101
rect 26332 11160 26384 11212
rect 28908 11203 28960 11212
rect 28908 11169 28917 11203
rect 28917 11169 28951 11203
rect 28951 11169 28960 11203
rect 28908 11160 28960 11169
rect 29368 11160 29420 11212
rect 30288 11160 30340 11212
rect 26424 11135 26476 11144
rect 26424 11101 26433 11135
rect 26433 11101 26467 11135
rect 26467 11101 26476 11135
rect 26424 11092 26476 11101
rect 26884 11135 26936 11144
rect 26884 11101 26896 11135
rect 26896 11101 26930 11135
rect 26930 11101 26936 11135
rect 26884 11092 26936 11101
rect 28540 11092 28592 11144
rect 17040 10956 17092 11008
rect 19524 10956 19576 11008
rect 19708 10956 19760 11008
rect 21548 10956 21600 11008
rect 22284 10956 22336 11008
rect 28080 11024 28132 11076
rect 30012 11067 30064 11076
rect 30012 11033 30021 11067
rect 30021 11033 30055 11067
rect 30055 11033 30064 11067
rect 30012 11024 30064 11033
rect 24032 10956 24084 11008
rect 29276 10956 29328 11008
rect 4193 10854 4245 10906
rect 4257 10854 4309 10906
rect 4321 10854 4373 10906
rect 4385 10854 4437 10906
rect 4449 10854 4501 10906
rect 11783 10854 11835 10906
rect 11847 10854 11899 10906
rect 11911 10854 11963 10906
rect 11975 10854 12027 10906
rect 12039 10854 12091 10906
rect 19373 10854 19425 10906
rect 19437 10854 19489 10906
rect 19501 10854 19553 10906
rect 19565 10854 19617 10906
rect 19629 10854 19681 10906
rect 26963 10854 27015 10906
rect 27027 10854 27079 10906
rect 27091 10854 27143 10906
rect 27155 10854 27207 10906
rect 27219 10854 27271 10906
rect 1308 10616 1360 10668
rect 2136 10616 2188 10668
rect 4620 10752 4672 10804
rect 3148 10616 3200 10668
rect 3700 10616 3752 10668
rect 5540 10659 5592 10668
rect 5540 10625 5549 10659
rect 5549 10625 5583 10659
rect 5583 10625 5592 10659
rect 5540 10616 5592 10625
rect 5816 10616 5868 10668
rect 6736 10616 6788 10668
rect 7840 10616 7892 10668
rect 1676 10412 1728 10464
rect 2964 10455 3016 10464
rect 2964 10421 2973 10455
rect 2973 10421 3007 10455
rect 3007 10421 3016 10455
rect 2964 10412 3016 10421
rect 4068 10548 4120 10600
rect 4620 10548 4672 10600
rect 6092 10548 6144 10600
rect 6276 10591 6328 10600
rect 6276 10557 6285 10591
rect 6285 10557 6319 10591
rect 6319 10557 6328 10591
rect 6276 10548 6328 10557
rect 6920 10548 6972 10600
rect 9680 10684 9732 10736
rect 11704 10795 11756 10804
rect 11704 10761 11713 10795
rect 11713 10761 11747 10795
rect 11747 10761 11756 10795
rect 11704 10752 11756 10761
rect 12992 10752 13044 10804
rect 15200 10752 15252 10804
rect 16396 10752 16448 10804
rect 16948 10752 17000 10804
rect 17868 10752 17920 10804
rect 9588 10616 9640 10668
rect 9864 10616 9916 10668
rect 10876 10616 10928 10668
rect 11244 10616 11296 10668
rect 12348 10684 12400 10736
rect 7380 10480 7432 10532
rect 8208 10480 8260 10532
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 9404 10480 9456 10532
rect 10232 10548 10284 10600
rect 13176 10684 13228 10736
rect 13360 10684 13412 10736
rect 20536 10752 20588 10804
rect 20720 10795 20772 10804
rect 20720 10761 20729 10795
rect 20729 10761 20763 10795
rect 20763 10761 20772 10795
rect 20720 10752 20772 10761
rect 12532 10548 12584 10600
rect 12624 10591 12676 10600
rect 12624 10557 12633 10591
rect 12633 10557 12667 10591
rect 12667 10557 12676 10591
rect 12624 10548 12676 10557
rect 14648 10616 14700 10668
rect 16580 10616 16632 10668
rect 13544 10591 13596 10600
rect 13544 10557 13553 10591
rect 13553 10557 13587 10591
rect 13587 10557 13596 10591
rect 13544 10548 13596 10557
rect 13820 10548 13872 10600
rect 15200 10548 15252 10600
rect 18144 10616 18196 10668
rect 18880 10616 18932 10668
rect 19340 10616 19392 10668
rect 22284 10752 22336 10804
rect 22652 10752 22704 10804
rect 24860 10752 24912 10804
rect 25136 10752 25188 10804
rect 25688 10752 25740 10804
rect 22744 10727 22796 10736
rect 22744 10693 22753 10727
rect 22753 10693 22787 10727
rect 22787 10693 22796 10727
rect 22744 10684 22796 10693
rect 18604 10548 18656 10600
rect 19248 10548 19300 10600
rect 19708 10548 19760 10600
rect 21548 10548 21600 10600
rect 21824 10616 21876 10668
rect 28264 10616 28316 10668
rect 3516 10412 3568 10464
rect 5632 10412 5684 10464
rect 6000 10455 6052 10464
rect 6000 10421 6015 10455
rect 6015 10421 6049 10455
rect 6049 10421 6052 10455
rect 6000 10412 6052 10421
rect 7656 10412 7708 10464
rect 10140 10412 10192 10464
rect 10876 10412 10928 10464
rect 24032 10591 24084 10600
rect 24032 10557 24041 10591
rect 24041 10557 24075 10591
rect 24075 10557 24084 10591
rect 24032 10548 24084 10557
rect 25320 10591 25372 10600
rect 25320 10557 25329 10591
rect 25329 10557 25363 10591
rect 25363 10557 25372 10591
rect 25320 10548 25372 10557
rect 25688 10548 25740 10600
rect 28540 10548 28592 10600
rect 29920 10752 29972 10804
rect 30288 10727 30340 10736
rect 30288 10693 30297 10727
rect 30297 10693 30331 10727
rect 30331 10693 30340 10727
rect 30288 10684 30340 10693
rect 29368 10616 29420 10668
rect 29460 10548 29512 10600
rect 26056 10480 26108 10532
rect 12164 10412 12216 10464
rect 12532 10412 12584 10464
rect 12900 10455 12952 10464
rect 12900 10421 12909 10455
rect 12909 10421 12943 10455
rect 12943 10421 12952 10455
rect 12900 10412 12952 10421
rect 13820 10412 13872 10464
rect 13912 10412 13964 10464
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 18788 10412 18840 10464
rect 19156 10455 19208 10464
rect 19156 10421 19171 10455
rect 19171 10421 19205 10455
rect 19205 10421 19208 10455
rect 19156 10412 19208 10421
rect 22468 10412 22520 10464
rect 22652 10412 22704 10464
rect 24124 10412 24176 10464
rect 24492 10412 24544 10464
rect 26240 10412 26292 10464
rect 26884 10480 26936 10532
rect 30472 10480 30524 10532
rect 29000 10412 29052 10464
rect 29736 10455 29788 10464
rect 29736 10421 29745 10455
rect 29745 10421 29779 10455
rect 29779 10421 29788 10455
rect 29736 10412 29788 10421
rect 7988 10310 8040 10362
rect 8052 10310 8104 10362
rect 8116 10310 8168 10362
rect 8180 10310 8232 10362
rect 8244 10310 8296 10362
rect 15578 10310 15630 10362
rect 15642 10310 15694 10362
rect 15706 10310 15758 10362
rect 15770 10310 15822 10362
rect 15834 10310 15886 10362
rect 23168 10310 23220 10362
rect 23232 10310 23284 10362
rect 23296 10310 23348 10362
rect 23360 10310 23412 10362
rect 23424 10310 23476 10362
rect 30758 10310 30810 10362
rect 30822 10310 30874 10362
rect 30886 10310 30938 10362
rect 30950 10310 31002 10362
rect 31014 10310 31066 10362
rect 940 10072 992 10124
rect 1308 10208 1360 10260
rect 1400 10208 1452 10260
rect 1676 10208 1728 10260
rect 3240 10208 3292 10260
rect 3884 10208 3936 10260
rect 5172 10208 5224 10260
rect 6920 10251 6972 10260
rect 6920 10217 6935 10251
rect 6935 10217 6969 10251
rect 6969 10217 6972 10251
rect 6920 10208 6972 10217
rect 8944 10208 8996 10260
rect 5356 10140 5408 10192
rect 6552 10140 6604 10192
rect 10140 10140 10192 10192
rect 11060 10140 11112 10192
rect 12624 10208 12676 10260
rect 16488 10208 16540 10260
rect 17132 10208 17184 10260
rect 18788 10208 18840 10260
rect 19248 10251 19300 10260
rect 19248 10217 19257 10251
rect 19257 10217 19291 10251
rect 19291 10217 19300 10251
rect 19248 10208 19300 10217
rect 20904 10208 20956 10260
rect 22008 10208 22060 10260
rect 22652 10208 22704 10260
rect 24032 10208 24084 10260
rect 24768 10208 24820 10260
rect 26700 10208 26752 10260
rect 26884 10251 26936 10260
rect 26884 10217 26899 10251
rect 26899 10217 26933 10251
rect 26933 10217 26936 10251
rect 26884 10208 26936 10217
rect 29920 10208 29972 10260
rect 1676 10004 1728 10056
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 2964 10004 3016 10056
rect 3240 10047 3292 10056
rect 3240 10013 3249 10047
rect 3249 10013 3283 10047
rect 3283 10013 3292 10047
rect 3240 10004 3292 10013
rect 3700 10047 3752 10056
rect 3700 10013 3712 10047
rect 3712 10013 3746 10047
rect 3746 10013 3752 10047
rect 3700 10004 3752 10013
rect 4160 10004 4212 10056
rect 5724 10004 5776 10056
rect 7288 10072 7340 10124
rect 6000 10004 6052 10056
rect 6828 10004 6880 10056
rect 7104 10004 7156 10056
rect 7564 10004 7616 10056
rect 9036 10047 9088 10056
rect 9036 10013 9038 10047
rect 9038 10013 9088 10047
rect 3056 9911 3108 9920
rect 3056 9877 3065 9911
rect 3065 9877 3099 9911
rect 3099 9877 3108 9911
rect 3056 9868 3108 9877
rect 3700 9868 3752 9920
rect 8484 9868 8536 9920
rect 8576 9868 8628 9920
rect 9036 10004 9088 10013
rect 10508 10072 10560 10124
rect 10692 10072 10744 10124
rect 10876 10004 10928 10056
rect 11336 10047 11388 10056
rect 11336 10013 11338 10047
rect 11338 10013 11388 10047
rect 11336 10004 11388 10013
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 13268 10183 13320 10192
rect 13268 10149 13277 10183
rect 13277 10149 13311 10183
rect 13311 10149 13320 10183
rect 13268 10140 13320 10149
rect 16396 10140 16448 10192
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 13912 10047 13964 10056
rect 13912 10013 13914 10047
rect 13914 10013 13964 10047
rect 13912 10004 13964 10013
rect 14372 10072 14424 10124
rect 15200 10072 15252 10124
rect 16672 10072 16724 10124
rect 17316 10140 17368 10192
rect 19984 10140 20036 10192
rect 20996 10140 21048 10192
rect 21272 10140 21324 10192
rect 17040 10072 17092 10124
rect 20260 10072 20312 10124
rect 21088 10072 21140 10124
rect 17960 10047 18012 10056
rect 17960 10013 17969 10047
rect 17969 10013 18003 10047
rect 18003 10013 18012 10047
rect 17960 10004 18012 10013
rect 18052 10004 18104 10056
rect 17132 9936 17184 9988
rect 21272 10047 21324 10056
rect 21272 10013 21281 10047
rect 21281 10013 21315 10047
rect 21315 10013 21324 10047
rect 21272 10004 21324 10013
rect 21732 10047 21784 10056
rect 21732 10013 21744 10047
rect 21744 10013 21778 10047
rect 21778 10013 21784 10047
rect 21732 10004 21784 10013
rect 21916 10004 21968 10056
rect 23756 10072 23808 10124
rect 24492 10115 24544 10124
rect 24492 10081 24494 10115
rect 24494 10081 24544 10115
rect 24492 10072 24544 10081
rect 24124 10047 24176 10056
rect 9496 9868 9548 9920
rect 11152 9868 11204 9920
rect 12348 9868 12400 9920
rect 12900 9868 12952 9920
rect 15292 9868 15344 9920
rect 15476 9868 15528 9920
rect 17960 9868 18012 9920
rect 20996 9911 21048 9920
rect 20996 9877 21005 9911
rect 21005 9877 21039 9911
rect 21039 9877 21048 9911
rect 20996 9868 21048 9877
rect 24124 10013 24133 10047
rect 24133 10013 24167 10047
rect 24167 10013 24176 10047
rect 24124 10004 24176 10013
rect 24952 10072 25004 10124
rect 24676 10004 24728 10056
rect 26424 10047 26476 10056
rect 26424 10013 26433 10047
rect 26433 10013 26467 10047
rect 26467 10013 26476 10047
rect 26424 10004 26476 10013
rect 29184 10072 29236 10124
rect 28264 10004 28316 10056
rect 28816 10004 28868 10056
rect 24676 9868 24728 9920
rect 28448 9911 28500 9920
rect 28448 9877 28457 9911
rect 28457 9877 28491 9911
rect 28491 9877 28500 9911
rect 28448 9868 28500 9877
rect 30012 9911 30064 9920
rect 30012 9877 30021 9911
rect 30021 9877 30055 9911
rect 30055 9877 30064 9911
rect 30012 9868 30064 9877
rect 30104 9868 30156 9920
rect 4193 9766 4245 9818
rect 4257 9766 4309 9818
rect 4321 9766 4373 9818
rect 4385 9766 4437 9818
rect 4449 9766 4501 9818
rect 11783 9766 11835 9818
rect 11847 9766 11899 9818
rect 11911 9766 11963 9818
rect 11975 9766 12027 9818
rect 12039 9766 12091 9818
rect 19373 9766 19425 9818
rect 19437 9766 19489 9818
rect 19501 9766 19553 9818
rect 19565 9766 19617 9818
rect 19629 9766 19681 9818
rect 26963 9766 27015 9818
rect 27027 9766 27079 9818
rect 27091 9766 27143 9818
rect 27155 9766 27207 9818
rect 27219 9766 27271 9818
rect 1124 9664 1176 9716
rect 1768 9664 1820 9716
rect 1860 9664 1912 9716
rect 5448 9664 5500 9716
rect 5816 9664 5868 9716
rect 940 9571 992 9580
rect 940 9537 949 9571
rect 949 9537 983 9571
rect 983 9537 992 9571
rect 940 9528 992 9537
rect 1584 9460 1636 9512
rect 1400 9367 1452 9376
rect 1400 9333 1415 9367
rect 1415 9333 1449 9367
rect 1449 9333 1452 9367
rect 1400 9324 1452 9333
rect 3056 9528 3108 9580
rect 3884 9528 3936 9580
rect 4712 9528 4764 9580
rect 5264 9528 5316 9580
rect 7288 9664 7340 9716
rect 8484 9664 8536 9716
rect 8760 9664 8812 9716
rect 10692 9664 10744 9716
rect 10968 9664 11020 9716
rect 11704 9664 11756 9716
rect 11888 9664 11940 9716
rect 3240 9460 3292 9512
rect 3608 9460 3660 9512
rect 6552 9571 6604 9580
rect 6552 9537 6564 9571
rect 6564 9537 6598 9571
rect 6598 9537 6604 9571
rect 6552 9528 6604 9537
rect 8392 9528 8444 9580
rect 8576 9571 8628 9580
rect 8576 9537 8585 9571
rect 8585 9537 8619 9571
rect 8619 9537 8628 9571
rect 8576 9528 8628 9537
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 4988 9392 5040 9444
rect 3700 9324 3752 9376
rect 3976 9324 4028 9376
rect 4712 9324 4764 9376
rect 5632 9324 5684 9376
rect 6736 9460 6788 9512
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 10784 9528 10836 9537
rect 9312 9503 9364 9512
rect 9312 9469 9321 9503
rect 9321 9469 9355 9503
rect 9355 9469 9364 9503
rect 9312 9460 9364 9469
rect 9404 9460 9456 9512
rect 11244 9571 11296 9580
rect 11244 9537 11256 9571
rect 11256 9537 11290 9571
rect 11290 9537 11296 9571
rect 11244 9528 11296 9537
rect 11336 9528 11388 9580
rect 13084 9528 13136 9580
rect 13544 9571 13596 9580
rect 13544 9537 13553 9571
rect 13553 9537 13587 9571
rect 13587 9537 13596 9571
rect 13544 9528 13596 9537
rect 13820 9528 13872 9580
rect 15016 9528 15068 9580
rect 11520 9503 11572 9512
rect 11520 9469 11529 9503
rect 11529 9469 11563 9503
rect 11563 9469 11572 9503
rect 11520 9460 11572 9469
rect 11612 9460 11664 9512
rect 17224 9664 17276 9716
rect 17592 9664 17644 9716
rect 18052 9664 18104 9716
rect 18604 9664 18656 9716
rect 24032 9664 24084 9716
rect 24124 9664 24176 9716
rect 22560 9596 22612 9648
rect 16764 9503 16816 9512
rect 16764 9469 16766 9503
rect 16766 9469 16816 9503
rect 6460 9324 6512 9376
rect 6920 9324 6972 9376
rect 7748 9324 7800 9376
rect 8944 9324 8996 9376
rect 9036 9367 9088 9376
rect 9036 9333 9051 9367
rect 9051 9333 9085 9367
rect 9085 9333 9088 9367
rect 9036 9324 9088 9333
rect 9588 9324 9640 9376
rect 10784 9324 10836 9376
rect 12440 9324 12492 9376
rect 13912 9324 13964 9376
rect 15016 9324 15068 9376
rect 16120 9367 16172 9376
rect 16120 9333 16129 9367
rect 16129 9333 16163 9367
rect 16163 9333 16172 9367
rect 16120 9324 16172 9333
rect 16304 9324 16356 9376
rect 16764 9460 16816 9469
rect 19248 9528 19300 9580
rect 19432 9571 19484 9580
rect 19432 9537 19441 9571
rect 19441 9537 19475 9571
rect 19475 9537 19484 9571
rect 19432 9528 19484 9537
rect 20812 9571 20864 9580
rect 20812 9537 20821 9571
rect 20821 9537 20855 9571
rect 20855 9537 20864 9571
rect 20812 9528 20864 9537
rect 21732 9528 21784 9580
rect 17040 9460 17092 9512
rect 17132 9503 17184 9512
rect 17132 9469 17141 9503
rect 17141 9469 17175 9503
rect 17175 9469 17184 9503
rect 17132 9460 17184 9469
rect 18696 9503 18748 9512
rect 18696 9469 18705 9503
rect 18705 9469 18739 9503
rect 18739 9469 18748 9503
rect 18696 9460 18748 9469
rect 20996 9460 21048 9512
rect 21640 9503 21692 9512
rect 21640 9469 21649 9503
rect 21649 9469 21683 9503
rect 21683 9469 21692 9503
rect 21640 9460 21692 9469
rect 21916 9460 21968 9512
rect 23756 9460 23808 9512
rect 24124 9528 24176 9580
rect 25688 9707 25740 9716
rect 25688 9673 25697 9707
rect 25697 9673 25731 9707
rect 25731 9673 25740 9707
rect 25688 9664 25740 9673
rect 28264 9707 28316 9716
rect 28264 9673 28273 9707
rect 28273 9673 28307 9707
rect 28307 9673 28316 9707
rect 28264 9664 28316 9673
rect 26240 9528 26292 9580
rect 24492 9460 24544 9512
rect 25688 9460 25740 9512
rect 26700 9528 26752 9580
rect 28816 9596 28868 9648
rect 26792 9503 26844 9512
rect 26792 9469 26801 9503
rect 26801 9469 26835 9503
rect 26835 9469 26844 9503
rect 26792 9460 26844 9469
rect 29000 9528 29052 9580
rect 16672 9324 16724 9376
rect 16856 9324 16908 9376
rect 17592 9324 17644 9376
rect 17776 9324 17828 9376
rect 19064 9324 19116 9376
rect 23020 9324 23072 9376
rect 23664 9324 23716 9376
rect 23940 9392 23992 9444
rect 25872 9392 25924 9444
rect 24216 9324 24268 9376
rect 24492 9324 24544 9376
rect 29736 9596 29788 9648
rect 29184 9460 29236 9512
rect 30472 9503 30524 9512
rect 30472 9469 30481 9503
rect 30481 9469 30515 9503
rect 30515 9469 30524 9503
rect 30472 9460 30524 9469
rect 27896 9367 27948 9376
rect 27896 9333 27905 9367
rect 27905 9333 27939 9367
rect 27939 9333 27948 9367
rect 27896 9324 27948 9333
rect 28540 9367 28592 9376
rect 28540 9333 28549 9367
rect 28549 9333 28583 9367
rect 28583 9333 28592 9367
rect 28540 9324 28592 9333
rect 30288 9367 30340 9376
rect 30288 9333 30297 9367
rect 30297 9333 30331 9367
rect 30331 9333 30340 9367
rect 30288 9324 30340 9333
rect 7988 9222 8040 9274
rect 8052 9222 8104 9274
rect 8116 9222 8168 9274
rect 8180 9222 8232 9274
rect 8244 9222 8296 9274
rect 15578 9222 15630 9274
rect 15642 9222 15694 9274
rect 15706 9222 15758 9274
rect 15770 9222 15822 9274
rect 15834 9222 15886 9274
rect 23168 9222 23220 9274
rect 23232 9222 23284 9274
rect 23296 9222 23348 9274
rect 23360 9222 23412 9274
rect 23424 9222 23476 9274
rect 30758 9222 30810 9274
rect 30822 9222 30874 9274
rect 30886 9222 30938 9274
rect 30950 9222 31002 9274
rect 31014 9222 31066 9274
rect 2964 9120 3016 9172
rect 3976 9120 4028 9172
rect 5264 9052 5316 9104
rect 5908 9052 5960 9104
rect 6736 9120 6788 9172
rect 7196 9120 7248 9172
rect 848 8916 900 8968
rect 1400 8959 1452 8968
rect 1400 8925 1402 8959
rect 1402 8925 1452 8959
rect 1400 8916 1452 8925
rect 1768 8959 1820 8968
rect 1768 8925 1777 8959
rect 1777 8925 1811 8959
rect 1811 8925 1820 8959
rect 1768 8916 1820 8925
rect 940 8780 992 8832
rect 2412 8780 2464 8832
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 6184 8984 6236 9036
rect 6368 9027 6420 9036
rect 6368 8993 6377 9027
rect 6377 8993 6411 9027
rect 6411 8993 6420 9027
rect 6368 8984 6420 8993
rect 6460 8984 6512 9036
rect 6736 9027 6788 9036
rect 6736 8993 6745 9027
rect 6745 8993 6779 9027
rect 6779 8993 6788 9027
rect 6736 8984 6788 8993
rect 7288 8984 7340 9036
rect 7472 9027 7524 9036
rect 7472 8993 7481 9027
rect 7481 8993 7515 9027
rect 7515 8993 7524 9027
rect 7472 8984 7524 8993
rect 9312 9120 9364 9172
rect 9404 9163 9456 9172
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 10324 9163 10376 9172
rect 10324 9129 10333 9163
rect 10333 9129 10367 9163
rect 10367 9129 10376 9163
rect 10324 9120 10376 9129
rect 11520 9120 11572 9172
rect 14740 9120 14792 9172
rect 16856 9120 16908 9172
rect 17592 9120 17644 9172
rect 19432 9120 19484 9172
rect 21640 9120 21692 9172
rect 12716 9052 12768 9104
rect 15200 9052 15252 9104
rect 15568 9052 15620 9104
rect 10416 8984 10468 9036
rect 10600 8984 10652 9036
rect 11336 9027 11388 9036
rect 11336 8993 11338 9027
rect 11338 8993 11388 9027
rect 5264 8848 5316 8900
rect 6828 8916 6880 8968
rect 6920 8959 6972 8968
rect 6920 8925 6929 8959
rect 6929 8925 6963 8959
rect 6963 8925 6972 8959
rect 6920 8916 6972 8925
rect 7380 8916 7432 8968
rect 7748 8916 7800 8968
rect 8024 8959 8076 8968
rect 8024 8925 8036 8959
rect 8036 8925 8070 8959
rect 8070 8925 8076 8959
rect 8024 8916 8076 8925
rect 8208 8916 8260 8968
rect 10048 8916 10100 8968
rect 10324 8916 10376 8968
rect 11336 8984 11388 8993
rect 11612 8984 11664 9036
rect 13084 8984 13136 9036
rect 13912 9027 13964 9036
rect 13912 8993 13914 9027
rect 13914 8993 13964 9027
rect 13912 8984 13964 8993
rect 14924 8984 14976 9036
rect 11152 8916 11204 8968
rect 11520 8916 11572 8968
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 16672 9052 16724 9104
rect 14096 8916 14148 8968
rect 15844 8916 15896 8968
rect 16764 9027 16816 9036
rect 16764 8993 16773 9027
rect 16773 8993 16807 9027
rect 16807 8993 16816 9027
rect 16764 8984 16816 8993
rect 19064 9052 19116 9104
rect 20996 9052 21048 9104
rect 21824 9052 21876 9104
rect 17960 8984 18012 9036
rect 19248 9027 19300 9036
rect 19248 8993 19257 9027
rect 19257 8993 19291 9027
rect 19291 8993 19300 9027
rect 19248 8984 19300 8993
rect 20168 8984 20220 9036
rect 16488 8916 16540 8968
rect 17132 8916 17184 8968
rect 17408 8916 17460 8968
rect 17776 8916 17828 8968
rect 18420 8916 18472 8968
rect 19800 8916 19852 8968
rect 5356 8780 5408 8832
rect 5448 8823 5500 8832
rect 5448 8789 5457 8823
rect 5457 8789 5491 8823
rect 5491 8789 5500 8823
rect 5448 8780 5500 8789
rect 6184 8823 6236 8832
rect 6184 8789 6193 8823
rect 6193 8789 6227 8823
rect 6227 8789 6236 8823
rect 6184 8780 6236 8789
rect 6460 8823 6512 8832
rect 6460 8789 6469 8823
rect 6469 8789 6503 8823
rect 6503 8789 6512 8823
rect 6460 8780 6512 8789
rect 10232 8848 10284 8900
rect 10416 8848 10468 8900
rect 10876 8780 10928 8832
rect 11336 8780 11388 8832
rect 12808 8823 12860 8832
rect 12808 8789 12817 8823
rect 12817 8789 12851 8823
rect 12851 8789 12860 8823
rect 12808 8780 12860 8789
rect 13360 8823 13412 8832
rect 13360 8789 13369 8823
rect 13369 8789 13403 8823
rect 13403 8789 13412 8823
rect 13360 8780 13412 8789
rect 13728 8780 13780 8832
rect 18328 8848 18380 8900
rect 18972 8848 19024 8900
rect 20904 8984 20956 9036
rect 22836 9027 22888 9036
rect 22836 8993 22845 9027
rect 22845 8993 22879 9027
rect 22879 8993 22888 9027
rect 22836 8984 22888 8993
rect 23940 9120 23992 9172
rect 25688 9163 25740 9172
rect 25688 9129 25697 9163
rect 25697 9129 25731 9163
rect 25731 9129 25740 9163
rect 25688 9120 25740 9129
rect 26792 9120 26844 9172
rect 26884 9163 26936 9172
rect 26884 9129 26899 9163
rect 26899 9129 26933 9163
rect 26933 9129 26936 9163
rect 26884 9120 26936 9129
rect 27896 9120 27948 9172
rect 28540 9120 28592 9172
rect 31116 9120 31168 9172
rect 23020 9052 23072 9104
rect 24860 9052 24912 9104
rect 23664 9027 23716 9036
rect 23664 8993 23673 9027
rect 23673 8993 23707 9027
rect 23707 8993 23716 9027
rect 23664 8984 23716 8993
rect 23756 8984 23808 9036
rect 25780 8984 25832 9036
rect 25964 8984 26016 9036
rect 26148 9027 26200 9036
rect 26148 8993 26157 9027
rect 26157 8993 26191 9027
rect 26191 8993 26200 9027
rect 26148 8984 26200 8993
rect 26424 9027 26476 9036
rect 26424 8993 26433 9027
rect 26433 8993 26467 9027
rect 26467 8993 26476 9027
rect 26424 8984 26476 8993
rect 26700 8984 26752 9036
rect 20536 8916 20588 8968
rect 22744 8916 22796 8968
rect 23572 8916 23624 8968
rect 23848 8916 23900 8968
rect 28172 8848 28224 8900
rect 30012 8984 30064 9036
rect 15200 8780 15252 8832
rect 16120 8823 16172 8832
rect 16120 8789 16129 8823
rect 16129 8789 16163 8823
rect 16163 8789 16172 8823
rect 16120 8780 16172 8789
rect 16672 8780 16724 8832
rect 17776 8780 17828 8832
rect 18788 8780 18840 8832
rect 22192 8780 22244 8832
rect 24492 8780 24544 8832
rect 24952 8823 25004 8832
rect 24952 8789 24961 8823
rect 24961 8789 24995 8823
rect 24995 8789 25004 8823
rect 24952 8780 25004 8789
rect 26884 8780 26936 8832
rect 27528 8780 27580 8832
rect 27896 8780 27948 8832
rect 28264 8823 28316 8832
rect 28264 8789 28273 8823
rect 28273 8789 28307 8823
rect 28307 8789 28316 8823
rect 28264 8780 28316 8789
rect 4193 8678 4245 8730
rect 4257 8678 4309 8730
rect 4321 8678 4373 8730
rect 4385 8678 4437 8730
rect 4449 8678 4501 8730
rect 11783 8678 11835 8730
rect 11847 8678 11899 8730
rect 11911 8678 11963 8730
rect 11975 8678 12027 8730
rect 12039 8678 12091 8730
rect 19373 8678 19425 8730
rect 19437 8678 19489 8730
rect 19501 8678 19553 8730
rect 19565 8678 19617 8730
rect 19629 8678 19681 8730
rect 26963 8678 27015 8730
rect 27027 8678 27079 8730
rect 27091 8678 27143 8730
rect 27155 8678 27207 8730
rect 27219 8678 27271 8730
rect 2044 8576 2096 8628
rect 2964 8576 3016 8628
rect 2412 8508 2464 8560
rect 5172 8551 5224 8560
rect 5172 8517 5181 8551
rect 5181 8517 5215 8551
rect 5215 8517 5224 8551
rect 5172 8508 5224 8517
rect 7104 8576 7156 8628
rect 7564 8576 7616 8628
rect 8944 8576 8996 8628
rect 3148 8440 3200 8492
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 3976 8440 4028 8492
rect 5264 8440 5316 8492
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 5724 8440 5776 8492
rect 6368 8440 6420 8492
rect 7012 8440 7064 8492
rect 11520 8619 11572 8628
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 11612 8576 11664 8628
rect 848 8372 900 8424
rect 2964 8372 3016 8424
rect 2780 8304 2832 8356
rect 3608 8372 3660 8424
rect 5448 8304 5500 8356
rect 7104 8372 7156 8424
rect 7656 8372 7708 8424
rect 10692 8440 10744 8492
rect 11152 8440 11204 8492
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 14188 8440 14240 8492
rect 15476 8440 15528 8492
rect 18144 8576 18196 8628
rect 18236 8619 18288 8628
rect 18236 8585 18245 8619
rect 18245 8585 18279 8619
rect 18279 8585 18288 8619
rect 18236 8576 18288 8585
rect 21548 8576 21600 8628
rect 21732 8576 21784 8628
rect 22836 8576 22888 8628
rect 8208 8415 8260 8424
rect 8208 8381 8217 8415
rect 8217 8381 8251 8415
rect 8251 8381 8260 8415
rect 8208 8372 8260 8381
rect 1400 8279 1452 8288
rect 1400 8245 1415 8279
rect 1415 8245 1449 8279
rect 1449 8245 1452 8279
rect 1400 8236 1452 8245
rect 6000 8279 6052 8288
rect 6000 8245 6015 8279
rect 6015 8245 6049 8279
rect 6049 8245 6052 8279
rect 6000 8236 6052 8245
rect 6368 8236 6420 8288
rect 6920 8236 6972 8288
rect 7288 8304 7340 8356
rect 7840 8304 7892 8356
rect 8668 8372 8720 8424
rect 9404 8372 9456 8424
rect 9496 8415 9548 8424
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 9588 8372 9640 8424
rect 10600 8372 10652 8424
rect 12624 8415 12676 8424
rect 12624 8381 12633 8415
rect 12633 8381 12667 8415
rect 12667 8381 12676 8415
rect 12624 8372 12676 8381
rect 12716 8372 12768 8424
rect 13084 8372 13136 8424
rect 15568 8372 15620 8424
rect 7104 8236 7156 8288
rect 9128 8236 9180 8288
rect 10968 8304 11020 8356
rect 11244 8304 11296 8356
rect 12164 8304 12216 8356
rect 13820 8236 13872 8288
rect 15844 8236 15896 8288
rect 16212 8236 16264 8288
rect 17224 8372 17276 8424
rect 17776 8236 17828 8288
rect 17960 8440 18012 8492
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 19064 8483 19116 8492
rect 19064 8449 19066 8483
rect 19066 8449 19116 8483
rect 19064 8440 19116 8449
rect 23756 8508 23808 8560
rect 18788 8372 18840 8424
rect 19708 8372 19760 8424
rect 20720 8372 20772 8424
rect 20812 8372 20864 8424
rect 20444 8304 20496 8356
rect 21732 8372 21784 8424
rect 24492 8440 24544 8492
rect 25320 8576 25372 8628
rect 26332 8619 26384 8628
rect 26332 8585 26341 8619
rect 26341 8585 26375 8619
rect 26375 8585 26384 8619
rect 26332 8576 26384 8585
rect 26516 8576 26568 8628
rect 27620 8576 27672 8628
rect 27804 8576 27856 8628
rect 28632 8576 28684 8628
rect 29276 8576 29328 8628
rect 30196 8576 30248 8628
rect 25872 8551 25924 8560
rect 25872 8517 25881 8551
rect 25881 8517 25915 8551
rect 25915 8517 25924 8551
rect 25872 8508 25924 8517
rect 29644 8508 29696 8560
rect 23940 8372 23992 8424
rect 24216 8415 24268 8424
rect 24216 8381 24218 8415
rect 24218 8381 24268 8415
rect 24216 8372 24268 8381
rect 24676 8372 24728 8424
rect 25964 8372 26016 8424
rect 23664 8304 23716 8356
rect 23756 8304 23808 8356
rect 25872 8236 25924 8288
rect 26884 8440 26936 8492
rect 28080 8440 28132 8492
rect 26424 8304 26476 8356
rect 27436 8415 27488 8424
rect 27436 8381 27445 8415
rect 27445 8381 27479 8415
rect 27479 8381 27488 8415
rect 27436 8372 27488 8381
rect 29368 8440 29420 8492
rect 28356 8372 28408 8424
rect 29092 8415 29144 8424
rect 29092 8381 29101 8415
rect 29101 8381 29135 8415
rect 29135 8381 29144 8415
rect 29092 8372 29144 8381
rect 29092 8236 29144 8288
rect 7988 8134 8040 8186
rect 8052 8134 8104 8186
rect 8116 8134 8168 8186
rect 8180 8134 8232 8186
rect 8244 8134 8296 8186
rect 15578 8134 15630 8186
rect 15642 8134 15694 8186
rect 15706 8134 15758 8186
rect 15770 8134 15822 8186
rect 15834 8134 15886 8186
rect 23168 8134 23220 8186
rect 23232 8134 23284 8186
rect 23296 8134 23348 8186
rect 23360 8134 23412 8186
rect 23424 8134 23476 8186
rect 30758 8134 30810 8186
rect 30822 8134 30874 8186
rect 30886 8134 30938 8186
rect 30950 8134 31002 8186
rect 31014 8134 31066 8186
rect 5172 8032 5224 8084
rect 5448 8075 5500 8084
rect 5448 8041 5457 8075
rect 5457 8041 5491 8075
rect 5491 8041 5500 8075
rect 5448 8032 5500 8041
rect 5724 8032 5776 8084
rect 3332 7896 3384 7948
rect 4804 7896 4856 7948
rect 5356 7964 5408 8016
rect 10508 7964 10560 8016
rect 5908 7896 5960 7948
rect 6000 7939 6052 7948
rect 6000 7905 6009 7939
rect 6009 7905 6043 7939
rect 6043 7905 6052 7939
rect 6000 7896 6052 7905
rect 8392 7939 8444 7948
rect 848 7828 900 7880
rect 1400 7871 1452 7880
rect 1400 7837 1402 7871
rect 1402 7837 1452 7871
rect 1400 7828 1452 7837
rect 1676 7828 1728 7880
rect 2596 7828 2648 7880
rect 3424 7828 3476 7880
rect 3608 7871 3660 7880
rect 3608 7837 3610 7871
rect 3610 7837 3660 7871
rect 3608 7828 3660 7837
rect 8392 7905 8401 7939
rect 8401 7905 8435 7939
rect 8435 7905 8444 7939
rect 8392 7896 8444 7905
rect 5908 7760 5960 7812
rect 6368 7828 6420 7880
rect 6736 7828 6788 7880
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 8760 7871 8812 7880
rect 8760 7837 8762 7871
rect 8762 7837 8812 7871
rect 8760 7828 8812 7837
rect 9312 7828 9364 7880
rect 10600 7803 10652 7812
rect 10600 7769 10609 7803
rect 10609 7769 10643 7803
rect 10643 7769 10652 7803
rect 10600 7760 10652 7769
rect 11244 7828 11296 7880
rect 12256 8032 12308 8084
rect 13452 8075 13504 8084
rect 13452 8041 13461 8075
rect 13461 8041 13495 8075
rect 13495 8041 13504 8075
rect 13452 8032 13504 8041
rect 13820 8032 13872 8084
rect 14096 8032 14148 8084
rect 14556 8032 14608 8084
rect 16120 8032 16172 8084
rect 16212 8032 16264 8084
rect 11704 7896 11756 7948
rect 16028 7964 16080 8016
rect 17500 8007 17552 8016
rect 17500 7973 17509 8007
rect 17509 7973 17543 8007
rect 17543 7973 17552 8007
rect 17500 7964 17552 7973
rect 18144 8032 18196 8084
rect 19892 8075 19944 8084
rect 19892 8041 19901 8075
rect 19901 8041 19935 8075
rect 19935 8041 19944 8075
rect 19892 8032 19944 8041
rect 20444 8075 20496 8084
rect 20444 8041 20453 8075
rect 20453 8041 20487 8075
rect 20487 8041 20496 8075
rect 20444 8032 20496 8041
rect 21456 8032 21508 8084
rect 23572 8075 23624 8084
rect 23572 8041 23581 8075
rect 23581 8041 23615 8075
rect 23615 8041 23624 8075
rect 23572 8032 23624 8041
rect 14556 7939 14608 7948
rect 14556 7905 14565 7939
rect 14565 7905 14599 7939
rect 14599 7905 14608 7939
rect 14556 7896 14608 7905
rect 16396 7939 16448 7948
rect 16396 7905 16405 7939
rect 16405 7905 16439 7939
rect 16439 7905 16448 7939
rect 16396 7896 16448 7905
rect 17592 7896 17644 7948
rect 17776 7896 17828 7948
rect 2964 7692 3016 7744
rect 5172 7692 5224 7744
rect 6552 7692 6604 7744
rect 9772 7692 9824 7744
rect 10232 7735 10284 7744
rect 10232 7701 10241 7735
rect 10241 7701 10275 7735
rect 10275 7701 10284 7735
rect 10232 7692 10284 7701
rect 13176 7692 13228 7744
rect 13820 7871 13872 7880
rect 13820 7837 13829 7871
rect 13829 7837 13863 7871
rect 13863 7837 13872 7871
rect 13820 7828 13872 7837
rect 15292 7828 15344 7880
rect 16764 7828 16816 7880
rect 17960 7828 18012 7880
rect 20904 7896 20956 7948
rect 21456 7939 21508 7948
rect 21456 7905 21475 7939
rect 21475 7905 21508 7939
rect 18788 7871 18840 7880
rect 18788 7837 18797 7871
rect 18797 7837 18831 7871
rect 18831 7837 18840 7871
rect 18788 7828 18840 7837
rect 16120 7760 16172 7812
rect 21456 7896 21508 7905
rect 21640 7896 21692 7948
rect 22560 7896 22612 7948
rect 21180 7760 21232 7812
rect 21456 7760 21508 7812
rect 21732 7828 21784 7880
rect 21916 7871 21968 7880
rect 21916 7837 21918 7871
rect 21918 7837 21968 7871
rect 21916 7828 21968 7837
rect 22008 7828 22060 7880
rect 23664 7828 23716 7880
rect 24492 7871 24544 7880
rect 24492 7837 24494 7871
rect 24494 7837 24544 7871
rect 24492 7828 24544 7837
rect 26608 7896 26660 7948
rect 27620 7896 27672 7948
rect 28172 8032 28224 8084
rect 28632 8032 28684 8084
rect 28908 8032 28960 8084
rect 30196 8032 30248 8084
rect 27896 7964 27948 8016
rect 28448 7896 28500 7948
rect 30104 7896 30156 7948
rect 26792 7828 26844 7880
rect 27804 7871 27856 7880
rect 27804 7837 27813 7871
rect 27813 7837 27847 7871
rect 27847 7837 27856 7871
rect 27804 7828 27856 7837
rect 29000 7828 29052 7880
rect 29552 7828 29604 7880
rect 15292 7692 15344 7744
rect 16488 7692 16540 7744
rect 16764 7692 16816 7744
rect 16948 7692 17000 7744
rect 18604 7692 18656 7744
rect 20812 7692 20864 7744
rect 21548 7692 21600 7744
rect 21732 7692 21784 7744
rect 24676 7692 24728 7744
rect 24768 7692 24820 7744
rect 27436 7692 27488 7744
rect 27528 7735 27580 7744
rect 27528 7701 27537 7735
rect 27537 7701 27571 7735
rect 27571 7701 27580 7735
rect 27528 7692 27580 7701
rect 28448 7692 28500 7744
rect 28632 7692 28684 7744
rect 30104 7735 30156 7744
rect 30104 7701 30113 7735
rect 30113 7701 30147 7735
rect 30147 7701 30156 7735
rect 30104 7692 30156 7701
rect 4193 7590 4245 7642
rect 4257 7590 4309 7642
rect 4321 7590 4373 7642
rect 4385 7590 4437 7642
rect 4449 7590 4501 7642
rect 11783 7590 11835 7642
rect 11847 7590 11899 7642
rect 11911 7590 11963 7642
rect 11975 7590 12027 7642
rect 12039 7590 12091 7642
rect 19373 7590 19425 7642
rect 19437 7590 19489 7642
rect 19501 7590 19553 7642
rect 19565 7590 19617 7642
rect 19629 7590 19681 7642
rect 26963 7590 27015 7642
rect 27027 7590 27079 7642
rect 27091 7590 27143 7642
rect 27155 7590 27207 7642
rect 27219 7590 27271 7642
rect 4712 7488 4764 7540
rect 848 7284 900 7336
rect 2412 7284 2464 7336
rect 4068 7352 4120 7404
rect 6460 7488 6512 7540
rect 6920 7488 6972 7540
rect 5356 7463 5408 7472
rect 5356 7429 5365 7463
rect 5365 7429 5399 7463
rect 5399 7429 5408 7463
rect 5356 7420 5408 7429
rect 7196 7420 7248 7472
rect 7472 7420 7524 7472
rect 5908 7352 5960 7404
rect 6276 7352 6328 7404
rect 2872 7284 2924 7336
rect 5724 7327 5776 7336
rect 5724 7293 5733 7327
rect 5733 7293 5767 7327
rect 5767 7293 5776 7327
rect 5724 7284 5776 7293
rect 8392 7352 8444 7404
rect 15108 7488 15160 7540
rect 6460 7327 6512 7336
rect 6460 7293 6469 7327
rect 6469 7293 6503 7327
rect 6503 7293 6512 7327
rect 6460 7284 6512 7293
rect 6828 7284 6880 7336
rect 8116 7327 8168 7336
rect 8116 7293 8125 7327
rect 8125 7293 8159 7327
rect 8159 7293 8168 7327
rect 8116 7284 8168 7293
rect 8760 7284 8812 7336
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 10416 7284 10468 7336
rect 10968 7284 11020 7336
rect 11244 7327 11296 7336
rect 11244 7293 11253 7327
rect 11253 7293 11287 7327
rect 11287 7293 11296 7327
rect 11244 7284 11296 7293
rect 11336 7284 11388 7336
rect 12348 7352 12400 7404
rect 12256 7284 12308 7336
rect 13820 7352 13872 7404
rect 14004 7352 14056 7404
rect 1400 7191 1452 7200
rect 1400 7157 1415 7191
rect 1415 7157 1449 7191
rect 1449 7157 1452 7191
rect 1400 7148 1452 7157
rect 2136 7148 2188 7200
rect 3240 7191 3292 7200
rect 3240 7157 3249 7191
rect 3249 7157 3283 7191
rect 3283 7157 3292 7191
rect 3240 7148 3292 7157
rect 6000 7148 6052 7200
rect 6368 7148 6420 7200
rect 7564 7191 7616 7200
rect 7564 7157 7573 7191
rect 7573 7157 7607 7191
rect 7607 7157 7616 7191
rect 7564 7148 7616 7157
rect 8392 7148 8444 7200
rect 12716 7216 12768 7268
rect 14280 7327 14332 7336
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 15200 7352 15252 7404
rect 16580 7352 16632 7404
rect 16764 7327 16816 7336
rect 16764 7293 16773 7327
rect 16773 7293 16807 7327
rect 16807 7293 16816 7327
rect 16764 7284 16816 7293
rect 17776 7488 17828 7540
rect 18604 7488 18656 7540
rect 19800 7488 19852 7540
rect 21364 7488 21416 7540
rect 21824 7488 21876 7540
rect 23756 7488 23808 7540
rect 25136 7488 25188 7540
rect 25872 7463 25924 7472
rect 25872 7429 25881 7463
rect 25881 7429 25915 7463
rect 25915 7429 25924 7463
rect 25872 7420 25924 7429
rect 28448 7531 28500 7540
rect 28448 7497 28457 7531
rect 28457 7497 28491 7531
rect 28491 7497 28500 7531
rect 28448 7488 28500 7497
rect 28724 7420 28776 7472
rect 17500 7352 17552 7404
rect 17868 7284 17920 7336
rect 18144 7284 18196 7336
rect 11336 7148 11388 7200
rect 11704 7191 11756 7200
rect 11704 7157 11719 7191
rect 11719 7157 11753 7191
rect 11753 7157 11756 7191
rect 18236 7216 18288 7268
rect 11704 7148 11756 7157
rect 14096 7148 14148 7200
rect 14740 7148 14792 7200
rect 15200 7148 15252 7200
rect 16304 7148 16356 7200
rect 17040 7191 17092 7200
rect 17040 7157 17049 7191
rect 17049 7157 17083 7191
rect 17083 7157 17092 7191
rect 17040 7148 17092 7157
rect 17132 7148 17184 7200
rect 17408 7148 17460 7200
rect 18604 7284 18656 7336
rect 21732 7352 21784 7404
rect 22100 7352 22152 7404
rect 22192 7352 22244 7404
rect 24584 7352 24636 7404
rect 24676 7352 24728 7404
rect 20812 7284 20864 7336
rect 21456 7284 21508 7336
rect 20168 7216 20220 7268
rect 21180 7216 21232 7268
rect 23480 7284 23532 7336
rect 23664 7284 23716 7336
rect 23572 7216 23624 7268
rect 24768 7327 24820 7336
rect 24768 7293 24777 7327
rect 24777 7293 24811 7327
rect 24811 7293 24820 7327
rect 24768 7284 24820 7293
rect 26240 7327 26292 7336
rect 26240 7293 26249 7327
rect 26249 7293 26283 7327
rect 26283 7293 26292 7327
rect 26240 7284 26292 7293
rect 20720 7148 20772 7200
rect 21916 7148 21968 7200
rect 24492 7191 24544 7200
rect 24492 7157 24507 7191
rect 24507 7157 24541 7191
rect 24541 7157 24544 7191
rect 26792 7284 26844 7336
rect 26976 7327 27028 7336
rect 26976 7293 26985 7327
rect 26985 7293 27019 7327
rect 27019 7293 27028 7327
rect 26976 7284 27028 7293
rect 27436 7284 27488 7336
rect 29092 7284 29144 7336
rect 29184 7327 29236 7336
rect 29184 7293 29193 7327
rect 29193 7293 29227 7327
rect 29227 7293 29236 7327
rect 29184 7284 29236 7293
rect 29368 7284 29420 7336
rect 24492 7148 24544 7157
rect 29000 7191 29052 7200
rect 29000 7157 29009 7191
rect 29009 7157 29043 7191
rect 29043 7157 29052 7191
rect 29000 7148 29052 7157
rect 29736 7148 29788 7200
rect 7988 7046 8040 7098
rect 8052 7046 8104 7098
rect 8116 7046 8168 7098
rect 8180 7046 8232 7098
rect 8244 7046 8296 7098
rect 15578 7046 15630 7098
rect 15642 7046 15694 7098
rect 15706 7046 15758 7098
rect 15770 7046 15822 7098
rect 15834 7046 15886 7098
rect 23168 7046 23220 7098
rect 23232 7046 23284 7098
rect 23296 7046 23348 7098
rect 23360 7046 23412 7098
rect 23424 7046 23476 7098
rect 30758 7046 30810 7098
rect 30822 7046 30874 7098
rect 30886 7046 30938 7098
rect 30950 7046 31002 7098
rect 31014 7046 31066 7098
rect 848 6740 900 6792
rect 3240 6944 3292 6996
rect 4896 6944 4948 6996
rect 6276 6944 6328 6996
rect 9404 6944 9456 6996
rect 10324 6944 10376 6996
rect 4804 6876 4856 6928
rect 1400 6783 1452 6792
rect 1400 6749 1402 6783
rect 1402 6749 1452 6783
rect 1400 6740 1452 6749
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 1768 6604 1820 6656
rect 2504 6604 2556 6656
rect 2872 6647 2924 6656
rect 2872 6613 2881 6647
rect 2881 6613 2915 6647
rect 2915 6613 2924 6647
rect 2872 6604 2924 6613
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 3608 6783 3660 6792
rect 3608 6749 3610 6783
rect 3610 6749 3660 6783
rect 3608 6740 3660 6749
rect 5356 6808 5408 6860
rect 8392 6876 8444 6928
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4712 6672 4764 6724
rect 5724 6672 5776 6724
rect 6000 6740 6052 6792
rect 6368 6740 6420 6792
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 7564 6740 7616 6792
rect 8484 6808 8536 6860
rect 8760 6783 8812 6792
rect 8760 6749 8762 6783
rect 8762 6749 8812 6783
rect 8760 6740 8812 6749
rect 9128 6783 9180 6792
rect 9128 6749 9137 6783
rect 9137 6749 9171 6783
rect 9171 6749 9180 6783
rect 9128 6740 9180 6749
rect 9496 6740 9548 6792
rect 10232 6740 10284 6792
rect 11336 6944 11388 6996
rect 12072 6944 12124 6996
rect 13176 6987 13228 6996
rect 13176 6953 13185 6987
rect 13185 6953 13219 6987
rect 13219 6953 13228 6987
rect 13176 6944 13228 6953
rect 14096 6944 14148 6996
rect 14648 6944 14700 6996
rect 11704 6851 11756 6860
rect 11704 6817 11706 6851
rect 11706 6817 11756 6851
rect 11704 6808 11756 6817
rect 11152 6740 11204 6792
rect 11520 6740 11572 6792
rect 12072 6783 12124 6792
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 12072 6740 12124 6749
rect 13544 6851 13596 6860
rect 13544 6817 13553 6851
rect 13553 6817 13587 6851
rect 13587 6817 13596 6851
rect 13544 6808 13596 6817
rect 13728 6808 13780 6860
rect 16120 6987 16172 6996
rect 16120 6953 16129 6987
rect 16129 6953 16163 6987
rect 16163 6953 16172 6987
rect 16120 6944 16172 6953
rect 17500 6987 17552 6996
rect 17500 6953 17509 6987
rect 17509 6953 17543 6987
rect 17543 6953 17552 6987
rect 17500 6944 17552 6953
rect 17776 6944 17828 6996
rect 16488 6808 16540 6860
rect 16580 6808 16632 6860
rect 16764 6808 16816 6860
rect 17132 6808 17184 6860
rect 12808 6740 12860 6792
rect 13820 6783 13872 6792
rect 13820 6749 13829 6783
rect 13829 6749 13863 6783
rect 13863 6749 13872 6783
rect 13820 6740 13872 6749
rect 14464 6740 14516 6792
rect 17316 6808 17368 6860
rect 18144 6944 18196 6996
rect 20904 6944 20956 6996
rect 22008 6944 22060 6996
rect 23664 6944 23716 6996
rect 26240 6944 26292 6996
rect 26976 6944 27028 6996
rect 27896 6944 27948 6996
rect 17868 6740 17920 6792
rect 18236 6740 18288 6792
rect 19248 6808 19300 6860
rect 26700 6876 26752 6928
rect 27436 6876 27488 6928
rect 18604 6740 18656 6792
rect 18696 6740 18748 6792
rect 5080 6647 5132 6656
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 5448 6647 5500 6656
rect 5448 6613 5457 6647
rect 5457 6613 5491 6647
rect 5491 6613 5500 6647
rect 5448 6604 5500 6613
rect 5816 6604 5868 6656
rect 6276 6604 6328 6656
rect 7656 6647 7708 6656
rect 7656 6613 7665 6647
rect 7665 6613 7699 6647
rect 7699 6613 7708 6647
rect 7656 6604 7708 6613
rect 9220 6604 9272 6656
rect 9588 6604 9640 6656
rect 11244 6672 11296 6724
rect 15476 6672 15528 6724
rect 19708 6672 19760 6724
rect 21272 6808 21324 6860
rect 21548 6808 21600 6860
rect 24124 6808 24176 6860
rect 21180 6740 21232 6792
rect 21364 6740 21416 6792
rect 21916 6740 21968 6792
rect 23388 6740 23440 6792
rect 24032 6783 24084 6792
rect 24032 6749 24049 6783
rect 24049 6749 24083 6783
rect 24083 6749 24084 6783
rect 24032 6740 24084 6749
rect 24492 6783 24544 6792
rect 24492 6749 24504 6783
rect 24504 6749 24538 6783
rect 24538 6749 24544 6783
rect 24492 6740 24544 6749
rect 24676 6740 24728 6792
rect 25964 6740 26016 6792
rect 30288 6808 30340 6860
rect 27804 6783 27856 6792
rect 27804 6749 27813 6783
rect 27813 6749 27847 6783
rect 27847 6749 27856 6783
rect 27804 6740 27856 6749
rect 27988 6740 28040 6792
rect 28264 6783 28316 6792
rect 28264 6749 28276 6783
rect 28276 6749 28310 6783
rect 28310 6749 28316 6783
rect 28264 6740 28316 6749
rect 9864 6604 9916 6656
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 10600 6604 10652 6613
rect 11060 6647 11112 6656
rect 11060 6613 11069 6647
rect 11069 6613 11103 6647
rect 11103 6613 11112 6647
rect 11060 6604 11112 6613
rect 11336 6604 11388 6656
rect 13360 6604 13412 6656
rect 13728 6647 13780 6656
rect 13728 6613 13737 6647
rect 13737 6613 13771 6647
rect 13771 6613 13780 6647
rect 13728 6604 13780 6613
rect 14464 6604 14516 6656
rect 16580 6647 16632 6656
rect 16580 6613 16589 6647
rect 16589 6613 16623 6647
rect 16623 6613 16632 6647
rect 16580 6604 16632 6613
rect 16672 6604 16724 6656
rect 17132 6647 17184 6656
rect 17132 6613 17141 6647
rect 17141 6613 17175 6647
rect 17175 6613 17184 6647
rect 17132 6604 17184 6613
rect 17224 6647 17276 6656
rect 17224 6613 17233 6647
rect 17233 6613 17267 6647
rect 17267 6613 17276 6647
rect 17224 6604 17276 6613
rect 17776 6604 17828 6656
rect 18604 6604 18656 6656
rect 20260 6647 20312 6656
rect 20260 6613 20269 6647
rect 20269 6613 20303 6647
rect 20303 6613 20312 6647
rect 20260 6604 20312 6613
rect 20536 6647 20588 6656
rect 20536 6613 20545 6647
rect 20545 6613 20579 6647
rect 20579 6613 20588 6647
rect 20536 6604 20588 6613
rect 21180 6604 21232 6656
rect 21548 6604 21600 6656
rect 21732 6604 21784 6656
rect 25228 6604 25280 6656
rect 25872 6604 25924 6656
rect 26056 6647 26108 6656
rect 26056 6613 26065 6647
rect 26065 6613 26099 6647
rect 26099 6613 26108 6647
rect 26056 6604 26108 6613
rect 27344 6672 27396 6724
rect 4193 6502 4245 6554
rect 4257 6502 4309 6554
rect 4321 6502 4373 6554
rect 4385 6502 4437 6554
rect 4449 6502 4501 6554
rect 11783 6502 11835 6554
rect 11847 6502 11899 6554
rect 11911 6502 11963 6554
rect 11975 6502 12027 6554
rect 12039 6502 12091 6554
rect 19373 6502 19425 6554
rect 19437 6502 19489 6554
rect 19501 6502 19553 6554
rect 19565 6502 19617 6554
rect 19629 6502 19681 6554
rect 26963 6502 27015 6554
rect 27027 6502 27079 6554
rect 27091 6502 27143 6554
rect 27155 6502 27207 6554
rect 27219 6502 27271 6554
rect 5080 6400 5132 6452
rect 5356 6400 5408 6452
rect 11060 6400 11112 6452
rect 11152 6400 11204 6452
rect 14556 6400 14608 6452
rect 16212 6443 16264 6452
rect 16212 6409 16221 6443
rect 16221 6409 16255 6443
rect 16255 6409 16264 6443
rect 16212 6400 16264 6409
rect 2596 6264 2648 6316
rect 848 6196 900 6248
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 2044 6196 2096 6248
rect 7380 6375 7432 6384
rect 7380 6341 7389 6375
rect 7389 6341 7423 6375
rect 7423 6341 7432 6375
rect 7380 6332 7432 6341
rect 8392 6332 8444 6384
rect 5724 6264 5776 6316
rect 5908 6307 5960 6316
rect 5908 6273 5910 6307
rect 5910 6273 5960 6307
rect 5908 6264 5960 6273
rect 6092 6264 6144 6316
rect 6184 6264 6236 6316
rect 8576 6264 8628 6316
rect 9036 6264 9088 6316
rect 11612 6307 11664 6316
rect 3148 6196 3200 6248
rect 3884 6196 3936 6248
rect 8392 6239 8444 6248
rect 8392 6205 8401 6239
rect 8401 6205 8435 6239
rect 8435 6205 8444 6239
rect 8392 6196 8444 6205
rect 8484 6196 8536 6248
rect 1400 6103 1452 6112
rect 1400 6069 1415 6103
rect 1415 6069 1449 6103
rect 1449 6069 1452 6103
rect 1400 6060 1452 6069
rect 2780 6103 2832 6112
rect 2780 6069 2789 6103
rect 2789 6069 2823 6103
rect 2823 6069 2832 6103
rect 2780 6060 2832 6069
rect 3240 6060 3292 6112
rect 3700 6060 3752 6112
rect 5080 6103 5132 6112
rect 5080 6069 5089 6103
rect 5089 6069 5123 6103
rect 5123 6069 5132 6103
rect 5080 6060 5132 6069
rect 8668 6060 8720 6112
rect 9588 6060 9640 6112
rect 10876 6196 10928 6248
rect 11060 6239 11112 6248
rect 11060 6205 11069 6239
rect 11069 6205 11103 6239
rect 11103 6205 11112 6239
rect 11060 6196 11112 6205
rect 11244 6239 11296 6248
rect 11244 6205 11253 6239
rect 11253 6205 11287 6239
rect 11287 6205 11296 6239
rect 11244 6196 11296 6205
rect 11612 6273 11614 6307
rect 11614 6273 11664 6307
rect 11612 6264 11664 6273
rect 12440 6264 12492 6316
rect 13820 6264 13872 6316
rect 14740 6307 14792 6316
rect 14740 6273 14742 6307
rect 14742 6273 14792 6307
rect 14740 6264 14792 6273
rect 15016 6264 15068 6316
rect 16304 6264 16356 6316
rect 13360 6196 13412 6248
rect 14096 6196 14148 6248
rect 10048 6060 10100 6112
rect 13636 6128 13688 6180
rect 16672 6196 16724 6248
rect 18696 6400 18748 6452
rect 20260 6400 20312 6452
rect 21272 6400 21324 6452
rect 18236 6332 18288 6384
rect 24768 6400 24820 6452
rect 25228 6400 25280 6452
rect 29644 6400 29696 6452
rect 23572 6332 23624 6384
rect 21548 6264 21600 6316
rect 23480 6264 23532 6316
rect 17592 6196 17644 6248
rect 17960 6239 18012 6248
rect 17960 6205 17969 6239
rect 17969 6205 18003 6239
rect 18003 6205 18012 6239
rect 17960 6196 18012 6205
rect 18236 6239 18288 6248
rect 18236 6205 18245 6239
rect 18245 6205 18279 6239
rect 18279 6205 18288 6239
rect 18236 6196 18288 6205
rect 18328 6239 18380 6248
rect 18328 6205 18337 6239
rect 18337 6205 18371 6239
rect 18371 6205 18380 6239
rect 18328 6196 18380 6205
rect 18696 6239 18748 6248
rect 18696 6205 18705 6239
rect 18705 6205 18739 6239
rect 18739 6205 18748 6239
rect 18696 6196 18748 6205
rect 18788 6196 18840 6248
rect 18972 6196 19024 6248
rect 21272 6196 21324 6248
rect 26332 6264 26384 6316
rect 27528 6264 27580 6316
rect 28080 6264 28132 6316
rect 23756 6196 23808 6248
rect 23940 6196 23992 6248
rect 24676 6196 24728 6248
rect 24860 6196 24912 6248
rect 18604 6128 18656 6180
rect 24124 6128 24176 6180
rect 26148 6171 26200 6180
rect 26148 6137 26157 6171
rect 26157 6137 26191 6171
rect 26191 6137 26200 6171
rect 26148 6128 26200 6137
rect 26516 6128 26568 6180
rect 26700 6239 26752 6248
rect 26700 6205 26709 6239
rect 26709 6205 26743 6239
rect 26743 6205 26752 6239
rect 26700 6196 26752 6205
rect 26792 6196 26844 6248
rect 29276 6196 29328 6248
rect 13452 6060 13504 6112
rect 13544 6103 13596 6112
rect 13544 6069 13553 6103
rect 13553 6069 13587 6103
rect 13587 6069 13596 6103
rect 13544 6060 13596 6069
rect 14464 6060 14516 6112
rect 16856 6060 16908 6112
rect 16948 6103 17000 6112
rect 16948 6069 16957 6103
rect 16957 6069 16991 6103
rect 16991 6069 17000 6103
rect 16948 6060 17000 6069
rect 17040 6060 17092 6112
rect 17224 6103 17276 6112
rect 17224 6069 17233 6103
rect 17233 6069 17267 6103
rect 17267 6069 17276 6103
rect 17224 6060 17276 6069
rect 17684 6103 17736 6112
rect 17684 6069 17693 6103
rect 17693 6069 17727 6103
rect 17727 6069 17736 6103
rect 17684 6060 17736 6069
rect 18512 6103 18564 6112
rect 18512 6069 18521 6103
rect 18521 6069 18555 6103
rect 18555 6069 18564 6103
rect 18512 6060 18564 6069
rect 18788 6060 18840 6112
rect 21548 6060 21600 6112
rect 22928 6060 22980 6112
rect 24768 6060 24820 6112
rect 26700 6060 26752 6112
rect 28356 6128 28408 6180
rect 27252 6060 27304 6112
rect 27344 6060 27396 6112
rect 7988 5958 8040 6010
rect 8052 5958 8104 6010
rect 8116 5958 8168 6010
rect 8180 5958 8232 6010
rect 8244 5958 8296 6010
rect 15578 5958 15630 6010
rect 15642 5958 15694 6010
rect 15706 5958 15758 6010
rect 15770 5958 15822 6010
rect 15834 5958 15886 6010
rect 23168 5958 23220 6010
rect 23232 5958 23284 6010
rect 23296 5958 23348 6010
rect 23360 5958 23412 6010
rect 23424 5958 23476 6010
rect 30758 5958 30810 6010
rect 30822 5958 30874 6010
rect 30886 5958 30938 6010
rect 30950 5958 31002 6010
rect 31014 5958 31066 6010
rect 1216 5856 1268 5908
rect 1584 5856 1636 5908
rect 2044 5856 2096 5908
rect 1032 5720 1084 5772
rect 1216 5763 1268 5772
rect 1216 5729 1225 5763
rect 1225 5729 1259 5763
rect 1259 5729 1268 5763
rect 1216 5720 1268 5729
rect 1308 5763 1360 5772
rect 1308 5729 1317 5763
rect 1317 5729 1351 5763
rect 1351 5729 1360 5763
rect 1308 5720 1360 5729
rect 2872 5856 2924 5908
rect 3792 5856 3844 5908
rect 5540 5856 5592 5908
rect 6460 5856 6512 5908
rect 8668 5856 8720 5908
rect 3516 5788 3568 5840
rect 5356 5788 5408 5840
rect 13452 5856 13504 5908
rect 16764 5856 16816 5908
rect 17040 5856 17092 5908
rect 20904 5856 20956 5908
rect 21548 5856 21600 5908
rect 23940 5899 23992 5908
rect 23940 5865 23955 5899
rect 23955 5865 23989 5899
rect 23989 5865 23992 5899
rect 23940 5856 23992 5865
rect 24860 5856 24912 5908
rect 25964 5899 26016 5908
rect 25964 5865 25973 5899
rect 25973 5865 26007 5899
rect 26007 5865 26016 5899
rect 25964 5856 26016 5865
rect 2872 5720 2924 5772
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 3332 5652 3384 5704
rect 4068 5652 4120 5704
rect 5448 5720 5500 5772
rect 7840 5720 7892 5772
rect 10416 5763 10468 5772
rect 10416 5729 10433 5763
rect 10433 5729 10467 5763
rect 10467 5729 10468 5763
rect 10416 5720 10468 5729
rect 5448 5584 5500 5636
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 5816 5695 5868 5704
rect 5816 5661 5825 5695
rect 5825 5661 5859 5695
rect 5859 5661 5868 5695
rect 5816 5652 5868 5661
rect 6184 5695 6236 5704
rect 6184 5661 6186 5695
rect 6186 5661 6236 5695
rect 6184 5652 6236 5661
rect 6276 5695 6328 5704
rect 6276 5661 6288 5695
rect 6288 5661 6322 5695
rect 6322 5661 6328 5695
rect 6276 5652 6328 5661
rect 6460 5652 6512 5704
rect 8300 5652 8352 5704
rect 8760 5695 8812 5704
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 10324 5652 10376 5704
rect 11244 5763 11296 5772
rect 11244 5729 11253 5763
rect 11253 5729 11287 5763
rect 11287 5729 11296 5763
rect 11244 5720 11296 5729
rect 14464 5720 14516 5772
rect 7656 5559 7708 5568
rect 7656 5525 7665 5559
rect 7665 5525 7699 5559
rect 7699 5525 7708 5559
rect 7656 5516 7708 5525
rect 8760 5516 8812 5568
rect 8944 5516 8996 5568
rect 11244 5584 11296 5636
rect 11612 5695 11664 5704
rect 11612 5661 11621 5695
rect 11621 5661 11655 5695
rect 11655 5661 11664 5695
rect 11612 5652 11664 5661
rect 11796 5652 11848 5704
rect 12164 5652 12216 5704
rect 14004 5652 14056 5704
rect 14188 5695 14240 5704
rect 14188 5661 14190 5695
rect 14190 5661 14240 5695
rect 14188 5652 14240 5661
rect 14280 5695 14332 5704
rect 14280 5661 14292 5695
rect 14292 5661 14326 5695
rect 14326 5661 14332 5695
rect 14280 5652 14332 5661
rect 16212 5695 16264 5704
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16212 5652 16264 5661
rect 16580 5695 16632 5704
rect 16580 5661 16582 5695
rect 16582 5661 16632 5695
rect 16580 5652 16632 5661
rect 16856 5720 16908 5772
rect 18788 5695 18840 5704
rect 18788 5661 18790 5695
rect 18790 5661 18840 5695
rect 10232 5559 10284 5568
rect 10232 5525 10241 5559
rect 10241 5525 10275 5559
rect 10275 5525 10284 5559
rect 10232 5516 10284 5525
rect 10784 5516 10836 5568
rect 11152 5516 11204 5568
rect 13728 5584 13780 5636
rect 14280 5516 14332 5568
rect 15384 5516 15436 5568
rect 17132 5516 17184 5568
rect 18788 5652 18840 5661
rect 27252 5856 27304 5908
rect 21272 5695 21324 5704
rect 21272 5661 21281 5695
rect 21281 5661 21315 5695
rect 21315 5661 21324 5695
rect 21272 5652 21324 5661
rect 21732 5695 21784 5704
rect 21732 5661 21744 5695
rect 21744 5661 21778 5695
rect 21778 5661 21784 5695
rect 21732 5652 21784 5661
rect 23664 5652 23716 5704
rect 24676 5720 24728 5772
rect 24952 5720 25004 5772
rect 25688 5720 25740 5772
rect 26516 5788 26568 5840
rect 29460 5856 29512 5908
rect 24216 5695 24268 5704
rect 24216 5661 24225 5695
rect 24225 5661 24259 5695
rect 24259 5661 24268 5695
rect 24216 5652 24268 5661
rect 26240 5720 26292 5772
rect 27988 5720 28040 5772
rect 25964 5652 26016 5704
rect 26884 5695 26936 5704
rect 26884 5661 26896 5695
rect 26896 5661 26930 5695
rect 26930 5661 26936 5695
rect 26884 5652 26936 5661
rect 27896 5584 27948 5636
rect 18696 5516 18748 5568
rect 21732 5516 21784 5568
rect 23388 5516 23440 5568
rect 24216 5516 24268 5568
rect 27804 5516 27856 5568
rect 29184 5559 29236 5568
rect 29184 5525 29193 5559
rect 29193 5525 29227 5559
rect 29227 5525 29236 5559
rect 29184 5516 29236 5525
rect 29460 5559 29512 5568
rect 29460 5525 29469 5559
rect 29469 5525 29503 5559
rect 29503 5525 29512 5559
rect 29460 5516 29512 5525
rect 4193 5414 4245 5466
rect 4257 5414 4309 5466
rect 4321 5414 4373 5466
rect 4385 5414 4437 5466
rect 4449 5414 4501 5466
rect 11783 5414 11835 5466
rect 11847 5414 11899 5466
rect 11911 5414 11963 5466
rect 11975 5414 12027 5466
rect 12039 5414 12091 5466
rect 19373 5414 19425 5466
rect 19437 5414 19489 5466
rect 19501 5414 19553 5466
rect 19565 5414 19617 5466
rect 19629 5414 19681 5466
rect 26963 5414 27015 5466
rect 27027 5414 27079 5466
rect 27091 5414 27143 5466
rect 27155 5414 27207 5466
rect 27219 5414 27271 5466
rect 1308 5312 1360 5364
rect 940 5219 992 5228
rect 940 5185 949 5219
rect 949 5185 983 5219
rect 983 5185 992 5219
rect 940 5176 992 5185
rect 2136 5176 2188 5228
rect 4068 5312 4120 5364
rect 6276 5312 6328 5364
rect 6368 5312 6420 5364
rect 6644 5312 6696 5364
rect 9312 5312 9364 5364
rect 9404 5312 9456 5364
rect 3700 5244 3752 5296
rect 7564 5244 7616 5296
rect 14372 5312 14424 5364
rect 20628 5312 20680 5364
rect 23112 5312 23164 5364
rect 24768 5312 24820 5364
rect 25412 5312 25464 5364
rect 26884 5312 26936 5364
rect 27068 5312 27120 5364
rect 28080 5312 28132 5364
rect 28540 5355 28592 5364
rect 28540 5321 28549 5355
rect 28549 5321 28583 5355
rect 28583 5321 28592 5355
rect 28540 5312 28592 5321
rect 13912 5244 13964 5296
rect 3148 5176 3200 5228
rect 3332 5176 3384 5228
rect 5080 5176 5132 5228
rect 5632 5176 5684 5228
rect 1584 5108 1636 5160
rect 1952 5108 2004 5160
rect 3792 5108 3844 5160
rect 4620 5151 4672 5160
rect 4620 5117 4629 5151
rect 4629 5117 4663 5151
rect 4663 5117 4672 5151
rect 4620 5108 4672 5117
rect 7656 5176 7708 5228
rect 3148 5040 3200 5092
rect 6920 5108 6972 5160
rect 9404 5176 9456 5228
rect 9680 5176 9732 5228
rect 9772 5219 9824 5226
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5174 9824 5185
rect 11152 5176 11204 5228
rect 7932 5108 7984 5160
rect 8760 5040 8812 5092
rect 6460 4972 6512 5024
rect 6828 4972 6880 5024
rect 7104 4972 7156 5024
rect 8392 4972 8444 5024
rect 8944 5108 8996 5160
rect 11520 5108 11572 5160
rect 11704 5219 11756 5228
rect 11704 5185 11716 5219
rect 11716 5185 11750 5219
rect 11750 5185 11756 5219
rect 11704 5176 11756 5185
rect 11888 5176 11940 5228
rect 14188 5176 14240 5228
rect 12256 5108 12308 5160
rect 14004 5151 14056 5160
rect 14004 5117 14013 5151
rect 14013 5117 14047 5151
rect 14047 5117 14056 5151
rect 14004 5108 14056 5117
rect 14556 5176 14608 5228
rect 16948 5219 17000 5228
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 20536 5176 20588 5228
rect 22008 5176 22060 5228
rect 16212 5151 16264 5160
rect 16212 5117 16221 5151
rect 16221 5117 16255 5151
rect 16255 5117 16264 5151
rect 16212 5108 16264 5117
rect 16580 5151 16632 5160
rect 16580 5117 16582 5151
rect 16582 5117 16632 5151
rect 16580 5108 16632 5117
rect 18696 5151 18748 5160
rect 18696 5117 18705 5151
rect 18705 5117 18739 5151
rect 18739 5117 18748 5151
rect 18696 5108 18748 5117
rect 9036 4972 9088 5024
rect 9680 4972 9732 5024
rect 10048 4972 10100 5024
rect 11520 4972 11572 5024
rect 11888 4972 11940 5024
rect 11980 4972 12032 5024
rect 13820 5040 13872 5092
rect 14096 5040 14148 5092
rect 13728 5015 13780 5024
rect 13728 4981 13737 5015
rect 13737 4981 13771 5015
rect 13771 4981 13780 5015
rect 13728 4972 13780 4981
rect 13912 4972 13964 5024
rect 21180 5108 21232 5160
rect 23388 5108 23440 5160
rect 23572 5151 23624 5160
rect 23572 5117 23581 5151
rect 23581 5117 23615 5151
rect 23615 5117 23624 5151
rect 23572 5108 23624 5117
rect 23664 5108 23716 5160
rect 24124 5176 24176 5228
rect 26424 5176 26476 5228
rect 29000 5176 29052 5228
rect 18788 4972 18840 5024
rect 20720 4972 20772 5024
rect 20904 4972 20956 5024
rect 21272 4972 21324 5024
rect 21548 4972 21600 5024
rect 22744 5015 22796 5024
rect 22744 4981 22753 5015
rect 22753 4981 22787 5015
rect 22787 4981 22796 5015
rect 22744 4972 22796 4981
rect 25964 5108 26016 5160
rect 23940 5040 23992 5092
rect 27528 5108 27580 5160
rect 23848 4972 23900 5024
rect 24124 4972 24176 5024
rect 26608 4972 26660 5024
rect 27068 4972 27120 5024
rect 28356 4972 28408 5024
rect 7988 4870 8040 4922
rect 8052 4870 8104 4922
rect 8116 4870 8168 4922
rect 8180 4870 8232 4922
rect 8244 4870 8296 4922
rect 15578 4870 15630 4922
rect 15642 4870 15694 4922
rect 15706 4870 15758 4922
rect 15770 4870 15822 4922
rect 15834 4870 15886 4922
rect 23168 4870 23220 4922
rect 23232 4870 23284 4922
rect 23296 4870 23348 4922
rect 23360 4870 23412 4922
rect 23424 4870 23476 4922
rect 30758 4870 30810 4922
rect 30822 4870 30874 4922
rect 30886 4870 30938 4922
rect 30950 4870 31002 4922
rect 31014 4870 31066 4922
rect 1492 4768 1544 4820
rect 3516 4768 3568 4820
rect 3792 4768 3844 4820
rect 7840 4811 7892 4820
rect 7840 4777 7849 4811
rect 7849 4777 7883 4811
rect 7883 4777 7892 4811
rect 7840 4768 7892 4777
rect 848 4675 900 4684
rect 848 4641 857 4675
rect 857 4641 891 4675
rect 891 4641 900 4675
rect 848 4632 900 4641
rect 1860 4632 1912 4684
rect 3332 4632 3384 4684
rect 3424 4675 3476 4684
rect 3424 4641 3433 4675
rect 3433 4641 3467 4675
rect 3467 4641 3476 4675
rect 3424 4632 3476 4641
rect 9496 4768 9548 4820
rect 9772 4768 9824 4820
rect 11152 4768 11204 4820
rect 11520 4768 11572 4820
rect 12256 4768 12308 4820
rect 14096 4768 14148 4820
rect 14188 4768 14240 4820
rect 16580 4768 16632 4820
rect 19340 4768 19392 4820
rect 19984 4768 20036 4820
rect 20168 4768 20220 4820
rect 1492 4564 1544 4616
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 1492 4428 1544 4480
rect 3240 4564 3292 4616
rect 4988 4632 5040 4684
rect 4068 4564 4120 4616
rect 5632 4496 5684 4548
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 3424 4428 3476 4480
rect 5816 4564 5868 4616
rect 6184 4564 6236 4616
rect 7196 4632 7248 4684
rect 9496 4632 9548 4684
rect 11244 4700 11296 4752
rect 11336 4632 11388 4684
rect 8300 4564 8352 4616
rect 8852 4564 8904 4616
rect 9036 4607 9088 4616
rect 9036 4573 9038 4607
rect 9038 4573 9088 4607
rect 9036 4564 9088 4573
rect 9220 4564 9272 4616
rect 11612 4675 11664 4684
rect 11612 4641 11621 4675
rect 11621 4641 11655 4675
rect 11655 4641 11664 4675
rect 11612 4632 11664 4641
rect 13728 4700 13780 4752
rect 18972 4700 19024 4752
rect 24492 4768 24544 4820
rect 26240 4768 26292 4820
rect 29184 4768 29236 4820
rect 13544 4632 13596 4684
rect 8484 4496 8536 4548
rect 11888 4564 11940 4616
rect 14004 4564 14056 4616
rect 14280 4607 14332 4616
rect 14280 4573 14292 4607
rect 14292 4573 14326 4607
rect 14326 4573 14332 4607
rect 14280 4564 14332 4573
rect 16212 4607 16264 4616
rect 16212 4573 16221 4607
rect 16221 4573 16255 4607
rect 16255 4573 16264 4607
rect 16212 4564 16264 4573
rect 17224 4632 17276 4684
rect 18052 4632 18104 4684
rect 18420 4675 18472 4684
rect 18420 4641 18429 4675
rect 18429 4641 18463 4675
rect 18463 4641 18472 4675
rect 18420 4632 18472 4641
rect 19064 4632 19116 4684
rect 18788 4564 18840 4616
rect 20444 4632 20496 4684
rect 20536 4632 20588 4684
rect 21916 4632 21968 4684
rect 27528 4700 27580 4752
rect 18880 4496 18932 4548
rect 20168 4564 20220 4616
rect 22560 4607 22612 4616
rect 22560 4573 22562 4607
rect 22562 4573 22612 4607
rect 22560 4564 22612 4573
rect 22744 4564 22796 4616
rect 22928 4675 22980 4684
rect 22928 4641 22937 4675
rect 22937 4641 22971 4675
rect 22971 4641 22980 4675
rect 22928 4632 22980 4641
rect 23572 4632 23624 4684
rect 27896 4632 27948 4684
rect 27988 4675 28040 4684
rect 27988 4641 27997 4675
rect 27997 4641 28031 4675
rect 28031 4641 28040 4675
rect 27988 4632 28040 4641
rect 30104 4632 30156 4684
rect 25228 4564 25280 4616
rect 28356 4607 28408 4616
rect 28356 4573 28358 4607
rect 28358 4573 28408 4607
rect 28356 4564 28408 4573
rect 28540 4564 28592 4616
rect 9864 4428 9916 4480
rect 12164 4428 12216 4480
rect 13820 4428 13872 4480
rect 17408 4428 17460 4480
rect 22192 4496 22244 4548
rect 25780 4496 25832 4548
rect 20996 4471 21048 4480
rect 20996 4437 21005 4471
rect 21005 4437 21039 4471
rect 21039 4437 21048 4471
rect 20996 4428 21048 4437
rect 21272 4471 21324 4480
rect 21272 4437 21281 4471
rect 21281 4437 21315 4471
rect 21315 4437 21324 4471
rect 21272 4428 21324 4437
rect 21548 4471 21600 4480
rect 21548 4437 21557 4471
rect 21557 4437 21591 4471
rect 21591 4437 21600 4471
rect 21548 4428 21600 4437
rect 21824 4471 21876 4480
rect 21824 4437 21833 4471
rect 21833 4437 21867 4471
rect 21867 4437 21876 4471
rect 21824 4428 21876 4437
rect 22008 4428 22060 4480
rect 23664 4428 23716 4480
rect 24768 4428 24820 4480
rect 25044 4471 25096 4480
rect 25044 4437 25053 4471
rect 25053 4437 25087 4471
rect 25087 4437 25096 4471
rect 25044 4428 25096 4437
rect 25964 4428 26016 4480
rect 26792 4428 26844 4480
rect 26884 4471 26936 4480
rect 26884 4437 26893 4471
rect 26893 4437 26927 4471
rect 26927 4437 26936 4471
rect 26884 4428 26936 4437
rect 4193 4326 4245 4378
rect 4257 4326 4309 4378
rect 4321 4326 4373 4378
rect 4385 4326 4437 4378
rect 4449 4326 4501 4378
rect 11783 4326 11835 4378
rect 11847 4326 11899 4378
rect 11911 4326 11963 4378
rect 11975 4326 12027 4378
rect 12039 4326 12091 4378
rect 19373 4326 19425 4378
rect 19437 4326 19489 4378
rect 19501 4326 19553 4378
rect 19565 4326 19617 4378
rect 19629 4326 19681 4378
rect 26963 4326 27015 4378
rect 27027 4326 27079 4378
rect 27091 4326 27143 4378
rect 27155 4326 27207 4378
rect 27219 4326 27271 4378
rect 1400 4224 1452 4276
rect 1860 4224 1912 4276
rect 940 4131 992 4140
rect 940 4097 949 4131
rect 949 4097 983 4131
rect 983 4097 992 4131
rect 940 4088 992 4097
rect 3240 4224 3292 4276
rect 6552 4224 6604 4276
rect 8300 4224 8352 4276
rect 9772 4224 9824 4276
rect 8392 4156 8444 4208
rect 1768 4020 1820 4072
rect 3608 4088 3660 4140
rect 4344 4088 4396 4140
rect 4528 4131 4580 4140
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 4528 4088 4580 4097
rect 5540 4088 5592 4140
rect 8576 4088 8628 4140
rect 8668 4131 8720 4140
rect 8668 4097 8677 4131
rect 8677 4097 8711 4131
rect 8711 4097 8720 4131
rect 8668 4088 8720 4097
rect 2780 4020 2832 4072
rect 3792 4063 3844 4072
rect 3792 4029 3801 4063
rect 3801 4029 3835 4063
rect 3835 4029 3844 4063
rect 3792 4020 3844 4029
rect 5816 4020 5868 4072
rect 6736 4063 6788 4072
rect 6736 4029 6745 4063
rect 6745 4029 6779 4063
rect 6779 4029 6788 4063
rect 6736 4020 6788 4029
rect 7472 4020 7524 4072
rect 5908 3995 5960 4004
rect 5908 3961 5917 3995
rect 5917 3961 5951 3995
rect 5951 3961 5960 3995
rect 5908 3952 5960 3961
rect 1676 3884 1728 3936
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 2780 3884 2832 3893
rect 3332 3884 3384 3936
rect 4528 3884 4580 3936
rect 6276 3884 6328 3936
rect 8944 4020 8996 4072
rect 9128 4063 9180 4072
rect 9128 4029 9137 4063
rect 9137 4029 9171 4063
rect 9171 4029 9180 4063
rect 9128 4020 9180 4029
rect 9864 4199 9916 4208
rect 9864 4165 9873 4199
rect 9873 4165 9907 4199
rect 9907 4165 9916 4199
rect 9864 4156 9916 4165
rect 10048 4156 10100 4208
rect 11704 4224 11756 4276
rect 17684 4224 17736 4276
rect 17776 4224 17828 4276
rect 20536 4224 20588 4276
rect 10324 4088 10376 4140
rect 10784 4088 10836 4140
rect 11244 4088 11296 4140
rect 11612 4088 11664 4140
rect 12072 4088 12124 4140
rect 12256 4088 12308 4140
rect 14464 4131 14516 4140
rect 14464 4097 14476 4131
rect 14476 4097 14510 4131
rect 14510 4097 14516 4131
rect 14464 4088 14516 4097
rect 21272 4224 21324 4276
rect 21456 4088 21508 4140
rect 21548 4088 21600 4140
rect 22008 4088 22060 4140
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 9404 3884 9456 3936
rect 10140 3952 10192 4004
rect 10416 4020 10468 4072
rect 11888 4020 11940 4072
rect 12716 4020 12768 4072
rect 13912 4063 13964 4072
rect 13912 4029 13921 4063
rect 13921 4029 13955 4063
rect 13955 4029 13964 4063
rect 13912 4020 13964 4029
rect 14004 4063 14056 4072
rect 14004 4029 14013 4063
rect 14013 4029 14047 4063
rect 14047 4029 14056 4063
rect 14004 4020 14056 4029
rect 14740 4063 14792 4072
rect 14740 4029 14749 4063
rect 14749 4029 14783 4063
rect 14783 4029 14792 4063
rect 14740 4020 14792 4029
rect 16212 4063 16264 4072
rect 16212 4029 16221 4063
rect 16221 4029 16255 4063
rect 16255 4029 16264 4063
rect 16212 4020 16264 4029
rect 12440 3952 12492 4004
rect 15476 3952 15528 4004
rect 18696 4063 18748 4072
rect 18696 4029 18705 4063
rect 18705 4029 18739 4063
rect 18739 4029 18748 4063
rect 18696 4020 18748 4029
rect 18972 4020 19024 4072
rect 20904 4063 20956 4072
rect 20904 4029 20913 4063
rect 20913 4029 20947 4063
rect 20947 4029 20956 4063
rect 20904 4020 20956 4029
rect 23572 4020 23624 4072
rect 23756 4020 23808 4072
rect 24216 4020 24268 4072
rect 26148 4088 26200 4140
rect 26516 4088 26568 4140
rect 26608 4088 26660 4140
rect 24584 4063 24636 4072
rect 24584 4029 24593 4063
rect 24593 4029 24627 4063
rect 24627 4029 24636 4063
rect 24584 4020 24636 4029
rect 24860 4063 24912 4072
rect 24860 4029 24869 4063
rect 24869 4029 24903 4063
rect 24903 4029 24912 4063
rect 24860 4020 24912 4029
rect 25964 4063 26016 4072
rect 25964 4029 25973 4063
rect 25973 4029 26007 4063
rect 26007 4029 26016 4063
rect 25964 4020 26016 4029
rect 27436 4020 27488 4072
rect 28172 4063 28224 4072
rect 28172 4029 28181 4063
rect 28181 4029 28215 4063
rect 28215 4029 28224 4063
rect 28172 4020 28224 4029
rect 29552 4088 29604 4140
rect 22560 3952 22612 4004
rect 10600 3927 10652 3936
rect 10600 3893 10615 3927
rect 10615 3893 10649 3927
rect 10649 3893 10652 3927
rect 10600 3884 10652 3893
rect 12072 3884 12124 3936
rect 13728 3927 13780 3936
rect 13728 3893 13737 3927
rect 13737 3893 13771 3927
rect 13771 3893 13780 3927
rect 13728 3884 13780 3893
rect 14280 3884 14332 3936
rect 16580 3884 16632 3936
rect 18788 3884 18840 3936
rect 22744 3927 22796 3936
rect 22744 3893 22753 3927
rect 22753 3893 22787 3927
rect 22787 3893 22796 3927
rect 22744 3884 22796 3893
rect 22928 3884 22980 3936
rect 24032 3884 24084 3936
rect 24124 3927 24176 3936
rect 24124 3893 24133 3927
rect 24133 3893 24167 3927
rect 24167 3893 24176 3927
rect 24124 3884 24176 3893
rect 24400 3927 24452 3936
rect 24400 3893 24409 3927
rect 24409 3893 24443 3927
rect 24443 3893 24452 3927
rect 24400 3884 24452 3893
rect 24676 3927 24728 3936
rect 24676 3893 24685 3927
rect 24685 3893 24719 3927
rect 24719 3893 24728 3927
rect 24676 3884 24728 3893
rect 25504 3927 25556 3936
rect 25504 3893 25513 3927
rect 25513 3893 25547 3927
rect 25547 3893 25556 3927
rect 25504 3884 25556 3893
rect 26424 3927 26476 3936
rect 26424 3893 26439 3927
rect 26439 3893 26473 3927
rect 26473 3893 26476 3927
rect 26424 3884 26476 3893
rect 26608 3884 26660 3936
rect 27528 3884 27580 3936
rect 28356 3927 28408 3936
rect 28356 3893 28365 3927
rect 28365 3893 28399 3927
rect 28399 3893 28408 3927
rect 28356 3884 28408 3893
rect 7988 3782 8040 3834
rect 8052 3782 8104 3834
rect 8116 3782 8168 3834
rect 8180 3782 8232 3834
rect 8244 3782 8296 3834
rect 15578 3782 15630 3834
rect 15642 3782 15694 3834
rect 15706 3782 15758 3834
rect 15770 3782 15822 3834
rect 15834 3782 15886 3834
rect 23168 3782 23220 3834
rect 23232 3782 23284 3834
rect 23296 3782 23348 3834
rect 23360 3782 23412 3834
rect 23424 3782 23476 3834
rect 30758 3782 30810 3834
rect 30822 3782 30874 3834
rect 30886 3782 30938 3834
rect 30950 3782 31002 3834
rect 31014 3782 31066 3834
rect 6736 3680 6788 3732
rect 6828 3680 6880 3732
rect 8668 3680 8720 3732
rect 9036 3680 9088 3732
rect 10600 3680 10652 3732
rect 2780 3612 2832 3664
rect 3608 3612 3660 3664
rect 1032 3476 1084 3528
rect 1676 3519 1728 3528
rect 1676 3485 1678 3519
rect 1678 3485 1728 3519
rect 1676 3476 1728 3485
rect 4068 3544 4120 3596
rect 5356 3544 5408 3596
rect 6460 3587 6512 3596
rect 6460 3553 6469 3587
rect 6469 3553 6503 3587
rect 6503 3553 6512 3587
rect 6460 3544 6512 3553
rect 10140 3612 10192 3664
rect 2044 3519 2096 3528
rect 2044 3485 2053 3519
rect 2053 3485 2087 3519
rect 2087 3485 2096 3519
rect 2044 3476 2096 3485
rect 3240 3476 3292 3528
rect 3700 3476 3752 3528
rect 4160 3476 4212 3528
rect 6276 3476 6328 3528
rect 7012 3476 7064 3528
rect 7564 3544 7616 3596
rect 8300 3476 8352 3528
rect 8852 3476 8904 3528
rect 9036 3519 9088 3528
rect 9036 3485 9038 3519
rect 9038 3485 9088 3519
rect 9036 3476 9088 3485
rect 9404 3587 9456 3596
rect 9404 3553 9413 3587
rect 9413 3553 9447 3587
rect 9447 3553 9456 3587
rect 9404 3544 9456 3553
rect 9680 3544 9732 3596
rect 10232 3544 10284 3596
rect 9312 3476 9364 3528
rect 9588 3476 9640 3528
rect 11888 3476 11940 3528
rect 5816 3408 5868 3460
rect 12072 3587 12124 3596
rect 12072 3553 12081 3587
rect 12081 3553 12115 3587
rect 12115 3553 12124 3587
rect 12072 3544 12124 3553
rect 14464 3680 14516 3732
rect 16212 3680 16264 3732
rect 16580 3612 16632 3664
rect 18972 3612 19024 3664
rect 13268 3544 13320 3596
rect 12256 3476 12308 3528
rect 12532 3519 12584 3528
rect 12532 3485 12544 3519
rect 12544 3485 12578 3519
rect 12578 3485 12584 3519
rect 12532 3476 12584 3485
rect 15292 3476 15344 3528
rect 16764 3519 16816 3528
rect 16764 3485 16773 3519
rect 16773 3485 16807 3519
rect 16807 3485 16816 3519
rect 16764 3476 16816 3485
rect 17132 3519 17184 3528
rect 17132 3485 17134 3519
rect 17134 3485 17184 3519
rect 17132 3476 17184 3485
rect 17224 3476 17276 3528
rect 20904 3612 20956 3664
rect 21640 3612 21692 3664
rect 25228 3612 25280 3664
rect 19340 3587 19392 3596
rect 19340 3553 19342 3587
rect 19342 3553 19392 3587
rect 19340 3544 19392 3553
rect 18420 3476 18472 3528
rect 18604 3476 18656 3528
rect 18880 3476 18932 3528
rect 20628 3476 20680 3528
rect 1584 3340 1636 3392
rect 1676 3340 1728 3392
rect 3700 3340 3752 3392
rect 4344 3340 4396 3392
rect 4620 3340 4672 3392
rect 6368 3340 6420 3392
rect 8944 3340 8996 3392
rect 11612 3340 11664 3392
rect 11704 3340 11756 3392
rect 12072 3408 12124 3460
rect 14096 3408 14148 3460
rect 22560 3587 22612 3596
rect 22560 3553 22562 3587
rect 22562 3553 22612 3587
rect 22560 3544 22612 3553
rect 22928 3587 22980 3596
rect 22928 3553 22937 3587
rect 22937 3553 22971 3587
rect 22971 3553 22980 3587
rect 22928 3544 22980 3553
rect 24768 3544 24820 3596
rect 25596 3544 25648 3596
rect 25872 3544 25924 3596
rect 28172 3680 28224 3732
rect 29000 3680 29052 3732
rect 27436 3544 27488 3596
rect 21916 3476 21968 3528
rect 22192 3519 22244 3528
rect 22192 3485 22201 3519
rect 22201 3485 22235 3519
rect 22235 3485 22244 3519
rect 22192 3476 22244 3485
rect 22744 3476 22796 3528
rect 12532 3340 12584 3392
rect 13636 3340 13688 3392
rect 14648 3340 14700 3392
rect 18972 3340 19024 3392
rect 21548 3340 21600 3392
rect 22100 3340 22152 3392
rect 23848 3340 23900 3392
rect 24216 3383 24268 3392
rect 24216 3349 24225 3383
rect 24225 3349 24259 3383
rect 24259 3349 24268 3383
rect 24216 3340 24268 3349
rect 24492 3340 24544 3392
rect 24952 3519 25004 3528
rect 24952 3485 24961 3519
rect 24961 3485 24995 3519
rect 24995 3485 25004 3519
rect 24952 3476 25004 3485
rect 26516 3476 26568 3528
rect 25596 3408 25648 3460
rect 25780 3451 25832 3460
rect 25780 3417 25789 3451
rect 25789 3417 25823 3451
rect 25823 3417 25832 3451
rect 25780 3408 25832 3417
rect 25228 3383 25280 3392
rect 25228 3349 25237 3383
rect 25237 3349 25271 3383
rect 25271 3349 25280 3383
rect 25228 3340 25280 3349
rect 25504 3383 25556 3392
rect 25504 3349 25513 3383
rect 25513 3349 25547 3383
rect 25547 3349 25556 3383
rect 25504 3340 25556 3349
rect 25872 3340 25924 3392
rect 27988 3544 28040 3596
rect 28632 3587 28684 3596
rect 28632 3553 28641 3587
rect 28641 3553 28675 3587
rect 28675 3553 28684 3587
rect 28632 3544 28684 3553
rect 28356 3519 28408 3528
rect 28356 3485 28368 3519
rect 28368 3485 28402 3519
rect 28402 3485 28408 3519
rect 28356 3476 28408 3485
rect 28448 3476 28500 3528
rect 29552 3408 29604 3460
rect 4193 3238 4245 3290
rect 4257 3238 4309 3290
rect 4321 3238 4373 3290
rect 4385 3238 4437 3290
rect 4449 3238 4501 3290
rect 11783 3238 11835 3290
rect 11847 3238 11899 3290
rect 11911 3238 11963 3290
rect 11975 3238 12027 3290
rect 12039 3238 12091 3290
rect 19373 3238 19425 3290
rect 19437 3238 19489 3290
rect 19501 3238 19553 3290
rect 19565 3238 19617 3290
rect 19629 3238 19681 3290
rect 26963 3238 27015 3290
rect 27027 3238 27079 3290
rect 27091 3238 27143 3290
rect 27155 3238 27207 3290
rect 27219 3238 27271 3290
rect 1584 3136 1636 3188
rect 3056 3136 3108 3188
rect 3240 3136 3292 3188
rect 3332 3136 3384 3188
rect 6368 3136 6420 3188
rect 940 3043 992 3052
rect 940 3009 949 3043
rect 949 3009 983 3043
rect 983 3009 992 3043
rect 940 3000 992 3009
rect 2964 3000 3016 3052
rect 1676 2975 1728 2984
rect 1676 2941 1685 2975
rect 1685 2941 1719 2975
rect 1719 2941 1728 2975
rect 1676 2932 1728 2941
rect 3608 3068 3660 3120
rect 5264 3000 5316 3052
rect 5816 3000 5868 3052
rect 9680 3136 9732 3188
rect 9864 3136 9916 3188
rect 9588 3000 9640 3052
rect 3700 2932 3752 2984
rect 1768 2796 1820 2848
rect 1952 2796 2004 2848
rect 6460 2932 6512 2984
rect 6184 2864 6236 2916
rect 4160 2796 4212 2848
rect 6920 2796 6972 2848
rect 8852 2932 8904 2984
rect 9312 2932 9364 2984
rect 11704 3136 11756 3188
rect 14740 3136 14792 3188
rect 16580 3136 16632 3188
rect 17132 3136 17184 3188
rect 11796 3000 11848 3052
rect 11244 2975 11296 2984
rect 11244 2941 11253 2975
rect 11253 2941 11287 2975
rect 11287 2941 11296 2975
rect 11244 2932 11296 2941
rect 21548 3136 21600 3188
rect 22100 3136 22152 3188
rect 28172 3068 28224 3120
rect 21456 3000 21508 3052
rect 21824 3000 21876 3052
rect 24492 3000 24544 3052
rect 13636 2932 13688 2984
rect 14096 2975 14148 2984
rect 14096 2941 14105 2975
rect 14105 2941 14139 2975
rect 14139 2941 14148 2975
rect 14096 2932 14148 2941
rect 14188 2932 14240 2984
rect 14832 2975 14884 2984
rect 14832 2941 14841 2975
rect 14841 2941 14875 2975
rect 14875 2941 14884 2975
rect 14832 2932 14884 2941
rect 16672 2975 16724 2984
rect 16672 2941 16674 2975
rect 16674 2941 16724 2975
rect 16672 2932 16724 2941
rect 17040 2975 17092 2984
rect 17040 2941 17049 2975
rect 17049 2941 17083 2975
rect 17083 2941 17092 2975
rect 17040 2932 17092 2941
rect 18512 2932 18564 2984
rect 18696 2975 18748 2984
rect 18696 2941 18705 2975
rect 18705 2941 18739 2975
rect 18739 2941 18748 2975
rect 18696 2932 18748 2941
rect 18972 2932 19024 2984
rect 20904 2975 20956 2984
rect 20904 2941 20913 2975
rect 20913 2941 20947 2975
rect 20947 2941 20956 2975
rect 20904 2932 20956 2941
rect 25964 3000 26016 3052
rect 26424 3043 26476 3052
rect 26424 3009 26426 3043
rect 26426 3009 26476 3043
rect 26424 3000 26476 3009
rect 22008 2932 22060 2984
rect 23848 2975 23900 2984
rect 23848 2941 23857 2975
rect 23857 2941 23891 2975
rect 23891 2941 23900 2975
rect 23848 2932 23900 2941
rect 25780 2932 25832 2984
rect 26700 3000 26752 3052
rect 26976 3000 27028 3052
rect 29092 3000 29144 3052
rect 29276 2975 29328 2984
rect 29276 2941 29285 2975
rect 29285 2941 29319 2975
rect 29319 2941 29328 2975
rect 29276 2932 29328 2941
rect 16212 2864 16264 2916
rect 8392 2796 8444 2848
rect 9036 2796 9088 2848
rect 11980 2796 12032 2848
rect 12256 2796 12308 2848
rect 18788 2796 18840 2848
rect 25964 2907 26016 2916
rect 25964 2873 25973 2907
rect 25973 2873 26007 2907
rect 26007 2873 26016 2907
rect 25964 2864 26016 2873
rect 24124 2796 24176 2848
rect 26792 2796 26844 2848
rect 7988 2694 8040 2746
rect 8052 2694 8104 2746
rect 8116 2694 8168 2746
rect 8180 2694 8232 2746
rect 8244 2694 8296 2746
rect 15578 2694 15630 2746
rect 15642 2694 15694 2746
rect 15706 2694 15758 2746
rect 15770 2694 15822 2746
rect 15834 2694 15886 2746
rect 23168 2694 23220 2746
rect 23232 2694 23284 2746
rect 23296 2694 23348 2746
rect 23360 2694 23412 2746
rect 23424 2694 23476 2746
rect 30758 2694 30810 2746
rect 30822 2694 30874 2746
rect 30886 2694 30938 2746
rect 30950 2694 31002 2746
rect 31014 2694 31066 2746
rect 2044 2592 2096 2644
rect 1860 2456 1912 2508
rect 1676 2388 1728 2440
rect 4068 2592 4120 2644
rect 4620 2592 4672 2644
rect 6184 2592 6236 2644
rect 6644 2592 6696 2644
rect 7012 2592 7064 2644
rect 9036 2592 9088 2644
rect 9312 2592 9364 2644
rect 10048 2592 10100 2644
rect 11520 2592 11572 2644
rect 15292 2592 15344 2644
rect 16580 2592 16632 2644
rect 17224 2592 17276 2644
rect 21640 2592 21692 2644
rect 22008 2592 22060 2644
rect 23848 2635 23900 2644
rect 23848 2601 23857 2635
rect 23857 2601 23891 2635
rect 23891 2601 23900 2635
rect 23848 2592 23900 2601
rect 24216 2592 24268 2644
rect 25780 2592 25832 2644
rect 28448 2635 28500 2644
rect 28448 2601 28463 2635
rect 28463 2601 28497 2635
rect 28497 2601 28500 2635
rect 28448 2592 28500 2601
rect 29368 2592 29420 2644
rect 8668 2524 8720 2576
rect 7656 2456 7708 2508
rect 8760 2456 8812 2508
rect 3424 2388 3476 2440
rect 3792 2388 3844 2440
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 4068 2388 4120 2440
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 6276 2431 6328 2440
rect 6276 2397 6288 2431
rect 6288 2397 6322 2431
rect 6322 2397 6328 2431
rect 6276 2388 6328 2397
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 9312 2456 9364 2508
rect 9404 2499 9456 2508
rect 9404 2465 9413 2499
rect 9413 2465 9447 2499
rect 9447 2465 9456 2499
rect 9404 2456 9456 2465
rect 11244 2456 11296 2508
rect 20536 2567 20588 2576
rect 20536 2533 20545 2567
rect 20545 2533 20579 2567
rect 20579 2533 20588 2567
rect 20536 2524 20588 2533
rect 9128 2431 9180 2440
rect 9128 2397 9140 2431
rect 9140 2397 9174 2431
rect 9174 2397 9180 2431
rect 9128 2388 9180 2397
rect 11796 2388 11848 2440
rect 11980 2431 12032 2440
rect 11980 2397 11982 2431
rect 11982 2397 12032 2431
rect 11980 2388 12032 2397
rect 12164 2388 12216 2440
rect 14004 2388 14056 2440
rect 14188 2431 14240 2440
rect 14188 2397 14190 2431
rect 14190 2397 14240 2431
rect 14188 2388 14240 2397
rect 16120 2456 16172 2508
rect 18420 2499 18472 2508
rect 18420 2465 18429 2499
rect 18429 2465 18463 2499
rect 18463 2465 18472 2499
rect 18420 2456 18472 2465
rect 18788 2499 18840 2508
rect 18788 2465 18790 2499
rect 18790 2465 18840 2499
rect 18788 2456 18840 2465
rect 19248 2456 19300 2508
rect 14556 2431 14608 2440
rect 14556 2397 14565 2431
rect 14565 2397 14599 2431
rect 14599 2397 14608 2431
rect 14556 2388 14608 2397
rect 3516 2252 3568 2304
rect 5356 2252 5408 2304
rect 12164 2252 12216 2304
rect 13544 2252 13596 2304
rect 16488 2252 16540 2304
rect 19156 2431 19208 2440
rect 19156 2397 19165 2431
rect 19165 2397 19199 2431
rect 19199 2397 19208 2431
rect 19156 2388 19208 2397
rect 20904 2456 20956 2508
rect 22744 2456 22796 2508
rect 24032 2456 24084 2508
rect 21456 2388 21508 2440
rect 21824 2388 21876 2440
rect 22836 2388 22888 2440
rect 22928 2388 22980 2440
rect 24400 2388 24452 2440
rect 25228 2456 25280 2508
rect 26240 2456 26292 2508
rect 27436 2524 27488 2576
rect 24952 2388 25004 2440
rect 26056 2388 26108 2440
rect 26332 2388 26384 2440
rect 27252 2456 27304 2508
rect 21088 2320 21140 2372
rect 20628 2252 20680 2304
rect 20812 2252 20864 2304
rect 23664 2320 23716 2372
rect 23940 2252 23992 2304
rect 24584 2252 24636 2304
rect 26792 2388 26844 2440
rect 27436 2388 27488 2440
rect 27988 2499 28040 2508
rect 27988 2465 27997 2499
rect 27997 2465 28031 2499
rect 28031 2465 28040 2499
rect 27988 2456 28040 2465
rect 27620 2388 27672 2440
rect 28724 2499 28776 2508
rect 28724 2465 28733 2499
rect 28733 2465 28767 2499
rect 28767 2465 28776 2499
rect 28724 2456 28776 2465
rect 29092 2388 29144 2440
rect 29460 2388 29512 2440
rect 25596 2252 25648 2304
rect 26056 2252 26108 2304
rect 29368 2252 29420 2304
rect 4193 2150 4245 2202
rect 4257 2150 4309 2202
rect 4321 2150 4373 2202
rect 4385 2150 4437 2202
rect 4449 2150 4501 2202
rect 11783 2150 11835 2202
rect 11847 2150 11899 2202
rect 11911 2150 11963 2202
rect 11975 2150 12027 2202
rect 12039 2150 12091 2202
rect 19373 2150 19425 2202
rect 19437 2150 19489 2202
rect 19501 2150 19553 2202
rect 19565 2150 19617 2202
rect 19629 2150 19681 2202
rect 26963 2150 27015 2202
rect 27027 2150 27079 2202
rect 27091 2150 27143 2202
rect 27155 2150 27207 2202
rect 27219 2150 27271 2202
rect 1676 2048 1728 2100
rect 2320 1912 2372 1964
rect 3884 2048 3936 2100
rect 3976 2048 4028 2100
rect 9864 2048 9916 2100
rect 11980 2048 12032 2100
rect 13544 2048 13596 2100
rect 14832 2048 14884 2100
rect 17040 2048 17092 2100
rect 19156 2048 19208 2100
rect 3884 1955 3936 1964
rect 940 1887 992 1896
rect 940 1853 949 1887
rect 949 1853 983 1887
rect 983 1853 992 1887
rect 940 1844 992 1853
rect 1584 1844 1636 1896
rect 2596 1844 2648 1896
rect 3056 1819 3108 1828
rect 3056 1785 3065 1819
rect 3065 1785 3099 1819
rect 3099 1785 3108 1819
rect 3056 1776 3108 1785
rect 1400 1751 1452 1760
rect 1400 1717 1415 1751
rect 1415 1717 1449 1751
rect 1449 1717 1452 1751
rect 1400 1708 1452 1717
rect 2044 1708 2096 1760
rect 3516 1887 3568 1896
rect 3516 1853 3525 1887
rect 3525 1853 3559 1887
rect 3559 1853 3568 1887
rect 3516 1844 3568 1853
rect 3884 1921 3886 1955
rect 3886 1921 3936 1955
rect 3884 1912 3936 1921
rect 4068 1912 4120 1964
rect 5448 1912 5500 1964
rect 6460 1912 6512 1964
rect 4988 1776 5040 1828
rect 6000 1844 6052 1896
rect 6644 1912 6696 1964
rect 6828 1955 6880 1964
rect 6828 1921 6837 1955
rect 6837 1921 6871 1955
rect 6871 1921 6880 1955
rect 6828 1912 6880 1921
rect 9680 1912 9732 1964
rect 9864 1912 9916 1964
rect 11244 1980 11296 2032
rect 23020 1980 23072 2032
rect 28172 2091 28224 2100
rect 28172 2057 28181 2091
rect 28181 2057 28215 2091
rect 28215 2057 28224 2091
rect 28172 2048 28224 2057
rect 29184 2091 29236 2100
rect 29184 2057 29193 2091
rect 29193 2057 29227 2091
rect 29227 2057 29236 2091
rect 29184 2048 29236 2057
rect 29644 2048 29696 2100
rect 16120 1955 16172 1964
rect 16120 1921 16129 1955
rect 16129 1921 16163 1955
rect 16163 1921 16172 1955
rect 16120 1912 16172 1921
rect 8760 1844 8812 1896
rect 8852 1844 8904 1896
rect 9312 1844 9364 1896
rect 11336 1844 11388 1896
rect 11612 1844 11664 1896
rect 11980 1887 12032 1896
rect 11980 1853 11989 1887
rect 11989 1853 12023 1887
rect 12023 1853 12032 1887
rect 11980 1844 12032 1853
rect 12440 1844 12492 1896
rect 13912 1887 13964 1896
rect 13912 1853 13921 1887
rect 13921 1853 13955 1887
rect 13955 1853 13964 1887
rect 13912 1844 13964 1853
rect 13544 1776 13596 1828
rect 19248 1912 19300 1964
rect 20720 1912 20772 1964
rect 21456 1912 21508 1964
rect 23112 1912 23164 1964
rect 23756 1980 23808 2032
rect 16856 1887 16908 1896
rect 16856 1853 16865 1887
rect 16865 1853 16899 1887
rect 16899 1853 16908 1887
rect 16856 1844 16908 1853
rect 6000 1751 6052 1760
rect 6000 1717 6009 1751
rect 6009 1717 6043 1751
rect 6043 1717 6052 1751
rect 6000 1708 6052 1717
rect 6920 1708 6972 1760
rect 9036 1708 9088 1760
rect 9680 1708 9732 1760
rect 10416 1708 10468 1760
rect 11704 1751 11756 1760
rect 11704 1717 11719 1751
rect 11719 1717 11753 1751
rect 11753 1717 11756 1751
rect 11704 1708 11756 1717
rect 14188 1708 14240 1760
rect 16580 1751 16632 1760
rect 16580 1717 16595 1751
rect 16595 1717 16629 1751
rect 16629 1717 16632 1751
rect 18696 1887 18748 1896
rect 18696 1853 18705 1887
rect 18705 1853 18739 1887
rect 18739 1853 18748 1887
rect 18696 1844 18748 1853
rect 18788 1844 18840 1896
rect 19432 1887 19484 1896
rect 19432 1853 19441 1887
rect 19441 1853 19475 1887
rect 19475 1853 19484 1887
rect 19432 1844 19484 1853
rect 20904 1887 20956 1896
rect 20904 1853 20913 1887
rect 20913 1853 20947 1887
rect 20947 1853 20956 1887
rect 20904 1844 20956 1853
rect 23664 1912 23716 1964
rect 23848 1887 23900 1896
rect 23848 1853 23857 1887
rect 23857 1853 23891 1887
rect 23891 1853 23900 1887
rect 23848 1844 23900 1853
rect 22652 1776 22704 1828
rect 24492 1912 24544 1964
rect 27712 1912 27764 1964
rect 28816 1912 28868 1964
rect 25780 1844 25832 1896
rect 16580 1708 16632 1717
rect 21916 1708 21968 1760
rect 23112 1708 23164 1760
rect 24124 1708 24176 1760
rect 24492 1708 24544 1760
rect 26424 1844 26476 1896
rect 26976 1844 27028 1896
rect 26332 1776 26384 1828
rect 26056 1751 26108 1760
rect 26056 1717 26065 1751
rect 26065 1717 26099 1751
rect 26099 1717 26108 1751
rect 26056 1708 26108 1717
rect 26424 1708 26476 1760
rect 29000 1887 29052 1896
rect 29000 1853 29018 1887
rect 29018 1853 29052 1887
rect 29000 1844 29052 1853
rect 28724 1751 28776 1760
rect 28724 1717 28733 1751
rect 28733 1717 28767 1751
rect 28767 1717 28776 1751
rect 28724 1708 28776 1717
rect 7988 1606 8040 1658
rect 8052 1606 8104 1658
rect 8116 1606 8168 1658
rect 8180 1606 8232 1658
rect 8244 1606 8296 1658
rect 15578 1606 15630 1658
rect 15642 1606 15694 1658
rect 15706 1606 15758 1658
rect 15770 1606 15822 1658
rect 15834 1606 15886 1658
rect 23168 1606 23220 1658
rect 23232 1606 23284 1658
rect 23296 1606 23348 1658
rect 23360 1606 23412 1658
rect 23424 1606 23476 1658
rect 30758 1606 30810 1658
rect 30822 1606 30874 1658
rect 30886 1606 30938 1658
rect 30950 1606 31002 1658
rect 31014 1606 31066 1658
rect 1124 1504 1176 1556
rect 1216 1504 1268 1556
rect 2320 1436 2372 1488
rect 2596 1504 2648 1556
rect 3148 1547 3200 1556
rect 3148 1513 3157 1547
rect 3157 1513 3191 1547
rect 3191 1513 3200 1547
rect 3148 1504 3200 1513
rect 4712 1504 4764 1556
rect 5356 1504 5408 1556
rect 1032 1411 1084 1420
rect 1032 1377 1041 1411
rect 1041 1377 1075 1411
rect 1075 1377 1084 1411
rect 1032 1368 1084 1377
rect 2044 1368 2096 1420
rect 3332 1436 3384 1488
rect 5816 1436 5868 1488
rect 3240 1232 3292 1284
rect 2228 1164 2280 1216
rect 2688 1207 2740 1216
rect 2688 1173 2697 1207
rect 2697 1173 2731 1207
rect 2731 1173 2740 1207
rect 2688 1164 2740 1173
rect 3516 1343 3568 1352
rect 3516 1309 3525 1343
rect 3525 1309 3559 1343
rect 3559 1309 3568 1343
rect 3516 1300 3568 1309
rect 3884 1343 3936 1352
rect 3884 1309 3886 1343
rect 3886 1309 3936 1343
rect 3884 1300 3936 1309
rect 3976 1343 4028 1352
rect 3976 1309 3988 1343
rect 3988 1309 4022 1343
rect 4022 1309 4028 1343
rect 3976 1300 4028 1309
rect 4252 1343 4304 1352
rect 4252 1309 4261 1343
rect 4261 1309 4295 1343
rect 4295 1309 4304 1343
rect 4252 1300 4304 1309
rect 6276 1436 6328 1488
rect 6460 1411 6512 1420
rect 6460 1377 6469 1411
rect 6469 1377 6503 1411
rect 6503 1377 6512 1411
rect 6460 1368 6512 1377
rect 6920 1547 6972 1556
rect 6920 1513 6935 1547
rect 6935 1513 6969 1547
rect 6969 1513 6972 1547
rect 6920 1504 6972 1513
rect 9128 1504 9180 1556
rect 8208 1436 8260 1488
rect 11520 1504 11572 1556
rect 11704 1504 11756 1556
rect 12256 1504 12308 1556
rect 14372 1504 14424 1556
rect 16580 1504 16632 1556
rect 18788 1504 18840 1556
rect 19432 1504 19484 1556
rect 21548 1504 21600 1556
rect 26884 1504 26936 1556
rect 27436 1504 27488 1556
rect 10416 1436 10468 1488
rect 11612 1411 11664 1420
rect 11612 1377 11621 1411
rect 11621 1377 11655 1411
rect 11655 1377 11664 1411
rect 11612 1368 11664 1377
rect 6920 1343 6972 1352
rect 6920 1309 6932 1343
rect 6932 1309 6966 1343
rect 6966 1309 6972 1343
rect 6920 1300 6972 1309
rect 8576 1300 8628 1352
rect 8852 1300 8904 1352
rect 9036 1343 9088 1352
rect 9036 1309 9038 1343
rect 9038 1309 9088 1343
rect 9036 1300 9088 1309
rect 9312 1300 9364 1352
rect 11888 1368 11940 1420
rect 13820 1343 13872 1352
rect 13820 1309 13829 1343
rect 13829 1309 13863 1343
rect 13863 1309 13872 1343
rect 13820 1300 13872 1309
rect 14188 1343 14240 1352
rect 14188 1309 14190 1343
rect 14190 1309 14240 1343
rect 14188 1300 14240 1309
rect 16120 1368 16172 1420
rect 14372 1300 14424 1352
rect 16948 1343 17000 1352
rect 16948 1309 16957 1343
rect 16957 1309 16991 1343
rect 16991 1309 17000 1343
rect 16948 1300 17000 1309
rect 17040 1300 17092 1352
rect 3976 1164 4028 1216
rect 4068 1164 4120 1216
rect 7656 1164 7708 1216
rect 12072 1164 12124 1216
rect 12164 1164 12216 1216
rect 14556 1164 14608 1216
rect 18604 1300 18656 1352
rect 20812 1411 20864 1420
rect 20812 1377 20821 1411
rect 20821 1377 20855 1411
rect 20855 1377 20864 1411
rect 20812 1368 20864 1377
rect 21088 1411 21140 1420
rect 21088 1377 21097 1411
rect 21097 1377 21131 1411
rect 21131 1377 21140 1411
rect 21088 1368 21140 1377
rect 20996 1300 21048 1352
rect 23572 1436 23624 1488
rect 24952 1436 25004 1488
rect 25780 1479 25832 1488
rect 25780 1445 25789 1479
rect 25789 1445 25823 1479
rect 25823 1445 25832 1479
rect 25780 1436 25832 1445
rect 24860 1368 24912 1420
rect 26516 1436 26568 1488
rect 25964 1368 26016 1420
rect 20628 1207 20680 1216
rect 20628 1173 20637 1207
rect 20637 1173 20671 1207
rect 20671 1173 20680 1207
rect 20628 1164 20680 1173
rect 20904 1232 20956 1284
rect 23664 1300 23716 1352
rect 23940 1343 23992 1352
rect 23940 1309 23952 1343
rect 23952 1309 23986 1343
rect 23986 1309 23992 1343
rect 23940 1300 23992 1309
rect 24124 1300 24176 1352
rect 25412 1300 25464 1352
rect 23020 1164 23072 1216
rect 23388 1164 23440 1216
rect 24032 1164 24084 1216
rect 25688 1232 25740 1284
rect 26608 1300 26660 1352
rect 26976 1300 27028 1352
rect 27988 1504 28040 1556
rect 28356 1504 28408 1556
rect 29368 1504 29420 1556
rect 28632 1368 28684 1420
rect 29000 1368 29052 1420
rect 29368 1368 29420 1420
rect 25320 1207 25372 1216
rect 25320 1173 25329 1207
rect 25329 1173 25363 1207
rect 25363 1173 25372 1207
rect 25320 1164 25372 1173
rect 26148 1164 26200 1216
rect 26976 1164 27028 1216
rect 28632 1207 28684 1216
rect 28632 1173 28641 1207
rect 28641 1173 28675 1207
rect 28675 1173 28684 1207
rect 28632 1164 28684 1173
rect 29368 1207 29420 1216
rect 29368 1173 29377 1207
rect 29377 1173 29411 1207
rect 29411 1173 29420 1207
rect 29368 1164 29420 1173
rect 4193 1062 4245 1114
rect 4257 1062 4309 1114
rect 4321 1062 4373 1114
rect 4385 1062 4437 1114
rect 4449 1062 4501 1114
rect 11783 1062 11835 1114
rect 11847 1062 11899 1114
rect 11911 1062 11963 1114
rect 11975 1062 12027 1114
rect 12039 1062 12091 1114
rect 19373 1062 19425 1114
rect 19437 1062 19489 1114
rect 19501 1062 19553 1114
rect 19565 1062 19617 1114
rect 19629 1062 19681 1114
rect 26963 1062 27015 1114
rect 27027 1062 27079 1114
rect 27091 1062 27143 1114
rect 27155 1062 27207 1114
rect 27219 1062 27271 1114
rect 6920 960 6972 1012
rect 7656 1003 7708 1012
rect 7656 969 7665 1003
rect 7665 969 7699 1003
rect 7699 969 7708 1003
rect 7656 960 7708 969
rect 9312 960 9364 1012
rect 10600 1003 10652 1012
rect 10600 969 10609 1003
rect 10609 969 10643 1003
rect 10643 969 10652 1003
rect 10600 960 10652 969
rect 12164 960 12216 1012
rect 12348 960 12400 1012
rect 940 867 992 876
rect 940 833 949 867
rect 949 833 983 867
rect 983 833 992 867
rect 940 824 992 833
rect 1676 867 1728 876
rect 1676 833 1685 867
rect 1685 833 1719 867
rect 1719 833 1728 867
rect 1676 824 1728 833
rect 5172 892 5224 944
rect 13360 960 13412 1012
rect 13544 1003 13596 1012
rect 13544 969 13553 1003
rect 13553 969 13587 1003
rect 13587 969 13596 1003
rect 13544 960 13596 969
rect 16856 960 16908 1012
rect 16948 960 17000 1012
rect 16212 892 16264 944
rect 17960 892 18012 944
rect 20444 960 20496 1012
rect 6276 865 6328 876
rect 6276 831 6288 865
rect 6288 831 6322 865
rect 6322 831 6328 865
rect 6276 824 6328 831
rect 6644 824 6696 876
rect 3608 756 3660 808
rect 4988 799 5040 808
rect 4988 765 4997 799
rect 4997 765 5031 799
rect 5031 765 5040 799
rect 4988 756 5040 765
rect 5632 799 5684 808
rect 5632 765 5641 799
rect 5641 765 5675 799
rect 5675 765 5684 799
rect 5632 756 5684 765
rect 5816 799 5868 808
rect 5816 765 5825 799
rect 5825 765 5859 799
rect 5859 765 5868 799
rect 5816 756 5868 765
rect 7840 756 7892 808
rect 8392 867 8444 876
rect 8392 833 8401 867
rect 8401 833 8435 867
rect 8435 833 8444 867
rect 8392 824 8444 833
rect 10508 824 10560 876
rect 9036 756 9088 808
rect 11612 824 11664 876
rect 12072 824 12124 876
rect 11152 799 11204 808
rect 11152 765 11161 799
rect 11161 765 11195 799
rect 11195 765 11204 799
rect 11152 756 11204 765
rect 11888 756 11940 808
rect 12256 756 12308 808
rect 1400 663 1452 672
rect 1400 629 1415 663
rect 1415 629 1449 663
rect 1449 629 1452 663
rect 1400 620 1452 629
rect 1676 620 1728 672
rect 5356 663 5408 672
rect 5356 629 5365 663
rect 5365 629 5399 663
rect 5399 629 5408 663
rect 5356 620 5408 629
rect 5448 663 5500 672
rect 5448 629 5457 663
rect 5457 629 5491 663
rect 5491 629 5500 663
rect 5448 620 5500 629
rect 7564 620 7616 672
rect 8300 620 8352 672
rect 9128 620 9180 672
rect 11336 620 11388 672
rect 12072 620 12124 672
rect 12256 620 12308 672
rect 14372 824 14424 876
rect 17040 824 17092 876
rect 18788 824 18840 876
rect 13728 799 13780 808
rect 13728 765 13729 799
rect 13729 765 13763 799
rect 13763 765 13780 799
rect 13728 756 13780 765
rect 13820 799 13872 808
rect 13820 765 13829 799
rect 13829 765 13863 799
rect 13863 765 13872 799
rect 13820 756 13872 765
rect 14464 756 14516 808
rect 15016 756 15068 808
rect 16304 799 16356 808
rect 16304 765 16313 799
rect 16313 765 16347 799
rect 16347 765 16356 799
rect 16304 756 16356 765
rect 16396 799 16448 808
rect 16396 765 16405 799
rect 16405 765 16439 799
rect 16439 765 16448 799
rect 16396 756 16448 765
rect 25320 960 25372 1012
rect 25412 960 25464 1012
rect 28540 1003 28592 1012
rect 28540 969 28549 1003
rect 28549 969 28583 1003
rect 28583 969 28592 1003
rect 28540 960 28592 969
rect 20904 892 20956 944
rect 25504 892 25556 944
rect 26148 892 26200 944
rect 20812 824 20864 876
rect 21548 867 21600 876
rect 21548 833 21557 867
rect 21557 833 21591 867
rect 21591 833 21600 867
rect 21548 824 21600 833
rect 16488 688 16540 740
rect 13636 620 13688 672
rect 18236 663 18288 672
rect 18236 629 18245 663
rect 18245 629 18279 663
rect 18279 629 18288 663
rect 18236 620 18288 629
rect 18420 688 18472 740
rect 21272 756 21324 808
rect 20444 688 20496 740
rect 21640 756 21692 808
rect 23020 756 23072 808
rect 23572 824 23624 876
rect 24584 867 24636 876
rect 24584 833 24593 867
rect 24593 833 24627 867
rect 24627 833 24636 867
rect 24584 824 24636 833
rect 25228 824 25280 876
rect 26424 824 26476 876
rect 26884 824 26936 876
rect 23664 799 23716 808
rect 23664 765 23673 799
rect 23673 765 23707 799
rect 23707 765 23716 799
rect 23664 756 23716 765
rect 23848 799 23900 808
rect 23848 765 23857 799
rect 23857 765 23891 799
rect 23891 765 23900 799
rect 23848 756 23900 765
rect 20536 620 20588 672
rect 20812 663 20864 672
rect 20812 629 20821 663
rect 20821 629 20855 663
rect 20855 629 20864 663
rect 20812 620 20864 629
rect 23756 688 23808 740
rect 24492 756 24544 808
rect 26608 799 26660 808
rect 26608 765 26617 799
rect 26617 765 26651 799
rect 26651 765 26660 799
rect 26608 756 26660 765
rect 26792 756 26844 808
rect 27344 824 27396 876
rect 27528 756 27580 808
rect 29460 756 29512 808
rect 24124 620 24176 672
rect 25688 663 25740 672
rect 25688 629 25697 663
rect 25697 629 25731 663
rect 25731 629 25740 663
rect 25688 620 25740 629
rect 26056 663 26108 672
rect 26056 629 26065 663
rect 26065 629 26099 663
rect 26099 629 26108 663
rect 26056 620 26108 629
rect 7988 518 8040 570
rect 8052 518 8104 570
rect 8116 518 8168 570
rect 8180 518 8232 570
rect 8244 518 8296 570
rect 15578 518 15630 570
rect 15642 518 15694 570
rect 15706 518 15758 570
rect 15770 518 15822 570
rect 15834 518 15886 570
rect 23168 518 23220 570
rect 23232 518 23284 570
rect 23296 518 23348 570
rect 23360 518 23412 570
rect 23424 518 23476 570
rect 30758 518 30810 570
rect 30822 518 30874 570
rect 30886 518 30938 570
rect 30950 518 31002 570
rect 31014 518 31066 570
rect 3976 416 4028 468
rect 6920 416 6972 468
rect 7564 416 7616 468
rect 7840 416 7892 468
rect 20720 416 20772 468
rect 23756 416 23808 468
rect 25596 416 25648 468
rect 13636 348 13688 400
rect 14464 348 14516 400
rect 18604 348 18656 400
rect 23020 348 23072 400
rect 25872 348 25924 400
rect 5448 280 5500 332
rect 11520 280 11572 332
rect 11612 280 11664 332
rect 13728 280 13780 332
rect 13820 280 13872 332
rect 18512 280 18564 332
rect 22836 280 22888 332
rect 26056 280 26108 332
rect 6000 212 6052 264
rect 9036 212 9088 264
rect 12348 212 12400 264
rect 21272 212 21324 264
rect 28632 212 28684 264
rect 5080 144 5132 196
rect 5356 144 5408 196
rect 15384 144 15436 196
rect 18788 144 18840 196
rect 28356 144 28408 196
rect 9128 76 9180 128
rect 22744 76 22796 128
rect 5816 8 5868 60
rect 16396 8 16448 60
rect 18420 8 18472 60
rect 18604 8 18656 60
rect 19708 8 19760 60
rect 26792 8 26844 60
<< metal2 >>
rect 1952 22296 2004 22302
rect 8852 22296 8904 22302
rect 1952 22238 2004 22244
rect 8850 22264 8852 22273
rect 9680 22296 9732 22302
rect 8904 22264 8906 22273
rect 1674 21584 1730 21593
rect 1674 21519 1730 21528
rect 1688 21486 1716 21519
rect 1676 21480 1728 21486
rect 1676 21422 1728 21428
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 1412 21010 1440 21286
rect 1964 21078 1992 22238
rect 4068 22228 4120 22234
rect 9678 22264 9680 22273
rect 18788 22296 18840 22302
rect 9732 22264 9734 22273
rect 8850 22199 8906 22208
rect 9128 22228 9180 22234
rect 4068 22170 4120 22176
rect 12636 22234 12940 22250
rect 23572 22296 23624 22302
rect 18788 22238 18840 22244
rect 21638 22264 21694 22273
rect 9678 22199 9734 22208
rect 9772 22228 9824 22234
rect 9128 22170 9180 22176
rect 9772 22170 9824 22176
rect 12636 22228 12952 22234
rect 12636 22222 12900 22228
rect 3056 22160 3108 22166
rect 3056 22102 3108 22108
rect 2136 21888 2188 21894
rect 2136 21830 2188 21836
rect 2504 21888 2556 21894
rect 2504 21830 2556 21836
rect 2148 21078 2176 21830
rect 1952 21072 2004 21078
rect 1952 21014 2004 21020
rect 2136 21072 2188 21078
rect 2136 21014 2188 21020
rect 1124 21004 1176 21010
rect 1124 20946 1176 20952
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 848 19848 900 19854
rect 848 19790 900 19796
rect 860 19378 888 19790
rect 848 19372 900 19378
rect 848 19314 900 19320
rect 860 18698 888 19314
rect 1030 18864 1086 18873
rect 1136 18834 1164 20946
rect 1216 20392 1268 20398
rect 1584 20392 1636 20398
rect 1216 20334 1268 20340
rect 1582 20360 1584 20369
rect 1636 20360 1638 20369
rect 1228 18902 1256 20334
rect 1582 20295 1638 20304
rect 1308 20256 1360 20262
rect 1308 20198 1360 20204
rect 1320 18902 1348 20198
rect 1400 20052 1452 20058
rect 1400 19994 1452 20000
rect 1412 19174 1440 19994
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1596 19417 1624 19790
rect 1582 19408 1638 19417
rect 1582 19343 1638 19352
rect 2044 19372 2096 19378
rect 2044 19314 2096 19320
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1400 19168 1452 19174
rect 1400 19110 1452 19116
rect 1216 18896 1268 18902
rect 1216 18838 1268 18844
rect 1308 18896 1360 18902
rect 1308 18838 1360 18844
rect 1030 18799 1032 18808
rect 1084 18799 1086 18808
rect 1124 18828 1176 18834
rect 1032 18770 1084 18776
rect 1124 18770 1176 18776
rect 848 18692 900 18698
rect 848 18634 900 18640
rect 860 18290 888 18634
rect 848 18284 900 18290
rect 848 18226 900 18232
rect 860 17746 888 18226
rect 1412 18086 1440 19110
rect 1584 18760 1636 18766
rect 1582 18728 1584 18737
rect 1636 18728 1638 18737
rect 1582 18663 1638 18672
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 1412 17882 1440 18022
rect 1400 17876 1452 17882
rect 1400 17818 1452 17824
rect 848 17740 900 17746
rect 848 17682 900 17688
rect 1674 17640 1730 17649
rect 1674 17575 1730 17584
rect 1308 17128 1360 17134
rect 1308 17070 1360 17076
rect 940 16652 992 16658
rect 860 16612 940 16640
rect 860 9058 888 16612
rect 940 16594 992 16600
rect 1320 16046 1348 17070
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15366 1348 15982
rect 1412 15910 1440 16934
rect 1688 16590 1716 17575
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1412 15706 1440 15846
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 940 15360 992 15366
rect 940 15302 992 15308
rect 1308 15360 1360 15366
rect 1308 15302 1360 15308
rect 952 11354 980 15302
rect 1320 15026 1348 15302
rect 1308 15020 1360 15026
rect 1308 14962 1360 14968
rect 1412 14822 1440 15642
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1688 15162 1716 15438
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1964 15065 1992 19246
rect 2056 16250 2084 19314
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 2424 18426 2452 18702
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2412 18216 2464 18222
rect 2412 18158 2464 18164
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 2042 16144 2098 16153
rect 2042 16079 2098 16088
rect 1950 15056 2006 15065
rect 1950 14991 2006 15000
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 1398 14512 1454 14521
rect 1124 14476 1176 14482
rect 1398 14447 1400 14456
rect 1124 14418 1176 14424
rect 1452 14447 1454 14456
rect 1400 14418 1452 14424
rect 1136 14074 1164 14418
rect 2056 14414 2084 16079
rect 2148 15473 2176 17070
rect 2424 16522 2452 18158
rect 2412 16516 2464 16522
rect 2412 16458 2464 16464
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2134 15464 2190 15473
rect 2134 15399 2190 15408
rect 1492 14408 1544 14414
rect 1492 14350 1544 14356
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 1124 14068 1176 14074
rect 1124 14010 1176 14016
rect 1136 13326 1164 14010
rect 1216 13864 1268 13870
rect 1216 13806 1268 13812
rect 1124 13320 1176 13326
rect 1124 13262 1176 13268
rect 1032 13184 1084 13190
rect 1032 13126 1084 13132
rect 1044 12442 1072 13126
rect 1032 12436 1084 12442
rect 1032 12378 1084 12384
rect 940 11348 992 11354
rect 940 11290 992 11296
rect 940 10124 992 10130
rect 940 10066 992 10072
rect 952 9586 980 10066
rect 1136 10010 1164 13262
rect 1228 11694 1256 13806
rect 1400 13728 1452 13734
rect 1400 13670 1452 13676
rect 1308 13320 1360 13326
rect 1308 13262 1360 13268
rect 1320 12850 1348 13262
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 1320 12238 1348 12786
rect 1308 12232 1360 12238
rect 1308 12174 1360 12180
rect 1216 11688 1268 11694
rect 1216 11630 1268 11636
rect 1044 9982 1164 10010
rect 940 9580 992 9586
rect 940 9522 992 9528
rect 1044 9489 1072 9982
rect 1124 9716 1176 9722
rect 1124 9658 1176 9664
rect 1030 9480 1086 9489
rect 1030 9415 1086 9424
rect 860 9030 980 9058
rect 848 8968 900 8974
rect 848 8910 900 8916
rect 860 8430 888 8910
rect 952 8838 980 9030
rect 940 8832 992 8838
rect 940 8774 992 8780
rect 848 8424 900 8430
rect 848 8366 900 8372
rect 860 7886 888 8366
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 860 7342 888 7822
rect 848 7336 900 7342
rect 848 7278 900 7284
rect 860 6798 888 7278
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 860 6254 888 6734
rect 848 6248 900 6254
rect 848 6190 900 6196
rect 860 4690 888 6190
rect 1044 5778 1072 9415
rect 1032 5772 1084 5778
rect 1032 5714 1084 5720
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 848 4684 900 4690
rect 848 4626 900 4632
rect 952 4146 980 5170
rect 940 4140 992 4146
rect 940 4082 992 4088
rect 952 3058 980 4082
rect 1030 3904 1086 3913
rect 1030 3839 1086 3848
rect 1044 3534 1072 3839
rect 1032 3528 1084 3534
rect 1032 3470 1084 3476
rect 940 3052 992 3058
rect 940 2994 992 3000
rect 940 1896 992 1902
rect 940 1838 992 1844
rect 952 882 980 1838
rect 1044 1426 1072 3470
rect 1136 1562 1164 9658
rect 1228 5914 1256 11630
rect 1320 11098 1348 12174
rect 1412 11558 1440 13670
rect 1504 13326 1532 14350
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1688 12986 1716 13806
rect 1780 13530 1808 14350
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1676 12640 1728 12646
rect 1780 12628 1808 13466
rect 1728 12600 1808 12628
rect 1676 12582 1728 12588
rect 1688 12238 1716 12582
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1964 12238 1992 12378
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1860 12232 1912 12238
rect 1860 12174 1912 12180
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1400 11144 1452 11150
rect 1398 11112 1400 11121
rect 1452 11112 1454 11121
rect 1320 11070 1398 11098
rect 1320 10674 1348 11070
rect 1398 11047 1454 11056
rect 1308 10668 1360 10674
rect 1308 10610 1360 10616
rect 1320 10266 1348 10610
rect 1308 10260 1360 10266
rect 1308 10202 1360 10208
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 1412 9382 1440 10202
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1412 8294 1440 8910
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 7886 1440 8230
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7206 1440 7822
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1412 6798 1440 7142
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6118 1440 6734
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1216 5908 1268 5914
rect 1216 5850 1268 5856
rect 1216 5772 1268 5778
rect 1216 5714 1268 5720
rect 1308 5772 1360 5778
rect 1308 5714 1360 5720
rect 1228 1562 1256 5714
rect 1320 5370 1348 5714
rect 1308 5364 1360 5370
rect 1308 5306 1360 5312
rect 1412 4282 1440 6054
rect 1504 4826 1532 11698
rect 1596 9518 1624 12038
rect 1688 11393 1716 12174
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1780 11694 1808 12038
rect 1768 11688 1820 11694
rect 1768 11630 1820 11636
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1674 11384 1730 11393
rect 1674 11319 1730 11328
rect 1688 11150 1716 11319
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1688 10470 1716 11086
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10266 1716 10406
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1674 10160 1730 10169
rect 1780 10146 1808 11494
rect 1872 11014 1900 12174
rect 2056 11370 2084 13874
rect 2134 13696 2190 13705
rect 2134 13631 2190 13640
rect 2148 12782 2176 13631
rect 2136 12776 2188 12782
rect 2136 12718 2188 12724
rect 2240 12617 2268 14350
rect 2226 12608 2282 12617
rect 2226 12543 2282 12552
rect 1964 11342 2084 11370
rect 2136 11348 2188 11354
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1964 10452 1992 11342
rect 2136 11290 2188 11296
rect 2148 11218 2176 11290
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2134 10704 2190 10713
rect 2134 10639 2136 10648
rect 2188 10639 2190 10648
rect 2136 10610 2188 10616
rect 1964 10424 2084 10452
rect 1780 10118 1992 10146
rect 1674 10095 1730 10104
rect 1688 10062 1716 10095
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1780 9722 1808 9998
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1676 7880 1728 7886
rect 1780 7857 1808 8910
rect 1676 7822 1728 7828
rect 1766 7848 1822 7857
rect 1688 7732 1716 7822
rect 1766 7783 1822 7792
rect 1688 7704 1808 7732
rect 1674 7304 1730 7313
rect 1674 7239 1730 7248
rect 1688 6254 1716 7239
rect 1780 7041 1808 7704
rect 1766 7032 1822 7041
rect 1766 6967 1822 6976
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1780 6662 1808 6734
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1872 6474 1900 9658
rect 1964 7528 1992 10118
rect 2056 8634 2084 10424
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1964 7500 2084 7528
rect 1950 7440 2006 7449
rect 1950 7375 2006 7384
rect 1780 6446 1900 6474
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1596 5166 1624 5850
rect 1584 5160 1636 5166
rect 1636 5108 1716 5114
rect 1584 5102 1716 5108
rect 1596 5086 1716 5102
rect 1492 4820 1544 4826
rect 1492 4762 1544 4768
rect 1582 4720 1638 4729
rect 1582 4655 1638 4664
rect 1596 4622 1624 4655
rect 1492 4616 1544 4622
rect 1492 4558 1544 4564
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1504 4486 1532 4558
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1400 4276 1452 4282
rect 1400 4218 1452 4224
rect 1688 3942 1716 5086
rect 1780 4078 1808 6446
rect 1964 5166 1992 7375
rect 2056 6254 2084 7500
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 2056 5914 2084 6190
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 2042 5808 2098 5817
rect 2042 5743 2098 5752
rect 2056 5710 2084 5743
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2148 5234 2176 7142
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 1860 4684 1912 4690
rect 1860 4626 1912 4632
rect 1872 4282 1900 4626
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1676 3936 1728 3942
rect 1728 3896 1808 3924
rect 1676 3878 1728 3884
rect 1676 3528 1728 3534
rect 1780 3505 1808 3896
rect 2042 3632 2098 3641
rect 2042 3567 2098 3576
rect 2056 3534 2084 3567
rect 2044 3528 2096 3534
rect 1676 3470 1728 3476
rect 1766 3496 1822 3505
rect 1688 3398 1716 3470
rect 2044 3470 2096 3476
rect 1766 3431 1822 3440
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1596 3194 1624 3334
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1674 3088 1730 3097
rect 1674 3023 1730 3032
rect 1688 2990 1716 3023
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1780 2854 1808 3431
rect 1768 2848 1820 2854
rect 1398 2816 1454 2825
rect 1768 2790 1820 2796
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 1398 2751 1454 2760
rect 1412 1766 1440 2751
rect 1858 2680 1914 2689
rect 1858 2615 1914 2624
rect 1872 2514 1900 2615
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 1676 2440 1728 2446
rect 1676 2382 1728 2388
rect 1688 2106 1716 2382
rect 1676 2100 1728 2106
rect 1676 2042 1728 2048
rect 1584 1896 1636 1902
rect 1964 1884 1992 2790
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 2056 2009 2084 2586
rect 2042 2000 2098 2009
rect 2332 1970 2360 16390
rect 2516 16046 2544 21830
rect 2780 21684 2832 21690
rect 2780 21626 2832 21632
rect 2792 20942 2820 21626
rect 2964 21004 3016 21010
rect 2964 20946 3016 20952
rect 2780 20936 2832 20942
rect 2780 20878 2832 20884
rect 2792 20584 2820 20878
rect 2976 20754 3004 20946
rect 3068 20942 3096 22102
rect 3792 21888 3844 21894
rect 3792 21830 3844 21836
rect 3424 21548 3476 21554
rect 3424 21490 3476 21496
rect 3240 21480 3292 21486
rect 3240 21422 3292 21428
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 2976 20726 3188 20754
rect 2792 20556 3004 20584
rect 2780 20460 2832 20466
rect 2780 20402 2832 20408
rect 2792 17882 2820 20402
rect 2976 19854 3004 20556
rect 2964 19848 3016 19854
rect 2964 19790 3016 19796
rect 3160 19836 3188 20726
rect 3252 19938 3280 21422
rect 3436 20058 3464 21490
rect 3516 21344 3568 21350
rect 3516 21286 3568 21292
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 3252 19910 3372 19938
rect 3240 19848 3292 19854
rect 3160 19808 3240 19836
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2884 17338 2912 19654
rect 2976 19378 3004 19790
rect 2964 19372 3016 19378
rect 2964 19314 3016 19320
rect 3160 19310 3188 19808
rect 3240 19790 3292 19796
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 2964 18760 3016 18766
rect 2964 18702 3016 18708
rect 2976 18426 3004 18702
rect 2964 18420 3016 18426
rect 2964 18362 3016 18368
rect 3148 18284 3200 18290
rect 3148 18226 3200 18232
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2424 11937 2452 15438
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 2410 11928 2466 11937
rect 2410 11863 2466 11872
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2424 8566 2452 8774
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2042 1935 2098 1944
rect 2320 1964 2372 1970
rect 2320 1906 2372 1912
rect 1636 1856 1992 1884
rect 1584 1838 1636 1844
rect 1400 1760 1452 1766
rect 1400 1702 1452 1708
rect 2044 1760 2096 1766
rect 2044 1702 2096 1708
rect 1124 1556 1176 1562
rect 1124 1498 1176 1504
rect 1216 1556 1268 1562
rect 1216 1498 1268 1504
rect 1032 1420 1084 1426
rect 1032 1362 1084 1368
rect 940 876 992 882
rect 940 818 992 824
rect 1412 678 1440 1702
rect 2056 1426 2084 1702
rect 2424 1578 2452 7278
rect 2516 6662 2544 13806
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2608 7886 2636 12582
rect 2700 12209 2728 14894
rect 2792 14074 2820 16526
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2884 12434 2912 16730
rect 2976 15162 3004 17682
rect 3160 15706 3188 18226
rect 3252 18222 3280 19314
rect 3344 18426 3372 19910
rect 3528 18834 3556 21286
rect 3804 21010 3832 21830
rect 3974 21584 4030 21593
rect 3974 21519 4030 21528
rect 3988 21486 4016 21519
rect 3976 21480 4028 21486
rect 3976 21422 4028 21428
rect 3792 21004 3844 21010
rect 3792 20946 3844 20952
rect 3700 20936 3752 20942
rect 3700 20878 3752 20884
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3620 19854 3648 20198
rect 3712 19854 3740 20878
rect 4080 20806 4108 22170
rect 7194 22128 7250 22137
rect 5264 22092 5316 22098
rect 7194 22063 7250 22072
rect 5264 22034 5316 22040
rect 4193 21788 4501 21797
rect 4193 21786 4199 21788
rect 4255 21786 4279 21788
rect 4335 21786 4359 21788
rect 4415 21786 4439 21788
rect 4495 21786 4501 21788
rect 4255 21734 4257 21786
rect 4437 21734 4439 21786
rect 4193 21732 4199 21734
rect 4255 21732 4279 21734
rect 4335 21732 4359 21734
rect 4415 21732 4439 21734
rect 4495 21732 4501 21734
rect 4193 21723 4501 21732
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 4193 20700 4501 20709
rect 4193 20698 4199 20700
rect 4255 20698 4279 20700
rect 4335 20698 4359 20700
rect 4415 20698 4439 20700
rect 4495 20698 4501 20700
rect 4255 20646 4257 20698
rect 4437 20646 4439 20698
rect 4193 20644 4199 20646
rect 4255 20644 4279 20646
rect 4335 20644 4359 20646
rect 4415 20644 4439 20646
rect 4495 20644 4501 20646
rect 4193 20635 4501 20644
rect 4540 20466 4568 20742
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 4620 20460 4672 20466
rect 4620 20402 4672 20408
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 4264 20058 4292 20198
rect 4252 20052 4304 20058
rect 4252 19994 4304 20000
rect 3608 19848 3660 19854
rect 3608 19790 3660 19796
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 4193 19612 4501 19621
rect 4193 19610 4199 19612
rect 4255 19610 4279 19612
rect 4335 19610 4359 19612
rect 4415 19610 4439 19612
rect 4495 19610 4501 19612
rect 4255 19558 4257 19610
rect 4437 19558 4439 19610
rect 4193 19556 4199 19558
rect 4255 19556 4279 19558
rect 4335 19556 4359 19558
rect 4415 19556 4439 19558
rect 4495 19556 4501 19558
rect 4193 19547 4501 19556
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 3896 19145 3924 19246
rect 3882 19136 3938 19145
rect 3882 19071 3938 19080
rect 3516 18828 3568 18834
rect 3792 18828 3844 18834
rect 3516 18770 3568 18776
rect 3712 18788 3792 18816
rect 3712 18737 3740 18788
rect 3792 18770 3844 18776
rect 3698 18728 3754 18737
rect 3698 18663 3754 18672
rect 3332 18420 3384 18426
rect 3332 18362 3384 18368
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3344 18086 3372 18362
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3528 17882 3556 18362
rect 3606 17912 3662 17921
rect 3516 17876 3568 17882
rect 3606 17847 3662 17856
rect 3516 17818 3568 17824
rect 3620 17746 3648 17847
rect 3608 17740 3660 17746
rect 3608 17682 3660 17688
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 3252 14634 3280 16526
rect 3344 16046 3372 17138
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3330 14648 3386 14657
rect 3252 14606 3330 14634
rect 3330 14583 3386 14592
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3146 13424 3202 13433
rect 3146 13359 3148 13368
rect 3200 13359 3202 13368
rect 3148 13330 3200 13336
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3068 12753 3096 12786
rect 3054 12744 3110 12753
rect 3054 12679 3110 12688
rect 3160 12434 3188 12922
rect 2792 12406 2912 12434
rect 3068 12406 3188 12434
rect 2686 12200 2742 12209
rect 2686 12135 2742 12144
rect 2792 8362 2820 12406
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2884 9081 2912 12242
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2976 10062 3004 10406
rect 3068 10282 3096 12406
rect 3252 11830 3280 14350
rect 3436 14074 3464 17614
rect 3712 17134 3740 18663
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3896 18222 3924 18566
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3896 17678 3924 18158
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3804 17338 3832 17478
rect 3896 17338 3924 17614
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3528 15994 3556 16526
rect 3528 15966 3648 15994
rect 3620 15910 3648 15966
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3514 15600 3570 15609
rect 3620 15570 3648 15846
rect 3514 15535 3570 15544
rect 3608 15564 3660 15570
rect 3528 15026 3556 15535
rect 3608 15506 3660 15512
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3712 14958 3740 17070
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3896 15910 3924 16526
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 15502 3924 15846
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 15026 3832 15302
rect 3792 15020 3844 15026
rect 3792 14962 3844 14968
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3896 14822 3924 15438
rect 3988 15065 4016 19246
rect 4264 18970 4292 19246
rect 4632 19009 4660 20402
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 4724 19242 4752 20334
rect 4712 19236 4764 19242
rect 4712 19178 4764 19184
rect 4618 19000 4674 19009
rect 4252 18964 4304 18970
rect 4618 18935 4674 18944
rect 4252 18906 4304 18912
rect 4724 18902 4752 19178
rect 4620 18896 4672 18902
rect 4620 18838 4672 18844
rect 4712 18896 4764 18902
rect 4816 18873 4844 21422
rect 5276 21078 5304 22034
rect 7208 21962 7236 22063
rect 7196 21956 7248 21962
rect 7196 21898 7248 21904
rect 8760 21888 8812 21894
rect 8760 21830 8812 21836
rect 8852 21888 8904 21894
rect 8852 21830 8904 21836
rect 5814 21720 5870 21729
rect 5814 21655 5870 21664
rect 8208 21684 8260 21690
rect 5540 21616 5592 21622
rect 5540 21558 5592 21564
rect 5552 21486 5580 21558
rect 5540 21480 5592 21486
rect 5540 21422 5592 21428
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5264 21072 5316 21078
rect 5264 21014 5316 21020
rect 4988 21004 5040 21010
rect 4988 20946 5040 20952
rect 4712 18838 4764 18844
rect 4802 18864 4858 18873
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 4080 18290 4108 18566
rect 4193 18524 4501 18533
rect 4193 18522 4199 18524
rect 4255 18522 4279 18524
rect 4335 18522 4359 18524
rect 4415 18522 4439 18524
rect 4495 18522 4501 18524
rect 4255 18470 4257 18522
rect 4437 18470 4439 18522
rect 4193 18468 4199 18470
rect 4255 18468 4279 18470
rect 4335 18468 4359 18470
rect 4415 18468 4439 18470
rect 4495 18468 4501 18470
rect 4193 18459 4501 18468
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 4264 17882 4292 18226
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4356 17746 4384 18226
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 4080 17218 4108 17614
rect 4193 17436 4501 17445
rect 4193 17434 4199 17436
rect 4255 17434 4279 17436
rect 4335 17434 4359 17436
rect 4415 17434 4439 17436
rect 4495 17434 4501 17436
rect 4255 17382 4257 17434
rect 4437 17382 4439 17434
rect 4193 17380 4199 17382
rect 4255 17380 4279 17382
rect 4335 17380 4359 17382
rect 4415 17380 4439 17382
rect 4495 17380 4501 17382
rect 4193 17371 4501 17380
rect 4080 17190 4200 17218
rect 4172 16794 4200 17190
rect 4540 16998 4568 17818
rect 4528 16992 4580 16998
rect 4528 16934 4580 16940
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4193 16348 4501 16357
rect 4193 16346 4199 16348
rect 4255 16346 4279 16348
rect 4335 16346 4359 16348
rect 4415 16346 4439 16348
rect 4495 16346 4501 16348
rect 4255 16294 4257 16346
rect 4437 16294 4439 16346
rect 4193 16292 4199 16294
rect 4255 16292 4279 16294
rect 4335 16292 4359 16294
rect 4415 16292 4439 16294
rect 4495 16292 4501 16294
rect 4193 16283 4501 16292
rect 4632 16250 4660 18838
rect 4802 18799 4858 18808
rect 4816 18136 4844 18799
rect 5000 18578 5028 20946
rect 5276 20806 5304 21014
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 5080 19712 5132 19718
rect 5080 19654 5132 19660
rect 5092 19514 5120 19654
rect 5170 19544 5226 19553
rect 5080 19508 5132 19514
rect 5170 19479 5226 19488
rect 5080 19450 5132 19456
rect 5184 19174 5212 19479
rect 5172 19168 5224 19174
rect 5172 19110 5224 19116
rect 5000 18550 5212 18578
rect 5078 18456 5134 18465
rect 5078 18391 5134 18400
rect 4724 18108 4844 18136
rect 4986 18184 5042 18193
rect 4986 18119 5042 18128
rect 4724 16969 4752 18108
rect 4894 18048 4950 18057
rect 4816 18006 4894 18034
rect 4710 16960 4766 16969
rect 4710 16895 4766 16904
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4724 16250 4752 16730
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4712 16244 4764 16250
rect 4712 16186 4764 16192
rect 4264 15570 4292 16186
rect 4436 16040 4488 16046
rect 4434 16008 4436 16017
rect 4528 16040 4580 16046
rect 4488 16008 4490 16017
rect 4528 15982 4580 15988
rect 4434 15943 4490 15952
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 4356 15366 4384 15506
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4193 15260 4501 15269
rect 4193 15258 4199 15260
rect 4255 15258 4279 15260
rect 4335 15258 4359 15260
rect 4415 15258 4439 15260
rect 4495 15258 4501 15260
rect 4255 15206 4257 15258
rect 4437 15206 4439 15258
rect 4193 15204 4199 15206
rect 4255 15204 4279 15206
rect 4335 15204 4359 15206
rect 4415 15204 4439 15206
rect 4495 15204 4501 15206
rect 4193 15195 4501 15204
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 3974 15056 4030 15065
rect 3974 14991 4030 15000
rect 4160 14952 4212 14958
rect 4080 14912 4160 14940
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 4080 14618 4108 14912
rect 4160 14894 4212 14900
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4264 14482 4292 15098
rect 4540 14618 4568 15982
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4620 14544 4672 14550
rect 4434 14512 4490 14521
rect 4252 14476 4304 14482
rect 4620 14486 4672 14492
rect 4434 14447 4436 14456
rect 4252 14418 4304 14424
rect 4488 14447 4490 14456
rect 4436 14418 4488 14424
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3332 13320 3384 13326
rect 3330 13288 3332 13297
rect 3384 13288 3386 13297
rect 3330 13223 3386 13232
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3344 12850 3372 13126
rect 3528 12986 3556 14214
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3514 12880 3570 12889
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3424 12844 3476 12850
rect 3514 12815 3570 12824
rect 3424 12786 3476 12792
rect 3344 12238 3372 12786
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 3344 11694 3372 12174
rect 3436 11744 3464 12786
rect 3528 12782 3556 12815
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3436 11716 3556 11744
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3238 11112 3294 11121
rect 3238 11047 3240 11056
rect 3292 11047 3294 11056
rect 3240 11018 3292 11024
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10674 3188 10950
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3238 10432 3294 10441
rect 3238 10367 3294 10376
rect 3146 10296 3202 10305
rect 3068 10254 3146 10282
rect 3252 10266 3280 10367
rect 3146 10231 3202 10240
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 3240 10056 3292 10062
rect 3344 10044 3372 11630
rect 3424 11620 3476 11626
rect 3424 11562 3476 11568
rect 3292 10016 3372 10044
rect 3240 9998 3292 10004
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 3068 9586 3096 9862
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3252 9518 3280 9998
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 9178 3004 9318
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2870 9072 2926 9081
rect 2870 9007 2926 9016
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2884 7342 2912 9007
rect 3252 8974 3280 9454
rect 3148 8968 3200 8974
rect 3146 8936 3148 8945
rect 3240 8968 3292 8974
rect 3200 8936 3202 8945
rect 3240 8910 3292 8916
rect 3146 8871 3202 8880
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2976 8430 3004 8570
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 2964 8424 3016 8430
rect 2964 8366 3016 8372
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2594 6760 2650 6769
rect 2594 6695 2650 6704
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2608 6322 2636 6695
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2594 5264 2650 5273
rect 2594 5199 2650 5208
rect 2608 1902 2636 5199
rect 2686 4992 2742 5001
rect 2686 4927 2742 4936
rect 2700 2802 2728 4927
rect 2792 4078 2820 6054
rect 2884 5914 2912 6598
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2884 5001 2912 5714
rect 2870 4992 2926 5001
rect 2870 4927 2926 4936
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2792 3670 2820 3878
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2976 3058 3004 7686
rect 3160 7177 3188 8434
rect 3344 7954 3372 8434
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3240 7200 3292 7206
rect 3146 7168 3202 7177
rect 3240 7142 3292 7148
rect 3146 7103 3202 7112
rect 3252 7002 3280 7142
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 3160 5234 3188 6190
rect 3252 6118 3280 6734
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3344 5710 3372 7890
rect 3436 7886 3464 11562
rect 3528 11529 3556 11716
rect 3514 11520 3570 11529
rect 3514 11455 3570 11464
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3528 5953 3556 10406
rect 3620 9518 3648 13942
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3712 11121 3740 11698
rect 3698 11112 3754 11121
rect 3698 11047 3754 11056
rect 3804 11014 3832 14214
rect 4080 14056 4108 14214
rect 4193 14172 4501 14181
rect 4193 14170 4199 14172
rect 4255 14170 4279 14172
rect 4335 14170 4359 14172
rect 4415 14170 4439 14172
rect 4495 14170 4501 14172
rect 4255 14118 4257 14170
rect 4437 14118 4439 14170
rect 4193 14116 4199 14118
rect 4255 14116 4279 14118
rect 4335 14116 4359 14118
rect 4415 14116 4439 14118
rect 4495 14116 4501 14118
rect 4193 14107 4501 14116
rect 4080 14028 4200 14056
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 3896 13190 3924 13806
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3988 13530 4016 13670
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3896 11762 3924 12922
rect 3988 12646 4016 13466
rect 4172 13240 4200 14028
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4080 13212 4200 13240
rect 4080 12968 4108 13212
rect 4264 13190 4292 13806
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4193 13084 4501 13093
rect 4193 13082 4199 13084
rect 4255 13082 4279 13084
rect 4335 13082 4359 13084
rect 4415 13082 4439 13084
rect 4495 13082 4501 13084
rect 4255 13030 4257 13082
rect 4437 13030 4439 13082
rect 4193 13028 4199 13030
rect 4255 13028 4279 13030
rect 4335 13028 4359 13030
rect 4415 13028 4439 13030
rect 4495 13028 4501 13030
rect 4193 13019 4501 13028
rect 4080 12940 4200 12968
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3988 12442 4016 12582
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3988 11558 4016 12378
rect 4172 12306 4200 12940
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4264 12753 4292 12786
rect 4250 12744 4306 12753
rect 4250 12679 4306 12688
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4193 11996 4501 12005
rect 4193 11994 4199 11996
rect 4255 11994 4279 11996
rect 4335 11994 4359 11996
rect 4415 11994 4439 11996
rect 4495 11994 4501 11996
rect 4255 11942 4257 11994
rect 4437 11942 4439 11994
rect 4193 11940 4199 11942
rect 4255 11940 4279 11942
rect 4335 11940 4359 11942
rect 4415 11940 4439 11942
rect 4495 11940 4501 11942
rect 4193 11931 4501 11940
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3884 11280 3936 11286
rect 3882 11248 3884 11257
rect 3936 11248 3938 11257
rect 3882 11183 3938 11192
rect 3988 11150 4016 11494
rect 4448 11286 4476 11834
rect 4540 11354 4568 13874
rect 4632 12782 4660 14486
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4620 11280 4672 11286
rect 4620 11222 4672 11228
rect 3976 11144 4028 11150
rect 4632 11132 4660 11222
rect 3976 11086 4028 11092
rect 4540 11104 4660 11132
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3700 10668 3752 10674
rect 3752 10628 3924 10656
rect 3700 10610 3752 10616
rect 3896 10266 3924 10628
rect 3988 10441 4016 11086
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10690 4108 10950
rect 4193 10908 4501 10917
rect 4193 10906 4199 10908
rect 4255 10906 4279 10908
rect 4335 10906 4359 10908
rect 4415 10906 4439 10908
rect 4495 10906 4501 10908
rect 4255 10854 4257 10906
rect 4437 10854 4439 10906
rect 4193 10852 4199 10854
rect 4255 10852 4279 10854
rect 4335 10852 4359 10854
rect 4415 10852 4439 10854
rect 4495 10852 4501 10854
rect 4193 10843 4501 10852
rect 4080 10662 4200 10690
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3974 10432 4030 10441
rect 3974 10367 4030 10376
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3712 9926 3740 9998
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3608 9512 3660 9518
rect 3608 9454 3660 9460
rect 3700 9376 3752 9382
rect 3896 9364 3924 9522
rect 3988 9382 4016 10367
rect 4080 10033 4108 10542
rect 4172 10062 4200 10662
rect 4540 10588 4568 11104
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4632 10810 4660 10950
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4620 10600 4672 10606
rect 4540 10560 4620 10588
rect 4620 10542 4672 10548
rect 4160 10056 4212 10062
rect 4066 10024 4122 10033
rect 4160 9998 4212 10004
rect 4066 9959 4122 9968
rect 4066 9888 4122 9897
rect 4066 9823 4122 9832
rect 3752 9336 3924 9364
rect 3976 9376 4028 9382
rect 3700 9318 3752 9324
rect 3976 9318 4028 9324
rect 3988 9178 4016 9318
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3974 8528 4030 8537
rect 3974 8463 3976 8472
rect 4028 8463 4030 8472
rect 3976 8434 4028 8440
rect 3608 8424 3660 8430
rect 4080 8378 4108 9823
rect 4193 9820 4501 9829
rect 4193 9818 4199 9820
rect 4255 9818 4279 9820
rect 4335 9818 4359 9820
rect 4415 9818 4439 9820
rect 4495 9818 4501 9820
rect 4255 9766 4257 9818
rect 4437 9766 4439 9818
rect 4193 9764 4199 9766
rect 4255 9764 4279 9766
rect 4335 9764 4359 9766
rect 4415 9764 4439 9766
rect 4495 9764 4501 9766
rect 4193 9755 4501 9764
rect 4724 9586 4752 15302
rect 4816 12628 4844 18006
rect 4894 17983 4950 17992
rect 4896 17740 4948 17746
rect 4896 17682 4948 17688
rect 4908 16794 4936 17682
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 4894 16688 4950 16697
rect 4894 16623 4950 16632
rect 4908 15366 4936 16623
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 5000 14498 5028 18119
rect 5092 15201 5120 18391
rect 5184 17796 5212 18550
rect 5276 17898 5304 19790
rect 5368 19310 5396 19790
rect 5356 19304 5408 19310
rect 5356 19246 5408 19252
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 5368 18601 5396 18770
rect 5354 18592 5410 18601
rect 5354 18527 5410 18536
rect 5354 18320 5410 18329
rect 5354 18255 5356 18264
rect 5408 18255 5410 18264
rect 5356 18226 5408 18232
rect 5276 17870 5396 17898
rect 5184 17768 5304 17796
rect 5368 17785 5396 17870
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5078 15192 5134 15201
rect 5078 15127 5134 15136
rect 5184 14793 5212 17614
rect 5276 17082 5304 17768
rect 5354 17776 5410 17785
rect 5354 17711 5410 17720
rect 5460 17202 5488 21286
rect 5828 21078 5856 21655
rect 8208 21626 8260 21632
rect 8220 21486 8248 21626
rect 5908 21480 5960 21486
rect 8208 21480 8260 21486
rect 6826 21448 6882 21457
rect 5908 21422 5960 21428
rect 5816 21072 5868 21078
rect 5816 21014 5868 21020
rect 5722 20904 5778 20913
rect 5722 20839 5778 20848
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5552 17218 5580 18702
rect 5644 18465 5672 19858
rect 5630 18456 5686 18465
rect 5736 18426 5764 20839
rect 5816 20800 5868 20806
rect 5814 20768 5816 20777
rect 5868 20768 5870 20777
rect 5814 20703 5870 20712
rect 5920 19854 5948 21422
rect 6196 21406 6826 21434
rect 6196 21350 6224 21406
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6276 21344 6328 21350
rect 6276 21286 6328 21292
rect 6182 21176 6238 21185
rect 6182 21111 6238 21120
rect 6196 21026 6224 21111
rect 6104 21010 6224 21026
rect 6000 21004 6052 21010
rect 6000 20946 6052 20952
rect 6092 21004 6224 21010
rect 6144 20998 6224 21004
rect 6092 20946 6144 20952
rect 6012 20097 6040 20946
rect 5998 20088 6054 20097
rect 5998 20023 6054 20032
rect 6000 19984 6052 19990
rect 5998 19952 6000 19961
rect 6052 19952 6054 19961
rect 6104 19938 6132 20946
rect 6184 20392 6236 20398
rect 6182 20360 6184 20369
rect 6236 20360 6238 20369
rect 6182 20295 6238 20304
rect 6184 20256 6236 20262
rect 6288 20210 6316 21286
rect 6236 20204 6316 20210
rect 6184 20198 6316 20204
rect 6196 20182 6316 20198
rect 6104 19910 6224 19938
rect 5998 19887 6054 19896
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6104 19514 6132 19790
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 6104 19378 6132 19450
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 6196 18714 6224 19910
rect 6288 19854 6316 20182
rect 6276 19848 6328 19854
rect 6276 19790 6328 19796
rect 6288 19174 6316 19790
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 6288 18970 6316 19110
rect 6276 18964 6328 18970
rect 6276 18906 6328 18912
rect 6380 18850 6408 21406
rect 8208 21422 8260 21428
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 6826 21383 6882 21392
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 6656 20466 6684 21286
rect 7194 21176 7250 21185
rect 7194 21111 7250 21120
rect 7208 21078 7236 21111
rect 7196 21072 7248 21078
rect 7196 21014 7248 21020
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 7286 20632 7342 20641
rect 7286 20567 7288 20576
rect 7340 20567 7342 20576
rect 7288 20538 7340 20544
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 6644 19848 6696 19854
rect 6840 19825 6868 20402
rect 6644 19790 6696 19796
rect 6826 19816 6882 19825
rect 6656 19417 6684 19790
rect 6826 19751 6882 19760
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 6642 19408 6698 19417
rect 6642 19343 6698 19352
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6288 18822 6592 18850
rect 6288 18766 6316 18822
rect 6012 18686 6224 18714
rect 6276 18760 6328 18766
rect 6276 18702 6328 18708
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 5630 18391 5686 18400
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5644 17814 5672 18226
rect 5632 17808 5684 17814
rect 5632 17750 5684 17756
rect 5448 17196 5500 17202
rect 5552 17190 5948 17218
rect 5448 17138 5500 17144
rect 5276 17054 5580 17082
rect 5262 16960 5318 16969
rect 5318 16918 5488 16946
rect 5262 16895 5318 16904
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 5170 14784 5226 14793
rect 5170 14719 5226 14728
rect 5080 14612 5132 14618
rect 5276 14600 5304 15914
rect 5354 15056 5410 15065
rect 5354 14991 5410 15000
rect 5132 14572 5304 14600
rect 5080 14554 5132 14560
rect 4908 14470 5028 14498
rect 5172 14476 5224 14482
rect 4908 13569 4936 14470
rect 5092 14436 5172 14464
rect 5092 13870 5120 14436
rect 5172 14418 5224 14424
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 4894 13560 4950 13569
rect 4894 13495 4950 13504
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4896 12640 4948 12646
rect 4816 12600 4896 12628
rect 4896 12582 4948 12588
rect 5092 12238 5120 13262
rect 5276 12753 5304 14418
rect 5368 13326 5396 14991
rect 5460 14482 5488 16918
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5446 13424 5502 13433
rect 5552 13410 5580 17054
rect 5632 17060 5684 17066
rect 5632 17002 5684 17008
rect 5816 17060 5868 17066
rect 5816 17002 5868 17008
rect 5644 15638 5672 17002
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 5632 15632 5684 15638
rect 5632 15574 5684 15580
rect 5736 14278 5764 16594
rect 5828 16590 5856 17002
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5814 15056 5870 15065
rect 5814 14991 5870 15000
rect 5828 14550 5856 14991
rect 5816 14544 5868 14550
rect 5816 14486 5868 14492
rect 5920 14278 5948 17190
rect 6012 16436 6040 18686
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 6104 18222 6132 18566
rect 6380 18426 6408 18702
rect 6368 18420 6420 18426
rect 6368 18362 6420 18368
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 6472 18306 6500 18362
rect 6288 18278 6500 18306
rect 6092 18216 6144 18222
rect 6144 18176 6224 18204
rect 6092 18158 6144 18164
rect 6196 18086 6224 18176
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6196 17678 6224 18022
rect 6288 17746 6316 18278
rect 6564 18170 6592 18822
rect 6472 18142 6592 18170
rect 6472 18086 6500 18142
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6550 18048 6606 18057
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6196 17134 6224 17614
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6196 16590 6224 16934
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 6012 16408 6224 16436
rect 6092 16040 6144 16046
rect 6092 15982 6144 15988
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 6012 15337 6040 15438
rect 6104 15434 6132 15982
rect 6092 15428 6144 15434
rect 6092 15370 6144 15376
rect 5998 15328 6054 15337
rect 5998 15263 6054 15272
rect 6104 14958 6132 15370
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 5724 14272 5776 14278
rect 5630 14240 5686 14249
rect 5724 14214 5776 14220
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5630 14175 5686 14184
rect 5644 13462 5672 14175
rect 5722 14104 5778 14113
rect 5828 14074 5856 14214
rect 5722 14039 5724 14048
rect 5776 14039 5778 14048
rect 5816 14068 5868 14074
rect 5724 14010 5776 14016
rect 5816 14010 5868 14016
rect 6104 13870 6132 14894
rect 6196 14657 6224 16408
rect 6288 15026 6316 16526
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6380 14770 6408 17682
rect 6472 17134 6500 18022
rect 6550 17983 6606 17992
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6458 16280 6514 16289
rect 6458 16215 6514 16224
rect 6472 16114 6500 16215
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6472 15638 6500 15846
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 6472 14822 6500 15574
rect 6288 14742 6408 14770
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6182 14648 6238 14657
rect 6182 14583 6238 14592
rect 6196 14482 6224 14583
rect 6184 14476 6236 14482
rect 6184 14418 6236 14424
rect 6288 14414 6316 14742
rect 6366 14512 6422 14521
rect 6366 14447 6422 14456
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6288 13462 6316 14350
rect 6380 14346 6408 14447
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6472 13938 6500 14758
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6564 13530 6592 17983
rect 6656 16590 6684 19246
rect 6736 18216 6788 18222
rect 6840 18193 6868 19654
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7392 18601 7420 19246
rect 7378 18592 7434 18601
rect 7378 18527 7434 18536
rect 6736 18158 6788 18164
rect 6826 18184 6882 18193
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6748 14521 6776 18158
rect 6826 18119 6882 18128
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6840 17678 6868 18022
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 6828 17128 6880 17134
rect 6826 17096 6828 17105
rect 6880 17096 6882 17105
rect 6826 17031 6882 17040
rect 7024 16794 7052 17614
rect 7208 17338 7236 17614
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6840 14618 6868 14894
rect 6932 14822 6960 16730
rect 7288 16448 7340 16454
rect 7484 16425 7512 20742
rect 7576 20262 7604 21354
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7564 20256 7616 20262
rect 7564 20198 7616 20204
rect 7668 19378 7696 20878
rect 7748 20800 7800 20806
rect 7748 20742 7800 20748
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7562 19272 7618 19281
rect 7562 19207 7618 19216
rect 7576 18698 7604 19207
rect 7656 18896 7708 18902
rect 7656 18838 7708 18844
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 7288 16390 7340 16396
rect 7470 16416 7526 16425
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7208 15065 7236 15438
rect 7194 15056 7250 15065
rect 7194 14991 7250 15000
rect 7300 14958 7328 16390
rect 7470 16351 7526 16360
rect 7668 15201 7696 18838
rect 7760 18834 7788 20742
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7746 17912 7802 17921
rect 7746 17847 7802 17856
rect 7760 17513 7788 17847
rect 7852 17649 7880 21286
rect 7988 21244 8296 21253
rect 7988 21242 7994 21244
rect 8050 21242 8074 21244
rect 8130 21242 8154 21244
rect 8210 21242 8234 21244
rect 8290 21242 8296 21244
rect 8050 21190 8052 21242
rect 8232 21190 8234 21242
rect 7988 21188 7994 21190
rect 8050 21188 8074 21190
rect 8130 21188 8154 21190
rect 8210 21188 8234 21190
rect 8290 21188 8296 21190
rect 7988 21179 8296 21188
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 7944 20602 7972 21082
rect 8022 21040 8078 21049
rect 8022 20975 8024 20984
rect 8076 20975 8078 20984
rect 8024 20946 8076 20952
rect 8300 20936 8352 20942
rect 8404 20890 8432 21422
rect 8484 21344 8536 21350
rect 8484 21286 8536 21292
rect 8574 21312 8630 21321
rect 8352 20884 8432 20890
rect 8300 20878 8432 20884
rect 8312 20862 8432 20878
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 8404 20369 8432 20862
rect 8496 20777 8524 21286
rect 8574 21247 8630 21256
rect 8588 21146 8616 21247
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8680 20942 8708 21422
rect 8772 21146 8800 21830
rect 8864 21729 8892 21830
rect 8850 21720 8906 21729
rect 8850 21655 8906 21664
rect 9140 21554 9168 22170
rect 9588 22092 9640 22098
rect 9588 22034 9640 22040
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 9496 21548 9548 21554
rect 9496 21490 9548 21496
rect 8760 21140 8812 21146
rect 8760 21082 8812 21088
rect 8668 20936 8720 20942
rect 8852 20936 8904 20942
rect 8668 20878 8720 20884
rect 8850 20904 8852 20913
rect 8904 20904 8906 20913
rect 8482 20768 8538 20777
rect 8482 20703 8538 20712
rect 8390 20360 8446 20369
rect 8390 20295 8392 20304
rect 8444 20295 8446 20304
rect 8392 20266 8444 20272
rect 7988 20156 8296 20165
rect 7988 20154 7994 20156
rect 8050 20154 8074 20156
rect 8130 20154 8154 20156
rect 8210 20154 8234 20156
rect 8290 20154 8296 20156
rect 8050 20102 8052 20154
rect 8232 20102 8234 20154
rect 7988 20100 7994 20102
rect 8050 20100 8074 20102
rect 8130 20100 8154 20102
rect 8210 20100 8234 20102
rect 8290 20100 8296 20102
rect 7988 20091 8296 20100
rect 8404 19922 8432 20266
rect 8482 20088 8538 20097
rect 8482 20023 8538 20032
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8312 19802 8340 19858
rect 8496 19802 8524 20023
rect 8312 19774 8524 19802
rect 8680 19802 8708 20878
rect 8850 20839 8906 20848
rect 8850 20632 8906 20641
rect 8956 20618 8984 21490
rect 9404 21480 9456 21486
rect 9404 21422 9456 21428
rect 8906 20590 8984 20618
rect 8850 20567 8906 20576
rect 9416 20482 9444 21422
rect 8852 20460 8904 20466
rect 8852 20402 8904 20408
rect 9140 20454 9444 20482
rect 8864 20210 8892 20402
rect 9140 20398 9168 20454
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 9312 20256 9364 20262
rect 8864 20182 9168 20210
rect 9312 20198 9364 20204
rect 8944 20052 8996 20058
rect 8772 20012 8944 20040
rect 8772 19802 8800 20012
rect 8944 19994 8996 20000
rect 8850 19952 8906 19961
rect 8906 19910 8984 19938
rect 8850 19887 8906 19896
rect 8680 19774 8892 19802
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8312 19514 8340 19654
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 7988 19068 8296 19077
rect 7988 19066 7994 19068
rect 8050 19066 8074 19068
rect 8130 19066 8154 19068
rect 8210 19066 8234 19068
rect 8290 19066 8296 19068
rect 8050 19014 8052 19066
rect 8232 19014 8234 19066
rect 7988 19012 7994 19014
rect 8050 19012 8074 19014
rect 8130 19012 8154 19014
rect 8210 19012 8234 19014
rect 8290 19012 8296 19014
rect 7988 19003 8296 19012
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8312 18714 8340 18770
rect 8404 18766 8432 19246
rect 8484 19236 8536 19242
rect 8484 19178 8536 19184
rect 8496 18766 8524 19178
rect 8588 18986 8616 19314
rect 8864 19258 8892 19774
rect 8956 19378 8984 19910
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8772 19230 9076 19258
rect 8772 19174 8800 19230
rect 9048 19174 9076 19230
rect 8760 19168 8812 19174
rect 8852 19168 8904 19174
rect 8760 19110 8812 19116
rect 8850 19136 8852 19145
rect 9036 19168 9088 19174
rect 8904 19136 8906 19145
rect 9036 19110 9088 19116
rect 8850 19071 8906 19080
rect 8588 18958 8800 18986
rect 8772 18902 8800 18958
rect 8760 18896 8812 18902
rect 8760 18838 8812 18844
rect 8128 18686 8340 18714
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8128 18601 8156 18686
rect 8208 18624 8260 18630
rect 8114 18592 8170 18601
rect 8298 18592 8354 18601
rect 8260 18572 8298 18578
rect 8208 18566 8298 18572
rect 8220 18550 8298 18566
rect 8114 18527 8170 18536
rect 8298 18527 8354 18536
rect 8404 18290 8432 18702
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 7988 17980 8296 17989
rect 7988 17978 7994 17980
rect 8050 17978 8074 17980
rect 8130 17978 8154 17980
rect 8210 17978 8234 17980
rect 8290 17978 8296 17980
rect 8050 17926 8052 17978
rect 8232 17926 8234 17978
rect 7988 17924 7994 17926
rect 8050 17924 8074 17926
rect 8130 17924 8154 17926
rect 8210 17924 8234 17926
rect 8290 17924 8296 17926
rect 7988 17915 8296 17924
rect 8404 17882 8432 18022
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8496 17746 8524 18090
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8588 17678 8616 18226
rect 8666 18048 8722 18057
rect 8666 17983 8722 17992
rect 8576 17672 8628 17678
rect 7838 17640 7894 17649
rect 8576 17614 8628 17620
rect 7838 17575 7894 17584
rect 7746 17504 7802 17513
rect 7746 17439 7802 17448
rect 8588 17270 8616 17614
rect 8392 17264 8444 17270
rect 8392 17206 8444 17212
rect 8576 17264 8628 17270
rect 8576 17206 8628 17212
rect 7988 16892 8296 16901
rect 7988 16890 7994 16892
rect 8050 16890 8074 16892
rect 8130 16890 8154 16892
rect 8210 16890 8234 16892
rect 8290 16890 8296 16892
rect 8050 16838 8052 16890
rect 8232 16838 8234 16890
rect 7988 16836 7994 16838
rect 8050 16836 8074 16838
rect 8130 16836 8154 16838
rect 8210 16836 8234 16838
rect 8290 16836 8296 16838
rect 7988 16827 8296 16836
rect 8404 16833 8432 17206
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8390 16824 8446 16833
rect 8390 16759 8446 16768
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 7988 15804 8296 15813
rect 7988 15802 7994 15804
rect 8050 15802 8074 15804
rect 8130 15802 8154 15804
rect 8210 15802 8234 15804
rect 8290 15802 8296 15804
rect 8050 15750 8052 15802
rect 8232 15750 8234 15802
rect 7988 15748 7994 15750
rect 8050 15748 8074 15750
rect 8130 15748 8154 15750
rect 8210 15748 8234 15750
rect 8290 15748 8296 15750
rect 7988 15739 8296 15748
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 7746 15328 7802 15337
rect 7746 15263 7802 15272
rect 7654 15192 7710 15201
rect 7654 15127 7710 15136
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 7102 14784 7158 14793
rect 7102 14719 7158 14728
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6734 14512 6790 14521
rect 6644 14476 6696 14482
rect 6734 14447 6790 14456
rect 6644 14418 6696 14424
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 5502 13382 5580 13410
rect 5632 13456 5684 13462
rect 5632 13398 5684 13404
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 5446 13359 5502 13368
rect 6656 13326 6684 14418
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5262 12744 5318 12753
rect 5262 12679 5318 12688
rect 5276 12442 5304 12679
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5368 11898 5396 12786
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4816 11354 4844 11630
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4193 8732 4501 8741
rect 4193 8730 4199 8732
rect 4255 8730 4279 8732
rect 4335 8730 4359 8732
rect 4415 8730 4439 8732
rect 4495 8730 4501 8732
rect 4255 8678 4257 8730
rect 4437 8678 4439 8730
rect 4193 8676 4199 8678
rect 4255 8676 4279 8678
rect 4335 8676 4359 8678
rect 4415 8676 4439 8678
rect 4495 8676 4501 8678
rect 4193 8667 4501 8676
rect 3608 8366 3660 8372
rect 3620 7886 3648 8366
rect 3896 8350 4108 8378
rect 3608 7880 3660 7886
rect 3660 7840 3832 7868
rect 3608 7822 3660 7828
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3514 5944 3570 5953
rect 3514 5879 3570 5888
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3344 5234 3372 5646
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3160 5098 3188 5170
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 3054 3768 3110 3777
rect 3054 3703 3110 3712
rect 3068 3194 3096 3703
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 2700 2774 2820 2802
rect 2596 1896 2648 1902
rect 2792 1884 2820 2774
rect 2596 1838 2648 1844
rect 2700 1856 2820 1884
rect 2240 1550 2452 1578
rect 2596 1556 2648 1562
rect 2044 1420 2096 1426
rect 2044 1362 2096 1368
rect 2240 1222 2268 1550
rect 2596 1498 2648 1504
rect 2320 1488 2372 1494
rect 2608 1442 2636 1498
rect 2372 1436 2636 1442
rect 2320 1430 2636 1436
rect 2332 1414 2636 1430
rect 2700 1222 2728 1856
rect 3056 1828 3108 1834
rect 3056 1770 3108 1776
rect 3068 1601 3096 1770
rect 3054 1592 3110 1601
rect 3160 1562 3188 5034
rect 3344 4690 3372 5170
rect 3528 4826 3556 5782
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3240 4616 3292 4622
rect 3238 4584 3240 4593
rect 3292 4584 3294 4593
rect 3238 4519 3294 4528
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3252 4282 3280 4422
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3344 4026 3372 4626
rect 3436 4486 3464 4626
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3620 4146 3648 6734
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3712 5302 3740 6054
rect 3804 5914 3832 7840
rect 3896 6254 3924 8350
rect 4066 7984 4122 7993
rect 4066 7919 4122 7928
rect 4080 7410 4108 7919
rect 4724 7834 4752 9318
rect 4816 7954 4844 10950
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4724 7806 4844 7834
rect 4193 7644 4501 7653
rect 4193 7642 4199 7644
rect 4255 7642 4279 7644
rect 4335 7642 4359 7644
rect 4415 7642 4439 7644
rect 4495 7642 4501 7644
rect 4255 7590 4257 7642
rect 4437 7590 4439 7642
rect 4193 7588 4199 7590
rect 4255 7588 4279 7590
rect 4335 7588 4359 7590
rect 4415 7588 4439 7590
rect 4495 7588 4501 7590
rect 4193 7579 4501 7588
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3700 5296 3752 5302
rect 3700 5238 3752 5244
rect 3804 5166 3832 5850
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3804 4826 3832 5102
rect 3792 4820 3844 4826
rect 3712 4780 3792 4808
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3252 3998 3372 4026
rect 3252 3534 3280 3998
rect 3332 3936 3384 3942
rect 3332 3878 3384 3884
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3252 3194 3280 3470
rect 3344 3194 3372 3878
rect 3608 3664 3660 3670
rect 3608 3606 3660 3612
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3252 2496 3280 3130
rect 3620 3126 3648 3606
rect 3712 3534 3740 4780
rect 3792 4762 3844 4768
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3712 3398 3740 3470
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3608 3120 3660 3126
rect 3608 3062 3660 3068
rect 3712 2990 3740 3334
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3804 2689 3832 4014
rect 3988 2774 4016 6734
rect 4724 6730 4752 7482
rect 4816 6934 4844 7806
rect 4908 7002 4936 11494
rect 5000 9674 5028 11834
rect 5644 11694 5672 12718
rect 5724 12436 5776 12442
rect 5724 12378 5776 12384
rect 5632 11688 5684 11694
rect 5446 11656 5502 11665
rect 5446 11591 5502 11600
rect 5552 11648 5632 11676
rect 5078 11384 5134 11393
rect 5078 11319 5134 11328
rect 5092 11286 5120 11319
rect 5080 11280 5132 11286
rect 5080 11222 5132 11228
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5000 9646 5120 9674
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 4193 6556 4501 6565
rect 4193 6554 4199 6556
rect 4255 6554 4279 6556
rect 4335 6554 4359 6556
rect 4415 6554 4439 6556
rect 4495 6554 4501 6556
rect 4255 6502 4257 6554
rect 4437 6502 4439 6554
rect 4193 6500 4199 6502
rect 4255 6500 4279 6502
rect 4335 6500 4359 6502
rect 4415 6500 4439 6502
rect 4495 6500 4501 6502
rect 4193 6491 4501 6500
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4080 5370 4108 5646
rect 4816 5545 4844 6870
rect 4802 5536 4858 5545
rect 4193 5468 4501 5477
rect 4802 5471 4858 5480
rect 4193 5466 4199 5468
rect 4255 5466 4279 5468
rect 4335 5466 4359 5468
rect 4415 5466 4439 5468
rect 4495 5466 4501 5468
rect 4255 5414 4257 5466
rect 4437 5414 4439 5466
rect 4193 5412 4199 5414
rect 4255 5412 4279 5414
rect 4335 5412 4359 5414
rect 4415 5412 4439 5414
rect 4495 5412 4501 5414
rect 4193 5403 4501 5412
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4068 4616 4120 4622
rect 4066 4584 4068 4593
rect 4120 4584 4122 4593
rect 4066 4519 4122 4528
rect 4193 4380 4501 4389
rect 4193 4378 4199 4380
rect 4255 4378 4279 4380
rect 4335 4378 4359 4380
rect 4415 4378 4439 4380
rect 4495 4378 4501 4380
rect 4255 4326 4257 4378
rect 4437 4326 4439 4378
rect 4193 4324 4199 4326
rect 4255 4324 4279 4326
rect 4335 4324 4359 4326
rect 4415 4324 4439 4326
rect 4495 4324 4501 4326
rect 4193 4315 4501 4324
rect 4526 4176 4582 4185
rect 4344 4140 4396 4146
rect 4526 4111 4528 4120
rect 4344 4082 4396 4088
rect 4580 4111 4582 4120
rect 4528 4082 4580 4088
rect 4158 3768 4214 3777
rect 4158 3703 4214 3712
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 3896 2746 4016 2774
rect 3790 2680 3846 2689
rect 3790 2615 3846 2624
rect 3252 2468 3372 2496
rect 3238 2408 3294 2417
rect 3238 2343 3294 2352
rect 3054 1527 3110 1536
rect 3148 1556 3200 1562
rect 3148 1498 3200 1504
rect 3252 1290 3280 2343
rect 3344 1494 3372 2468
rect 3424 2440 3476 2446
rect 3792 2440 3844 2446
rect 3476 2388 3648 2394
rect 3424 2382 3648 2388
rect 3792 2382 3844 2388
rect 3436 2366 3648 2382
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3528 1902 3556 2246
rect 3516 1896 3568 1902
rect 3516 1838 3568 1844
rect 3332 1488 3384 1494
rect 3332 1430 3384 1436
rect 3528 1358 3556 1838
rect 3516 1352 3568 1358
rect 3516 1294 3568 1300
rect 3240 1284 3292 1290
rect 3240 1226 3292 1232
rect 2228 1216 2280 1222
rect 2228 1158 2280 1164
rect 2688 1216 2740 1222
rect 2688 1158 2740 1164
rect 1676 876 1728 882
rect 1676 818 1728 824
rect 1688 678 1716 818
rect 3620 814 3648 2366
rect 3608 808 3660 814
rect 3608 750 3660 756
rect 1400 672 1452 678
rect 1400 614 1452 620
rect 1676 672 1728 678
rect 1676 614 1728 620
rect 3804 105 3832 2382
rect 3896 2106 3924 2746
rect 4080 2650 4108 3538
rect 4172 3534 4200 3703
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4356 3398 4384 4082
rect 4632 4026 4660 5102
rect 4632 3998 4752 4026
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4193 3292 4501 3301
rect 4193 3290 4199 3292
rect 4255 3290 4279 3292
rect 4335 3290 4359 3292
rect 4415 3290 4439 3292
rect 4495 3290 4501 3292
rect 4255 3238 4257 3290
rect 4437 3238 4439 3290
rect 4193 3236 4199 3238
rect 4255 3236 4279 3238
rect 4335 3236 4359 3238
rect 4415 3236 4439 3238
rect 4495 3236 4501 3238
rect 4193 3227 4501 3236
rect 4160 2848 4212 2854
rect 4158 2816 4160 2825
rect 4212 2816 4214 2825
rect 4158 2751 4214 2760
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 3976 2440 4028 2446
rect 3974 2408 3976 2417
rect 4068 2440 4120 2446
rect 4028 2408 4030 2417
rect 4068 2382 4120 2388
rect 3974 2343 4030 2352
rect 4080 2258 4108 2382
rect 3988 2230 4108 2258
rect 3988 2106 4016 2230
rect 4193 2204 4501 2213
rect 4193 2202 4199 2204
rect 4255 2202 4279 2204
rect 4335 2202 4359 2204
rect 4415 2202 4439 2204
rect 4495 2202 4501 2204
rect 4255 2150 4257 2202
rect 4437 2150 4439 2202
rect 4193 2148 4199 2150
rect 4255 2148 4279 2150
rect 4335 2148 4359 2150
rect 4415 2148 4439 2150
rect 4495 2148 4501 2150
rect 4193 2139 4501 2148
rect 3884 2100 3936 2106
rect 3884 2042 3936 2048
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 3884 1964 3936 1970
rect 3988 1952 4016 2042
rect 4540 2009 4568 3878
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4632 2650 4660 3334
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4526 2000 4582 2009
rect 3936 1924 4016 1952
rect 4068 1964 4120 1970
rect 3884 1906 3936 1912
rect 4526 1935 4582 1944
rect 4068 1906 4120 1912
rect 3896 1358 3924 1906
rect 3884 1352 3936 1358
rect 3884 1294 3936 1300
rect 3976 1352 4028 1358
rect 3976 1294 4028 1300
rect 3988 1222 4016 1294
rect 4080 1222 4108 1906
rect 4540 1465 4568 1935
rect 4724 1562 4752 3998
rect 4816 2774 4844 5471
rect 5000 4690 5028 9386
rect 5092 8106 5120 9646
rect 5184 8566 5212 10202
rect 5368 10198 5396 11154
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5460 9722 5488 11591
rect 5552 10674 5580 11648
rect 5632 11630 5684 11636
rect 5736 11354 5764 12378
rect 5920 11937 5948 13126
rect 6288 12866 6316 13126
rect 6104 12838 6316 12866
rect 6104 12442 6132 12838
rect 6184 12776 6236 12782
rect 6380 12764 6408 13194
rect 6236 12736 6408 12764
rect 6184 12718 6236 12724
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 6380 12306 6408 12736
rect 6458 12472 6514 12481
rect 6514 12416 6592 12434
rect 6458 12407 6592 12416
rect 6472 12406 6592 12407
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 5906 11928 5962 11937
rect 5906 11863 5962 11872
rect 6012 11778 6040 12038
rect 6104 11898 6132 12038
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6012 11762 6132 11778
rect 5908 11756 5960 11762
rect 6012 11756 6144 11762
rect 6012 11750 6092 11756
rect 5908 11698 5960 11704
rect 6092 11698 6144 11704
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5828 11558 5856 11630
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5448 9716 5500 9722
rect 5448 9658 5500 9664
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5276 9489 5304 9522
rect 5262 9480 5318 9489
rect 5262 9415 5318 9424
rect 5264 9104 5316 9110
rect 5262 9072 5264 9081
rect 5316 9072 5318 9081
rect 5262 9007 5318 9016
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5276 8498 5304 8842
rect 5356 8832 5408 8838
rect 5448 8832 5500 8838
rect 5356 8774 5408 8780
rect 5446 8800 5448 8809
rect 5500 8800 5502 8809
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5092 8090 5212 8106
rect 5092 8084 5224 8090
rect 5092 8078 5172 8084
rect 5172 8026 5224 8032
rect 5368 8022 5396 8774
rect 5446 8735 5502 8744
rect 5552 8498 5580 10610
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5644 9697 5672 10406
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5630 9688 5686 9697
rect 5630 9623 5686 9632
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5460 8090 5488 8298
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 6458 5120 6598
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5092 5234 5120 6054
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4816 2746 5028 2774
rect 5000 1834 5028 2746
rect 5078 2680 5134 2689
rect 5078 2615 5134 2624
rect 4988 1828 5040 1834
rect 4988 1770 5040 1776
rect 4712 1556 4764 1562
rect 4712 1498 4764 1504
rect 4526 1456 4582 1465
rect 4526 1391 4582 1400
rect 4252 1352 4304 1358
rect 4250 1320 4252 1329
rect 4304 1320 4306 1329
rect 4250 1255 4306 1264
rect 3976 1216 4028 1222
rect 3976 1158 4028 1164
rect 4068 1216 4120 1222
rect 4068 1158 4120 1164
rect 3988 474 4016 1158
rect 4193 1116 4501 1125
rect 4193 1114 4199 1116
rect 4255 1114 4279 1116
rect 4335 1114 4359 1116
rect 4415 1114 4439 1116
rect 4495 1114 4501 1116
rect 4255 1062 4257 1114
rect 4437 1062 4439 1114
rect 4193 1060 4199 1062
rect 4255 1060 4279 1062
rect 4335 1060 4359 1062
rect 4415 1060 4439 1062
rect 4495 1060 4501 1062
rect 4193 1051 4501 1060
rect 4988 808 5040 814
rect 4986 776 4988 785
rect 5040 776 5042 785
rect 4986 711 5042 720
rect 3976 468 4028 474
rect 3976 410 4028 416
rect 5092 202 5120 2615
rect 5184 950 5212 7686
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5368 6866 5396 7414
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5262 6216 5318 6225
rect 5262 6151 5318 6160
rect 5276 3058 5304 6151
rect 5368 5846 5396 6394
rect 5356 5840 5408 5846
rect 5356 5782 5408 5788
rect 5460 5778 5488 6598
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5552 5658 5580 5850
rect 5460 5642 5580 5658
rect 5448 5636 5580 5642
rect 5500 5630 5580 5636
rect 5448 5578 5500 5584
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5446 4584 5502 4593
rect 5446 4519 5502 4528
rect 5354 4040 5410 4049
rect 5354 3975 5410 3984
rect 5368 3602 5396 3975
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 5368 1562 5396 2246
rect 5460 1970 5488 4519
rect 5552 4146 5580 5510
rect 5644 5234 5672 9318
rect 5736 8498 5764 9998
rect 5828 9722 5856 10610
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5814 9480 5870 9489
rect 5814 9415 5870 9424
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5722 8392 5778 8401
rect 5722 8327 5778 8336
rect 5736 8090 5764 8327
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5736 6730 5764 7278
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5736 6322 5764 6666
rect 5828 6662 5856 9415
rect 5920 9110 5948 11698
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 6182 11520 6238 11529
rect 6012 11150 6040 11494
rect 6182 11455 6238 11464
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6012 10470 6040 11086
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 6012 10062 6040 10406
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 6012 8294 6040 9998
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 5906 8120 5962 8129
rect 5906 8055 5962 8064
rect 5920 7954 5948 8055
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5920 7410 5948 7754
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6012 7290 6040 7890
rect 5920 7262 6040 7290
rect 5920 6905 5948 7262
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 5906 6896 5962 6905
rect 5906 6831 5962 6840
rect 6012 6798 6040 7142
rect 6000 6792 6052 6798
rect 5920 6752 6000 6780
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5920 6322 5948 6752
rect 6000 6734 6052 6740
rect 6104 6610 6132 10542
rect 6196 9042 6224 11455
rect 6380 11218 6408 12242
rect 6564 11370 6592 12406
rect 6748 12102 6776 14282
rect 6840 13394 6868 14350
rect 7010 14104 7066 14113
rect 6920 14068 6972 14074
rect 7010 14039 7012 14048
rect 6920 14010 6972 14016
rect 7064 14039 7066 14048
rect 7012 14010 7064 14016
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6840 12238 6868 12378
rect 6932 12238 6960 14010
rect 7116 13297 7144 14719
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7208 13326 7236 14350
rect 7300 14249 7328 14350
rect 7286 14240 7342 14249
rect 7286 14175 7342 14184
rect 7196 13320 7248 13326
rect 7102 13288 7158 13297
rect 7196 13262 7248 13268
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7102 13223 7158 13232
rect 7208 12782 7236 13262
rect 7300 12986 7328 13262
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7208 12442 7236 12718
rect 7484 12646 7512 13126
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7378 12472 7434 12481
rect 7196 12436 7248 12442
rect 7472 12436 7524 12442
rect 7434 12416 7472 12434
rect 7378 12407 7472 12416
rect 7392 12406 7472 12407
rect 7196 12378 7248 12384
rect 7472 12378 7524 12384
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6564 11342 6684 11370
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6012 6582 6132 6610
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5722 5944 5778 5953
rect 5778 5902 5856 5930
rect 5722 5879 5778 5888
rect 5828 5710 5856 5902
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5828 4622 5856 5646
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5448 1964 5500 1970
rect 5448 1906 5500 1912
rect 5356 1556 5408 1562
rect 5356 1498 5408 1504
rect 5644 1193 5672 4490
rect 5828 4078 5856 4558
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5828 3466 5856 4014
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5828 3058 5856 3402
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5828 2446 5856 2994
rect 5920 2961 5948 3946
rect 5906 2952 5962 2961
rect 5906 2887 5962 2896
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5828 1494 5856 2382
rect 6012 1902 6040 6582
rect 6090 6352 6146 6361
rect 6196 6322 6224 8774
rect 6288 8401 6316 10542
rect 6380 10169 6408 11018
rect 6366 10160 6422 10169
rect 6366 10095 6422 10104
rect 6472 9382 6500 11154
rect 6656 10282 6684 11342
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6748 10674 6776 11154
rect 6840 11132 6868 12174
rect 7576 11898 7604 14350
rect 7760 14074 7788 15263
rect 7944 15094 7972 15574
rect 8404 15570 8432 15846
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8312 15162 8340 15302
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 7932 15088 7984 15094
rect 7932 15030 7984 15036
rect 8496 14958 8524 17070
rect 8576 16788 8628 16794
rect 8680 16776 8708 17983
rect 8772 17814 8800 18226
rect 8864 18086 8892 19071
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 8852 18080 8904 18086
rect 8852 18022 8904 18028
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8864 17678 8892 18022
rect 8852 17672 8904 17678
rect 8852 17614 8904 17620
rect 8956 17490 8984 18770
rect 9036 18760 9088 18766
rect 9140 18748 9168 20182
rect 9218 20088 9274 20097
rect 9218 20023 9220 20032
rect 9272 20023 9274 20032
rect 9220 19994 9272 20000
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9232 18850 9260 19790
rect 9324 18970 9352 20198
rect 9508 19553 9536 21490
rect 9494 19544 9550 19553
rect 9494 19479 9550 19488
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 9232 18822 9352 18850
rect 9088 18720 9168 18748
rect 9036 18702 9088 18708
rect 9140 18290 9168 18720
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 8628 16748 8708 16776
rect 8772 17462 8984 17490
rect 8576 16730 8628 16736
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 8680 16046 8708 16594
rect 8668 16040 8720 16046
rect 8668 15982 8720 15988
rect 8680 15366 8708 15982
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8574 15056 8630 15065
rect 8574 14991 8630 15000
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 7988 14716 8296 14725
rect 7988 14714 7994 14716
rect 8050 14714 8074 14716
rect 8130 14714 8154 14716
rect 8210 14714 8234 14716
rect 8290 14714 8296 14716
rect 8050 14662 8052 14714
rect 8232 14662 8234 14714
rect 7988 14660 7994 14662
rect 8050 14660 8074 14662
rect 8130 14660 8154 14662
rect 8210 14660 8234 14662
rect 8290 14660 8296 14662
rect 7988 14651 8296 14660
rect 8496 14482 8524 14894
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7988 13628 8296 13637
rect 7988 13626 7994 13628
rect 8050 13626 8074 13628
rect 8130 13626 8154 13628
rect 8210 13626 8234 13628
rect 8290 13626 8296 13628
rect 8050 13574 8052 13626
rect 8232 13574 8234 13626
rect 7988 13572 7994 13574
rect 8050 13572 8074 13574
rect 8130 13572 8154 13574
rect 8210 13572 8234 13574
rect 8290 13572 8296 13574
rect 7654 13560 7710 13569
rect 7988 13563 8296 13572
rect 7654 13495 7710 13504
rect 7668 12986 7696 13495
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 8496 12714 8524 14418
rect 8588 14414 8616 14991
rect 8680 14958 8708 15302
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8772 14482 8800 17462
rect 9048 16998 9076 17614
rect 9232 17542 9260 17614
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9324 17354 9352 18822
rect 9402 17640 9458 17649
rect 9402 17575 9458 17584
rect 9140 17326 9352 17354
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8850 16280 8906 16289
rect 8850 16215 8906 16224
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8772 13530 8800 14214
rect 8864 14006 8892 16215
rect 8956 16130 8984 16526
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 9048 16289 9076 16390
rect 9034 16280 9090 16289
rect 9034 16215 9090 16224
rect 8956 16102 9076 16130
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 8956 14074 8984 15982
rect 9048 15910 9076 16102
rect 9036 15904 9088 15910
rect 9036 15846 9088 15852
rect 9048 15502 9076 15846
rect 9036 15496 9088 15502
rect 9140 15473 9168 17326
rect 9218 17232 9274 17241
rect 9416 17202 9444 17575
rect 9218 17167 9274 17176
rect 9404 17196 9456 17202
rect 9232 15502 9260 17167
rect 9404 17138 9456 17144
rect 9310 16824 9366 16833
rect 9366 16782 9444 16810
rect 9310 16759 9366 16768
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9220 15496 9272 15502
rect 9036 15438 9088 15444
rect 9126 15464 9182 15473
rect 9048 15026 9076 15438
rect 9220 15438 9272 15444
rect 9126 15399 9182 15408
rect 9218 15056 9274 15065
rect 9036 15020 9088 15026
rect 9218 14991 9220 15000
rect 9036 14962 9088 14968
rect 9272 14991 9274 15000
rect 9220 14962 9272 14968
rect 9048 14618 9076 14962
rect 9218 14920 9274 14929
rect 9218 14855 9274 14864
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 9232 14074 9260 14855
rect 9324 14074 9352 16594
rect 9416 14958 9444 16782
rect 9508 16538 9536 19314
rect 9600 19310 9628 22034
rect 9680 21004 9732 21010
rect 9680 20946 9732 20952
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 9692 18601 9720 20946
rect 9784 19961 9812 22170
rect 12636 22114 12664 22222
rect 12900 22170 12952 22176
rect 18512 22228 18564 22234
rect 18512 22170 18564 22176
rect 12452 22098 12664 22114
rect 12808 22160 12860 22166
rect 12808 22102 12860 22108
rect 12440 22092 12664 22098
rect 12492 22086 12664 22092
rect 12440 22034 12492 22040
rect 12624 22024 12676 22030
rect 10322 21992 10378 22001
rect 12438 21992 12494 22001
rect 10378 21950 10456 21978
rect 10322 21927 10378 21936
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 9770 19952 9826 19961
rect 9770 19887 9826 19896
rect 9772 18624 9824 18630
rect 9678 18592 9734 18601
rect 9772 18566 9824 18572
rect 9678 18527 9734 18536
rect 9678 18456 9734 18465
rect 9678 18391 9734 18400
rect 9692 17134 9720 18391
rect 9784 17649 9812 18566
rect 9862 17776 9918 17785
rect 9918 17734 9996 17762
rect 9862 17711 9918 17720
rect 9770 17640 9826 17649
rect 9770 17575 9826 17584
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9772 16584 9824 16590
rect 9508 16510 9628 16538
rect 9772 16526 9824 16532
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9508 15609 9536 16390
rect 9494 15600 9550 15609
rect 9494 15535 9550 15544
rect 9496 15496 9548 15502
rect 9496 15438 9548 15444
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 8852 14000 8904 14006
rect 9508 13954 9536 15438
rect 8852 13942 8904 13948
rect 9416 13926 9536 13954
rect 9416 13870 9444 13926
rect 8944 13864 8996 13870
rect 9404 13864 9456 13870
rect 8996 13824 9404 13852
rect 8944 13806 8996 13812
rect 9600 13818 9628 16510
rect 9784 16250 9812 16526
rect 9862 16280 9918 16289
rect 9772 16244 9824 16250
rect 9862 16215 9918 16224
rect 9772 16186 9824 16192
rect 9784 14482 9812 16186
rect 9876 16046 9904 16215
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9692 14113 9720 14282
rect 9678 14104 9734 14113
rect 9678 14039 9734 14048
rect 9404 13806 9456 13812
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 7988 12540 8296 12549
rect 7988 12538 7994 12540
rect 8050 12538 8074 12540
rect 8130 12538 8154 12540
rect 8210 12538 8234 12540
rect 8290 12538 8296 12540
rect 8050 12486 8052 12538
rect 8232 12486 8234 12538
rect 7988 12484 7994 12486
rect 8050 12484 8074 12486
rect 8130 12484 8154 12486
rect 8210 12484 8234 12486
rect 8290 12484 8296 12486
rect 7988 12475 8296 12484
rect 8588 12442 8616 12582
rect 8772 12442 8800 12718
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7380 11824 7432 11830
rect 7380 11766 7432 11772
rect 7012 11552 7064 11558
rect 7392 11529 7420 11766
rect 7944 11694 7972 12378
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11694 8248 12038
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8680 11676 8708 12174
rect 8864 11762 8892 13126
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8760 11688 8812 11694
rect 8680 11648 8760 11676
rect 7748 11552 7800 11558
rect 7012 11494 7064 11500
rect 7378 11520 7434 11529
rect 6920 11144 6972 11150
rect 6840 11104 6920 11132
rect 6920 11086 6972 11092
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6656 10254 6776 10282
rect 6932 10266 6960 10542
rect 6552 10192 6604 10198
rect 6604 10152 6684 10180
rect 6552 10134 6604 10140
rect 6550 9888 6606 9897
rect 6550 9823 6606 9832
rect 6564 9586 6592 9823
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6472 9042 6500 9318
rect 6656 9058 6684 10152
rect 6748 9518 6776 10254
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6748 9178 6776 9454
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6840 9058 6868 9998
rect 6932 9382 6960 10202
rect 7024 9897 7052 11494
rect 7748 11494 7800 11500
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 7378 11455 7434 11464
rect 7760 11218 7788 11494
rect 7988 11452 8296 11461
rect 7988 11450 7994 11452
rect 8050 11450 8074 11452
rect 8130 11450 8154 11452
rect 8210 11450 8234 11452
rect 8290 11450 8296 11452
rect 8050 11398 8052 11450
rect 8232 11398 8234 11450
rect 7988 11396 7994 11398
rect 8050 11396 8074 11398
rect 8130 11396 8154 11398
rect 8210 11396 8234 11398
rect 8290 11396 8296 11398
rect 7988 11387 8296 11396
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 7392 10146 7420 10474
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7300 10130 7420 10146
rect 7288 10124 7420 10130
rect 7340 10118 7420 10124
rect 7288 10066 7340 10072
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7010 9888 7066 9897
rect 7010 9823 7066 9832
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6656 9042 6776 9058
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6460 9036 6512 9042
rect 6656 9036 6788 9042
rect 6656 9030 6736 9036
rect 6460 8978 6512 8984
rect 6840 9030 7052 9058
rect 6736 8978 6788 8984
rect 6380 8498 6408 8978
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6274 8392 6330 8401
rect 6274 8327 6330 8336
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6380 7886 6408 8230
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6288 7002 6316 7346
rect 6380 7206 6408 7822
rect 6472 7546 6500 8774
rect 6748 8106 6776 8978
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6656 8078 6776 8106
rect 6550 7984 6606 7993
rect 6550 7919 6606 7928
rect 6564 7750 6592 7919
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6090 6287 6092 6296
rect 6144 6287 6146 6296
rect 6184 6316 6236 6322
rect 6092 6258 6144 6264
rect 6184 6258 6236 6264
rect 6288 5794 6316 6598
rect 6196 5766 6316 5794
rect 6196 5710 6224 5766
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6276 5704 6328 5710
rect 6380 5681 6408 6734
rect 6472 5914 6500 7278
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6460 5704 6512 5710
rect 6276 5646 6328 5652
rect 6366 5672 6422 5681
rect 6196 4622 6224 5646
rect 6288 5370 6316 5646
rect 6460 5646 6512 5652
rect 6366 5607 6422 5616
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6196 3924 6224 4558
rect 6276 3936 6328 3942
rect 6196 3896 6276 3924
rect 6196 2922 6224 3896
rect 6276 3878 6328 3884
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6184 2916 6236 2922
rect 6184 2858 6236 2864
rect 6196 2650 6224 2858
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6288 2446 6316 3470
rect 6380 3398 6408 5306
rect 6472 5030 6500 5646
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6472 3602 6500 4966
rect 6564 4282 6592 6734
rect 6656 5370 6684 8078
rect 6734 7984 6790 7993
rect 6734 7919 6790 7928
rect 6748 7886 6776 7919
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6840 7342 6868 8910
rect 6932 8294 6960 8910
rect 7024 8498 7052 9030
rect 7116 8634 7144 9998
rect 7392 9738 7420 10118
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7300 9722 7420 9738
rect 7288 9716 7420 9722
rect 7340 9710 7420 9716
rect 7288 9658 7340 9664
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 7104 8424 7156 8430
rect 7024 8372 7104 8378
rect 7024 8366 7156 8372
rect 7024 8350 7144 8366
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6918 8120 6974 8129
rect 7024 8106 7052 8350
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 6974 8078 7052 8106
rect 6918 8055 6974 8064
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6932 7546 6960 7822
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6920 5160 6972 5166
rect 6656 5108 6920 5114
rect 6656 5102 6972 5108
rect 6656 5086 6960 5102
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 6368 3392 6420 3398
rect 6368 3334 6420 3340
rect 6380 3194 6408 3334
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6472 2990 6500 3538
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 6472 1970 6500 2926
rect 6656 2774 6684 5086
rect 7116 5030 7144 8230
rect 7208 7478 7236 9114
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7300 8362 7328 8978
rect 7392 8974 7420 9710
rect 7470 9072 7526 9081
rect 7470 9007 7472 9016
rect 7524 9007 7526 9016
rect 7472 8978 7524 8984
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7484 8072 7512 8978
rect 7576 8634 7604 9998
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7668 8430 7696 10406
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7760 8974 7788 9318
rect 7852 9058 7880 10610
rect 8220 10538 8248 11290
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 7988 10364 8296 10373
rect 7988 10362 7994 10364
rect 8050 10362 8074 10364
rect 8130 10362 8154 10364
rect 8210 10362 8234 10364
rect 8290 10362 8296 10364
rect 8050 10310 8052 10362
rect 8232 10310 8234 10362
rect 7988 10308 7994 10310
rect 8050 10308 8074 10310
rect 8130 10308 8154 10310
rect 8210 10308 8234 10310
rect 8290 10308 8296 10310
rect 7988 10299 8296 10308
rect 8404 9586 8432 11494
rect 8588 11218 8616 11630
rect 8680 11354 8708 11648
rect 8760 11630 8812 11636
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 11393 8892 11494
rect 8850 11384 8906 11393
rect 8668 11348 8720 11354
rect 8850 11319 8906 11328
rect 8668 11290 8720 11296
rect 8956 11218 8984 13806
rect 9416 13530 9444 13806
rect 9508 13790 9628 13818
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9324 13190 9352 13398
rect 9508 13190 9536 13790
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9324 12782 9352 12922
rect 9128 12776 9180 12782
rect 9126 12744 9128 12753
rect 9312 12776 9364 12782
rect 9180 12744 9182 12753
rect 9312 12718 9364 12724
rect 9126 12679 9182 12688
rect 9600 12646 9628 13670
rect 9692 12782 9720 13806
rect 9784 13326 9812 14418
rect 9876 14385 9904 14554
rect 9862 14376 9918 14385
rect 9862 14311 9918 14320
rect 9968 13954 9996 17734
rect 10060 16726 10088 21286
rect 10322 20632 10378 20641
rect 10322 20567 10324 20576
rect 10376 20567 10378 20576
rect 10324 20538 10376 20544
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10244 19514 10272 20402
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10244 18154 10272 19178
rect 10322 19000 10378 19009
rect 10322 18935 10378 18944
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10048 16720 10100 16726
rect 10048 16662 10100 16668
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 9876 13926 9996 13954
rect 9876 13530 9904 13926
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9864 13388 9916 13394
rect 9968 13376 9996 13806
rect 9916 13348 9996 13376
rect 9864 13330 9916 13336
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9048 12238 9076 12582
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 9048 11558 9076 12174
rect 9126 11928 9182 11937
rect 9126 11863 9182 11872
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8588 10554 8616 11154
rect 9140 11014 9168 11863
rect 9692 11608 9720 12718
rect 9600 11580 9720 11608
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 8944 10600 8996 10606
rect 8588 10526 8708 10554
rect 8944 10542 8996 10548
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8496 9722 8524 9862
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8588 9586 8616 9862
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 7988 9276 8296 9285
rect 7988 9274 7994 9276
rect 8050 9274 8074 9276
rect 8130 9274 8154 9276
rect 8210 9274 8234 9276
rect 8290 9274 8296 9276
rect 8050 9222 8052 9274
rect 8232 9222 8234 9274
rect 7988 9220 7994 9222
rect 8050 9220 8074 9222
rect 8130 9220 8154 9222
rect 8210 9220 8234 9222
rect 8290 9220 8296 9222
rect 7988 9211 8296 9220
rect 7852 9030 8064 9058
rect 8036 8974 8064 9030
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8220 8430 8248 8910
rect 8680 8430 8708 10526
rect 8956 10266 8984 10542
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 8760 9716 8812 9722
rect 8812 9664 8892 9674
rect 8760 9658 8892 9664
rect 8772 9646 8892 9658
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 7300 8044 7512 8072
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 7194 6896 7250 6905
rect 7300 6882 7328 8044
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7378 7032 7434 7041
rect 7378 6967 7434 6976
rect 7250 6854 7328 6882
rect 7194 6831 7250 6840
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6748 3738 6776 4014
rect 6840 3738 6868 4966
rect 7208 4690 7236 6831
rect 7392 6390 7420 6967
rect 7380 6384 7432 6390
rect 7380 6326 7432 6332
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7208 3913 7236 4626
rect 7484 4078 7512 7414
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7654 7168 7710 7177
rect 7576 6798 7604 7142
rect 7654 7103 7710 7112
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7668 6662 7696 7103
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7852 5896 7880 8298
rect 7988 8188 8296 8197
rect 7988 8186 7994 8188
rect 8050 8186 8074 8188
rect 8130 8186 8154 8188
rect 8210 8186 8234 8188
rect 8290 8186 8296 8188
rect 8050 8134 8052 8186
rect 8232 8134 8234 8186
rect 7988 8132 7994 8134
rect 8050 8132 8074 8134
rect 8130 8132 8154 8134
rect 8210 8132 8234 8134
rect 8290 8132 8296 8134
rect 7988 8123 8296 8132
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8114 7576 8170 7585
rect 8114 7511 8170 7520
rect 8128 7342 8156 7511
rect 8404 7410 8432 7890
rect 8680 7721 8708 8366
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8666 7712 8722 7721
rect 8666 7647 8722 7656
rect 8392 7404 8444 7410
rect 8444 7364 8524 7392
rect 8392 7346 8444 7352
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 7988 7100 8296 7109
rect 7988 7098 7994 7100
rect 8050 7098 8074 7100
rect 8130 7098 8154 7100
rect 8210 7098 8234 7100
rect 8290 7098 8296 7100
rect 8050 7046 8052 7098
rect 8232 7046 8234 7098
rect 7988 7044 7994 7046
rect 8050 7044 8074 7046
rect 8130 7044 8154 7046
rect 8210 7044 8234 7046
rect 8290 7044 8296 7046
rect 7988 7035 8296 7044
rect 8404 6934 8432 7142
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 8496 6866 8524 7364
rect 8772 7342 8800 7822
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8392 6384 8444 6390
rect 8496 6372 8524 6802
rect 8772 6798 8800 7278
rect 8760 6792 8812 6798
rect 8760 6734 8812 6740
rect 8864 6440 8892 9646
rect 9048 9382 9076 9998
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 8956 8634 8984 9318
rect 9140 9081 9168 10950
rect 9416 10538 9444 11494
rect 9600 11354 9628 11580
rect 9784 11506 9812 13262
rect 9876 12753 9904 13330
rect 10060 13308 10088 16458
rect 10152 15366 10180 17682
rect 10244 16697 10272 18090
rect 10230 16688 10286 16697
rect 10230 16623 10286 16632
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 10336 14958 10364 18935
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10322 14648 10378 14657
rect 10322 14583 10378 14592
rect 10336 14550 10364 14583
rect 10324 14544 10376 14550
rect 10324 14486 10376 14492
rect 10138 14104 10194 14113
rect 10138 14039 10194 14048
rect 10152 13938 10180 14039
rect 10428 13954 10456 21950
rect 12624 21966 12676 21972
rect 12438 21927 12494 21936
rect 11783 21788 12091 21797
rect 11783 21786 11789 21788
rect 11845 21786 11869 21788
rect 11925 21786 11949 21788
rect 12005 21786 12029 21788
rect 12085 21786 12091 21788
rect 11845 21734 11847 21786
rect 12027 21734 12029 21786
rect 11783 21732 11789 21734
rect 11845 21732 11869 21734
rect 11925 21732 11949 21734
rect 12005 21732 12029 21734
rect 12085 21732 12091 21734
rect 11783 21723 12091 21732
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 10968 21480 11020 21486
rect 11060 21480 11112 21486
rect 10968 21422 11020 21428
rect 11058 21448 11060 21457
rect 11612 21480 11664 21486
rect 11112 21448 11114 21457
rect 10600 21344 10652 21350
rect 10600 21286 10652 21292
rect 10612 21146 10640 21286
rect 10600 21140 10652 21146
rect 10704 21128 10732 21422
rect 10888 21321 10916 21422
rect 10874 21312 10930 21321
rect 10874 21247 10930 21256
rect 10704 21100 10916 21128
rect 10600 21082 10652 21088
rect 10784 21004 10836 21010
rect 10784 20946 10836 20952
rect 10508 20936 10560 20942
rect 10796 20913 10824 20946
rect 10888 20924 10916 21100
rect 10980 21078 11008 21422
rect 11612 21422 11664 21428
rect 11058 21383 11114 21392
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 10968 21072 11020 21078
rect 10968 21014 11020 21020
rect 11060 21072 11112 21078
rect 11060 21014 11112 21020
rect 11072 20924 11100 21014
rect 10782 20904 10838 20913
rect 10508 20878 10560 20884
rect 10520 20602 10548 20878
rect 10704 20862 10782 20890
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 10508 18828 10560 18834
rect 10508 18770 10560 18776
rect 10520 17338 10548 18770
rect 10612 18204 10640 20198
rect 10704 18426 10732 20862
rect 10782 20839 10838 20848
rect 10888 20896 11100 20924
rect 10888 20369 10916 20896
rect 11244 20868 11296 20874
rect 11244 20810 11296 20816
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 10980 20466 11008 20742
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 10874 20360 10930 20369
rect 11072 20346 11100 20402
rect 10874 20295 10930 20304
rect 10980 20318 11100 20346
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10796 18698 10824 19654
rect 10876 19236 10928 19242
rect 10876 19178 10928 19184
rect 10888 19009 10916 19178
rect 10874 19000 10930 19009
rect 10874 18935 10930 18944
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10784 18692 10836 18698
rect 10784 18634 10836 18640
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10784 18216 10836 18222
rect 10612 18176 10784 18204
rect 10784 18158 10836 18164
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10506 16008 10562 16017
rect 10506 15943 10562 15952
rect 10520 15910 10548 15943
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10612 14482 10640 17070
rect 10690 16416 10746 16425
rect 10690 16351 10746 16360
rect 10704 16017 10732 16351
rect 10690 16008 10746 16017
rect 10690 15943 10746 15952
rect 10796 14618 10824 18158
rect 10888 17338 10916 18702
rect 10980 17746 11008 20318
rect 11164 20058 11192 20742
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11058 19680 11114 19689
rect 11114 19638 11192 19666
rect 11058 19615 11114 19624
rect 11060 19304 11112 19310
rect 11058 19272 11060 19281
rect 11112 19272 11114 19281
rect 11058 19207 11114 19216
rect 11164 18834 11192 19638
rect 11256 19514 11284 20810
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11244 18828 11296 18834
rect 11244 18770 11296 18776
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 11072 17513 11100 18566
rect 11256 17785 11284 18770
rect 11348 18290 11376 21286
rect 11520 21140 11572 21146
rect 11520 21082 11572 21088
rect 11532 21010 11560 21082
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11440 18766 11468 20198
rect 11428 18760 11480 18766
rect 11428 18702 11480 18708
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11440 18086 11468 18702
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11242 17776 11298 17785
rect 11152 17740 11204 17746
rect 11242 17711 11298 17720
rect 11152 17682 11204 17688
rect 11058 17504 11114 17513
rect 11058 17439 11114 17448
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10876 17060 10928 17066
rect 10876 17002 10928 17008
rect 10888 15162 10916 17002
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10980 16182 11008 16730
rect 11072 16182 11100 17439
rect 11164 16590 11192 17682
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 10968 15496 11020 15502
rect 11072 15484 11100 16118
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11020 15456 11100 15484
rect 10968 15438 11020 15444
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 11072 14958 11100 15302
rect 10876 14952 10928 14958
rect 11060 14952 11112 14958
rect 10876 14894 10928 14900
rect 10980 14912 11060 14940
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10888 14482 10916 14894
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10704 14278 10732 14418
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10140 13932 10192 13938
rect 10428 13926 10548 13954
rect 10140 13874 10192 13880
rect 10416 13864 10468 13870
rect 9968 13280 10088 13308
rect 10336 13824 10416 13852
rect 9862 12744 9918 12753
rect 9862 12679 9918 12688
rect 9692 11478 9812 11506
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9508 11014 9536 11154
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9508 9926 9536 10950
rect 9600 10674 9628 11290
rect 9692 10742 9720 11478
rect 9770 11384 9826 11393
rect 9770 11319 9826 11328
rect 9784 11121 9812 11319
rect 9864 11144 9916 11150
rect 9770 11112 9826 11121
rect 9864 11086 9916 11092
rect 9770 11047 9826 11056
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9876 10674 9904 11086
rect 9968 10713 9996 13280
rect 10336 13274 10364 13824
rect 10416 13806 10468 13812
rect 10414 13696 10470 13705
rect 10414 13631 10470 13640
rect 10152 13246 10364 13274
rect 10428 13258 10456 13631
rect 10416 13252 10468 13258
rect 10046 13016 10102 13025
rect 10046 12951 10048 12960
rect 10100 12951 10102 12960
rect 10048 12922 10100 12928
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10060 12442 10088 12786
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10152 11082 10180 13246
rect 10416 13194 10468 13200
rect 10520 13190 10548 13926
rect 10704 13734 10732 14214
rect 10874 13832 10930 13841
rect 10874 13767 10930 13776
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10782 13696 10838 13705
rect 10782 13631 10838 13640
rect 10796 13444 10824 13631
rect 10888 13530 10916 13767
rect 10980 13530 11008 14912
rect 11060 14894 11112 14900
rect 11164 13546 11192 15846
rect 11256 14385 11284 17711
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11532 17202 11560 17614
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11428 16720 11480 16726
rect 11426 16688 11428 16697
rect 11480 16688 11482 16697
rect 11532 16658 11560 17138
rect 11426 16623 11482 16632
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11428 16516 11480 16522
rect 11428 16458 11480 16464
rect 11336 15632 11388 15638
rect 11440 15609 11468 16458
rect 11532 16114 11560 16594
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11532 15638 11560 16050
rect 11520 15632 11572 15638
rect 11336 15574 11388 15580
rect 11426 15600 11482 15609
rect 11348 14958 11376 15574
rect 11520 15574 11572 15580
rect 11426 15535 11482 15544
rect 11518 15192 11574 15201
rect 11518 15127 11574 15136
rect 11336 14952 11388 14958
rect 11388 14900 11468 14906
rect 11336 14894 11468 14900
rect 11348 14878 11468 14894
rect 11336 14816 11388 14822
rect 11334 14784 11336 14793
rect 11388 14784 11390 14793
rect 11334 14719 11390 14728
rect 11440 14482 11468 14878
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11336 14408 11388 14414
rect 11242 14376 11298 14385
rect 11336 14350 11388 14356
rect 11426 14376 11482 14385
rect 11242 14311 11298 14320
rect 11242 14240 11298 14249
rect 11242 14175 11298 14184
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 11072 13518 11192 13546
rect 10704 13416 10824 13444
rect 10704 13258 10732 13416
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10244 12968 10272 13126
rect 10244 12940 10548 12968
rect 10520 12850 10548 12940
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10508 12844 10560 12850
rect 10508 12786 10560 12792
rect 10428 12238 10456 12786
rect 10796 12442 10824 13262
rect 10980 12753 11008 13466
rect 11072 13258 11100 13518
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11060 13252 11112 13258
rect 11060 13194 11112 13200
rect 10966 12744 11022 12753
rect 11164 12714 11192 13330
rect 11256 12918 11284 14175
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 10966 12679 11022 12688
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 11058 12608 11114 12617
rect 11058 12543 11114 12552
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10508 11212 10560 11218
rect 10244 11172 10508 11200
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 9954 10704 10010 10713
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9864 10668 9916 10674
rect 10244 10690 10272 11172
rect 10784 11212 10836 11218
rect 10508 11154 10560 11160
rect 10704 11172 10784 11200
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 9954 10639 10010 10648
rect 10060 10662 10272 10690
rect 9864 10610 9916 10616
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9324 9178 9352 9454
rect 9416 9178 9444 9454
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9126 9072 9182 9081
rect 9126 9007 9182 9016
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 9508 8430 9536 9862
rect 10060 9625 10088 10662
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10140 10464 10192 10470
rect 10140 10406 10192 10412
rect 10152 10198 10180 10406
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 10046 9616 10102 9625
rect 10046 9551 10102 9560
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 8430 9628 9318
rect 10060 8974 10088 9551
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10244 8906 10272 10542
rect 10520 10130 10548 11018
rect 10704 10452 10732 11172
rect 10784 11154 10836 11160
rect 10888 10674 10916 12242
rect 11072 11286 11100 12543
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10612 10424 10732 10452
rect 10876 10464 10928 10470
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10336 9081 10364 9114
rect 10322 9072 10378 9081
rect 10612 9042 10640 10424
rect 10876 10406 10928 10412
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10704 9722 10732 10066
rect 10888 10062 10916 10406
rect 10876 10056 10928 10062
rect 10796 10016 10876 10044
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10796 9586 10824 10016
rect 10876 9998 10928 10004
rect 10980 9874 11008 11018
rect 11072 10198 11100 11018
rect 11164 10452 11192 12650
rect 11348 12442 11376 14350
rect 11426 14311 11482 14320
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11440 11778 11468 14311
rect 11532 13870 11560 15127
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11520 13728 11572 13734
rect 11518 13696 11520 13705
rect 11572 13696 11574 13705
rect 11518 13631 11574 13640
rect 11532 13462 11560 13631
rect 11624 13530 11652 21422
rect 12452 21146 12480 21927
rect 12532 21888 12584 21894
rect 12532 21830 12584 21836
rect 12544 21690 12572 21830
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12636 21554 12664 21966
rect 12820 21690 12848 22102
rect 16120 21956 16172 21962
rect 16120 21898 16172 21904
rect 18420 21956 18472 21962
rect 18420 21898 18472 21904
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 13740 21554 13768 21830
rect 16132 21690 16160 21898
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16120 21684 16172 21690
rect 16120 21626 16172 21632
rect 16684 21622 16712 21830
rect 13912 21616 13964 21622
rect 16672 21616 16724 21622
rect 13912 21558 13964 21564
rect 15198 21584 15254 21593
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13176 21344 13228 21350
rect 12714 21312 12770 21321
rect 13176 21286 13228 21292
rect 12714 21247 12770 21256
rect 12348 21140 12400 21146
rect 12348 21082 12400 21088
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12360 21026 12388 21082
rect 12360 20998 12480 21026
rect 11796 20936 11848 20942
rect 11702 20904 11758 20913
rect 11758 20884 11796 20890
rect 11758 20878 11848 20884
rect 11758 20862 11836 20878
rect 11702 20839 11758 20848
rect 11783 20700 12091 20709
rect 11783 20698 11789 20700
rect 11845 20698 11869 20700
rect 11925 20698 11949 20700
rect 12005 20698 12029 20700
rect 12085 20698 12091 20700
rect 11845 20646 11847 20698
rect 12027 20646 12029 20698
rect 11783 20644 11789 20646
rect 11845 20644 11869 20646
rect 11925 20644 11949 20646
rect 12005 20644 12029 20646
rect 12085 20644 12091 20646
rect 11783 20635 12091 20644
rect 11704 20392 11756 20398
rect 11704 20334 11756 20340
rect 11978 20360 12034 20369
rect 11716 19990 11744 20334
rect 11978 20295 12034 20304
rect 11796 20256 11848 20262
rect 11796 20198 11848 20204
rect 11704 19984 11756 19990
rect 11704 19926 11756 19932
rect 11808 19922 11836 20198
rect 11796 19916 11848 19922
rect 11796 19858 11848 19864
rect 11992 19854 12020 20295
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11992 19700 12020 19790
rect 11716 19672 12020 19700
rect 11716 19334 11744 19672
rect 11783 19612 12091 19621
rect 11783 19610 11789 19612
rect 11845 19610 11869 19612
rect 11925 19610 11949 19612
rect 12005 19610 12029 19612
rect 12085 19610 12091 19612
rect 11845 19558 11847 19610
rect 12027 19558 12029 19610
rect 11783 19556 11789 19558
rect 11845 19556 11869 19558
rect 11925 19556 11949 19558
rect 12005 19556 12029 19558
rect 12085 19556 12091 19558
rect 11783 19547 12091 19556
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 11992 19360 12020 19450
rect 12176 19378 12204 20198
rect 12452 20058 12480 20998
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12544 20505 12572 20538
rect 12530 20496 12586 20505
rect 12530 20431 12586 20440
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12268 19530 12296 19994
rect 12268 19514 12388 19530
rect 12268 19508 12400 19514
rect 12268 19502 12348 19508
rect 12348 19450 12400 19456
rect 12164 19372 12216 19378
rect 11716 19310 11928 19334
rect 11992 19332 12112 19360
rect 11716 19306 11940 19310
rect 11888 19304 11940 19306
rect 11888 19246 11940 19252
rect 12084 18850 12112 19332
rect 12164 19314 12216 19320
rect 12452 19258 12480 19994
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12360 19230 12480 19258
rect 12360 19174 12388 19230
rect 12452 19174 12480 19230
rect 12348 19168 12400 19174
rect 12348 19110 12400 19116
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12084 18822 12296 18850
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 11716 17678 11744 18702
rect 11783 18524 12091 18533
rect 11783 18522 11789 18524
rect 11845 18522 11869 18524
rect 11925 18522 11949 18524
rect 12005 18522 12029 18524
rect 12085 18522 12091 18524
rect 11845 18470 11847 18522
rect 12027 18470 12029 18522
rect 11783 18468 11789 18470
rect 11845 18468 11869 18470
rect 11925 18468 11949 18470
rect 12005 18468 12029 18470
rect 12085 18468 12091 18470
rect 11783 18459 12091 18468
rect 12176 17678 12204 18702
rect 12268 18358 12296 18822
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 11783 17436 12091 17445
rect 11783 17434 11789 17436
rect 11845 17434 11869 17436
rect 11925 17434 11949 17436
rect 12005 17434 12029 17436
rect 12085 17434 12091 17436
rect 11845 17382 11847 17434
rect 12027 17382 12029 17434
rect 11783 17380 11789 17382
rect 11845 17380 11869 17382
rect 11925 17380 11949 17382
rect 12005 17380 12029 17382
rect 12085 17380 12091 17382
rect 11783 17371 12091 17380
rect 12072 16992 12124 16998
rect 12176 16980 12204 17614
rect 12124 16952 12204 16980
rect 12072 16934 12124 16940
rect 11980 16584 12032 16590
rect 12176 16572 12204 16952
rect 12032 16544 12204 16572
rect 11980 16526 12032 16532
rect 11783 16348 12091 16357
rect 11783 16346 11789 16348
rect 11845 16346 11869 16348
rect 11925 16346 11949 16348
rect 12005 16346 12029 16348
rect 12085 16346 12091 16348
rect 11845 16294 11847 16346
rect 12027 16294 12029 16346
rect 11783 16292 11789 16294
rect 11845 16292 11869 16294
rect 11925 16292 11949 16294
rect 12005 16292 12029 16294
rect 12085 16292 12091 16294
rect 11783 16283 12091 16292
rect 11704 16108 11756 16114
rect 11756 16068 11836 16096
rect 11704 16050 11756 16056
rect 11808 15745 11836 16068
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 12072 15904 12124 15910
rect 12176 15892 12204 16544
rect 12124 15864 12204 15892
rect 12072 15846 12124 15852
rect 11794 15736 11850 15745
rect 11794 15671 11850 15680
rect 11900 15570 11928 15846
rect 12268 15586 12296 18294
rect 12346 18184 12402 18193
rect 12346 18119 12402 18128
rect 12360 17882 12388 18119
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12360 16590 12388 16730
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 11888 15564 11940 15570
rect 11716 15524 11888 15552
rect 11716 14822 11744 15524
rect 11888 15506 11940 15512
rect 12176 15558 12296 15586
rect 12176 15366 12204 15558
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 11783 15260 12091 15269
rect 11783 15258 11789 15260
rect 11845 15258 11869 15260
rect 11925 15258 11949 15260
rect 12005 15258 12029 15260
rect 12085 15258 12091 15260
rect 11845 15206 11847 15258
rect 12027 15206 12029 15258
rect 11783 15204 11789 15206
rect 11845 15204 11869 15206
rect 11925 15204 11949 15206
rect 12005 15204 12029 15206
rect 12085 15204 12091 15206
rect 11783 15195 12091 15204
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11808 15026 11836 15098
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11704 14816 11756 14822
rect 12176 14770 12204 15302
rect 11704 14758 11756 14764
rect 11716 14396 11744 14758
rect 12084 14742 12204 14770
rect 11796 14408 11848 14414
rect 11716 14368 11796 14396
rect 11716 14006 11744 14368
rect 11796 14350 11848 14356
rect 12084 14260 12112 14742
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 12084 14232 12148 14260
rect 11783 14172 12091 14181
rect 11783 14170 11789 14172
rect 11845 14170 11869 14172
rect 11925 14170 11949 14172
rect 12005 14170 12029 14172
rect 12085 14170 12091 14172
rect 11845 14118 11847 14170
rect 12027 14118 12029 14170
rect 11783 14116 11789 14118
rect 11845 14116 11869 14118
rect 11925 14116 11949 14118
rect 12005 14116 12029 14118
rect 12085 14116 12091 14118
rect 11783 14107 12091 14116
rect 12120 14056 12148 14232
rect 11992 14028 12148 14056
rect 11704 14000 11756 14006
rect 11704 13942 11756 13948
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11886 13832 11942 13841
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11520 13456 11572 13462
rect 11716 13410 11744 13466
rect 11520 13398 11572 13404
rect 11624 13382 11744 13410
rect 11518 13288 11574 13297
rect 11518 13223 11520 13232
rect 11572 13223 11574 13232
rect 11520 13194 11572 13200
rect 11624 12782 11652 13382
rect 11808 13172 11836 13806
rect 11886 13767 11942 13776
rect 11900 13462 11928 13767
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 11992 13394 12020 14028
rect 12072 13932 12124 13938
rect 12176 13920 12204 14554
rect 12268 14278 12296 15438
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12360 14074 12388 14214
rect 12452 14074 12480 14894
rect 12544 14074 12572 18702
rect 12636 18426 12664 19790
rect 12728 19553 12756 21247
rect 13188 20602 13216 21286
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 12992 20324 13044 20330
rect 12992 20266 13044 20272
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12820 19718 12848 19790
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12714 19544 12770 19553
rect 13004 19514 13032 20266
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 12714 19479 12770 19488
rect 12992 19508 13044 19514
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12728 16130 12756 19479
rect 12992 19450 13044 19456
rect 13096 19310 13124 19654
rect 13084 19304 13136 19310
rect 12898 19272 12954 19281
rect 13084 19246 13136 19252
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 12898 19207 12954 19216
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12820 16697 12848 16730
rect 12806 16688 12862 16697
rect 12806 16623 12862 16632
rect 12728 16102 12848 16130
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12636 14793 12664 14894
rect 12622 14784 12678 14793
rect 12622 14719 12678 14728
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12124 13892 12204 13920
rect 12072 13874 12124 13880
rect 12636 13870 12664 14418
rect 12728 14006 12756 15982
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12070 13560 12126 13569
rect 12070 13495 12126 13504
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11886 13288 11942 13297
rect 11886 13223 11942 13232
rect 11900 13190 11928 13223
rect 11716 13144 11836 13172
rect 11888 13184 11940 13190
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11612 12368 11664 12374
rect 11716 12356 11744 13144
rect 11992 13172 12020 13330
rect 12084 13297 12112 13495
rect 12532 13456 12584 13462
rect 12532 13398 12584 13404
rect 12440 13320 12492 13326
rect 12070 13288 12126 13297
rect 12440 13262 12492 13268
rect 12070 13223 12126 13232
rect 12256 13184 12308 13190
rect 11992 13144 12204 13172
rect 11888 13126 11940 13132
rect 11783 13084 12091 13093
rect 11783 13082 11789 13084
rect 11845 13082 11869 13084
rect 11925 13082 11949 13084
rect 12005 13082 12029 13084
rect 12085 13082 12091 13084
rect 11845 13030 11847 13082
rect 12027 13030 12029 13082
rect 11783 13028 11789 13030
rect 11845 13028 11869 13030
rect 11925 13028 11949 13030
rect 12005 13028 12029 13030
rect 12085 13028 12091 13030
rect 11783 13019 12091 13028
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11980 12776 12032 12782
rect 11978 12744 11980 12753
rect 12032 12744 12034 12753
rect 11978 12679 12034 12688
rect 11978 12472 12034 12481
rect 11978 12407 11980 12416
rect 12032 12407 12034 12416
rect 11980 12378 12032 12384
rect 11796 12368 11848 12374
rect 11716 12328 11796 12356
rect 11612 12310 11664 12316
rect 11796 12310 11848 12316
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11532 11898 11560 12038
rect 11624 11898 11652 12310
rect 12084 12306 12112 12854
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 11783 11996 12091 12005
rect 11783 11994 11789 11996
rect 11845 11994 11869 11996
rect 11925 11994 11949 11996
rect 12005 11994 12029 11996
rect 12085 11994 12091 11996
rect 11845 11942 11847 11994
rect 12027 11942 12029 11994
rect 11783 11940 11789 11942
rect 11845 11940 11869 11942
rect 11925 11940 11949 11942
rect 12005 11940 12029 11942
rect 12085 11940 12091 11942
rect 11783 11931 12091 11940
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11348 11750 11468 11778
rect 11532 11762 11928 11778
rect 11520 11756 11928 11762
rect 11244 11688 11296 11694
rect 11244 11630 11296 11636
rect 11256 11014 11284 11630
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11256 10674 11284 10950
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11348 10577 11376 11750
rect 11572 11750 11928 11756
rect 11520 11698 11572 11704
rect 11900 11694 11928 11750
rect 11612 11688 11664 11694
rect 11426 11656 11482 11665
rect 11426 11591 11482 11600
rect 11610 11656 11612 11665
rect 11796 11688 11848 11694
rect 11664 11656 11666 11665
rect 11610 11591 11666 11600
rect 11716 11648 11796 11676
rect 11440 11014 11468 11591
rect 11428 11008 11480 11014
rect 11520 11008 11572 11014
rect 11428 10950 11480 10956
rect 11518 10976 11520 10985
rect 11572 10976 11574 10985
rect 11518 10911 11574 10920
rect 11716 10810 11744 11648
rect 11796 11630 11848 11636
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 12070 11384 12126 11393
rect 12070 11319 12072 11328
rect 12124 11319 12126 11328
rect 12072 11290 12124 11296
rect 12176 11234 12204 13144
rect 12256 13126 12308 13132
rect 12268 12850 12296 13126
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12360 12782 12388 12922
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12256 12640 12308 12646
rect 12256 12582 12308 12588
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12268 11642 12296 12582
rect 12360 11762 12388 12582
rect 12452 12288 12480 13262
rect 12544 12424 12572 13398
rect 12636 12617 12664 13806
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12728 13530 12756 13738
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12820 13138 12848 16102
rect 12912 13870 12940 19207
rect 13188 18970 13216 19246
rect 13176 18964 13228 18970
rect 13176 18906 13228 18912
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 13004 15065 13032 18566
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 13096 16250 13124 16934
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13096 15706 13124 15846
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13188 15586 13216 17002
rect 13096 15558 13216 15586
rect 12990 15056 13046 15065
rect 12990 14991 13046 15000
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12728 13110 12848 13138
rect 12728 12986 12756 13110
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12622 12608 12678 12617
rect 12622 12543 12678 12552
rect 12820 12442 12848 12922
rect 12808 12436 12860 12442
rect 12544 12396 12756 12424
rect 12532 12300 12584 12306
rect 12452 12260 12532 12288
rect 12452 11762 12480 12260
rect 12532 12242 12584 12248
rect 12728 11898 12756 12396
rect 12808 12378 12860 12384
rect 12912 12102 12940 13806
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 13004 12986 13032 13262
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 13096 12866 13124 15558
rect 13280 14770 13308 21490
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 13372 20369 13400 21286
rect 13544 21004 13596 21010
rect 13544 20946 13596 20952
rect 13358 20360 13414 20369
rect 13358 20295 13414 20304
rect 13372 19334 13400 20295
rect 13556 20058 13584 20946
rect 13820 20528 13872 20534
rect 13818 20496 13820 20505
rect 13872 20496 13874 20505
rect 13818 20431 13874 20440
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13372 19310 13584 19334
rect 13372 19306 13596 19310
rect 13544 19304 13596 19306
rect 13544 19246 13596 19252
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13464 17542 13492 18906
rect 13740 18290 13768 19926
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13544 18216 13596 18222
rect 13544 18158 13596 18164
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13464 15706 13492 17138
rect 13452 15700 13504 15706
rect 13452 15642 13504 15648
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13188 14742 13308 14770
rect 13188 14482 13216 14742
rect 13266 14648 13322 14657
rect 13372 14618 13400 15302
rect 13452 14884 13504 14890
rect 13452 14826 13504 14832
rect 13266 14583 13322 14592
rect 13360 14612 13412 14618
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13280 13682 13308 14583
rect 13360 14554 13412 14560
rect 13280 13654 13400 13682
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13280 13326 13308 13466
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13372 13025 13400 13654
rect 13358 13016 13414 13025
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13280 12974 13358 13002
rect 13004 12838 13124 12866
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12268 11614 12388 11642
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12268 11354 12296 11494
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12084 11206 12204 11234
rect 12084 10996 12112 11206
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12084 10968 12148 10996
rect 11783 10908 12091 10917
rect 11783 10906 11789 10908
rect 11845 10906 11869 10908
rect 11925 10906 11949 10908
rect 12005 10906 12029 10908
rect 12085 10906 12091 10908
rect 11845 10854 11847 10906
rect 12027 10854 12029 10906
rect 11783 10852 11789 10854
rect 11845 10852 11869 10854
rect 11925 10852 11949 10854
rect 12005 10852 12029 10854
rect 12085 10852 12091 10854
rect 11783 10843 12091 10852
rect 11704 10804 11756 10810
rect 12120 10792 12148 10968
rect 11704 10746 11756 10752
rect 12084 10764 12148 10792
rect 11334 10568 11390 10577
rect 11334 10503 11390 10512
rect 11164 10424 11652 10452
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 10888 9846 11008 9874
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10782 9480 10838 9489
rect 10782 9415 10838 9424
rect 10796 9382 10824 9415
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10888 9160 10916 9846
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 10704 9132 10916 9160
rect 10322 9007 10378 9016
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 9862 8800 9918 8809
rect 9918 8758 9996 8786
rect 9862 8735 9918 8744
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 6798 9168 8230
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9232 6662 9260 7278
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 8864 6412 9260 6440
rect 8444 6344 8524 6372
rect 8392 6326 8444 6332
rect 8576 6316 8628 6322
rect 9036 6316 9088 6322
rect 8576 6258 8628 6264
rect 8864 6276 9036 6304
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 7988 6012 8296 6021
rect 7988 6010 7994 6012
rect 8050 6010 8074 6012
rect 8130 6010 8154 6012
rect 8210 6010 8234 6012
rect 8290 6010 8296 6012
rect 8050 5958 8052 6010
rect 8232 5958 8234 6010
rect 7988 5956 7994 5958
rect 8050 5956 8074 5958
rect 8130 5956 8154 5958
rect 8210 5956 8234 5958
rect 8290 5956 8296 5958
rect 7988 5947 8296 5956
rect 7852 5868 7972 5896
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7194 3904 7250 3913
rect 7194 3839 7250 3848
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6840 2938 6868 3674
rect 7576 3602 7604 5238
rect 7668 5234 7696 5510
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7852 4826 7880 5714
rect 7944 5166 7972 5868
rect 8300 5704 8352 5710
rect 8404 5692 8432 6190
rect 8352 5664 8432 5692
rect 8300 5646 8352 5652
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 7988 4924 8296 4933
rect 7988 4922 7994 4924
rect 8050 4922 8074 4924
rect 8130 4922 8154 4924
rect 8210 4922 8234 4924
rect 8290 4922 8296 4924
rect 8050 4870 8052 4922
rect 8232 4870 8234 4922
rect 7988 4868 7994 4870
rect 8050 4868 8074 4870
rect 8130 4868 8154 4870
rect 8210 4868 8234 4870
rect 8290 4868 8296 4870
rect 7988 4859 8296 4868
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 4282 8340 4558
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8404 4214 8432 4966
rect 8496 4554 8524 6190
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8392 4208 8444 4214
rect 8392 4150 8444 4156
rect 8588 4146 8616 6258
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8680 5914 8708 6054
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8680 4146 8708 5850
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8772 5574 8800 5646
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8760 5092 8812 5098
rect 8760 5034 8812 5040
rect 8772 5001 8800 5034
rect 8758 4992 8814 5001
rect 8758 4927 8814 4936
rect 8864 4842 8892 6276
rect 9036 6258 9088 6264
rect 9126 6080 9182 6089
rect 9126 6015 9182 6024
rect 8944 5568 8996 5574
rect 8942 5536 8944 5545
rect 8996 5536 8998 5545
rect 8942 5471 8998 5480
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 8772 4814 8892 4842
rect 8576 4140 8628 4146
rect 8576 4082 8628 4088
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 7988 3836 8296 3845
rect 7988 3834 7994 3836
rect 8050 3834 8074 3836
rect 8130 3834 8154 3836
rect 8210 3834 8234 3836
rect 8290 3834 8296 3836
rect 8050 3782 8052 3834
rect 8232 3782 8234 3834
rect 7988 3780 7994 3782
rect 8050 3780 8074 3782
rect 8130 3780 8154 3782
rect 8210 3780 8234 3782
rect 8290 3780 8296 3782
rect 7988 3771 8296 3780
rect 8680 3738 8708 4082
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8772 3618 8800 4814
rect 8852 4616 8904 4622
rect 8956 4604 8984 5102
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 9048 4622 9076 4966
rect 8904 4576 8984 4604
rect 9036 4616 9088 4622
rect 8852 4558 8904 4564
rect 9036 4558 9088 4564
rect 7564 3596 7616 3602
rect 7564 3538 7616 3544
rect 8588 3590 8800 3618
rect 7012 3528 7064 3534
rect 8300 3528 8352 3534
rect 7012 3470 7064 3476
rect 8298 3496 8300 3505
rect 8352 3496 8354 3505
rect 6840 2910 6960 2938
rect 6932 2854 6960 2910
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6656 2746 6868 2774
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6552 2440 6604 2446
rect 6550 2408 6552 2417
rect 6604 2408 6606 2417
rect 6550 2343 6606 2352
rect 6656 1970 6684 2586
rect 6840 1970 6868 2746
rect 6460 1964 6512 1970
rect 6460 1906 6512 1912
rect 6644 1964 6696 1970
rect 6644 1906 6696 1912
rect 6828 1964 6880 1970
rect 6828 1906 6880 1912
rect 6000 1896 6052 1902
rect 6000 1838 6052 1844
rect 6274 1864 6330 1873
rect 6274 1799 6330 1808
rect 6000 1760 6052 1766
rect 6000 1702 6052 1708
rect 5816 1488 5868 1494
rect 5816 1430 5868 1436
rect 5630 1184 5686 1193
rect 5630 1119 5686 1128
rect 5172 944 5224 950
rect 5172 886 5224 892
rect 5644 814 5672 1119
rect 5632 808 5684 814
rect 5632 750 5684 756
rect 5816 808 5868 814
rect 5816 750 5868 756
rect 5356 672 5408 678
rect 5356 614 5408 620
rect 5448 672 5500 678
rect 5448 614 5500 620
rect 5368 202 5396 614
rect 5460 338 5488 614
rect 5448 332 5500 338
rect 5448 274 5500 280
rect 5080 196 5132 202
rect 5080 138 5132 144
rect 5356 196 5408 202
rect 5356 138 5408 144
rect 3790 96 3846 105
rect 5828 66 5856 750
rect 6012 270 6040 1702
rect 6288 1494 6316 1799
rect 6276 1488 6328 1494
rect 6276 1430 6328 1436
rect 6472 1426 6500 1906
rect 6932 1766 6960 2790
rect 7024 2650 7052 3470
rect 8298 3431 8354 3440
rect 7654 3224 7710 3233
rect 7654 3159 7710 3168
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7668 2514 7696 3159
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 7988 2748 8296 2757
rect 7988 2746 7994 2748
rect 8050 2746 8074 2748
rect 8130 2746 8154 2748
rect 8210 2746 8234 2748
rect 8290 2746 8296 2748
rect 8050 2694 8052 2746
rect 8232 2694 8234 2746
rect 7988 2692 7994 2694
rect 8050 2692 8074 2694
rect 8130 2692 8154 2694
rect 8210 2692 8234 2694
rect 8290 2692 8296 2694
rect 7988 2683 8296 2692
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 6920 1760 6972 1766
rect 6920 1702 6972 1708
rect 6642 1592 6698 1601
rect 6932 1562 6960 1702
rect 7988 1660 8296 1669
rect 7988 1658 7994 1660
rect 8050 1658 8074 1660
rect 8130 1658 8154 1660
rect 8210 1658 8234 1660
rect 8290 1658 8296 1660
rect 8050 1606 8052 1658
rect 8232 1606 8234 1658
rect 7988 1604 7994 1606
rect 8050 1604 8074 1606
rect 8130 1604 8154 1606
rect 8210 1604 8234 1606
rect 8290 1604 8296 1606
rect 7988 1595 8296 1604
rect 6642 1527 6698 1536
rect 6920 1556 6972 1562
rect 6460 1420 6512 1426
rect 6460 1362 6512 1368
rect 6656 882 6684 1527
rect 6920 1498 6972 1504
rect 8208 1488 8260 1494
rect 8260 1448 8340 1476
rect 8208 1430 8260 1436
rect 6920 1352 6972 1358
rect 6920 1294 6972 1300
rect 6932 1018 6960 1294
rect 7656 1216 7708 1222
rect 7656 1158 7708 1164
rect 7668 1018 7696 1158
rect 6920 1012 6972 1018
rect 6920 954 6972 960
rect 7656 1012 7708 1018
rect 7656 954 7708 960
rect 6276 876 6328 882
rect 6276 818 6328 824
rect 6644 876 6696 882
rect 6644 818 6696 824
rect 6000 264 6052 270
rect 6288 241 6316 818
rect 7840 808 7892 814
rect 7840 750 7892 756
rect 7564 672 7616 678
rect 7564 614 7616 620
rect 7576 474 7604 614
rect 7852 474 7880 750
rect 8312 678 8340 1448
rect 8404 882 8432 2790
rect 8588 1358 8616 3590
rect 8864 3534 8892 4558
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8666 3360 8722 3369
rect 8666 3295 8722 3304
rect 8680 2825 8708 3295
rect 8864 2990 8892 3470
rect 8956 3398 8984 4014
rect 9048 3738 9076 4558
rect 9140 4078 9168 6015
rect 9232 5080 9260 6412
rect 9324 5370 9352 7822
rect 9416 7177 9444 8366
rect 9772 7744 9824 7750
rect 9586 7712 9642 7721
rect 9772 7686 9824 7692
rect 9586 7647 9642 7656
rect 9402 7168 9458 7177
rect 9402 7103 9458 7112
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9416 6905 9444 6938
rect 9402 6896 9458 6905
rect 9402 6831 9458 6840
rect 9496 6792 9548 6798
rect 9402 6760 9458 6769
rect 9458 6740 9496 6746
rect 9458 6734 9548 6740
rect 9458 6718 9536 6734
rect 9402 6695 9458 6704
rect 9600 6662 9628 7647
rect 9784 6769 9812 7686
rect 9770 6760 9826 6769
rect 9770 6695 9826 6704
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9416 5234 9444 5306
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9232 5052 9352 5080
rect 9218 4992 9274 5001
rect 9218 4927 9274 4936
rect 9232 4622 9260 4927
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9324 4026 9352 5052
rect 9496 4820 9548 4826
rect 9600 4808 9628 6054
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9772 5226 9824 5232
rect 9692 5030 9720 5170
rect 9772 5168 9824 5174
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9784 4826 9812 5168
rect 9548 4780 9628 4808
rect 9772 4820 9824 4826
rect 9496 4762 9548 4768
rect 9772 4762 9824 4768
rect 9402 4720 9458 4729
rect 9496 4684 9548 4690
rect 9458 4664 9496 4672
rect 9402 4655 9496 4664
rect 9416 4644 9496 4655
rect 9496 4626 9548 4632
rect 9876 4486 9904 6598
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9324 3998 9536 4026
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9048 3534 9076 3674
rect 9324 3534 9352 3878
rect 9416 3602 9444 3878
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8666 2816 8722 2825
rect 8956 2774 8984 3334
rect 9048 2854 9076 3470
rect 9508 3176 9536 3998
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9416 3148 9536 3176
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 8666 2751 8722 2760
rect 8680 2582 8708 2751
rect 8772 2746 8984 2774
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8772 2514 8800 2746
rect 9048 2650 9076 2790
rect 9324 2650 9352 2926
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 8772 1902 8800 2450
rect 8760 1896 8812 1902
rect 8760 1838 8812 1844
rect 8852 1896 8904 1902
rect 8852 1838 8904 1844
rect 8864 1358 8892 1838
rect 9048 1766 9076 2586
rect 9324 2514 9352 2586
rect 9416 2514 9444 3148
rect 9600 3058 9628 3470
rect 9692 3194 9720 3538
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9784 3097 9812 4218
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9876 3194 9904 4150
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9770 3088 9826 3097
rect 9588 3052 9640 3058
rect 9770 3023 9826 3032
rect 9588 2994 9640 3000
rect 9968 2774 9996 8758
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 6798 10272 7686
rect 10336 7002 10364 8910
rect 10428 8906 10456 8978
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10612 8430 10640 8978
rect 10704 8498 10732 9132
rect 10980 9058 11008 9658
rect 10888 9030 11008 9058
rect 10888 8838 10916 9030
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10690 8392 10746 8401
rect 10690 8327 10746 8336
rect 10968 8356 11020 8362
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10520 7585 10548 7958
rect 10598 7848 10654 7857
rect 10598 7783 10600 7792
rect 10652 7783 10654 7792
rect 10600 7754 10652 7760
rect 10506 7576 10562 7585
rect 10506 7511 10562 7520
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5030 10088 6054
rect 10428 5778 10456 7278
rect 10520 7041 10548 7511
rect 10506 7032 10562 7041
rect 10506 6967 10562 6976
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10048 4208 10100 4214
rect 10048 4150 10100 4156
rect 9692 2746 9996 2774
rect 9494 2544 9550 2553
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 9404 2508 9456 2514
rect 9494 2479 9550 2488
rect 9404 2450 9456 2456
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9036 1760 9088 1766
rect 9036 1702 9088 1708
rect 9048 1358 9076 1702
rect 9140 1562 9168 2382
rect 9324 1902 9352 2450
rect 9508 2281 9536 2479
rect 9494 2272 9550 2281
rect 9494 2207 9550 2216
rect 9494 2136 9550 2145
rect 9494 2071 9550 2080
rect 9312 1896 9364 1902
rect 9508 1850 9536 2071
rect 9692 1970 9720 2746
rect 10060 2650 10088 4150
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10152 3670 10180 3946
rect 10140 3664 10192 3670
rect 10140 3606 10192 3612
rect 10244 3602 10272 5510
rect 10336 4146 10364 5646
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10428 4078 10456 5714
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9864 2100 9916 2106
rect 9864 2042 9916 2048
rect 9876 1970 9904 2042
rect 9680 1964 9732 1970
rect 9680 1906 9732 1912
rect 9864 1964 9916 1970
rect 9864 1906 9916 1912
rect 9312 1838 9364 1844
rect 9416 1822 9720 1850
rect 9128 1556 9180 1562
rect 9128 1498 9180 1504
rect 8576 1352 8628 1358
rect 8576 1294 8628 1300
rect 8852 1352 8904 1358
rect 8852 1294 8904 1300
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 9312 1352 9364 1358
rect 9312 1294 9364 1300
rect 9324 1018 9352 1294
rect 9416 1193 9444 1822
rect 9692 1766 9720 1822
rect 9680 1760 9732 1766
rect 9680 1702 9732 1708
rect 10416 1760 10468 1766
rect 10416 1702 10468 1708
rect 10428 1494 10456 1702
rect 10416 1488 10468 1494
rect 10416 1430 10468 1436
rect 9402 1184 9458 1193
rect 9402 1119 9458 1128
rect 9312 1012 9364 1018
rect 9312 954 9364 960
rect 10520 882 10548 6967
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 6225 10640 6598
rect 10598 6216 10654 6225
rect 10598 6151 10654 6160
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3738 10640 3878
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10704 1873 10732 8327
rect 10968 8298 11020 8304
rect 10980 7342 11008 8298
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 11072 6746 11100 10134
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11164 9674 11192 9862
rect 11164 9646 11284 9674
rect 11256 9586 11284 9646
rect 11348 9586 11376 9998
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11336 9580 11388 9586
rect 11336 9522 11388 9528
rect 11348 9042 11376 9522
rect 11624 9518 11652 10424
rect 12084 10282 12112 10764
rect 12176 10470 12204 11086
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12084 10254 12204 10282
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11716 9722 11744 9998
rect 11783 9820 12091 9829
rect 11783 9818 11789 9820
rect 11845 9818 11869 9820
rect 11925 9818 11949 9820
rect 12005 9818 12029 9820
rect 12085 9818 12091 9820
rect 11845 9766 11847 9818
rect 12027 9766 12029 9818
rect 11783 9764 11789 9766
rect 11845 9764 11869 9766
rect 11925 9764 11949 9766
rect 12005 9764 12029 9766
rect 12085 9764 12091 9766
rect 11783 9755 12091 9764
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 11900 9625 11928 9658
rect 11886 9616 11942 9625
rect 11886 9551 11942 9560
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11532 9178 11560 9454
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11426 9072 11482 9081
rect 11336 9036 11388 9042
rect 11482 9042 11652 9058
rect 11482 9036 11664 9042
rect 11482 9030 11612 9036
rect 11426 9007 11482 9016
rect 11336 8978 11388 8984
rect 11612 8978 11664 8984
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11164 8498 11192 8910
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 11256 7886 11284 8298
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11256 7342 11284 7822
rect 11348 7342 11376 8774
rect 11532 8634 11560 8910
rect 11783 8732 12091 8741
rect 11783 8730 11789 8732
rect 11845 8730 11869 8732
rect 11925 8730 11949 8732
rect 12005 8730 12029 8732
rect 12085 8730 12091 8732
rect 11845 8678 11847 8730
rect 12027 8678 12029 8730
rect 11783 8676 11789 8678
rect 11845 8676 11869 8678
rect 11925 8676 11949 8678
rect 12005 8676 12029 8678
rect 12085 8676 12091 8678
rect 11783 8667 12091 8676
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11624 7449 11652 8570
rect 12176 8362 12204 10254
rect 12268 9489 12296 11290
rect 12360 11286 12388 11614
rect 12348 11280 12400 11286
rect 12348 11222 12400 11228
rect 12452 11150 12480 11698
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12360 10742 12388 11018
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12544 10470 12572 10542
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12254 9480 12310 9489
rect 12254 9415 12310 9424
rect 12164 8356 12216 8362
rect 12164 8298 12216 8304
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11610 7440 11666 7449
rect 11610 7375 11666 7384
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11336 7336 11388 7342
rect 11388 7296 11468 7324
rect 11336 7278 11388 7284
rect 10980 6718 11100 6746
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 10980 6338 11008 6718
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 6458 11100 6598
rect 11164 6458 11192 6734
rect 11256 6730 11284 7278
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 7002 11376 7142
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 11440 6882 11468 7296
rect 11716 7206 11744 7890
rect 11783 7644 12091 7653
rect 11783 7642 11789 7644
rect 11845 7642 11869 7644
rect 11925 7642 11949 7644
rect 12005 7642 12029 7644
rect 12085 7642 12091 7644
rect 11845 7590 11847 7642
rect 12027 7590 12029 7642
rect 11783 7588 11789 7590
rect 11845 7588 11869 7590
rect 11925 7588 11949 7590
rect 12005 7588 12029 7590
rect 12085 7588 12091 7590
rect 11783 7579 12091 7588
rect 12268 7342 12296 8026
rect 12360 7410 12388 9862
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11348 6854 11468 6882
rect 11716 6866 11744 7142
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 11704 6860 11756 6866
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 10980 6310 11100 6338
rect 11072 6254 11100 6310
rect 11256 6254 11284 6666
rect 11348 6662 11376 6854
rect 11704 6802 11756 6808
rect 11520 6792 11572 6798
rect 11440 6752 11520 6780
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 10876 6248 10928 6254
rect 10874 6216 10876 6225
rect 11060 6248 11112 6254
rect 10928 6216 10930 6225
rect 11060 6190 11112 6196
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 10874 6151 10930 6160
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11256 5642 11284 5714
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 10796 4146 10824 5510
rect 11164 5234 11192 5510
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11150 5128 11206 5137
rect 11150 5063 11206 5072
rect 11164 4826 11192 5063
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11256 4758 11284 5578
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11348 4690 11376 6598
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11440 4570 11468 6752
rect 11520 6734 11572 6740
rect 11612 6316 11664 6322
rect 11716 6304 11744 6802
rect 12084 6798 12112 6938
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11783 6556 12091 6565
rect 11783 6554 11789 6556
rect 11845 6554 11869 6556
rect 11925 6554 11949 6556
rect 12005 6554 12029 6556
rect 12085 6554 12091 6556
rect 11845 6502 11847 6554
rect 12027 6502 12029 6554
rect 11783 6500 11789 6502
rect 11845 6500 11869 6502
rect 11925 6500 11949 6502
rect 12005 6500 12029 6502
rect 12085 6500 12091 6502
rect 11783 6491 12091 6500
rect 12452 6322 12480 9318
rect 12544 7177 12572 10406
rect 12636 10266 12664 10542
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12728 9110 12756 11834
rect 13004 10810 13032 12838
rect 13188 12782 13216 12922
rect 13176 12776 13228 12782
rect 13096 12724 13176 12730
rect 13096 12718 13228 12724
rect 13096 12702 13216 12718
rect 13096 12481 13124 12702
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 13082 12472 13138 12481
rect 13082 12407 13138 12416
rect 13188 12306 13216 12582
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13174 12064 13230 12073
rect 13096 11830 13124 12038
rect 13174 11999 13230 12008
rect 13084 11824 13136 11830
rect 13084 11766 13136 11772
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 13188 10742 13216 11999
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 12898 10568 12954 10577
rect 12898 10503 12954 10512
rect 12912 10470 12940 10503
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 13280 10198 13308 12974
rect 13358 12951 13414 12960
rect 13464 12073 13492 14826
rect 13450 12064 13506 12073
rect 13450 11999 13506 12008
rect 13556 11914 13584 18158
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13648 17105 13676 17478
rect 13634 17096 13690 17105
rect 13634 17031 13690 17040
rect 13726 16824 13782 16833
rect 13726 16759 13782 16768
rect 13740 15434 13768 16759
rect 13832 16454 13860 18022
rect 13924 17746 13952 21558
rect 16672 21558 16724 21564
rect 17958 21584 18014 21593
rect 15198 21519 15254 21528
rect 17958 21519 18014 21528
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14016 18057 14044 18226
rect 14002 18048 14058 18057
rect 14002 17983 14058 17992
rect 13912 17740 13964 17746
rect 13912 17682 13964 17688
rect 13912 17536 13964 17542
rect 13912 17478 13964 17484
rect 13924 17338 13952 17478
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14004 17128 14056 17134
rect 13910 17096 13966 17105
rect 14004 17070 14056 17076
rect 13910 17031 13912 17040
rect 13964 17031 13966 17040
rect 13912 17002 13964 17008
rect 14016 16590 14044 17070
rect 14004 16584 14056 16590
rect 13910 16552 13966 16561
rect 14004 16526 14056 16532
rect 13910 16487 13966 16496
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13818 16280 13874 16289
rect 13818 16215 13874 16224
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13648 15026 13676 15302
rect 13832 15178 13860 16215
rect 13740 15150 13860 15178
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13740 14890 13768 15150
rect 13924 15094 13952 16487
rect 14016 15910 14044 16526
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 14016 15502 14044 15846
rect 14004 15496 14056 15502
rect 14004 15438 14056 15444
rect 13912 15088 13964 15094
rect 13912 15030 13964 15036
rect 14016 14890 14044 15438
rect 14108 15094 14136 21422
rect 14384 21026 14412 21422
rect 14660 21078 14688 21422
rect 15212 21146 15240 21519
rect 15936 21412 15988 21418
rect 15936 21354 15988 21360
rect 15578 21244 15886 21253
rect 15578 21242 15584 21244
rect 15640 21242 15664 21244
rect 15720 21242 15744 21244
rect 15800 21242 15824 21244
rect 15880 21242 15886 21244
rect 15640 21190 15642 21242
rect 15822 21190 15824 21242
rect 15578 21188 15584 21190
rect 15640 21188 15664 21190
rect 15720 21188 15744 21190
rect 15800 21188 15824 21190
rect 15880 21188 15886 21190
rect 15578 21179 15886 21188
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 14292 21010 14412 21026
rect 14648 21072 14700 21078
rect 14648 21014 14700 21020
rect 14280 21004 14412 21010
rect 14332 20998 14412 21004
rect 14280 20946 14332 20952
rect 14280 20528 14332 20534
rect 14280 20470 14332 20476
rect 14292 20398 14320 20470
rect 14280 20392 14332 20398
rect 14384 20346 14412 20998
rect 14660 20466 14688 21014
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14332 20340 14412 20346
rect 14280 20334 14412 20340
rect 14292 20318 14412 20334
rect 14384 19854 14412 20318
rect 14554 20360 14610 20369
rect 14554 20295 14610 20304
rect 14568 19922 14596 20295
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14384 19378 14412 19790
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14200 18970 14228 19110
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14200 17270 14228 18770
rect 14292 18329 14320 19246
rect 14370 19000 14426 19009
rect 14370 18935 14426 18944
rect 14384 18737 14412 18935
rect 14476 18766 14504 19450
rect 14660 18834 14688 20402
rect 14844 20330 14872 20946
rect 15108 20800 15160 20806
rect 15108 20742 15160 20748
rect 15292 20800 15344 20806
rect 15292 20742 15344 20748
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 14844 19922 14872 20266
rect 14832 19916 14884 19922
rect 15120 19904 15148 20742
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15212 20058 15240 20402
rect 15304 20330 15332 20742
rect 15948 20466 15976 21354
rect 17972 21146 18000 21519
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 18432 21010 18460 21898
rect 18524 21690 18552 22170
rect 18604 22160 18656 22166
rect 18604 22102 18656 22108
rect 18512 21684 18564 21690
rect 18512 21626 18564 21632
rect 18616 21486 18644 22102
rect 18800 21622 18828 22238
rect 22466 22264 22522 22273
rect 21638 22199 21694 22208
rect 22376 22228 22428 22234
rect 19246 22128 19302 22137
rect 19246 22063 19302 22072
rect 19260 21962 19288 22063
rect 19248 21956 19300 21962
rect 19248 21898 19300 21904
rect 21364 21888 21416 21894
rect 21364 21830 21416 21836
rect 19373 21788 19681 21797
rect 19373 21786 19379 21788
rect 19435 21786 19459 21788
rect 19515 21786 19539 21788
rect 19595 21786 19619 21788
rect 19675 21786 19681 21788
rect 19435 21734 19437 21786
rect 19617 21734 19619 21786
rect 19373 21732 19379 21734
rect 19435 21732 19459 21734
rect 19515 21732 19539 21734
rect 19595 21732 19619 21734
rect 19675 21732 19681 21734
rect 19373 21723 19681 21732
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18510 21040 18566 21049
rect 18144 21004 18196 21010
rect 18144 20946 18196 20952
rect 18420 21004 18472 21010
rect 18510 20975 18566 20984
rect 18420 20946 18472 20952
rect 16396 20936 16448 20942
rect 16396 20878 16448 20884
rect 16118 20496 16174 20505
rect 15936 20460 15988 20466
rect 16118 20431 16174 20440
rect 15936 20402 15988 20408
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15304 20058 15332 20266
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15578 20156 15886 20165
rect 15578 20154 15584 20156
rect 15640 20154 15664 20156
rect 15720 20154 15744 20156
rect 15800 20154 15824 20156
rect 15880 20154 15886 20156
rect 15640 20102 15642 20154
rect 15822 20102 15824 20154
rect 15578 20100 15584 20102
rect 15640 20100 15664 20102
rect 15720 20100 15744 20102
rect 15800 20100 15824 20102
rect 15880 20100 15886 20102
rect 15578 20091 15886 20100
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15568 19916 15620 19922
rect 14832 19858 14884 19864
rect 15028 19876 15568 19904
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 14464 18760 14516 18766
rect 14370 18728 14426 18737
rect 14464 18702 14516 18708
rect 14370 18663 14426 18672
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14278 18320 14334 18329
rect 14278 18255 14334 18264
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14292 17513 14320 17614
rect 14464 17536 14516 17542
rect 14278 17504 14334 17513
rect 14464 17478 14516 17484
rect 14278 17439 14334 17448
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14200 17082 14228 17206
rect 14200 17054 14412 17082
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14200 16590 14228 16934
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 14200 15910 14228 16526
rect 14384 16250 14412 17054
rect 14476 16658 14504 17478
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 14004 14884 14056 14890
rect 14004 14826 14056 14832
rect 13740 13954 13768 14826
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14002 14648 14058 14657
rect 14002 14583 14058 14592
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13924 14074 13952 14418
rect 14016 14414 14044 14583
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 14108 14006 14136 14758
rect 14292 14362 14320 14894
rect 14384 14822 14412 16186
rect 14476 15994 14504 16390
rect 14568 16114 14596 18566
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14476 15966 14596 15994
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14476 15570 14504 15846
rect 14568 15570 14596 15966
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14476 14414 14504 14894
rect 14200 14334 14320 14362
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14200 14278 14228 14334
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14096 14000 14148 14006
rect 13648 13926 13768 13954
rect 14016 13960 14096 13988
rect 13648 12986 13676 13926
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 13912 13796 13964 13802
rect 13912 13738 13964 13744
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13648 12442 13676 12786
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13464 11886 13584 11914
rect 13464 11665 13492 11886
rect 13544 11824 13596 11830
rect 13544 11766 13596 11772
rect 13556 11694 13584 11766
rect 13648 11694 13676 12378
rect 13740 12306 13768 13738
rect 13924 13462 13952 13738
rect 13912 13456 13964 13462
rect 13912 13398 13964 13404
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 13818 13016 13874 13025
rect 13818 12951 13874 12960
rect 13832 12782 13860 12951
rect 13924 12850 13952 13262
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 14016 12714 14044 13960
rect 14096 13942 14148 13948
rect 14200 13870 14228 14214
rect 14384 13977 14412 14350
rect 14370 13968 14426 13977
rect 14370 13903 14426 13912
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14188 13864 14240 13870
rect 14188 13806 14240 13812
rect 14108 12986 14136 13806
rect 14556 13728 14608 13734
rect 14278 13696 14334 13705
rect 14556 13670 14608 13676
rect 14278 13631 14334 13640
rect 14292 13530 14320 13631
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14292 12832 14320 13126
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14462 12880 14518 12889
rect 14108 12804 14320 12832
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 13818 12608 13874 12617
rect 13818 12543 13874 12552
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13544 11688 13596 11694
rect 13450 11656 13506 11665
rect 13360 11620 13412 11626
rect 13544 11630 13596 11636
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13450 11591 13506 11600
rect 13360 11562 13412 11568
rect 13372 10742 13400 11562
rect 13464 11540 13492 11591
rect 13464 11512 13584 11540
rect 13556 11150 13584 11512
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13832 10606 13860 12543
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13924 12102 13952 12242
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12912 8922 12940 9862
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13096 9042 13124 9522
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 12728 8894 12940 8922
rect 12728 8430 12756 8894
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12636 7857 12664 8366
rect 12622 7848 12678 7857
rect 12622 7783 12678 7792
rect 12728 7274 12756 8366
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12530 7168 12586 7177
rect 12530 7103 12586 7112
rect 11664 6276 11744 6304
rect 12440 6316 12492 6322
rect 11612 6258 11664 6264
rect 12440 6258 12492 6264
rect 11612 5704 11664 5710
rect 11796 5704 11848 5710
rect 11612 5646 11664 5652
rect 11716 5664 11796 5692
rect 11520 5160 11572 5166
rect 11624 5148 11652 5646
rect 11716 5352 11744 5664
rect 11796 5646 11848 5652
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 11783 5468 12091 5477
rect 11783 5466 11789 5468
rect 11845 5466 11869 5468
rect 11925 5466 11949 5468
rect 12005 5466 12029 5468
rect 12085 5466 12091 5468
rect 11845 5414 11847 5466
rect 12027 5414 12029 5466
rect 11783 5412 11789 5414
rect 11845 5412 11869 5414
rect 11925 5412 11949 5414
rect 12005 5412 12029 5414
rect 12085 5412 12091 5414
rect 11783 5403 12091 5412
rect 11716 5324 11928 5352
rect 11900 5234 11928 5324
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11572 5120 11652 5148
rect 11520 5102 11572 5108
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4826 11560 4966
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11624 4690 11652 5120
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11164 4542 11468 4570
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 11164 3233 11192 4542
rect 11624 4146 11652 4626
rect 11716 4282 11744 5170
rect 11900 5030 11928 5170
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11888 4616 11940 4622
rect 11992 4604 12020 4966
rect 11940 4576 12020 4604
rect 11888 4558 11940 4564
rect 12176 4486 12204 5646
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12268 4826 12296 5102
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 11783 4380 12091 4389
rect 11783 4378 11789 4380
rect 11845 4378 11869 4380
rect 11925 4378 11949 4380
rect 12005 4378 12029 4380
rect 12085 4378 12091 4380
rect 11845 4326 11847 4378
rect 12027 4326 12029 4378
rect 11783 4324 11789 4326
rect 11845 4324 11869 4326
rect 11925 4324 11949 4326
rect 12005 4324 12029 4326
rect 12085 4324 12091 4326
rect 11783 4315 12091 4324
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 12268 4146 12296 4762
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 11150 3224 11206 3233
rect 11150 3159 11206 3168
rect 10690 1864 10746 1873
rect 10690 1799 10746 1808
rect 10598 1592 10654 1601
rect 10598 1527 10654 1536
rect 10612 1018 10640 1527
rect 10600 1012 10652 1018
rect 10600 954 10652 960
rect 8392 876 8444 882
rect 8392 818 8444 824
rect 10508 876 10560 882
rect 10508 818 10560 824
rect 11164 814 11192 3159
rect 11256 2990 11284 4082
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11900 3534 11928 4014
rect 12084 3942 12112 4082
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 12084 3602 12112 3878
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 12268 3534 12296 4082
rect 12728 4078 12756 7210
rect 12820 6798 12848 8774
rect 13096 8430 13124 8978
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 13188 7002 13216 7686
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12440 4004 12492 4010
rect 12440 3946 12492 3952
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 12072 3460 12124 3466
rect 12124 3420 12204 3448
rect 12072 3402 12124 3408
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11624 3074 11652 3334
rect 11716 3194 11744 3334
rect 11783 3292 12091 3301
rect 11783 3290 11789 3292
rect 11845 3290 11869 3292
rect 11925 3290 11949 3292
rect 12005 3290 12029 3292
rect 12085 3290 12091 3292
rect 11845 3238 11847 3290
rect 12027 3238 12029 3290
rect 11783 3236 11789 3238
rect 11845 3236 11869 3238
rect 11925 3236 11949 3238
rect 12005 3236 12029 3238
rect 12085 3236 12091 3238
rect 11783 3227 12091 3236
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 12176 3097 12204 3420
rect 12162 3088 12218 3097
rect 11624 3058 11836 3074
rect 11624 3052 11848 3058
rect 11624 3046 11796 3052
rect 12162 3023 12218 3032
rect 11796 2994 11848 3000
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11256 2514 11284 2926
rect 12268 2854 12296 3470
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 12256 2848 12308 2854
rect 12256 2790 12308 2796
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11244 2508 11296 2514
rect 11296 2468 11376 2496
rect 11244 2450 11296 2456
rect 11244 2032 11296 2038
rect 11242 2000 11244 2009
rect 11296 2000 11298 2009
rect 11242 1935 11298 1944
rect 11348 1902 11376 2468
rect 11336 1896 11388 1902
rect 11336 1838 11388 1844
rect 11532 1562 11560 2586
rect 11992 2446 12020 2790
rect 11796 2440 11848 2446
rect 11716 2400 11796 2428
rect 11612 1896 11664 1902
rect 11612 1838 11664 1844
rect 11520 1556 11572 1562
rect 11520 1498 11572 1504
rect 11334 1456 11390 1465
rect 11624 1426 11652 1838
rect 11716 1766 11744 2400
rect 11796 2382 11848 2388
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 12176 2310 12204 2382
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 11783 2204 12091 2213
rect 11783 2202 11789 2204
rect 11845 2202 11869 2204
rect 11925 2202 11949 2204
rect 12005 2202 12029 2204
rect 12085 2202 12091 2204
rect 11845 2150 11847 2202
rect 12027 2150 12029 2202
rect 11783 2148 11789 2150
rect 11845 2148 11869 2150
rect 11925 2148 11949 2150
rect 12005 2148 12029 2150
rect 12085 2148 12091 2150
rect 11783 2139 12091 2148
rect 11980 2100 12032 2106
rect 11980 2042 12032 2048
rect 11992 2009 12020 2042
rect 11978 2000 12034 2009
rect 11978 1935 12034 1944
rect 12452 1902 12480 3946
rect 13280 3602 13308 10134
rect 13556 10130 13584 10542
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13556 9586 13584 10066
rect 13726 10024 13782 10033
rect 13726 9959 13782 9968
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13556 8974 13584 9522
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13372 6662 13400 8774
rect 13556 8498 13584 8910
rect 13740 8838 13768 9959
rect 13832 9586 13860 10406
rect 13924 10062 13952 10406
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13924 9382 13952 9998
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13924 9042 13952 9318
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 14108 8974 14136 12804
rect 14384 12434 14412 12854
rect 14568 12850 14596 13670
rect 14462 12815 14518 12824
rect 14556 12844 14608 12850
rect 14292 12406 14412 12434
rect 14292 11762 14320 12406
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 14200 8498 14228 11018
rect 14384 10130 14412 12038
rect 14476 11082 14504 12815
rect 14556 12786 14608 12792
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14568 11694 14596 12582
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14660 11098 14688 18158
rect 14830 17776 14886 17785
rect 14830 17711 14832 17720
rect 14884 17711 14886 17720
rect 14832 17682 14884 17688
rect 14924 17672 14976 17678
rect 14924 17614 14976 17620
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14844 16998 14872 17070
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 14936 16697 14964 17614
rect 14922 16688 14978 16697
rect 14922 16623 14978 16632
rect 15028 16289 15056 19876
rect 15568 19858 15620 19864
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15106 19408 15162 19417
rect 15106 19343 15162 19352
rect 15120 19242 15148 19343
rect 15304 19281 15332 19654
rect 15948 19378 15976 20198
rect 16132 20058 16160 20431
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 16408 19990 16436 20878
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 16212 19984 16264 19990
rect 16040 19932 16212 19938
rect 16396 19984 16448 19990
rect 16040 19926 16264 19932
rect 16316 19944 16396 19972
rect 16040 19910 16252 19926
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 15290 19272 15346 19281
rect 15108 19236 15160 19242
rect 15290 19207 15346 19216
rect 15108 19178 15160 19184
rect 15382 19136 15438 19145
rect 15382 19071 15438 19080
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15108 18080 15160 18086
rect 15108 18022 15160 18028
rect 15014 16280 15070 16289
rect 14832 16244 14884 16250
rect 15014 16215 15070 16224
rect 14832 16186 14884 16192
rect 14738 15736 14794 15745
rect 14738 15671 14794 15680
rect 14752 12628 14780 15671
rect 14844 15570 14872 16186
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 14830 14920 14886 14929
rect 14830 14855 14886 14864
rect 14844 12730 14872 14855
rect 14936 14822 14964 15846
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14936 14657 14964 14758
rect 14922 14648 14978 14657
rect 14922 14583 14978 14592
rect 14936 13734 14964 14583
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 15028 14278 15056 14418
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14936 13326 14964 13670
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 14936 12850 14964 13262
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14844 12702 14964 12730
rect 14832 12640 14884 12646
rect 14752 12600 14832 12628
rect 14832 12582 14884 12588
rect 14936 12442 14964 12702
rect 14924 12436 14976 12442
rect 15120 12434 15148 18022
rect 15304 15910 15332 18906
rect 15396 18698 15424 19071
rect 15578 19068 15886 19077
rect 15578 19066 15584 19068
rect 15640 19066 15664 19068
rect 15720 19066 15744 19068
rect 15800 19066 15824 19068
rect 15880 19066 15886 19068
rect 15640 19014 15642 19066
rect 15822 19014 15824 19066
rect 15578 19012 15584 19014
rect 15640 19012 15664 19014
rect 15720 19012 15744 19014
rect 15800 19012 15824 19014
rect 15880 19012 15886 19014
rect 15578 19003 15886 19012
rect 15948 18952 15976 19314
rect 16040 19310 16068 19910
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 15856 18924 15976 18952
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15856 18290 15884 18924
rect 16040 18834 16068 19246
rect 16028 18828 16080 18834
rect 16028 18770 16080 18776
rect 16132 18748 16160 19790
rect 16316 19786 16344 19944
rect 16396 19926 16448 19932
rect 16304 19780 16356 19786
rect 16304 19722 16356 19728
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 16224 18970 16252 19246
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16316 18766 16344 19722
rect 16394 19272 16450 19281
rect 16394 19207 16450 19216
rect 16212 18760 16264 18766
rect 16132 18720 16212 18748
rect 16212 18702 16264 18708
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 15568 18080 15620 18086
rect 15488 18040 15568 18068
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15212 13870 15240 14894
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15304 12730 15332 14894
rect 15396 14550 15424 15098
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15488 13512 15516 18040
rect 15568 18022 15620 18028
rect 15578 17980 15886 17989
rect 15578 17978 15584 17980
rect 15640 17978 15664 17980
rect 15720 17978 15744 17980
rect 15800 17978 15824 17980
rect 15880 17978 15886 17980
rect 15640 17926 15642 17978
rect 15822 17926 15824 17978
rect 15578 17924 15584 17926
rect 15640 17924 15664 17926
rect 15720 17924 15744 17926
rect 15800 17924 15824 17926
rect 15880 17924 15886 17926
rect 15578 17915 15886 17924
rect 16040 17882 16068 18226
rect 16224 18086 16252 18702
rect 16408 18222 16436 19207
rect 16500 18290 16528 20742
rect 17960 20324 18012 20330
rect 17960 20266 18012 20272
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 16868 19854 16896 20198
rect 16856 19848 16908 19854
rect 16856 19790 16908 19796
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 16868 19310 16896 19790
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16868 18766 16896 19246
rect 16856 18760 16908 18766
rect 16856 18702 16908 18708
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16028 17876 16080 17882
rect 16028 17818 16080 17824
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 15578 16892 15886 16901
rect 15578 16890 15584 16892
rect 15640 16890 15664 16892
rect 15720 16890 15744 16892
rect 15800 16890 15824 16892
rect 15880 16890 15886 16892
rect 15640 16838 15642 16890
rect 15822 16838 15824 16890
rect 15578 16836 15584 16838
rect 15640 16836 15664 16838
rect 15720 16836 15744 16838
rect 15800 16836 15824 16838
rect 15880 16836 15886 16838
rect 15578 16827 15886 16836
rect 15578 15804 15886 15813
rect 15578 15802 15584 15804
rect 15640 15802 15664 15804
rect 15720 15802 15744 15804
rect 15800 15802 15824 15804
rect 15880 15802 15886 15804
rect 15640 15750 15642 15802
rect 15822 15750 15824 15802
rect 15578 15748 15584 15750
rect 15640 15748 15664 15750
rect 15720 15748 15744 15750
rect 15800 15748 15824 15750
rect 15880 15748 15886 15750
rect 15578 15739 15886 15748
rect 15948 15706 15976 17070
rect 16316 16658 16344 17478
rect 16408 16794 16436 17682
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16500 17134 16528 17614
rect 16776 17610 16804 17818
rect 16868 17814 16896 18702
rect 17236 18426 17264 19790
rect 17512 18834 17540 20198
rect 17972 19922 18000 20266
rect 18050 19952 18106 19961
rect 17960 19916 18012 19922
rect 18050 19887 18106 19896
rect 17960 19858 18012 19864
rect 18064 19514 18092 19887
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 18156 19394 18184 20946
rect 18326 19544 18382 19553
rect 18326 19479 18382 19488
rect 18064 19366 18184 19394
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 16856 17808 16908 17814
rect 16856 17750 16908 17756
rect 17512 17678 17540 18362
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 16764 17604 16816 17610
rect 16764 17546 16816 17552
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 17040 17128 17092 17134
rect 17328 17116 17356 17614
rect 17092 17088 17356 17116
rect 17040 17070 17092 17076
rect 16396 16788 16448 16794
rect 16396 16730 16448 16736
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 16132 16114 16160 16390
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16500 16046 16528 17070
rect 16672 16992 16724 16998
rect 16578 16960 16634 16969
rect 16672 16934 16724 16940
rect 16578 16895 16634 16904
rect 16592 16794 16620 16895
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16488 16040 16540 16046
rect 16210 16008 16266 16017
rect 16578 16008 16634 16017
rect 16540 15988 16578 15994
rect 16488 15982 16578 15988
rect 16210 15943 16266 15952
rect 16500 15966 16578 15982
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 16118 15464 16174 15473
rect 16118 15399 16120 15408
rect 16172 15399 16174 15408
rect 16120 15370 16172 15376
rect 16224 15162 16252 15943
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16408 15502 16436 15642
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 16118 14920 16174 14929
rect 16118 14855 16174 14864
rect 15578 14716 15886 14725
rect 15578 14714 15584 14716
rect 15640 14714 15664 14716
rect 15720 14714 15744 14716
rect 15800 14714 15824 14716
rect 15880 14714 15886 14716
rect 15640 14662 15642 14714
rect 15822 14662 15824 14714
rect 15578 14660 15584 14662
rect 15640 14660 15664 14662
rect 15720 14660 15744 14662
rect 15800 14660 15824 14662
rect 15880 14660 15886 14662
rect 15578 14651 15886 14660
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 15578 13628 15886 13637
rect 15578 13626 15584 13628
rect 15640 13626 15664 13628
rect 15720 13626 15744 13628
rect 15800 13626 15824 13628
rect 15880 13626 15886 13628
rect 15640 13574 15642 13626
rect 15822 13574 15824 13626
rect 15578 13572 15584 13574
rect 15640 13572 15664 13574
rect 15720 13572 15744 13574
rect 15800 13572 15824 13574
rect 15880 13572 15886 13574
rect 15578 13563 15886 13572
rect 15488 13484 15608 13512
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15304 12702 15424 12730
rect 15396 12442 15424 12702
rect 14924 12378 14976 12384
rect 15028 12406 15148 12434
rect 15292 12436 15344 12442
rect 15028 12186 15056 12406
rect 15292 12378 15344 12384
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15304 12345 15332 12378
rect 15290 12336 15346 12345
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15200 12300 15252 12306
rect 15290 12271 15346 12280
rect 15200 12242 15252 12248
rect 14844 12158 15056 12186
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 11354 14780 12038
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14464 11076 14516 11082
rect 14660 11070 14780 11098
rect 14464 11018 14516 11024
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14660 10674 14688 10950
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14752 9178 14780 11070
rect 14740 9172 14792 9178
rect 14740 9114 14792 9120
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 8090 13860 8230
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 14096 8084 14148 8090
rect 14096 8026 14148 8032
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 13464 7993 13492 8026
rect 13450 7984 13506 7993
rect 13450 7919 13506 7928
rect 13820 7880 13872 7886
rect 13820 7822 13872 7828
rect 13832 7410 13860 7822
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 13726 6896 13782 6905
rect 13544 6860 13596 6866
rect 13726 6831 13728 6840
rect 13544 6802 13596 6808
rect 13780 6831 13782 6840
rect 13728 6802 13780 6808
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13372 6254 13400 6598
rect 13360 6248 13412 6254
rect 13556 6225 13584 6802
rect 13832 6798 13860 7346
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13360 6190 13412 6196
rect 13542 6216 13598 6225
rect 13542 6151 13598 6160
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13544 6112 13596 6118
rect 13544 6054 13596 6060
rect 13358 5944 13414 5953
rect 13464 5914 13492 6054
rect 13358 5879 13414 5888
rect 13452 5908 13504 5914
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12544 3398 12572 3470
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 11980 1896 12032 1902
rect 12440 1896 12492 1902
rect 11980 1838 12032 1844
rect 12346 1864 12402 1873
rect 11704 1760 11756 1766
rect 11704 1702 11756 1708
rect 11716 1562 11744 1702
rect 11992 1601 12020 1838
rect 12440 1838 12492 1844
rect 12346 1799 12402 1808
rect 11978 1592 12034 1601
rect 11704 1556 11756 1562
rect 12256 1556 12308 1562
rect 11978 1527 12034 1536
rect 11704 1498 11756 1504
rect 12084 1516 12256 1544
rect 11334 1391 11390 1400
rect 11612 1420 11664 1426
rect 9036 808 9088 814
rect 9036 750 9088 756
rect 11152 808 11204 814
rect 11152 750 11204 756
rect 8300 672 8352 678
rect 8300 614 8352 620
rect 7988 572 8296 581
rect 7988 570 7994 572
rect 8050 570 8074 572
rect 8130 570 8154 572
rect 8210 570 8234 572
rect 8290 570 8296 572
rect 8050 518 8052 570
rect 8232 518 8234 570
rect 7988 516 7994 518
rect 8050 516 8074 518
rect 8130 516 8154 518
rect 8210 516 8234 518
rect 8290 516 8296 518
rect 7988 507 8296 516
rect 6920 468 6972 474
rect 6920 410 6972 416
rect 7564 468 7616 474
rect 7564 410 7616 416
rect 7840 468 7892 474
rect 7840 410 7892 416
rect 6932 377 6960 410
rect 6918 368 6974 377
rect 6918 303 6974 312
rect 9048 270 9076 750
rect 11348 678 11376 1391
rect 11888 1420 11940 1426
rect 11612 1362 11664 1368
rect 11716 1380 11888 1408
rect 11716 1000 11744 1380
rect 11888 1362 11940 1368
rect 12084 1222 12112 1516
rect 12256 1498 12308 1504
rect 12072 1216 12124 1222
rect 12072 1158 12124 1164
rect 12164 1216 12216 1222
rect 12360 1170 12388 1799
rect 12164 1158 12216 1164
rect 11783 1116 12091 1125
rect 11783 1114 11789 1116
rect 11845 1114 11869 1116
rect 11925 1114 11949 1116
rect 12005 1114 12029 1116
rect 12085 1114 12091 1116
rect 11845 1062 11847 1114
rect 12027 1062 12029 1114
rect 11783 1060 11789 1062
rect 11845 1060 11869 1062
rect 11925 1060 11949 1062
rect 12005 1060 12029 1062
rect 12085 1060 12091 1062
rect 11783 1051 12091 1060
rect 12176 1018 12204 1158
rect 12268 1142 12388 1170
rect 11532 972 11744 1000
rect 12164 1012 12216 1018
rect 9128 672 9180 678
rect 9128 614 9180 620
rect 11336 672 11388 678
rect 11336 614 11388 620
rect 9036 264 9088 270
rect 6000 206 6052 212
rect 6274 232 6330 241
rect 9036 206 9088 212
rect 6274 167 6330 176
rect 9140 134 9168 614
rect 11532 338 11560 972
rect 12164 954 12216 960
rect 12070 912 12126 921
rect 11612 876 11664 882
rect 12070 847 12072 856
rect 11612 818 11664 824
rect 12124 847 12126 856
rect 12072 818 12124 824
rect 11624 338 11652 818
rect 12268 814 12296 1142
rect 13372 1018 13400 5879
rect 13452 5850 13504 5856
rect 13556 4690 13584 6054
rect 13648 5273 13676 6122
rect 13740 5817 13768 6598
rect 13832 6322 13860 6734
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 14016 6202 14044 7346
rect 14108 7206 14136 8026
rect 14568 7954 14596 8026
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14462 7576 14518 7585
rect 14292 7534 14462 7562
rect 14292 7342 14320 7534
rect 14462 7511 14518 7520
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14096 7200 14148 7206
rect 14292 7177 14320 7278
rect 14740 7200 14792 7206
rect 14096 7142 14148 7148
rect 14278 7168 14334 7177
rect 14108 7002 14136 7142
rect 14740 7142 14792 7148
rect 14278 7103 14334 7112
rect 14646 7032 14702 7041
rect 14096 6996 14148 7002
rect 14646 6967 14648 6976
rect 14096 6938 14148 6944
rect 14700 6967 14702 6976
rect 14648 6938 14700 6944
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14476 6662 14504 6734
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14096 6248 14148 6254
rect 13924 6196 14096 6202
rect 13924 6190 14148 6196
rect 13924 6174 14136 6190
rect 13726 5808 13782 5817
rect 13726 5743 13782 5752
rect 13924 5658 13952 6174
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5778 14504 6054
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 13740 5642 13952 5658
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14280 5704 14332 5710
rect 14332 5664 14412 5692
rect 14280 5646 14332 5652
rect 13728 5636 13952 5642
rect 13780 5630 13952 5636
rect 13728 5578 13780 5584
rect 13912 5296 13964 5302
rect 13634 5264 13690 5273
rect 13912 5238 13964 5244
rect 13634 5199 13690 5208
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13740 4758 13768 4966
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13832 4486 13860 5034
rect 13924 5030 13952 5238
rect 14016 5166 14044 5646
rect 14200 5234 14228 5646
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 14016 4622 14044 5102
rect 14096 5092 14148 5098
rect 14096 5034 14148 5040
rect 14108 4826 14136 5034
rect 14200 4826 14228 5170
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13910 4312 13966 4321
rect 13910 4247 13966 4256
rect 13924 4078 13952 4247
rect 14016 4078 14044 4558
rect 13912 4072 13964 4078
rect 13726 4040 13782 4049
rect 13912 4014 13964 4020
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 13726 3975 13782 3984
rect 13740 3942 13768 3975
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 14016 3618 14044 4014
rect 14200 3924 14228 4762
rect 14292 4622 14320 5510
rect 14384 5370 14412 5664
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14568 5234 14596 6394
rect 14752 6322 14780 7142
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14280 3936 14332 3942
rect 14200 3896 14280 3924
rect 14016 3590 14136 3618
rect 14108 3466 14136 3590
rect 14096 3460 14148 3466
rect 14096 3402 14148 3408
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 2990 13676 3334
rect 14108 2990 14136 3402
rect 14200 2990 14228 3896
rect 14280 3878 14332 3884
rect 14476 3738 14504 4082
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14648 3392 14700 3398
rect 14476 3352 14648 3380
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 14108 2774 14136 2926
rect 14016 2746 14136 2774
rect 14016 2446 14044 2746
rect 14200 2446 14228 2926
rect 14004 2440 14056 2446
rect 13924 2400 14004 2428
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13556 2106 13584 2246
rect 13544 2100 13596 2106
rect 13544 2042 13596 2048
rect 13924 1902 13952 2400
rect 14004 2382 14056 2388
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 13912 1896 13964 1902
rect 13912 1838 13964 1844
rect 13544 1828 13596 1834
rect 13544 1770 13596 1776
rect 13556 1018 13584 1770
rect 13820 1352 13872 1358
rect 13924 1340 13952 1838
rect 14200 1766 14228 2382
rect 14188 1760 14240 1766
rect 14188 1702 14240 1708
rect 14200 1358 14228 1702
rect 14372 1556 14424 1562
rect 14372 1498 14424 1504
rect 14384 1358 14412 1498
rect 13872 1312 13952 1340
rect 14188 1352 14240 1358
rect 13820 1294 13872 1300
rect 14188 1294 14240 1300
rect 14372 1352 14424 1358
rect 14372 1294 14424 1300
rect 12348 1012 12400 1018
rect 12348 954 12400 960
rect 13360 1012 13412 1018
rect 13360 954 13412 960
rect 13544 1012 13596 1018
rect 13544 954 13596 960
rect 11888 808 11940 814
rect 12256 808 12308 814
rect 11940 756 12020 762
rect 11888 750 12020 756
rect 12256 750 12308 756
rect 11900 734 12020 750
rect 11992 490 12020 734
rect 12072 672 12124 678
rect 12256 672 12308 678
rect 12124 649 12204 660
rect 12124 640 12218 649
rect 12124 632 12162 640
rect 12072 614 12124 620
rect 12256 614 12308 620
rect 12162 575 12218 584
rect 12268 490 12296 614
rect 11992 462 12296 490
rect 11520 332 11572 338
rect 11520 274 11572 280
rect 11612 332 11664 338
rect 11612 274 11664 280
rect 12360 270 12388 954
rect 14476 898 14504 3352
rect 14648 3334 14700 3340
rect 14752 3194 14780 4014
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14844 3074 14872 12158
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 15028 11937 15056 12038
rect 15014 11928 15070 11937
rect 15014 11863 15070 11872
rect 15120 11830 15148 12242
rect 15108 11824 15160 11830
rect 15108 11766 15160 11772
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14936 9042 14964 11018
rect 15028 9586 15056 11494
rect 15120 11354 15148 11630
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 15028 6322 15056 9318
rect 15120 7546 15148 11290
rect 15212 10810 15240 12242
rect 15488 11370 15516 13330
rect 15580 12730 15608 13484
rect 16040 13394 16068 14214
rect 16132 13394 16160 14855
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16408 14618 16436 14758
rect 16500 14618 16528 15966
rect 16578 15943 16634 15952
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 15752 13388 15804 13394
rect 16028 13388 16080 13394
rect 15804 13348 15884 13376
rect 15752 13330 15804 13336
rect 15856 13190 15884 13348
rect 16028 13330 16080 13336
rect 16120 13388 16172 13394
rect 16172 13348 16252 13376
rect 16120 13330 16172 13336
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15764 12850 15792 13126
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15580 12702 15976 12730
rect 15578 12540 15886 12549
rect 15578 12538 15584 12540
rect 15640 12538 15664 12540
rect 15720 12538 15744 12540
rect 15800 12538 15824 12540
rect 15880 12538 15886 12540
rect 15640 12486 15642 12538
rect 15822 12486 15824 12538
rect 15578 12484 15584 12486
rect 15640 12484 15664 12486
rect 15720 12484 15744 12486
rect 15800 12484 15824 12486
rect 15880 12484 15886 12486
rect 15578 12475 15886 12484
rect 15566 12200 15622 12209
rect 15566 12135 15568 12144
rect 15620 12135 15622 12144
rect 15568 12106 15620 12112
rect 15578 11452 15886 11461
rect 15578 11450 15584 11452
rect 15640 11450 15664 11452
rect 15720 11450 15744 11452
rect 15800 11450 15824 11452
rect 15880 11450 15886 11452
rect 15640 11398 15642 11450
rect 15822 11398 15824 11450
rect 15578 11396 15584 11398
rect 15640 11396 15664 11398
rect 15720 11396 15744 11398
rect 15800 11396 15824 11398
rect 15880 11396 15886 11398
rect 15578 11387 15886 11396
rect 15396 11342 15516 11370
rect 15396 11286 15424 11342
rect 15384 11280 15436 11286
rect 15384 11222 15436 11228
rect 15474 11248 15530 11257
rect 15474 11183 15476 11192
rect 15528 11183 15530 11192
rect 15476 11154 15528 11160
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15212 10130 15240 10542
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15212 9110 15240 10066
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15212 7410 15240 8774
rect 15304 7886 15332 9862
rect 15396 8378 15424 10406
rect 15578 10364 15886 10373
rect 15578 10362 15584 10364
rect 15640 10362 15664 10364
rect 15720 10362 15744 10364
rect 15800 10362 15824 10364
rect 15880 10362 15886 10364
rect 15640 10310 15642 10362
rect 15822 10310 15824 10362
rect 15578 10308 15584 10310
rect 15640 10308 15664 10310
rect 15720 10308 15744 10310
rect 15800 10308 15824 10310
rect 15880 10308 15886 10310
rect 15578 10299 15886 10308
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15488 8498 15516 9862
rect 15578 9276 15886 9285
rect 15578 9274 15584 9276
rect 15640 9274 15664 9276
rect 15720 9274 15744 9276
rect 15800 9274 15824 9276
rect 15880 9274 15886 9276
rect 15640 9222 15642 9274
rect 15822 9222 15824 9274
rect 15578 9220 15584 9222
rect 15640 9220 15664 9222
rect 15720 9220 15744 9222
rect 15800 9220 15824 9222
rect 15880 9220 15886 9222
rect 15578 9211 15886 9220
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15580 8430 15608 9046
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15568 8424 15620 8430
rect 15396 8350 15516 8378
rect 15568 8366 15620 8372
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 15212 5681 15240 7142
rect 15304 6361 15332 7686
rect 15488 6730 15516 8350
rect 15856 8294 15884 8910
rect 15948 8537 15976 12702
rect 16224 12322 16252 13348
rect 16316 12782 16344 14350
rect 16500 14278 16528 14554
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16500 13870 16528 14214
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16592 13530 16620 15506
rect 16684 14618 16712 16934
rect 16776 15910 16804 17070
rect 17040 16992 17092 16998
rect 16868 16952 17040 16980
rect 16868 16658 16896 16952
rect 17040 16934 17092 16940
rect 16946 16824 17002 16833
rect 17328 16794 17356 17088
rect 17788 16810 17816 19178
rect 18064 18970 18092 19366
rect 18340 19310 18368 19479
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 18064 18222 18092 18906
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 18156 18222 18184 18702
rect 18248 18358 18276 19246
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18340 18601 18368 19110
rect 18326 18592 18382 18601
rect 18326 18527 18382 18536
rect 18236 18352 18288 18358
rect 18236 18294 18288 18300
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 17866 17232 17922 17241
rect 17866 17167 17868 17176
rect 17920 17167 17922 17176
rect 17868 17138 17920 17144
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 17866 16824 17922 16833
rect 16946 16759 17002 16768
rect 17316 16788 17368 16794
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 16960 15586 16988 16759
rect 17788 16782 17866 16810
rect 18156 16794 18184 17070
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 17866 16759 17922 16768
rect 18144 16788 18196 16794
rect 17316 16730 17368 16736
rect 18144 16730 18196 16736
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17866 16552 17922 16561
rect 17132 16448 17184 16454
rect 17132 16390 17184 16396
rect 17144 15910 17172 16390
rect 17236 16046 17264 16526
rect 17866 16487 17922 16496
rect 17880 16114 17908 16487
rect 18248 16250 18276 16934
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17224 16040 17276 16046
rect 17222 16008 17224 16017
rect 17276 16008 17278 16017
rect 17222 15943 17278 15952
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17052 15638 17080 15846
rect 16776 15558 16988 15586
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16580 13524 16632 13530
rect 16776 13512 16804 15558
rect 16854 15464 16910 15473
rect 16854 15399 16856 15408
rect 16908 15399 16910 15408
rect 16856 15370 16908 15376
rect 16580 13466 16632 13472
rect 16684 13484 16804 13512
rect 16408 13258 16436 13466
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16304 12776 16356 12782
rect 16302 12744 16304 12753
rect 16356 12744 16358 12753
rect 16302 12679 16358 12688
rect 16028 12300 16080 12306
rect 16224 12294 16344 12322
rect 16408 12306 16436 13194
rect 16028 12242 16080 12248
rect 16040 11898 16068 12242
rect 16210 12064 16266 12073
rect 16316 12050 16344 12294
rect 16396 12300 16448 12306
rect 16396 12242 16448 12248
rect 16396 12164 16448 12170
rect 16396 12106 16448 12112
rect 16266 12022 16344 12050
rect 16210 11999 16266 12008
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16132 11354 16160 11494
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 15934 8528 15990 8537
rect 15934 8463 15990 8472
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15578 8188 15886 8197
rect 15578 8186 15584 8188
rect 15640 8186 15664 8188
rect 15720 8186 15744 8188
rect 15800 8186 15824 8188
rect 15880 8186 15886 8188
rect 15640 8134 15642 8186
rect 15822 8134 15824 8186
rect 15578 8132 15584 8134
rect 15640 8132 15664 8134
rect 15720 8132 15744 8134
rect 15800 8132 15824 8134
rect 15880 8132 15886 8134
rect 15578 8123 15886 8132
rect 16040 8022 16068 11154
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 16132 9217 16160 9318
rect 16118 9208 16174 9217
rect 16118 9143 16174 9152
rect 16224 8922 16252 11999
rect 16304 11824 16356 11830
rect 16408 11812 16436 12106
rect 16356 11784 16436 11812
rect 16304 11766 16356 11772
rect 16316 11354 16344 11766
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16396 10804 16448 10810
rect 16500 10792 16528 13330
rect 16592 12102 16620 13466
rect 16684 13190 16712 13484
rect 16762 13424 16818 13433
rect 16762 13359 16818 13368
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16776 12986 16804 13359
rect 16868 13138 16896 15370
rect 17052 14618 17080 15574
rect 17236 15502 17264 15943
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17144 15026 17172 15098
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17040 14612 17092 14618
rect 17092 14572 17172 14600
rect 17040 14554 17092 14560
rect 16946 14104 17002 14113
rect 16946 14039 17002 14048
rect 16960 13938 16988 14039
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17052 13394 17080 13806
rect 17144 13734 17172 14572
rect 17420 14414 17448 15302
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17144 13530 17172 13670
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 17408 13388 17460 13394
rect 17604 13376 17632 14894
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 17972 14618 18000 14826
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 18340 14482 18368 17818
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18156 14113 18184 14214
rect 18142 14104 18198 14113
rect 18142 14039 18198 14048
rect 17682 13968 17738 13977
rect 17682 13903 17738 13912
rect 17696 13530 17724 13903
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17460 13348 17632 13376
rect 17408 13330 17460 13336
rect 16946 13288 17002 13297
rect 17002 13246 17080 13274
rect 16946 13223 17002 13232
rect 16868 13110 16988 13138
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16868 12866 16896 12922
rect 16776 12838 16896 12866
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16776 11762 16804 12838
rect 16960 12646 16988 13110
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 17052 12442 17080 13246
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17604 12306 17632 13348
rect 17972 13297 18000 13806
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 17958 13288 18014 13297
rect 17958 13223 18014 13232
rect 18248 12850 18276 13670
rect 18524 13462 18552 20975
rect 18800 20466 18828 21558
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19800 21480 19852 21486
rect 19800 21422 19852 21428
rect 19156 21344 19208 21350
rect 19156 21286 19208 21292
rect 19062 20904 19118 20913
rect 18892 20862 19062 20890
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18708 18766 18736 19790
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18708 17746 18736 18702
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18694 17640 18750 17649
rect 18694 17575 18750 17584
rect 18708 17202 18736 17575
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18800 15706 18828 17478
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18892 15450 18920 20862
rect 19062 20839 19118 20848
rect 19168 18154 19196 21286
rect 19248 21072 19300 21078
rect 19246 21040 19248 21049
rect 19300 21040 19302 21049
rect 19246 20975 19302 20984
rect 19352 20788 19380 21422
rect 19444 21146 19472 21422
rect 19432 21140 19484 21146
rect 19432 21082 19484 21088
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19260 20760 19380 20788
rect 19260 20602 19288 20760
rect 19373 20700 19681 20709
rect 19373 20698 19379 20700
rect 19435 20698 19459 20700
rect 19515 20698 19539 20700
rect 19595 20698 19619 20700
rect 19675 20698 19681 20700
rect 19435 20646 19437 20698
rect 19617 20646 19619 20698
rect 19373 20644 19379 20646
rect 19435 20644 19459 20646
rect 19515 20644 19539 20646
rect 19595 20644 19619 20646
rect 19675 20644 19681 20646
rect 19373 20635 19681 20644
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19720 20466 19748 20878
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 19524 20324 19576 20330
rect 19524 20266 19576 20272
rect 19536 19802 19564 20266
rect 19812 20058 19840 21422
rect 19800 20052 19852 20058
rect 19800 19994 19852 20000
rect 19536 19774 19748 19802
rect 19904 19786 19932 21626
rect 20996 21344 21048 21350
rect 20996 21286 21048 21292
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 19373 19612 19681 19621
rect 19373 19610 19379 19612
rect 19435 19610 19459 19612
rect 19515 19610 19539 19612
rect 19595 19610 19619 19612
rect 19675 19610 19681 19612
rect 19435 19558 19437 19610
rect 19617 19558 19619 19610
rect 19373 19556 19379 19558
rect 19435 19556 19459 19558
rect 19515 19556 19539 19558
rect 19595 19556 19619 19558
rect 19675 19556 19681 19558
rect 19373 19547 19681 19556
rect 19373 18524 19681 18533
rect 19373 18522 19379 18524
rect 19435 18522 19459 18524
rect 19515 18522 19539 18524
rect 19595 18522 19619 18524
rect 19675 18522 19681 18524
rect 19435 18470 19437 18522
rect 19617 18470 19619 18522
rect 19373 18468 19379 18470
rect 19435 18468 19459 18470
rect 19515 18468 19539 18470
rect 19595 18468 19619 18470
rect 19675 18468 19681 18470
rect 19373 18459 19681 18468
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18984 17338 19012 17478
rect 19373 17436 19681 17445
rect 19373 17434 19379 17436
rect 19435 17434 19459 17436
rect 19515 17434 19539 17436
rect 19595 17434 19619 17436
rect 19675 17434 19681 17436
rect 19435 17382 19437 17434
rect 19617 17382 19619 17434
rect 19373 17380 19379 17382
rect 19435 17380 19459 17382
rect 19515 17380 19539 17382
rect 19595 17380 19619 17382
rect 19675 17380 19681 17382
rect 19373 17371 19681 17380
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 19720 17270 19748 19774
rect 19892 19780 19944 19786
rect 19892 19722 19944 19728
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19064 17264 19116 17270
rect 19064 17206 19116 17212
rect 19524 17264 19576 17270
rect 19524 17206 19576 17212
rect 19708 17264 19760 17270
rect 19708 17206 19760 17212
rect 19076 16726 19104 17206
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19064 16720 19116 16726
rect 19064 16662 19116 16668
rect 19352 16658 19380 17070
rect 19536 16697 19564 17206
rect 19522 16688 19578 16697
rect 19340 16652 19392 16658
rect 19812 16658 19840 18566
rect 19904 18358 19932 19722
rect 19996 18902 20024 21082
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20548 20058 20576 20742
rect 20732 20398 20760 20946
rect 21008 20806 21036 21286
rect 20996 20800 21048 20806
rect 20902 20768 20958 20777
rect 20996 20742 21048 20748
rect 20902 20703 20958 20712
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20628 19916 20680 19922
rect 20628 19858 20680 19864
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 19892 18352 19944 18358
rect 19892 18294 19944 18300
rect 19892 18148 19944 18154
rect 19892 18090 19944 18096
rect 19904 17746 19932 18090
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 19890 17504 19946 17513
rect 19890 17439 19946 17448
rect 19904 17066 19932 17439
rect 19996 17354 20024 18838
rect 20088 18154 20116 19110
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 18222 20300 18566
rect 20640 18290 20668 19858
rect 20732 19854 20760 20334
rect 20916 19922 20944 20703
rect 21100 20058 21128 21626
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 21284 21146 21312 21422
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21284 20398 21312 20878
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 21376 19718 21404 21830
rect 21652 21622 21680 22199
rect 23572 22238 23624 22244
rect 25964 22296 26016 22302
rect 25964 22238 26016 22244
rect 22466 22199 22468 22208
rect 22376 22170 22428 22176
rect 22520 22199 22522 22208
rect 22468 22170 22520 22176
rect 22282 21992 22338 22001
rect 22282 21927 22338 21936
rect 22296 21894 22324 21927
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 21640 21616 21692 21622
rect 22008 21616 22060 21622
rect 21640 21558 21692 21564
rect 22006 21584 22008 21593
rect 22060 21584 22062 21593
rect 21548 21548 21600 21554
rect 22006 21519 22062 21528
rect 21548 21490 21600 21496
rect 21456 21480 21508 21486
rect 21456 21422 21508 21428
rect 21468 20058 21496 21422
rect 21560 20262 21588 21490
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 21916 20800 21968 20806
rect 21916 20742 21968 20748
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 21560 19922 21588 19994
rect 21548 19916 21600 19922
rect 21548 19858 21600 19864
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21454 19544 21510 19553
rect 21454 19479 21510 19488
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 20824 18873 20852 19110
rect 20810 18864 20866 18873
rect 20810 18799 20866 18808
rect 21100 18737 21128 19110
rect 21086 18728 21142 18737
rect 21086 18663 21142 18672
rect 20628 18284 20680 18290
rect 20628 18226 20680 18232
rect 20260 18216 20312 18222
rect 20996 18216 21048 18222
rect 20260 18158 20312 18164
rect 20916 18176 20996 18204
rect 20076 18148 20128 18154
rect 20076 18090 20128 18096
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 20364 17746 20392 18022
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 19996 17326 20116 17354
rect 19892 17060 19944 17066
rect 19892 17002 19944 17008
rect 19984 17060 20036 17066
rect 19984 17002 20036 17008
rect 19904 16969 19932 17002
rect 19890 16960 19946 16969
rect 19890 16895 19946 16904
rect 19522 16623 19578 16632
rect 19800 16652 19852 16658
rect 19340 16594 19392 16600
rect 19800 16594 19852 16600
rect 19708 16448 19760 16454
rect 19708 16390 19760 16396
rect 19373 16348 19681 16357
rect 19373 16346 19379 16348
rect 19435 16346 19459 16348
rect 19515 16346 19539 16348
rect 19595 16346 19619 16348
rect 19675 16346 19681 16348
rect 19435 16294 19437 16346
rect 19617 16294 19619 16346
rect 19373 16292 19379 16294
rect 19435 16292 19459 16294
rect 19515 16292 19539 16294
rect 19595 16292 19619 16294
rect 19675 16292 19681 16294
rect 19373 16283 19681 16292
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 19248 15904 19300 15910
rect 19248 15846 19300 15852
rect 18800 15422 18920 15450
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18800 14958 18828 15422
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18788 14816 18840 14822
rect 18788 14758 18840 14764
rect 18800 14618 18828 14758
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18892 14074 18920 15302
rect 18984 14074 19012 15438
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18878 13968 18934 13977
rect 18878 13903 18934 13912
rect 18892 13870 18920 13903
rect 19168 13870 19196 14758
rect 19260 14521 19288 15846
rect 19444 15348 19472 15982
rect 19720 15586 19748 16390
rect 19800 16244 19852 16250
rect 19800 16186 19852 16192
rect 19628 15558 19748 15586
rect 19628 15502 19656 15558
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19444 15320 19748 15348
rect 19373 15260 19681 15269
rect 19373 15258 19379 15260
rect 19435 15258 19459 15260
rect 19515 15258 19539 15260
rect 19595 15258 19619 15260
rect 19675 15258 19681 15260
rect 19435 15206 19437 15258
rect 19617 15206 19619 15258
rect 19373 15204 19379 15206
rect 19435 15204 19459 15206
rect 19515 15204 19539 15206
rect 19595 15204 19619 15206
rect 19675 15204 19681 15206
rect 19373 15195 19681 15204
rect 19720 15144 19748 15320
rect 19628 15116 19748 15144
rect 19432 15088 19484 15094
rect 19432 15030 19484 15036
rect 19246 14512 19302 14521
rect 19444 14482 19472 15030
rect 19246 14447 19302 14456
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19444 14362 19472 14418
rect 19522 14376 19578 14385
rect 19260 14334 19380 14362
rect 19444 14334 19522 14362
rect 19260 13988 19288 14334
rect 19352 14260 19380 14334
rect 19522 14311 19578 14320
rect 19628 14260 19656 15116
rect 19708 14952 19760 14958
rect 19812 14940 19840 16186
rect 19996 16114 20024 17002
rect 20088 16454 20116 17326
rect 20364 17134 20392 17682
rect 20442 17640 20498 17649
rect 20442 17575 20498 17584
rect 20626 17640 20682 17649
rect 20626 17575 20682 17584
rect 20260 17128 20312 17134
rect 20260 17070 20312 17076
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20272 16969 20300 17070
rect 20258 16960 20314 16969
rect 20258 16895 20314 16904
rect 20364 16590 20392 17070
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 20364 16250 20392 16526
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20272 15162 20300 15982
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 20364 15706 20392 15846
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20364 15042 20392 15098
rect 19996 15026 20392 15042
rect 19984 15020 20392 15026
rect 20036 15014 20392 15020
rect 19984 14962 20036 14968
rect 19760 14912 19840 14940
rect 20352 14952 20404 14958
rect 19708 14894 19760 14900
rect 20352 14894 20404 14900
rect 19352 14232 19656 14260
rect 19373 14172 19681 14181
rect 19373 14170 19379 14172
rect 19435 14170 19459 14172
rect 19515 14170 19539 14172
rect 19595 14170 19619 14172
rect 19675 14170 19681 14172
rect 19435 14118 19437 14170
rect 19617 14118 19619 14170
rect 19373 14116 19379 14118
rect 19435 14116 19459 14118
rect 19515 14116 19539 14118
rect 19595 14116 19619 14118
rect 19675 14116 19681 14118
rect 19373 14107 19681 14116
rect 20364 14074 20392 14894
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 19260 13960 19380 13988
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 19156 13864 19208 13870
rect 19156 13806 19208 13812
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 18512 13456 18564 13462
rect 18512 13398 18564 13404
rect 18708 13394 18736 13670
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 18328 12708 18380 12714
rect 18328 12650 18380 12656
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17052 11762 17080 12038
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16684 11150 16712 11630
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16448 10764 16528 10792
rect 16396 10746 16448 10752
rect 16408 10198 16436 10746
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 16408 9897 16436 10134
rect 16394 9888 16450 9897
rect 16394 9823 16450 9832
rect 16500 9674 16528 10202
rect 16408 9646 16528 9674
rect 16408 9568 16436 9646
rect 16408 9540 16528 9568
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 9081 16344 9318
rect 16302 9072 16358 9081
rect 16302 9007 16358 9016
rect 16500 8974 16528 9540
rect 16488 8968 16540 8974
rect 16224 8894 16436 8922
rect 16488 8910 16540 8916
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16132 8090 16160 8774
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16224 8090 16252 8230
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16028 8016 16080 8022
rect 15934 7984 15990 7993
rect 16028 7958 16080 7964
rect 16408 7954 16436 8894
rect 15934 7919 15990 7928
rect 16396 7948 16448 7954
rect 15578 7100 15886 7109
rect 15578 7098 15584 7100
rect 15640 7098 15664 7100
rect 15720 7098 15744 7100
rect 15800 7098 15824 7100
rect 15880 7098 15886 7100
rect 15640 7046 15642 7098
rect 15822 7046 15824 7098
rect 15578 7044 15584 7046
rect 15640 7044 15664 7046
rect 15720 7044 15744 7046
rect 15800 7044 15824 7046
rect 15880 7044 15886 7046
rect 15578 7035 15886 7044
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15290 6352 15346 6361
rect 15290 6287 15346 6296
rect 15578 6012 15886 6021
rect 15578 6010 15584 6012
rect 15640 6010 15664 6012
rect 15720 6010 15744 6012
rect 15800 6010 15824 6012
rect 15880 6010 15886 6012
rect 15640 5958 15642 6010
rect 15822 5958 15824 6010
rect 15578 5956 15584 5958
rect 15640 5956 15664 5958
rect 15720 5956 15744 5958
rect 15800 5956 15824 5958
rect 15880 5956 15886 5958
rect 15578 5947 15886 5956
rect 15198 5672 15254 5681
rect 15198 5607 15254 5616
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 14752 3046 14872 3074
rect 14752 2825 14780 3046
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 14738 2816 14794 2825
rect 14738 2751 14794 2760
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14568 1222 14596 2382
rect 14844 2106 14872 2926
rect 15304 2650 15332 3470
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 14832 2100 14884 2106
rect 14832 2042 14884 2048
rect 15014 2000 15070 2009
rect 15014 1935 15070 1944
rect 14556 1216 14608 1222
rect 14556 1158 14608 1164
rect 14384 882 14504 898
rect 14372 876 14504 882
rect 14424 870 14504 876
rect 14372 818 14424 824
rect 15028 814 15056 1935
rect 13728 808 13780 814
rect 13728 750 13780 756
rect 13820 808 13872 814
rect 13820 750 13872 756
rect 14464 808 14516 814
rect 14464 750 14516 756
rect 15016 808 15068 814
rect 15016 750 15068 756
rect 13636 672 13688 678
rect 13636 614 13688 620
rect 13648 406 13676 614
rect 13636 400 13688 406
rect 13636 342 13688 348
rect 13740 338 13768 750
rect 13832 338 13860 750
rect 14476 649 14504 750
rect 14462 640 14518 649
rect 14462 575 14518 584
rect 14476 406 14504 575
rect 14464 400 14516 406
rect 14464 342 14516 348
rect 13728 332 13780 338
rect 13728 274 13780 280
rect 13820 332 13872 338
rect 13820 274 13872 280
rect 12348 264 12400 270
rect 12348 206 12400 212
rect 15396 202 15424 5510
rect 15578 4924 15886 4933
rect 15578 4922 15584 4924
rect 15640 4922 15664 4924
rect 15720 4922 15744 4924
rect 15800 4922 15824 4924
rect 15880 4922 15886 4924
rect 15640 4870 15642 4922
rect 15822 4870 15824 4922
rect 15578 4868 15584 4870
rect 15640 4868 15664 4870
rect 15720 4868 15744 4870
rect 15800 4868 15824 4870
rect 15880 4868 15886 4870
rect 15578 4859 15886 4868
rect 15474 4040 15530 4049
rect 15474 3975 15476 3984
rect 15528 3975 15530 3984
rect 15476 3946 15528 3952
rect 15578 3836 15886 3845
rect 15578 3834 15584 3836
rect 15640 3834 15664 3836
rect 15720 3834 15744 3836
rect 15800 3834 15824 3836
rect 15880 3834 15886 3836
rect 15640 3782 15642 3834
rect 15822 3782 15824 3834
rect 15578 3780 15584 3782
rect 15640 3780 15664 3782
rect 15720 3780 15744 3782
rect 15800 3780 15824 3782
rect 15880 3780 15886 3782
rect 15578 3771 15886 3780
rect 15948 3505 15976 7919
rect 16396 7890 16448 7896
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 16132 7002 16160 7754
rect 16500 7750 16528 8910
rect 16592 8401 16620 10610
rect 16684 10130 16712 11086
rect 16960 10810 16988 11698
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17144 11354 17172 11494
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 17052 10130 17080 10950
rect 17144 10266 17172 11290
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 17132 9988 17184 9994
rect 17132 9930 17184 9936
rect 17144 9518 17172 9930
rect 17236 9722 17264 12242
rect 18064 12238 18092 12650
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 18340 11694 18368 12650
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18708 12306 18736 12582
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18524 11898 18552 12174
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18892 11762 18920 12038
rect 18880 11756 18932 11762
rect 18880 11698 18932 11704
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17316 10192 17368 10198
rect 17316 10134 17368 10140
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17328 9674 17356 10134
rect 17592 9716 17644 9722
rect 17328 9646 17362 9674
rect 17644 9664 17724 9674
rect 17592 9658 17724 9664
rect 17604 9646 17724 9658
rect 17334 9602 17362 9646
rect 17328 9574 17362 9602
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 16672 9376 16724 9382
rect 16776 9353 16804 9454
rect 16856 9376 16908 9382
rect 16672 9318 16724 9324
rect 16762 9344 16818 9353
rect 16684 9110 16712 9318
rect 16856 9318 16908 9324
rect 16762 9279 16818 9288
rect 16868 9178 16896 9318
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16672 9104 16724 9110
rect 17052 9081 17080 9454
rect 17222 9344 17278 9353
rect 17144 9302 17222 9330
rect 16672 9046 16724 9052
rect 16762 9072 16818 9081
rect 16762 9007 16764 9016
rect 16816 9007 16818 9016
rect 17038 9072 17094 9081
rect 17038 9007 17094 9016
rect 16764 8978 16816 8984
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16578 8392 16634 8401
rect 16578 8327 16634 8336
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16394 7168 16450 7177
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 16210 6760 16266 6769
rect 16210 6695 16266 6704
rect 16224 6458 16252 6695
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16316 6322 16344 7142
rect 16394 7103 16450 7112
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16224 5166 16252 5646
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 16224 4622 16252 5102
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16224 4078 16252 4558
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16224 3738 16252 4014
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 15934 3496 15990 3505
rect 15934 3431 15990 3440
rect 16224 2922 16252 3674
rect 16408 2961 16436 7103
rect 16500 6866 16528 7686
rect 16578 7440 16634 7449
rect 16578 7375 16580 7384
rect 16632 7375 16634 7384
rect 16580 7346 16632 7352
rect 16578 6896 16634 6905
rect 16488 6860 16540 6866
rect 16578 6831 16580 6840
rect 16488 6802 16540 6808
rect 16632 6831 16634 6840
rect 16580 6802 16632 6808
rect 16500 5953 16528 6802
rect 16684 6746 16712 8774
rect 16776 7886 16804 8978
rect 17144 8974 17172 9302
rect 17222 9279 17278 9288
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16776 7342 16804 7686
rect 16960 7585 16988 7686
rect 16946 7576 17002 7585
rect 16946 7511 17002 7520
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16960 6882 16988 7511
rect 17038 7304 17094 7313
rect 17038 7239 17094 7248
rect 17052 7206 17080 7239
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17038 6896 17094 6905
rect 16764 6860 16816 6866
rect 16960 6854 17038 6882
rect 17144 6866 17172 7142
rect 17038 6831 17094 6840
rect 17132 6860 17184 6866
rect 16764 6802 16816 6808
rect 17132 6802 17184 6808
rect 16592 6718 16712 6746
rect 16592 6662 16620 6718
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16684 6254 16712 6598
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16486 5944 16542 5953
rect 16776 5914 16804 6802
rect 17130 6760 17186 6769
rect 17130 6695 17186 6704
rect 17144 6662 17172 6695
rect 17236 6662 17264 8366
rect 17328 6866 17356 9574
rect 17498 9480 17554 9489
rect 17498 9415 17554 9424
rect 17408 8968 17460 8974
rect 17406 8936 17408 8945
rect 17460 8936 17462 8945
rect 17406 8871 17462 8880
rect 17512 8022 17540 9415
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17604 9178 17632 9318
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17500 8016 17552 8022
rect 17500 7958 17552 7964
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17316 6860 17368 6866
rect 17316 6802 17368 6808
rect 17132 6656 17184 6662
rect 17132 6598 17184 6604
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 17040 6112 17092 6118
rect 17040 6054 17092 6060
rect 16486 5879 16542 5888
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16868 5778 16896 6054
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16592 5166 16620 5646
rect 16960 5234 16988 6054
rect 17052 5914 17080 6054
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17144 5574 17172 6598
rect 17224 6112 17276 6118
rect 17224 6054 17276 6060
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16592 4826 16620 5102
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16592 3942 16620 4762
rect 17236 4690 17264 6054
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16592 3670 16620 3878
rect 16580 3664 16632 3670
rect 16632 3612 16712 3618
rect 16580 3606 16712 3612
rect 16592 3590 16712 3606
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16592 3074 16620 3130
rect 16500 3046 16620 3074
rect 16394 2952 16450 2961
rect 16212 2916 16264 2922
rect 16394 2887 16450 2896
rect 16212 2858 16264 2864
rect 16224 2774 16252 2858
rect 15578 2748 15886 2757
rect 15578 2746 15584 2748
rect 15640 2746 15664 2748
rect 15720 2746 15744 2748
rect 15800 2746 15824 2748
rect 15880 2746 15886 2748
rect 15640 2694 15642 2746
rect 15822 2694 15824 2746
rect 15578 2692 15584 2694
rect 15640 2692 15664 2694
rect 15720 2692 15744 2694
rect 15800 2692 15824 2694
rect 15880 2692 15886 2694
rect 15578 2683 15886 2692
rect 16132 2746 16252 2774
rect 16132 2514 16160 2746
rect 16120 2508 16172 2514
rect 16120 2450 16172 2456
rect 16132 1970 16160 2450
rect 16500 2310 16528 3046
rect 16684 2990 16712 3590
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 17132 3528 17184 3534
rect 17224 3528 17276 3534
rect 17132 3470 17184 3476
rect 17222 3496 17224 3505
rect 17276 3496 17278 3505
rect 16672 2984 16724 2990
rect 16592 2932 16672 2938
rect 16592 2926 16724 2932
rect 16592 2910 16712 2926
rect 16592 2650 16620 2910
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16120 1964 16172 1970
rect 16120 1906 16172 1912
rect 15578 1660 15886 1669
rect 15578 1658 15584 1660
rect 15640 1658 15664 1660
rect 15720 1658 15744 1660
rect 15800 1658 15824 1660
rect 15880 1658 15886 1660
rect 15640 1606 15642 1658
rect 15822 1606 15824 1658
rect 15578 1604 15584 1606
rect 15640 1604 15664 1606
rect 15720 1604 15744 1606
rect 15800 1604 15824 1606
rect 15880 1604 15886 1606
rect 15578 1595 15886 1604
rect 16132 1426 16160 1906
rect 16592 1766 16620 2586
rect 16776 2281 16804 3470
rect 17144 3194 17172 3470
rect 17222 3431 17278 3440
rect 17132 3188 17184 3194
rect 17132 3130 17184 3136
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 16762 2272 16818 2281
rect 16762 2207 16818 2216
rect 17052 2106 17080 2926
rect 17144 2774 17172 3130
rect 17144 2746 17264 2774
rect 17236 2650 17264 2746
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17040 2100 17092 2106
rect 17040 2042 17092 2048
rect 16856 1896 16908 1902
rect 16856 1838 16908 1844
rect 16580 1760 16632 1766
rect 16580 1702 16632 1708
rect 16302 1592 16358 1601
rect 16592 1562 16620 1702
rect 16302 1527 16358 1536
rect 16580 1556 16632 1562
rect 16210 1456 16266 1465
rect 16120 1420 16172 1426
rect 16210 1391 16266 1400
rect 16120 1362 16172 1368
rect 16224 950 16252 1391
rect 16212 944 16264 950
rect 16212 886 16264 892
rect 16316 814 16344 1527
rect 16580 1498 16632 1504
rect 16868 1018 16896 1838
rect 17328 1578 17356 6802
rect 17420 4486 17448 7142
rect 17512 7002 17540 7346
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17604 6254 17632 7890
rect 17696 6780 17724 9646
rect 17776 9376 17828 9382
rect 17774 9344 17776 9353
rect 17828 9344 17830 9353
rect 17774 9279 17830 9288
rect 17774 9208 17830 9217
rect 17774 9143 17830 9152
rect 17788 8974 17816 9143
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17776 8832 17828 8838
rect 17880 8820 17908 10746
rect 18892 10713 18920 11698
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 18984 11354 19012 11630
rect 19168 11558 19196 12378
rect 19260 12306 19288 13670
rect 19352 13190 19380 13960
rect 20456 13954 20484 17575
rect 20640 17542 20668 17575
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20628 17128 20680 17134
rect 20628 17070 20680 17076
rect 20640 16726 20668 17070
rect 20628 16720 20680 16726
rect 20628 16662 20680 16668
rect 20640 14822 20668 16662
rect 20732 15570 20760 17478
rect 20916 16697 20944 18176
rect 20996 18158 21048 18164
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 21100 17542 21128 17682
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 21008 17134 21036 17478
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 20902 16688 20958 16697
rect 20902 16623 20958 16632
rect 21086 16688 21142 16697
rect 21086 16623 21088 16632
rect 21140 16623 21142 16632
rect 21088 16594 21140 16600
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21008 16114 21036 16390
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 21192 15065 21220 19246
rect 21364 19236 21416 19242
rect 21364 19178 21416 19184
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21284 15502 21312 16390
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21178 15056 21234 15065
rect 21178 14991 21234 15000
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21192 14414 21220 14758
rect 21284 14482 21312 15438
rect 21272 14476 21324 14482
rect 21272 14418 21324 14424
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20088 13926 20484 13954
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19800 13728 19852 13734
rect 19800 13670 19852 13676
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19373 13084 19681 13093
rect 19373 13082 19379 13084
rect 19435 13082 19459 13084
rect 19515 13082 19539 13084
rect 19595 13082 19619 13084
rect 19675 13082 19681 13084
rect 19435 13030 19437 13082
rect 19617 13030 19619 13082
rect 19373 13028 19379 13030
rect 19435 13028 19459 13030
rect 19515 13028 19539 13030
rect 19595 13028 19619 13030
rect 19675 13028 19681 13030
rect 19373 13019 19681 13028
rect 19812 12782 19840 13670
rect 19904 12850 19932 13806
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19996 13190 20024 13330
rect 20088 13297 20116 13926
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20074 13288 20130 13297
rect 20074 13223 20076 13232
rect 20128 13223 20130 13232
rect 20076 13194 20128 13200
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19373 11996 19681 12005
rect 19373 11994 19379 11996
rect 19435 11994 19459 11996
rect 19515 11994 19539 11996
rect 19595 11994 19619 11996
rect 19675 11994 19681 11996
rect 19435 11942 19437 11994
rect 19617 11942 19619 11994
rect 19373 11940 19379 11942
rect 19435 11940 19459 11942
rect 19515 11940 19539 11942
rect 19595 11940 19619 11942
rect 19675 11940 19681 11942
rect 19373 11931 19681 11940
rect 19432 11756 19484 11762
rect 19720 11744 19748 12582
rect 20180 12442 20208 13806
rect 20272 13734 20300 13806
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 20548 13394 20576 14282
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20260 13388 20312 13394
rect 20260 13330 20312 13336
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20272 12782 20300 13330
rect 20352 13184 20404 13190
rect 20404 13132 20484 13138
rect 20352 13126 20484 13132
rect 20364 13110 20484 13126
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20352 12776 20404 12782
rect 20352 12718 20404 12724
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20364 12238 20392 12718
rect 19800 12232 19852 12238
rect 19800 12174 19852 12180
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 19484 11716 19748 11744
rect 19432 11698 19484 11704
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 18972 11212 19024 11218
rect 18972 11154 19024 11160
rect 18878 10704 18934 10713
rect 18144 10668 18196 10674
rect 18878 10639 18880 10648
rect 18144 10610 18196 10616
rect 18932 10639 18934 10648
rect 18880 10610 18932 10616
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 17972 9926 18000 9998
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 18064 9722 18092 9998
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17828 8792 17908 8820
rect 17776 8774 17828 8780
rect 17972 8498 18000 8978
rect 18156 8786 18184 10610
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18616 9722 18644 10542
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18800 10266 18828 10406
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 18234 9072 18290 9081
rect 18234 9007 18290 9016
rect 18064 8758 18184 8786
rect 17960 8492 18012 8498
rect 17880 8452 17960 8480
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 17788 7954 17816 8230
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17788 7546 17816 7890
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17788 7002 17816 7482
rect 17880 7342 17908 8452
rect 17960 8434 18012 8440
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17868 6792 17920 6798
rect 17696 6752 17868 6780
rect 17868 6734 17920 6740
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17408 4480 17460 4486
rect 17408 4422 17460 4428
rect 17604 3097 17632 6190
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17696 4282 17724 6054
rect 17788 5137 17816 6598
rect 17774 5128 17830 5137
rect 17774 5063 17830 5072
rect 17774 4312 17830 4321
rect 17684 4276 17736 4282
rect 17880 4298 17908 6734
rect 17972 6254 18000 7822
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 17830 4270 17908 4298
rect 17774 4247 17776 4256
rect 17684 4218 17736 4224
rect 17828 4247 17830 4256
rect 17776 4218 17828 4224
rect 17590 3088 17646 3097
rect 17590 3023 17646 3032
rect 17406 1592 17462 1601
rect 17328 1550 17406 1578
rect 17406 1527 17462 1536
rect 16948 1352 17000 1358
rect 16948 1294 17000 1300
rect 17040 1352 17092 1358
rect 17040 1294 17092 1300
rect 16960 1018 16988 1294
rect 16856 1012 16908 1018
rect 16856 954 16908 960
rect 16948 1012 17000 1018
rect 16948 954 17000 960
rect 17052 882 17080 1294
rect 17972 950 18000 6190
rect 18064 4690 18092 8758
rect 18248 8634 18276 9007
rect 18420 8968 18472 8974
rect 18418 8936 18420 8945
rect 18472 8936 18474 8945
rect 18328 8900 18380 8906
rect 18418 8871 18474 8880
rect 18328 8842 18380 8848
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18156 8090 18184 8570
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18156 7342 18184 8026
rect 18340 7562 18368 8842
rect 18708 8498 18736 9454
rect 18984 8906 19012 11154
rect 19168 10470 19196 11494
rect 19812 11218 19840 12174
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19536 11014 19564 11154
rect 20456 11121 20484 13110
rect 20640 12986 20668 13806
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20628 12980 20680 12986
rect 20628 12922 20680 12928
rect 20812 12844 20864 12850
rect 20732 12804 20812 12832
rect 20442 11112 20498 11121
rect 20442 11047 20498 11056
rect 19524 11008 19576 11014
rect 19524 10950 19576 10956
rect 19708 11008 19760 11014
rect 19708 10950 19760 10956
rect 19373 10908 19681 10917
rect 19373 10906 19379 10908
rect 19435 10906 19459 10908
rect 19515 10906 19539 10908
rect 19595 10906 19619 10908
rect 19675 10906 19681 10908
rect 19435 10854 19437 10906
rect 19617 10854 19619 10906
rect 19373 10852 19379 10854
rect 19435 10852 19459 10854
rect 19515 10852 19539 10854
rect 19595 10852 19619 10854
rect 19675 10852 19681 10854
rect 19373 10843 19681 10852
rect 19338 10704 19394 10713
rect 19338 10639 19340 10648
rect 19392 10639 19394 10648
rect 19340 10610 19392 10616
rect 19720 10606 19748 10950
rect 20732 10810 20760 12804
rect 20812 12786 20864 12792
rect 20916 12782 20944 13670
rect 21284 13326 21312 14214
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 21100 12442 21128 12718
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 21192 12442 21220 12582
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 21180 12436 21232 12442
rect 21376 12434 21404 19178
rect 21468 15502 21496 19479
rect 21824 19304 21876 19310
rect 21824 19246 21876 19252
rect 21836 18834 21864 19246
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 21732 18624 21784 18630
rect 21732 18566 21784 18572
rect 21928 18578 21956 20742
rect 22020 19378 22048 21286
rect 22204 21146 22232 21422
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22204 19922 22232 20742
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22388 19666 22416 22170
rect 23584 22001 23612 22238
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23768 22114 23796 22170
rect 23676 22086 23796 22114
rect 23570 21992 23626 22001
rect 23296 21956 23348 21962
rect 23570 21927 23626 21936
rect 23296 21898 23348 21904
rect 22742 21584 22798 21593
rect 22742 21519 22798 21528
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22480 19854 22508 20198
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 22388 19638 22600 19666
rect 22468 19508 22520 19514
rect 22468 19450 22520 19456
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 22192 19168 22244 19174
rect 22192 19110 22244 19116
rect 22204 18970 22232 19110
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 22480 18766 22508 19450
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 22284 18624 22336 18630
rect 21744 18086 21772 18566
rect 21928 18550 22048 18578
rect 22284 18566 22336 18572
rect 21914 18456 21970 18465
rect 21914 18391 21970 18400
rect 21548 18080 21600 18086
rect 21732 18080 21784 18086
rect 21600 18040 21680 18068
rect 21548 18022 21600 18028
rect 21652 17746 21680 18040
rect 21732 18022 21784 18028
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21652 16590 21680 17682
rect 21732 17672 21784 17678
rect 21928 17660 21956 18391
rect 21784 17632 21956 17660
rect 21732 17614 21784 17620
rect 22020 17338 22048 18550
rect 22100 17740 22152 17746
rect 22100 17682 22152 17688
rect 22112 17649 22140 17682
rect 22098 17640 22154 17649
rect 22098 17575 22154 17584
rect 21916 17332 21968 17338
rect 21916 17274 21968 17280
rect 22008 17332 22060 17338
rect 22008 17274 22060 17280
rect 21928 16590 21956 17274
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21916 16584 21968 16590
rect 22204 16561 22232 16934
rect 21916 16526 21968 16532
rect 22190 16552 22246 16561
rect 21652 15502 21680 16526
rect 22190 16487 22246 16496
rect 22296 16114 22324 18566
rect 22284 16108 22336 16114
rect 22284 16050 22336 16056
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21640 15496 21692 15502
rect 22008 15496 22060 15502
rect 21640 15438 21692 15444
rect 21836 15444 22008 15450
rect 21836 15438 22060 15444
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21560 14618 21588 14758
rect 21652 14618 21680 15438
rect 21836 15422 22048 15438
rect 21548 14612 21600 14618
rect 21548 14554 21600 14560
rect 21640 14612 21692 14618
rect 21640 14554 21692 14560
rect 21730 13424 21786 13433
rect 21730 13359 21732 13368
rect 21784 13359 21786 13368
rect 21732 13330 21784 13336
rect 21640 13320 21692 13326
rect 21640 13262 21692 13268
rect 21652 13002 21680 13262
rect 21836 13190 21864 15422
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21928 14414 21956 15302
rect 22100 14884 22152 14890
rect 22100 14826 22152 14832
rect 22112 14618 22140 14826
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 21916 14408 21968 14414
rect 21916 14350 21968 14356
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 21824 13184 21876 13190
rect 21824 13126 21876 13132
rect 21916 13184 21968 13190
rect 22020 13138 22048 14350
rect 22284 13864 22336 13870
rect 22284 13806 22336 13812
rect 22296 13326 22324 13806
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22284 13320 22336 13326
rect 22284 13262 22336 13268
rect 21968 13132 22048 13138
rect 21916 13126 22048 13132
rect 21928 13110 22048 13126
rect 21652 12974 21864 13002
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21180 12378 21232 12384
rect 21284 12406 21404 12434
rect 21284 12186 21312 12406
rect 21364 12300 21416 12306
rect 21468 12288 21496 12582
rect 21548 12436 21600 12442
rect 21548 12378 21600 12384
rect 21560 12306 21588 12378
rect 21416 12260 21496 12288
rect 21548 12300 21600 12306
rect 21364 12242 21416 12248
rect 21548 12242 21600 12248
rect 21836 12238 21864 12974
rect 22204 12850 22232 13262
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22020 12442 22048 12786
rect 22008 12436 22060 12442
rect 22572 12434 22600 19638
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22664 18329 22692 18702
rect 22756 18426 22784 21519
rect 23308 21418 23336 21898
rect 23584 21486 23612 21927
rect 23676 21486 23704 22086
rect 25976 21622 26004 22238
rect 28724 22228 28776 22234
rect 28724 22170 28776 22176
rect 28080 22160 28132 22166
rect 28080 22102 28132 22108
rect 26608 21888 26660 21894
rect 26608 21830 26660 21836
rect 25964 21616 26016 21622
rect 24490 21584 24546 21593
rect 23756 21548 23808 21554
rect 23756 21490 23808 21496
rect 23940 21548 23992 21554
rect 23940 21490 23992 21496
rect 24032 21548 24084 21554
rect 24596 21554 25084 21570
rect 25964 21558 26016 21564
rect 24490 21519 24492 21528
rect 24032 21490 24084 21496
rect 24544 21519 24546 21528
rect 24584 21548 25084 21554
rect 24492 21490 24544 21496
rect 24636 21542 25084 21548
rect 24584 21490 24636 21496
rect 23572 21480 23624 21486
rect 23572 21422 23624 21428
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23296 21412 23348 21418
rect 23296 21354 23348 21360
rect 23168 21244 23476 21253
rect 23168 21242 23174 21244
rect 23230 21242 23254 21244
rect 23310 21242 23334 21244
rect 23390 21242 23414 21244
rect 23470 21242 23476 21244
rect 23230 21190 23232 21242
rect 23412 21190 23414 21242
rect 23168 21188 23174 21190
rect 23230 21188 23254 21190
rect 23310 21188 23334 21190
rect 23390 21188 23414 21190
rect 23470 21188 23476 21190
rect 23168 21179 23476 21188
rect 22836 21072 22888 21078
rect 22834 21040 22836 21049
rect 22888 21040 22890 21049
rect 22834 20975 22890 20984
rect 23112 21004 23164 21010
rect 23112 20946 23164 20952
rect 22926 20904 22982 20913
rect 22926 20839 22982 20848
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22650 18320 22706 18329
rect 22650 18255 22706 18264
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22652 17060 22704 17066
rect 22652 17002 22704 17008
rect 22664 16590 22692 17002
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22848 16522 22876 18226
rect 22940 18222 22968 20839
rect 23020 20596 23072 20602
rect 23020 20538 23072 20544
rect 23032 19514 23060 20538
rect 23124 20330 23152 20946
rect 23662 20768 23718 20777
rect 23662 20703 23718 20712
rect 23572 20528 23624 20534
rect 23572 20470 23624 20476
rect 23112 20324 23164 20330
rect 23112 20266 23164 20272
rect 23168 20156 23476 20165
rect 23168 20154 23174 20156
rect 23230 20154 23254 20156
rect 23310 20154 23334 20156
rect 23390 20154 23414 20156
rect 23470 20154 23476 20156
rect 23230 20102 23232 20154
rect 23412 20102 23414 20154
rect 23168 20100 23174 20102
rect 23230 20100 23254 20102
rect 23310 20100 23334 20102
rect 23390 20100 23414 20102
rect 23470 20100 23476 20102
rect 23168 20091 23476 20100
rect 23584 20097 23612 20470
rect 23570 20088 23626 20097
rect 23570 20023 23626 20032
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 23168 19068 23476 19077
rect 23168 19066 23174 19068
rect 23230 19066 23254 19068
rect 23310 19066 23334 19068
rect 23390 19066 23414 19068
rect 23470 19066 23476 19068
rect 23230 19014 23232 19066
rect 23412 19014 23414 19066
rect 23168 19012 23174 19014
rect 23230 19012 23254 19014
rect 23310 19012 23334 19014
rect 23390 19012 23414 19014
rect 23470 19012 23476 19014
rect 23168 19003 23476 19012
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23492 18630 23520 18906
rect 23584 18737 23612 19110
rect 23570 18728 23626 18737
rect 23570 18663 23626 18672
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23492 18426 23520 18566
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23676 18222 23704 20703
rect 23768 19310 23796 21490
rect 23848 21412 23900 21418
rect 23848 21354 23900 21360
rect 23860 19310 23888 21354
rect 23952 20058 23980 21490
rect 24044 21350 24072 21490
rect 25056 21486 25084 21542
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 25044 21480 25096 21486
rect 25044 21422 25096 21428
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 24768 20868 24820 20874
rect 24768 20810 24820 20816
rect 24308 20800 24360 20806
rect 24308 20742 24360 20748
rect 24124 20324 24176 20330
rect 24124 20266 24176 20272
rect 24136 20058 24164 20266
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 24320 19310 24348 20742
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 23756 19304 23808 19310
rect 23756 19246 23808 19252
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 24308 19304 24360 19310
rect 24308 19246 24360 19252
rect 24124 19236 24176 19242
rect 24124 19178 24176 19184
rect 23756 19168 23808 19174
rect 23756 19110 23808 19116
rect 23768 18426 23796 19110
rect 23848 18964 23900 18970
rect 23848 18906 23900 18912
rect 23756 18420 23808 18426
rect 23756 18362 23808 18368
rect 22928 18216 22980 18222
rect 23664 18216 23716 18222
rect 22928 18158 22980 18164
rect 23386 18184 23442 18193
rect 23664 18158 23716 18164
rect 23386 18119 23442 18128
rect 23400 18086 23428 18119
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23168 17980 23476 17989
rect 23168 17978 23174 17980
rect 23230 17978 23254 17980
rect 23310 17978 23334 17980
rect 23390 17978 23414 17980
rect 23470 17978 23476 17980
rect 23230 17926 23232 17978
rect 23412 17926 23414 17978
rect 23168 17924 23174 17926
rect 23230 17924 23254 17926
rect 23310 17924 23334 17926
rect 23390 17924 23414 17926
rect 23470 17924 23476 17926
rect 23168 17915 23476 17924
rect 23754 17912 23810 17921
rect 23584 17870 23754 17898
rect 23020 17604 23072 17610
rect 23020 17546 23072 17552
rect 22926 17368 22982 17377
rect 22926 17303 22982 17312
rect 22836 16516 22888 16522
rect 22836 16458 22888 16464
rect 22744 16448 22796 16454
rect 22664 16408 22744 16436
rect 22664 13410 22692 16408
rect 22744 16390 22796 16396
rect 22744 16040 22796 16046
rect 22744 15982 22796 15988
rect 22756 14822 22784 15982
rect 22940 15026 22968 17303
rect 23032 17270 23060 17546
rect 23112 17536 23164 17542
rect 23112 17478 23164 17484
rect 23020 17264 23072 17270
rect 23124 17241 23152 17478
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 23020 17206 23072 17212
rect 23110 17232 23166 17241
rect 23110 17167 23166 17176
rect 23112 17128 23164 17134
rect 23216 17116 23244 17274
rect 23584 17202 23612 17870
rect 23754 17847 23810 17856
rect 23756 17740 23808 17746
rect 23756 17682 23808 17688
rect 23662 17232 23718 17241
rect 23572 17196 23624 17202
rect 23662 17167 23718 17176
rect 23572 17138 23624 17144
rect 23164 17088 23244 17116
rect 23112 17070 23164 17076
rect 23020 17060 23072 17066
rect 23020 17002 23072 17008
rect 23032 16969 23060 17002
rect 23018 16960 23074 16969
rect 23676 16946 23704 17167
rect 23018 16895 23074 16904
rect 23584 16918 23704 16946
rect 23168 16892 23476 16901
rect 23168 16890 23174 16892
rect 23230 16890 23254 16892
rect 23310 16890 23334 16892
rect 23390 16890 23414 16892
rect 23470 16890 23476 16892
rect 23230 16838 23232 16890
rect 23412 16838 23414 16890
rect 23168 16836 23174 16838
rect 23230 16836 23254 16838
rect 23310 16836 23334 16838
rect 23390 16836 23414 16838
rect 23470 16836 23476 16838
rect 23168 16827 23476 16836
rect 23584 16674 23612 16918
rect 23492 16646 23612 16674
rect 23492 16046 23520 16646
rect 23768 16640 23796 17682
rect 23860 17134 23888 18906
rect 23938 18592 23994 18601
rect 23938 18527 23994 18536
rect 23952 18154 23980 18527
rect 23940 18148 23992 18154
rect 23940 18090 23992 18096
rect 24030 18048 24086 18057
rect 24030 17983 24086 17992
rect 24044 17746 24072 17983
rect 24136 17814 24164 19178
rect 24412 18970 24440 19790
rect 24688 19553 24716 19790
rect 24674 19544 24730 19553
rect 24674 19479 24730 19488
rect 24780 19334 24808 20810
rect 24872 20262 24900 21422
rect 25320 21344 25372 21350
rect 25320 21286 25372 21292
rect 25134 21176 25190 21185
rect 25332 21146 25360 21286
rect 25134 21111 25190 21120
rect 25320 21140 25372 21146
rect 25148 21010 25176 21111
rect 25320 21082 25372 21088
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 25148 20398 25176 20946
rect 25320 20528 25372 20534
rect 25320 20470 25372 20476
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 25148 20058 25176 20334
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 24584 19304 24636 19310
rect 24780 19306 24992 19334
rect 24584 19246 24636 19252
rect 24400 18964 24452 18970
rect 24400 18906 24452 18912
rect 24492 18964 24544 18970
rect 24492 18906 24544 18912
rect 24504 18850 24532 18906
rect 24412 18834 24532 18850
rect 24400 18828 24532 18834
rect 24452 18822 24532 18828
rect 24400 18770 24452 18776
rect 24320 18686 24532 18714
rect 24216 18284 24268 18290
rect 24216 18226 24268 18232
rect 24124 17808 24176 17814
rect 24124 17750 24176 17756
rect 24032 17740 24084 17746
rect 24032 17682 24084 17688
rect 24032 17604 24084 17610
rect 24032 17546 24084 17552
rect 23848 17128 23900 17134
rect 23848 17070 23900 17076
rect 23848 16992 23900 16998
rect 24044 16980 24072 17546
rect 24228 17513 24256 18226
rect 24320 18086 24348 18686
rect 24504 18630 24532 18686
rect 24400 18624 24452 18630
rect 24400 18566 24452 18572
rect 24492 18624 24544 18630
rect 24492 18566 24544 18572
rect 24308 18080 24360 18086
rect 24308 18022 24360 18028
rect 24412 18034 24440 18566
rect 24596 18358 24624 19246
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24858 18728 24914 18737
rect 24584 18352 24636 18358
rect 24584 18294 24636 18300
rect 24412 18006 24532 18034
rect 24306 17912 24362 17921
rect 24400 17876 24452 17882
rect 24362 17856 24400 17864
rect 24306 17847 24400 17856
rect 24320 17836 24400 17847
rect 24214 17504 24270 17513
rect 24214 17439 24270 17448
rect 24228 17134 24256 17439
rect 24216 17128 24268 17134
rect 24216 17070 24268 17076
rect 23900 16952 24072 16980
rect 23848 16934 23900 16940
rect 24044 16658 24072 16952
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 23940 16652 23992 16658
rect 23768 16612 23888 16640
rect 23860 16561 23888 16612
rect 23940 16594 23992 16600
rect 24032 16652 24084 16658
rect 24032 16594 24084 16600
rect 23846 16552 23902 16561
rect 23756 16516 23808 16522
rect 23952 16522 23980 16594
rect 23846 16487 23902 16496
rect 23940 16516 23992 16522
rect 23756 16458 23808 16464
rect 23940 16458 23992 16464
rect 23572 16448 23624 16454
rect 23572 16390 23624 16396
rect 23480 16040 23532 16046
rect 23480 15982 23532 15988
rect 23168 15804 23476 15813
rect 23168 15802 23174 15804
rect 23230 15802 23254 15804
rect 23310 15802 23334 15804
rect 23390 15802 23414 15804
rect 23470 15802 23476 15804
rect 23230 15750 23232 15802
rect 23412 15750 23414 15802
rect 23168 15748 23174 15750
rect 23230 15748 23254 15750
rect 23310 15748 23334 15750
rect 23390 15748 23414 15750
rect 23470 15748 23476 15750
rect 23168 15739 23476 15748
rect 23020 15632 23072 15638
rect 23480 15632 23532 15638
rect 23020 15574 23072 15580
rect 23386 15600 23442 15609
rect 22928 15020 22980 15026
rect 22928 14962 22980 14968
rect 22744 14816 22796 14822
rect 22744 14758 22796 14764
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 22940 14074 22968 14758
rect 23032 14074 23060 15574
rect 23480 15574 23532 15580
rect 23386 15535 23442 15544
rect 23400 15162 23428 15535
rect 23492 15162 23520 15574
rect 23584 15570 23612 16390
rect 23768 16114 23796 16458
rect 24044 16402 24072 16594
rect 23860 16374 24072 16402
rect 23756 16108 23808 16114
rect 23756 16050 23808 16056
rect 23664 16040 23716 16046
rect 23664 15982 23716 15988
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 23676 15502 23704 15982
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23388 15156 23440 15162
rect 23388 15098 23440 15104
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23676 15026 23704 15438
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23572 14952 23624 14958
rect 23572 14894 23624 14900
rect 23584 14793 23612 14894
rect 23570 14784 23626 14793
rect 23168 14716 23476 14725
rect 23570 14719 23626 14728
rect 23168 14714 23174 14716
rect 23230 14714 23254 14716
rect 23310 14714 23334 14716
rect 23390 14714 23414 14716
rect 23470 14714 23476 14716
rect 23230 14662 23232 14714
rect 23412 14662 23414 14714
rect 23168 14660 23174 14662
rect 23230 14660 23254 14662
rect 23310 14660 23334 14662
rect 23390 14660 23414 14662
rect 23470 14660 23476 14662
rect 23168 14651 23476 14660
rect 23676 14414 23704 14962
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 22928 14068 22980 14074
rect 22928 14010 22980 14016
rect 23020 14068 23072 14074
rect 23020 14010 23072 14016
rect 23572 14000 23624 14006
rect 23572 13942 23624 13948
rect 23020 13796 23072 13802
rect 23020 13738 23072 13744
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22742 13424 22798 13433
rect 22664 13382 22742 13410
rect 22742 13359 22798 13368
rect 22848 12782 22876 13670
rect 22928 12912 22980 12918
rect 22926 12880 22928 12889
rect 22980 12880 22982 12889
rect 22926 12815 22982 12824
rect 22836 12776 22888 12782
rect 22836 12718 22888 12724
rect 23032 12764 23060 13738
rect 23168 13628 23476 13637
rect 23168 13626 23174 13628
rect 23230 13626 23254 13628
rect 23310 13626 23334 13628
rect 23390 13626 23414 13628
rect 23470 13626 23476 13628
rect 23230 13574 23232 13626
rect 23412 13574 23414 13626
rect 23168 13572 23174 13574
rect 23230 13572 23254 13574
rect 23310 13572 23334 13574
rect 23390 13572 23414 13574
rect 23470 13572 23476 13574
rect 23168 13563 23476 13572
rect 23584 13394 23612 13942
rect 23768 13938 23796 16050
rect 23860 16046 23888 16374
rect 23848 16040 23900 16046
rect 23848 15982 23900 15988
rect 23848 15904 23900 15910
rect 23848 15846 23900 15852
rect 23860 15502 23888 15846
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 23860 15094 23888 15438
rect 23848 15088 23900 15094
rect 23848 15030 23900 15036
rect 23860 14482 23888 15030
rect 24136 14482 24164 16730
rect 24320 16590 24348 17836
rect 24400 17818 24452 17824
rect 24504 17762 24532 18006
rect 24412 17734 24532 17762
rect 24412 16674 24440 17734
rect 24492 17672 24544 17678
rect 24596 17660 24624 18294
rect 24688 18057 24716 18702
rect 24858 18663 24914 18672
rect 24872 18290 24900 18663
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24964 18170 24992 19306
rect 25136 19168 25188 19174
rect 25136 19110 25188 19116
rect 24872 18142 24992 18170
rect 24674 18048 24730 18057
rect 24674 17983 24730 17992
rect 24544 17632 24624 17660
rect 24768 17672 24820 17678
rect 24492 17614 24544 17620
rect 24872 17660 24900 18142
rect 25148 18086 25176 19110
rect 25332 18601 25360 20470
rect 25424 20398 25452 21490
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25872 21344 25924 21350
rect 25872 21286 25924 21292
rect 25700 20874 25728 21286
rect 25688 20868 25740 20874
rect 25688 20810 25740 20816
rect 25884 20806 25912 21286
rect 25872 20800 25924 20806
rect 25872 20742 25924 20748
rect 25976 20398 26004 21558
rect 26620 21486 26648 21830
rect 26963 21788 27271 21797
rect 26963 21786 26969 21788
rect 27025 21786 27049 21788
rect 27105 21786 27129 21788
rect 27185 21786 27209 21788
rect 27265 21786 27271 21788
rect 27025 21734 27027 21786
rect 27207 21734 27209 21786
rect 26963 21732 26969 21734
rect 27025 21732 27049 21734
rect 27105 21732 27129 21734
rect 27185 21732 27209 21734
rect 27265 21732 27271 21734
rect 26963 21723 27271 21732
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 26240 21480 26292 21486
rect 26240 21422 26292 21428
rect 26608 21480 26660 21486
rect 26608 21422 26660 21428
rect 26792 21480 26844 21486
rect 26792 21422 26844 21428
rect 26148 21412 26200 21418
rect 26148 21354 26200 21360
rect 26056 20936 26108 20942
rect 26056 20878 26108 20884
rect 25412 20392 25464 20398
rect 25412 20334 25464 20340
rect 25964 20392 26016 20398
rect 25964 20334 26016 20340
rect 25688 19304 25740 19310
rect 25688 19246 25740 19252
rect 25700 18970 25728 19246
rect 25688 18964 25740 18970
rect 25688 18906 25740 18912
rect 25318 18592 25374 18601
rect 25318 18527 25374 18536
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 25136 18080 25188 18086
rect 25136 18022 25188 18028
rect 24820 17632 24900 17660
rect 24768 17614 24820 17620
rect 24766 16688 24822 16697
rect 24412 16646 24624 16674
rect 24596 16590 24624 16646
rect 24688 16646 24766 16674
rect 24308 16584 24360 16590
rect 24584 16584 24636 16590
rect 24490 16552 24546 16561
rect 24308 16526 24360 16532
rect 24216 16108 24268 16114
rect 24216 16050 24268 16056
rect 24228 15586 24256 16050
rect 24320 15910 24348 16526
rect 24412 16510 24490 16538
rect 24412 16114 24440 16510
rect 24584 16526 24636 16532
rect 24490 16487 24546 16496
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24308 15904 24360 15910
rect 24308 15846 24360 15852
rect 24596 15706 24624 15982
rect 24584 15700 24636 15706
rect 24584 15642 24636 15648
rect 24228 15570 24348 15586
rect 24228 15564 24360 15570
rect 24228 15558 24308 15564
rect 24308 15506 24360 15512
rect 24688 15502 24716 16646
rect 24964 16658 24992 18022
rect 25148 17882 25176 18022
rect 25136 17876 25188 17882
rect 25136 17818 25188 17824
rect 25136 17060 25188 17066
rect 25136 17002 25188 17008
rect 24766 16623 24822 16632
rect 24952 16652 25004 16658
rect 24952 16594 25004 16600
rect 24766 16144 24822 16153
rect 24766 16079 24822 16088
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24490 15192 24546 15201
rect 24490 15127 24546 15136
rect 24504 14482 24532 15127
rect 24780 15026 24808 16079
rect 24950 15056 25006 15065
rect 24768 15020 24820 15026
rect 24950 14991 24952 15000
rect 24768 14962 24820 14968
rect 25004 14991 25006 15000
rect 24952 14962 25004 14968
rect 24676 14952 24728 14958
rect 24596 14912 24676 14940
rect 23848 14476 23900 14482
rect 23848 14418 23900 14424
rect 24124 14476 24176 14482
rect 24124 14418 24176 14424
rect 24492 14476 24544 14482
rect 24492 14418 24544 14424
rect 24596 14362 24624 14912
rect 24676 14894 24728 14900
rect 24320 14334 24624 14362
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24032 14272 24084 14278
rect 24032 14214 24084 14220
rect 23756 13932 23808 13938
rect 23756 13874 23808 13880
rect 24044 13462 24072 14214
rect 24320 13802 24348 14334
rect 24872 13938 24900 14350
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24400 13864 24452 13870
rect 24398 13832 24400 13841
rect 24452 13832 24454 13841
rect 24308 13796 24360 13802
rect 24398 13767 24454 13776
rect 24584 13796 24636 13802
rect 24308 13738 24360 13744
rect 24032 13456 24084 13462
rect 24032 13398 24084 13404
rect 24216 13456 24268 13462
rect 24216 13398 24268 13404
rect 24306 13424 24362 13433
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 24124 13320 24176 13326
rect 24124 13262 24176 13268
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23112 12776 23164 12782
rect 23032 12736 23112 12764
rect 22572 12406 22692 12434
rect 22008 12378 22060 12384
rect 21192 12158 21312 12186
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21192 12102 21220 12158
rect 21180 12096 21232 12102
rect 21180 12038 21232 12044
rect 21744 11898 21772 12174
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 19248 10600 19300 10606
rect 19248 10542 19300 10548
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19156 10464 19208 10470
rect 19156 10406 19208 10412
rect 19260 10266 19288 10542
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19984 10192 20036 10198
rect 19984 10134 20036 10140
rect 19373 9820 19681 9829
rect 19373 9818 19379 9820
rect 19435 9818 19459 9820
rect 19515 9818 19539 9820
rect 19595 9818 19619 9820
rect 19675 9818 19681 9820
rect 19435 9766 19437 9818
rect 19617 9766 19619 9818
rect 19373 9764 19379 9766
rect 19435 9764 19459 9766
rect 19515 9764 19539 9766
rect 19595 9764 19619 9766
rect 19675 9764 19681 9766
rect 19373 9755 19681 9764
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19076 9110 19104 9318
rect 19260 9160 19288 9522
rect 19444 9178 19472 9522
rect 19432 9172 19484 9178
rect 19260 9132 19380 9160
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 19352 9058 19380 9132
rect 19432 9114 19484 9120
rect 18972 8900 19024 8906
rect 18972 8842 19024 8848
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18800 8430 18828 8774
rect 19076 8498 19104 9046
rect 19248 9036 19300 9042
rect 19352 9030 19932 9058
rect 19248 8978 19300 8984
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 18788 8424 18840 8430
rect 18788 8366 18840 8372
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18248 7534 18460 7562
rect 18616 7546 18644 7686
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18156 7002 18184 7278
rect 18248 7274 18276 7534
rect 18326 7440 18382 7449
rect 18326 7375 18382 7384
rect 18236 7268 18288 7274
rect 18236 7210 18288 7216
rect 18144 6996 18196 7002
rect 18144 6938 18196 6944
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18248 6390 18276 6734
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 18248 6254 18276 6326
rect 18340 6254 18368 7375
rect 18236 6248 18288 6254
rect 18236 6190 18288 6196
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18432 4690 18460 7534
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18616 7342 18644 7482
rect 18694 7440 18750 7449
rect 18694 7375 18750 7384
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18708 7154 18736 7375
rect 18616 7126 18736 7154
rect 18616 6798 18644 7126
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18604 6656 18656 6662
rect 18604 6598 18656 6604
rect 18616 6186 18644 6598
rect 18708 6458 18736 6734
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18800 6254 18828 7822
rect 19260 6866 19288 8978
rect 19800 8968 19852 8974
rect 19800 8910 19852 8916
rect 19373 8732 19681 8741
rect 19373 8730 19379 8732
rect 19435 8730 19459 8732
rect 19515 8730 19539 8732
rect 19595 8730 19619 8732
rect 19675 8730 19681 8732
rect 19435 8678 19437 8730
rect 19617 8678 19619 8730
rect 19373 8676 19379 8678
rect 19435 8676 19459 8678
rect 19515 8676 19539 8678
rect 19595 8676 19619 8678
rect 19675 8676 19681 8678
rect 19373 8667 19681 8676
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19373 7644 19681 7653
rect 19373 7642 19379 7644
rect 19435 7642 19459 7644
rect 19515 7642 19539 7644
rect 19595 7642 19619 7644
rect 19675 7642 19681 7644
rect 19435 7590 19437 7642
rect 19617 7590 19619 7642
rect 19373 7588 19379 7590
rect 19435 7588 19459 7590
rect 19515 7588 19539 7590
rect 19595 7588 19619 7590
rect 19675 7588 19681 7590
rect 19373 7579 19681 7588
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19720 6730 19748 8366
rect 19812 7546 19840 8910
rect 19904 8090 19932 9030
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19373 6556 19681 6565
rect 19373 6554 19379 6556
rect 19435 6554 19459 6556
rect 19515 6554 19539 6556
rect 19595 6554 19619 6556
rect 19675 6554 19681 6556
rect 19435 6502 19437 6554
rect 19617 6502 19619 6554
rect 19373 6500 19379 6502
rect 19435 6500 19459 6502
rect 19515 6500 19539 6502
rect 19595 6500 19619 6502
rect 19675 6500 19681 6502
rect 19373 6491 19681 6500
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18788 6248 18840 6254
rect 18788 6190 18840 6196
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 18420 4684 18472 4690
rect 18420 4626 18472 4632
rect 18432 3534 18460 4626
rect 18524 3641 18552 6054
rect 18708 5574 18736 6190
rect 18788 6112 18840 6118
rect 18788 6054 18840 6060
rect 18800 5710 18828 6054
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18708 5166 18736 5510
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18708 4078 18736 5102
rect 18800 5030 18828 5646
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18878 4992 18934 5001
rect 18800 4622 18828 4966
rect 18878 4927 18934 4936
rect 18788 4616 18840 4622
rect 18788 4558 18840 4564
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18800 3942 18828 4558
rect 18892 4554 18920 4927
rect 18984 4758 19012 6190
rect 19373 5468 19681 5477
rect 19373 5466 19379 5468
rect 19435 5466 19459 5468
rect 19515 5466 19539 5468
rect 19595 5466 19619 5468
rect 19675 5466 19681 5468
rect 19435 5414 19437 5466
rect 19617 5414 19619 5466
rect 19373 5412 19379 5414
rect 19435 5412 19459 5414
rect 19515 5412 19539 5414
rect 19595 5412 19619 5414
rect 19675 5412 19681 5414
rect 19373 5403 19681 5412
rect 19996 4826 20024 10134
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20272 9058 20300 10066
rect 20180 9042 20300 9058
rect 20168 9036 20300 9042
rect 20220 9030 20300 9036
rect 20168 8978 20220 8984
rect 20548 8974 20576 10746
rect 20824 9586 20852 11086
rect 20916 10266 20944 11154
rect 21008 11150 21036 11766
rect 21088 11280 21140 11286
rect 21088 11222 21140 11228
rect 20996 11144 21048 11150
rect 20996 11086 21048 11092
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 21008 10198 21036 11086
rect 20996 10192 21048 10198
rect 20996 10134 21048 10140
rect 21100 10130 21128 11222
rect 21836 11218 21864 12174
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21928 11898 21956 12038
rect 21916 11892 21968 11898
rect 21916 11834 21968 11840
rect 21928 11762 21956 11834
rect 21916 11756 21968 11762
rect 21916 11698 21968 11704
rect 22020 11558 22048 12378
rect 22664 12102 22692 12406
rect 23032 12238 23060 12736
rect 23112 12718 23164 12724
rect 23168 12540 23476 12549
rect 23168 12538 23174 12540
rect 23230 12538 23254 12540
rect 23310 12538 23334 12540
rect 23390 12538 23414 12540
rect 23470 12538 23476 12540
rect 23230 12486 23232 12538
rect 23412 12486 23414 12538
rect 23168 12484 23174 12486
rect 23230 12484 23254 12486
rect 23310 12484 23334 12486
rect 23390 12484 23414 12486
rect 23470 12484 23476 12486
rect 23168 12475 23476 12484
rect 23388 12436 23440 12442
rect 23584 12424 23612 12922
rect 23768 12918 23796 13126
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 24136 12850 24164 13262
rect 23848 12844 23900 12850
rect 23848 12786 23900 12792
rect 24124 12844 24176 12850
rect 24124 12786 24176 12792
rect 23756 12776 23808 12782
rect 23756 12718 23808 12724
rect 23768 12617 23796 12718
rect 23754 12608 23810 12617
rect 23754 12543 23810 12552
rect 23440 12396 23612 12424
rect 23388 12378 23440 12384
rect 23860 12306 23888 12786
rect 24228 12646 24256 13398
rect 24412 13410 24440 13767
rect 24584 13738 24636 13744
rect 24362 13382 24440 13410
rect 24306 13359 24362 13368
rect 24124 12640 24176 12646
rect 24124 12582 24176 12588
rect 24216 12640 24268 12646
rect 24216 12582 24268 12588
rect 24136 12306 24164 12582
rect 24228 12442 24256 12582
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 24124 12300 24176 12306
rect 24124 12242 24176 12248
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 23940 12232 23992 12238
rect 23940 12174 23992 12180
rect 22652 12096 22704 12102
rect 22652 12038 22704 12044
rect 23952 11898 23980 12174
rect 23940 11892 23992 11898
rect 23940 11834 23992 11840
rect 24122 11792 24178 11801
rect 24122 11727 24124 11736
rect 24176 11727 24178 11736
rect 24124 11698 24176 11704
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 22296 11354 22324 11630
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 21824 11212 21876 11218
rect 21824 11154 21876 11160
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 21548 11008 21600 11014
rect 21548 10950 21600 10956
rect 21560 10606 21588 10950
rect 21824 10668 21876 10674
rect 21824 10610 21876 10616
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21272 10192 21324 10198
rect 21272 10134 21324 10140
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 21284 10062 21312 10134
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 21732 10056 21784 10062
rect 21732 9998 21784 10004
rect 20996 9920 21048 9926
rect 20996 9862 21048 9868
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 21008 9518 21036 9862
rect 21744 9704 21772 9998
rect 21560 9676 21772 9704
rect 20996 9512 21048 9518
rect 20996 9454 21048 9460
rect 21008 9110 21036 9454
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 20444 8356 20496 8362
rect 20444 8298 20496 8304
rect 20456 8090 20484 8298
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 20168 7268 20220 7274
rect 20168 7210 20220 7216
rect 20180 6769 20208 7210
rect 20732 7206 20760 8366
rect 20824 7750 20852 8366
rect 20916 7954 20944 8978
rect 21560 8634 21588 9676
rect 21732 9580 21784 9586
rect 21732 9522 21784 9528
rect 21640 9512 21692 9518
rect 21640 9454 21692 9460
rect 21652 9178 21680 9454
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21744 8634 21772 9522
rect 21836 9110 21864 10610
rect 22020 10266 22048 11154
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22296 10810 22324 10950
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22480 10470 22508 11290
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22008 10260 22060 10266
rect 21928 10220 22008 10248
rect 21928 10062 21956 10220
rect 22008 10202 22060 10208
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 22572 9654 22600 11086
rect 22664 10810 22692 11086
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22756 10742 22784 11630
rect 23168 11452 23476 11461
rect 23168 11450 23174 11452
rect 23230 11450 23254 11452
rect 23310 11450 23334 11452
rect 23390 11450 23414 11452
rect 23470 11450 23476 11452
rect 23230 11398 23232 11450
rect 23412 11398 23414 11450
rect 23168 11396 23174 11398
rect 23230 11396 23254 11398
rect 23310 11396 23334 11398
rect 23390 11396 23414 11398
rect 23470 11396 23476 11398
rect 23168 11387 23476 11396
rect 24032 11008 24084 11014
rect 24032 10950 24084 10956
rect 22744 10736 22796 10742
rect 22744 10678 22796 10684
rect 24044 10606 24072 10950
rect 24032 10600 24084 10606
rect 24032 10542 24084 10548
rect 22652 10464 22704 10470
rect 22652 10406 22704 10412
rect 24124 10464 24176 10470
rect 24124 10406 24176 10412
rect 22664 10266 22692 10406
rect 23168 10364 23476 10373
rect 23168 10362 23174 10364
rect 23230 10362 23254 10364
rect 23310 10362 23334 10364
rect 23390 10362 23414 10364
rect 23470 10362 23476 10364
rect 23230 10310 23232 10362
rect 23412 10310 23414 10362
rect 23168 10308 23174 10310
rect 23230 10308 23254 10310
rect 23310 10308 23334 10310
rect 23390 10308 23414 10310
rect 23470 10308 23476 10310
rect 23168 10299 23476 10308
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 23756 10124 23808 10130
rect 23756 10066 23808 10072
rect 22560 9648 22612 9654
rect 22560 9590 22612 9596
rect 23768 9518 23796 10066
rect 24044 9722 24072 10202
rect 24136 10062 24164 10406
rect 24124 10056 24176 10062
rect 24124 9998 24176 10004
rect 24136 9722 24164 9998
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 24124 9716 24176 9722
rect 24124 9658 24176 9664
rect 24124 9580 24176 9586
rect 24124 9522 24176 9528
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 23756 9512 23808 9518
rect 23756 9454 23808 9460
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 21928 8956 21956 9454
rect 23940 9444 23992 9450
rect 23940 9386 23992 9392
rect 23020 9376 23072 9382
rect 23020 9318 23072 9324
rect 23664 9376 23716 9382
rect 23664 9318 23716 9324
rect 23032 9110 23060 9318
rect 23168 9276 23476 9285
rect 23168 9274 23174 9276
rect 23230 9274 23254 9276
rect 23310 9274 23334 9276
rect 23390 9274 23414 9276
rect 23470 9274 23476 9276
rect 23230 9222 23232 9274
rect 23412 9222 23414 9274
rect 23168 9220 23174 9222
rect 23230 9220 23254 9222
rect 23310 9220 23334 9222
rect 23390 9220 23414 9222
rect 23470 9220 23476 9222
rect 23168 9211 23476 9220
rect 23020 9104 23072 9110
rect 22926 9072 22982 9081
rect 22848 9042 22926 9058
rect 22836 9036 22926 9042
rect 22888 9030 22926 9036
rect 23020 9046 23072 9052
rect 23676 9042 23704 9318
rect 23952 9178 23980 9386
rect 23940 9172 23992 9178
rect 23940 9114 23992 9120
rect 22926 9007 22982 9016
rect 23664 9036 23716 9042
rect 22836 8978 22888 8984
rect 23664 8978 23716 8984
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 21836 8928 21956 8956
rect 22744 8968 22796 8974
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21732 8424 21784 8430
rect 21732 8366 21784 8372
rect 21456 8084 21508 8090
rect 21508 8044 21680 8072
rect 21456 8026 21508 8032
rect 21652 7954 21680 8044
rect 20904 7948 20956 7954
rect 21456 7948 21508 7954
rect 20904 7890 20956 7896
rect 21376 7908 21456 7936
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20824 7342 20852 7686
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20916 7002 20944 7890
rect 21180 7812 21232 7818
rect 21180 7754 21232 7760
rect 21192 7274 21220 7754
rect 21376 7546 21404 7908
rect 21456 7890 21508 7896
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21744 7886 21772 8366
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21456 7812 21508 7818
rect 21456 7754 21508 7760
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21468 7342 21496 7754
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21732 7744 21784 7750
rect 21732 7686 21784 7692
rect 21456 7336 21508 7342
rect 21376 7296 21456 7324
rect 21180 7268 21232 7274
rect 21180 7210 21232 7216
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 20166 6760 20222 6769
rect 20166 6695 20222 6704
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20272 6458 20300 6598
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20548 5234 20576 6598
rect 20916 5914 20944 6938
rect 21192 6798 21220 7210
rect 21272 6860 21324 6866
rect 21272 6802 21324 6808
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19984 4820 20036 4826
rect 19984 4762 20036 4768
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 18880 4548 18932 4554
rect 18880 4490 18932 4496
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18510 3632 18566 3641
rect 18510 3567 18566 3576
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 18420 2508 18472 2514
rect 18524 2496 18552 2926
rect 18472 2468 18552 2496
rect 18420 2450 18472 2456
rect 18616 1986 18644 3470
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18524 1958 18644 1986
rect 17960 944 18012 950
rect 17960 886 18012 892
rect 17040 876 17092 882
rect 17040 818 17092 824
rect 16304 808 16356 814
rect 16304 750 16356 756
rect 16396 808 16448 814
rect 16396 750 16448 756
rect 15578 572 15886 581
rect 15578 570 15584 572
rect 15640 570 15664 572
rect 15720 570 15744 572
rect 15800 570 15824 572
rect 15880 570 15886 572
rect 15640 518 15642 570
rect 15822 518 15824 570
rect 15578 516 15584 518
rect 15640 516 15664 518
rect 15720 516 15744 518
rect 15800 516 15824 518
rect 15880 516 15886 518
rect 15578 507 15886 516
rect 15384 196 15436 202
rect 15384 138 15436 144
rect 9128 128 9180 134
rect 9128 70 9180 76
rect 16408 66 16436 750
rect 16488 740 16540 746
rect 16488 682 16540 688
rect 18420 740 18472 746
rect 18420 682 18472 688
rect 16500 649 16528 682
rect 18236 672 18288 678
rect 16486 640 16542 649
rect 18236 614 18288 620
rect 16486 575 16542 584
rect 18248 105 18276 614
rect 18234 96 18290 105
rect 3790 31 3846 40
rect 5816 60 5868 66
rect 5816 2 5868 8
rect 16396 60 16448 66
rect 18432 66 18460 682
rect 18524 338 18552 1958
rect 18708 1902 18736 2926
rect 18800 2854 18828 3878
rect 18892 3534 18920 4490
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 18984 3670 19012 4014
rect 18972 3664 19024 3670
rect 18972 3606 19024 3612
rect 18880 3528 18932 3534
rect 18880 3470 18932 3476
rect 18984 3398 19012 3606
rect 18972 3392 19024 3398
rect 18972 3334 19024 3340
rect 18984 2990 19012 3334
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 18788 2848 18840 2854
rect 18788 2790 18840 2796
rect 18800 2514 18828 2790
rect 19076 2774 19104 4626
rect 19352 4468 19380 4762
rect 20180 4622 20208 4762
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 20536 4684 20588 4690
rect 20536 4626 20588 4632
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 19260 4440 19380 4468
rect 19260 4264 19288 4440
rect 19373 4380 19681 4389
rect 19373 4378 19379 4380
rect 19435 4378 19459 4380
rect 19515 4378 19539 4380
rect 19595 4378 19619 4380
rect 19675 4378 19681 4380
rect 19435 4326 19437 4378
rect 19617 4326 19619 4378
rect 19373 4324 19379 4326
rect 19435 4324 19459 4326
rect 19515 4324 19539 4326
rect 19595 4324 19619 4326
rect 19675 4324 19681 4326
rect 19373 4315 19681 4324
rect 19260 4236 19380 4264
rect 19352 3602 19380 4236
rect 19340 3596 19392 3602
rect 19392 3556 19748 3584
rect 19340 3538 19392 3544
rect 19373 3292 19681 3301
rect 19373 3290 19379 3292
rect 19435 3290 19459 3292
rect 19515 3290 19539 3292
rect 19595 3290 19619 3292
rect 19675 3290 19681 3292
rect 19435 3238 19437 3290
rect 19617 3238 19619 3290
rect 19373 3236 19379 3238
rect 19435 3236 19459 3238
rect 19515 3236 19539 3238
rect 19595 3236 19619 3238
rect 19675 3236 19681 3238
rect 19373 3227 19681 3236
rect 19076 2746 19288 2774
rect 19260 2514 19288 2746
rect 18788 2508 18840 2514
rect 18788 2450 18840 2456
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 18800 1902 18828 2450
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 19168 2106 19196 2382
rect 19246 2272 19302 2281
rect 19246 2207 19302 2216
rect 19156 2100 19208 2106
rect 19156 2042 19208 2048
rect 19260 1970 19288 2207
rect 19373 2204 19681 2213
rect 19373 2202 19379 2204
rect 19435 2202 19459 2204
rect 19515 2202 19539 2204
rect 19595 2202 19619 2204
rect 19675 2202 19681 2204
rect 19435 2150 19437 2202
rect 19617 2150 19619 2202
rect 19373 2148 19379 2150
rect 19435 2148 19459 2150
rect 19515 2148 19539 2150
rect 19595 2148 19619 2150
rect 19675 2148 19681 2150
rect 19373 2139 19681 2148
rect 19248 1964 19300 1970
rect 19248 1906 19300 1912
rect 18696 1896 18748 1902
rect 18616 1856 18696 1884
rect 18616 1358 18644 1856
rect 18696 1838 18748 1844
rect 18788 1896 18840 1902
rect 18788 1838 18840 1844
rect 19432 1896 19484 1902
rect 19432 1838 19484 1844
rect 18800 1562 18828 1838
rect 19444 1562 19472 1838
rect 18788 1556 18840 1562
rect 18788 1498 18840 1504
rect 19432 1556 19484 1562
rect 19432 1498 19484 1504
rect 18604 1352 18656 1358
rect 18604 1294 18656 1300
rect 19373 1116 19681 1125
rect 19373 1114 19379 1116
rect 19435 1114 19459 1116
rect 19515 1114 19539 1116
rect 19595 1114 19619 1116
rect 19675 1114 19681 1116
rect 19435 1062 19437 1114
rect 19617 1062 19619 1114
rect 19373 1060 19379 1062
rect 19435 1060 19459 1062
rect 19515 1060 19539 1062
rect 19595 1060 19619 1062
rect 19675 1060 19681 1062
rect 19373 1051 19681 1060
rect 18788 876 18840 882
rect 18788 818 18840 824
rect 18604 400 18656 406
rect 18604 342 18656 348
rect 18512 332 18564 338
rect 18512 274 18564 280
rect 18616 66 18644 342
rect 18800 202 18828 818
rect 18878 640 18934 649
rect 18878 575 18934 584
rect 18788 196 18840 202
rect 18788 138 18840 144
rect 18892 105 18920 575
rect 18878 96 18934 105
rect 18234 31 18290 40
rect 18420 60 18472 66
rect 16396 2 16448 8
rect 18420 2 18472 8
rect 18604 60 18656 66
rect 19720 66 19748 3556
rect 20456 2961 20484 4626
rect 20548 4282 20576 4626
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20640 3534 20668 5306
rect 21192 5166 21220 6598
rect 21284 6458 21312 6802
rect 21376 6798 21404 7296
rect 21456 7278 21508 7284
rect 21560 6866 21588 7686
rect 21744 7562 21772 7686
rect 21652 7534 21772 7562
rect 21836 7546 21864 8928
rect 22744 8910 22796 8916
rect 23572 8968 23624 8974
rect 23572 8910 23624 8916
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 21916 7880 21968 7886
rect 22008 7880 22060 7886
rect 21916 7822 21968 7828
rect 22006 7848 22008 7857
rect 22060 7848 22062 7857
rect 21824 7540 21876 7546
rect 21548 6860 21600 6866
rect 21548 6802 21600 6808
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21560 6322 21588 6598
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 21272 6248 21324 6254
rect 21272 6190 21324 6196
rect 21284 5710 21312 6190
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 21560 5914 21588 6054
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 21284 5030 21312 5646
rect 21560 5030 21588 5850
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 21272 5024 21324 5030
rect 21548 5024 21600 5030
rect 21272 4966 21324 4972
rect 21468 4984 21548 5012
rect 20732 4049 20760 4966
rect 20916 4078 20944 4966
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 21272 4480 21324 4486
rect 21272 4422 21324 4428
rect 20904 4072 20956 4078
rect 20718 4040 20774 4049
rect 20904 4014 20956 4020
rect 20718 3975 20774 3984
rect 20916 3670 20944 4014
rect 20904 3664 20956 3670
rect 20904 3606 20956 3612
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20916 2990 20944 3606
rect 21008 3097 21036 4422
rect 21284 4282 21312 4422
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 21468 4146 21496 4984
rect 21548 4966 21600 4972
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21560 4146 21588 4422
rect 21456 4140 21508 4146
rect 21456 4082 21508 4088
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 20994 3088 21050 3097
rect 21468 3058 21496 4082
rect 21652 3670 21680 7534
rect 21824 7482 21876 7488
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 21744 6662 21772 7346
rect 21732 6656 21784 6662
rect 21732 6598 21784 6604
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 21744 5574 21772 5646
rect 21732 5568 21784 5574
rect 21732 5510 21784 5516
rect 21836 4672 21864 7482
rect 21928 7206 21956 7822
rect 22006 7783 22062 7792
rect 22204 7410 22232 8774
rect 22756 8616 22784 8910
rect 22836 8628 22888 8634
rect 22756 8588 22836 8616
rect 22836 8570 22888 8576
rect 23168 8188 23476 8197
rect 23168 8186 23174 8188
rect 23230 8186 23254 8188
rect 23310 8186 23334 8188
rect 23390 8186 23414 8188
rect 23470 8186 23476 8188
rect 23230 8134 23232 8186
rect 23412 8134 23414 8186
rect 23168 8132 23174 8134
rect 23230 8132 23254 8134
rect 23310 8132 23334 8134
rect 23390 8132 23414 8134
rect 23470 8132 23476 8134
rect 23168 8123 23476 8132
rect 23584 8090 23612 8910
rect 23768 8566 23796 8978
rect 23848 8968 23900 8974
rect 23848 8910 23900 8916
rect 23756 8560 23808 8566
rect 23756 8502 23808 8508
rect 23664 8356 23716 8362
rect 23664 8298 23716 8304
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 22558 7984 22614 7993
rect 22558 7919 22560 7928
rect 22612 7919 22614 7928
rect 22560 7890 22612 7896
rect 23676 7886 23704 8298
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 21928 6798 21956 7142
rect 22008 6996 22060 7002
rect 22008 6938 22060 6944
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 22020 5234 22048 6938
rect 22112 6338 22140 7346
rect 23676 7342 23704 7822
rect 23768 7546 23796 8298
rect 23756 7540 23808 7546
rect 23756 7482 23808 7488
rect 23480 7336 23532 7342
rect 23478 7304 23480 7313
rect 23664 7336 23716 7342
rect 23532 7304 23534 7313
rect 23664 7278 23716 7284
rect 23478 7239 23534 7248
rect 23572 7268 23624 7274
rect 23572 7210 23624 7216
rect 23168 7100 23476 7109
rect 23168 7098 23174 7100
rect 23230 7098 23254 7100
rect 23310 7098 23334 7100
rect 23390 7098 23414 7100
rect 23470 7098 23476 7100
rect 23230 7046 23232 7098
rect 23412 7046 23414 7098
rect 23168 7044 23174 7046
rect 23230 7044 23254 7046
rect 23310 7044 23334 7046
rect 23390 7044 23414 7046
rect 23470 7044 23476 7046
rect 23168 7035 23476 7044
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 22190 6352 22246 6361
rect 22112 6310 22190 6338
rect 22190 6287 22246 6296
rect 23400 6225 23428 6734
rect 23584 6474 23612 7210
rect 23676 7002 23704 7278
rect 23664 6996 23716 7002
rect 23664 6938 23716 6944
rect 23492 6446 23612 6474
rect 23492 6322 23520 6446
rect 23572 6384 23624 6390
rect 23572 6326 23624 6332
rect 23480 6316 23532 6322
rect 23480 6258 23532 6264
rect 23386 6216 23442 6225
rect 23386 6151 23442 6160
rect 22928 6112 22980 6118
rect 22928 6054 22980 6060
rect 22650 5944 22706 5953
rect 22650 5879 22706 5888
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 22664 4729 22692 5879
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22650 4720 22706 4729
rect 21916 4684 21968 4690
rect 21836 4644 21916 4672
rect 22650 4655 22706 4664
rect 21916 4626 21968 4632
rect 21824 4480 21876 4486
rect 21824 4422 21876 4428
rect 21640 3664 21692 3670
rect 21640 3606 21692 3612
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21560 3194 21588 3334
rect 21548 3188 21600 3194
rect 21548 3130 21600 3136
rect 21836 3058 21864 4422
rect 21928 3534 21956 4626
rect 22756 4622 22784 4966
rect 22940 4690 22968 6054
rect 23168 6012 23476 6021
rect 23168 6010 23174 6012
rect 23230 6010 23254 6012
rect 23310 6010 23334 6012
rect 23390 6010 23414 6012
rect 23470 6010 23476 6012
rect 23230 5958 23232 6010
rect 23412 5958 23414 6010
rect 23168 5956 23174 5958
rect 23230 5956 23254 5958
rect 23310 5956 23334 5958
rect 23390 5956 23414 5958
rect 23470 5956 23476 5958
rect 23168 5947 23476 5956
rect 23110 5672 23166 5681
rect 23110 5607 23166 5616
rect 23124 5370 23152 5607
rect 23388 5568 23440 5574
rect 23388 5510 23440 5516
rect 23112 5364 23164 5370
rect 23112 5306 23164 5312
rect 23400 5166 23428 5510
rect 23584 5166 23612 6326
rect 23756 6248 23808 6254
rect 23860 6236 23888 8910
rect 23952 8430 23980 9114
rect 23940 8424 23992 8430
rect 23940 8366 23992 8372
rect 24136 6866 24164 9522
rect 24216 9376 24268 9382
rect 24216 9318 24268 9324
rect 24228 8430 24256 9318
rect 24216 8424 24268 8430
rect 24216 8366 24268 8372
rect 24124 6860 24176 6866
rect 24124 6802 24176 6808
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 23808 6208 23888 6236
rect 23940 6248 23992 6254
rect 23756 6190 23808 6196
rect 24044 6202 24072 6734
rect 23992 6196 24072 6202
rect 23940 6190 24072 6196
rect 23664 5704 23716 5710
rect 23664 5646 23716 5652
rect 23676 5166 23704 5646
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 23572 5160 23624 5166
rect 23572 5102 23624 5108
rect 23664 5160 23716 5166
rect 23664 5102 23716 5108
rect 23168 4924 23476 4933
rect 23168 4922 23174 4924
rect 23230 4922 23254 4924
rect 23310 4922 23334 4924
rect 23390 4922 23414 4924
rect 23470 4922 23476 4924
rect 23230 4870 23232 4922
rect 23412 4870 23414 4922
rect 23168 4868 23174 4870
rect 23230 4868 23254 4870
rect 23310 4868 23334 4870
rect 23390 4868 23414 4870
rect 23470 4868 23476 4870
rect 23168 4859 23476 4868
rect 23584 4690 23612 5102
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 23572 4684 23624 4690
rect 23572 4626 23624 4632
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22192 4548 22244 4554
rect 22192 4490 22244 4496
rect 22008 4480 22060 4486
rect 22008 4422 22060 4428
rect 22020 4146 22048 4422
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 22204 3534 22232 4490
rect 22572 4010 22600 4558
rect 23664 4480 23716 4486
rect 23584 4440 23664 4468
rect 23584 4078 23612 4440
rect 23664 4422 23716 4428
rect 23768 4078 23796 6190
rect 23952 6174 24072 6190
rect 24044 5953 24072 6174
rect 24124 6180 24176 6186
rect 24124 6122 24176 6128
rect 24030 5944 24086 5953
rect 23940 5908 23992 5914
rect 24030 5879 24086 5888
rect 23940 5850 23992 5856
rect 23952 5098 23980 5850
rect 24136 5234 24164 6122
rect 24216 5704 24268 5710
rect 24216 5646 24268 5652
rect 24228 5574 24256 5646
rect 24216 5568 24268 5574
rect 24216 5510 24268 5516
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 23940 5092 23992 5098
rect 23940 5034 23992 5040
rect 23848 5024 23900 5030
rect 23848 4966 23900 4972
rect 24124 5024 24176 5030
rect 24124 4966 24176 4972
rect 23572 4072 23624 4078
rect 23572 4014 23624 4020
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 22560 4004 22612 4010
rect 22560 3946 22612 3952
rect 22572 3602 22600 3946
rect 22744 3936 22796 3942
rect 22744 3878 22796 3884
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 22560 3596 22612 3602
rect 22560 3538 22612 3544
rect 22756 3534 22784 3878
rect 22940 3602 22968 3878
rect 23168 3836 23476 3845
rect 23168 3834 23174 3836
rect 23230 3834 23254 3836
rect 23310 3834 23334 3836
rect 23390 3834 23414 3836
rect 23470 3834 23476 3836
rect 23230 3782 23232 3834
rect 23412 3782 23414 3834
rect 23168 3780 23174 3782
rect 23230 3780 23254 3782
rect 23310 3780 23334 3782
rect 23390 3780 23414 3782
rect 23470 3780 23476 3782
rect 23168 3771 23476 3780
rect 23570 3768 23626 3777
rect 23570 3703 23626 3712
rect 22928 3596 22980 3602
rect 22928 3538 22980 3544
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 22192 3528 22244 3534
rect 22192 3470 22244 3476
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 20994 3023 21050 3032
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 20904 2984 20956 2990
rect 20442 2952 20498 2961
rect 20904 2926 20956 2932
rect 20442 2887 20498 2896
rect 20534 2680 20590 2689
rect 20534 2615 20590 2624
rect 20548 2582 20576 2615
rect 20536 2576 20588 2582
rect 20536 2518 20588 2524
rect 20916 2514 20944 2926
rect 20904 2508 20956 2514
rect 20904 2450 20956 2456
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20534 1728 20590 1737
rect 20534 1663 20590 1672
rect 20444 1012 20496 1018
rect 20444 954 20496 960
rect 20456 746 20484 954
rect 20444 740 20496 746
rect 20444 682 20496 688
rect 20548 678 20576 1663
rect 20640 1222 20668 2246
rect 20720 1964 20772 1970
rect 20720 1906 20772 1912
rect 20628 1216 20680 1222
rect 20628 1158 20680 1164
rect 20732 1034 20760 1906
rect 20824 1426 20852 2246
rect 20916 1902 20944 2450
rect 21468 2446 21496 2994
rect 21822 2680 21878 2689
rect 21640 2644 21692 2650
rect 21822 2615 21878 2624
rect 21640 2586 21692 2592
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 21088 2372 21140 2378
rect 21088 2314 21140 2320
rect 21100 2281 21128 2314
rect 21086 2272 21142 2281
rect 21086 2207 21142 2216
rect 21468 1970 21496 2382
rect 21652 2145 21680 2586
rect 21836 2446 21864 2615
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 21638 2136 21694 2145
rect 21638 2071 21694 2080
rect 21456 1964 21508 1970
rect 21456 1906 21508 1912
rect 20904 1896 20956 1902
rect 20904 1838 20956 1844
rect 20916 1442 20944 1838
rect 20994 1592 21050 1601
rect 21050 1550 21128 1578
rect 20994 1527 21050 1536
rect 20812 1420 20864 1426
rect 20916 1414 21036 1442
rect 21100 1426 21128 1550
rect 21468 1544 21496 1906
rect 21548 1556 21600 1562
rect 21468 1516 21548 1544
rect 21548 1498 21600 1504
rect 20812 1362 20864 1368
rect 21008 1358 21036 1414
rect 21088 1420 21140 1426
rect 21088 1362 21140 1368
rect 20996 1352 21048 1358
rect 20996 1294 21048 1300
rect 20904 1284 20956 1290
rect 20904 1226 20956 1232
rect 20732 1006 20852 1034
rect 20824 882 20852 1006
rect 20916 950 20944 1226
rect 21546 1048 21602 1057
rect 21546 983 21602 992
rect 20904 944 20956 950
rect 20904 886 20956 892
rect 21560 882 21588 983
rect 20812 876 20864 882
rect 20812 818 20864 824
rect 21548 876 21600 882
rect 21548 818 21600 824
rect 21652 814 21680 2071
rect 21928 1766 21956 3470
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 22112 3194 22140 3334
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 22020 2650 22048 2926
rect 23168 2748 23476 2757
rect 23168 2746 23174 2748
rect 23230 2746 23254 2748
rect 23310 2746 23334 2748
rect 23390 2746 23414 2748
rect 23470 2746 23476 2748
rect 23230 2694 23232 2746
rect 23412 2694 23414 2746
rect 23168 2692 23174 2694
rect 23230 2692 23254 2694
rect 23310 2692 23334 2694
rect 23390 2692 23414 2694
rect 23470 2692 23476 2694
rect 23168 2683 23476 2692
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 22744 2508 22796 2514
rect 22744 2450 22796 2456
rect 22652 1828 22704 1834
rect 22652 1770 22704 1776
rect 21916 1760 21968 1766
rect 21916 1702 21968 1708
rect 22664 1601 22692 1770
rect 22650 1592 22706 1601
rect 22650 1527 22706 1536
rect 21272 808 21324 814
rect 21272 750 21324 756
rect 21640 808 21692 814
rect 21640 750 21692 756
rect 20536 672 20588 678
rect 20536 614 20588 620
rect 20812 672 20864 678
rect 20812 614 20864 620
rect 20824 513 20852 614
rect 20810 504 20866 513
rect 20720 468 20772 474
rect 20810 439 20866 448
rect 20720 410 20772 416
rect 20732 377 20760 410
rect 20718 368 20774 377
rect 20718 303 20774 312
rect 21284 270 21312 750
rect 21272 264 21324 270
rect 21272 206 21324 212
rect 22756 134 22784 2450
rect 22836 2440 22888 2446
rect 22836 2382 22888 2388
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 22848 338 22876 2382
rect 22940 1737 22968 2382
rect 23020 2032 23072 2038
rect 23020 1974 23072 1980
rect 22926 1728 22982 1737
rect 22926 1663 22982 1672
rect 23032 1222 23060 1974
rect 23112 1964 23164 1970
rect 23112 1906 23164 1912
rect 23124 1766 23152 1906
rect 23584 1873 23612 3703
rect 23664 2372 23716 2378
rect 23664 2314 23716 2320
rect 23676 1970 23704 2314
rect 23768 2038 23796 4014
rect 23860 3398 23888 4966
rect 24136 4536 24164 4966
rect 24320 4706 24348 13359
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 24492 13320 24544 13326
rect 24596 13308 24624 13738
rect 24676 13320 24728 13326
rect 24596 13280 24676 13308
rect 24492 13262 24544 13268
rect 24676 13262 24728 13268
rect 24412 12782 24440 13262
rect 24504 12986 24532 13262
rect 24492 12980 24544 12986
rect 24492 12922 24544 12928
rect 24490 12880 24546 12889
rect 24490 12815 24492 12824
rect 24544 12815 24546 12824
rect 24492 12786 24544 12792
rect 24400 12776 24452 12782
rect 24400 12718 24452 12724
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24688 11694 24716 11834
rect 24676 11688 24728 11694
rect 24676 11630 24728 11636
rect 24400 11620 24452 11626
rect 24400 11562 24452 11568
rect 24768 11620 24820 11626
rect 24768 11562 24820 11568
rect 24412 11150 24440 11562
rect 24780 11218 24808 11562
rect 24768 11212 24820 11218
rect 24768 11154 24820 11160
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24860 11144 24912 11150
rect 24860 11086 24912 11092
rect 24872 10810 24900 11086
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 24964 10690 24992 14962
rect 25148 10810 25176 17002
rect 25332 14770 25360 18527
rect 25412 18216 25464 18222
rect 25412 18158 25464 18164
rect 25424 17338 25452 18158
rect 25976 17762 26004 20334
rect 26068 19310 26096 20878
rect 26056 19304 26108 19310
rect 26056 19246 26108 19252
rect 25700 17734 26004 17762
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25410 14784 25466 14793
rect 25332 14742 25410 14770
rect 25410 14719 25466 14728
rect 25424 14618 25452 14719
rect 25412 14612 25464 14618
rect 25412 14554 25464 14560
rect 25700 13954 25728 17734
rect 25964 17672 26016 17678
rect 25778 17640 25834 17649
rect 25964 17614 26016 17620
rect 25778 17575 25834 17584
rect 25792 17134 25820 17575
rect 25976 17134 26004 17614
rect 25780 17128 25832 17134
rect 25780 17070 25832 17076
rect 25964 17128 26016 17134
rect 25964 17070 26016 17076
rect 25872 16652 25924 16658
rect 25872 16594 25924 16600
rect 25778 14512 25834 14521
rect 25778 14447 25834 14456
rect 25608 13926 25728 13954
rect 25608 13734 25636 13926
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 25320 13728 25372 13734
rect 25320 13670 25372 13676
rect 25596 13728 25648 13734
rect 25596 13670 25648 13676
rect 25332 13530 25360 13670
rect 25320 13524 25372 13530
rect 25320 13466 25372 13472
rect 25700 12986 25728 13806
rect 25688 12980 25740 12986
rect 25688 12922 25740 12928
rect 25792 12442 25820 14447
rect 25780 12436 25832 12442
rect 25780 12378 25832 12384
rect 25412 12300 25464 12306
rect 25412 12242 25464 12248
rect 25136 10804 25188 10810
rect 25136 10746 25188 10752
rect 24872 10662 24992 10690
rect 24492 10464 24544 10470
rect 24492 10406 24544 10412
rect 24504 10130 24532 10406
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24676 10056 24728 10062
rect 24676 9998 24728 10004
rect 24688 9926 24716 9998
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24492 9512 24544 9518
rect 24492 9454 24544 9460
rect 24504 9382 24532 9454
rect 24492 9376 24544 9382
rect 24492 9318 24544 9324
rect 24492 8832 24544 8838
rect 24492 8774 24544 8780
rect 24504 8498 24532 8774
rect 24492 8492 24544 8498
rect 24492 8434 24544 8440
rect 24676 8424 24728 8430
rect 24596 8384 24676 8412
rect 24492 7880 24544 7886
rect 24492 7822 24544 7828
rect 24504 7206 24532 7822
rect 24596 7410 24624 8384
rect 24676 8366 24728 8372
rect 24780 7750 24808 10202
rect 24872 9489 24900 10662
rect 25320 10600 25372 10606
rect 25320 10542 25372 10548
rect 24952 10124 25004 10130
rect 24952 10066 25004 10072
rect 24858 9480 24914 9489
rect 24858 9415 24914 9424
rect 24872 9110 24900 9415
rect 24860 9104 24912 9110
rect 24860 9046 24912 9052
rect 24964 8838 24992 10066
rect 24952 8832 25004 8838
rect 24952 8774 25004 8780
rect 25332 8634 25360 10542
rect 25320 8628 25372 8634
rect 25320 8570 25372 8576
rect 24676 7744 24728 7750
rect 24676 7686 24728 7692
rect 24768 7744 24820 7750
rect 24768 7686 24820 7692
rect 24688 7410 24716 7686
rect 25136 7540 25188 7546
rect 25136 7482 25188 7488
rect 25148 7449 25176 7482
rect 25134 7440 25190 7449
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 24676 7404 24728 7410
rect 25134 7375 25190 7384
rect 24676 7346 24728 7352
rect 24768 7336 24820 7342
rect 24768 7278 24820 7284
rect 24492 7200 24544 7206
rect 24492 7142 24544 7148
rect 24582 6896 24638 6905
rect 24582 6831 24638 6840
rect 24492 6792 24544 6798
rect 24492 6734 24544 6740
rect 24504 4826 24532 6734
rect 24492 4820 24544 4826
rect 24492 4762 24544 4768
rect 24044 4508 24164 4536
rect 24228 4678 24348 4706
rect 24044 3942 24072 4508
rect 24228 4078 24256 4678
rect 24596 4078 24624 6831
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24688 6338 24716 6734
rect 24780 6458 24808 7278
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 25240 6458 25268 6598
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 24688 6310 24808 6338
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 24688 5778 24716 6190
rect 24780 6118 24808 6310
rect 24860 6248 24912 6254
rect 24860 6190 24912 6196
rect 24768 6112 24820 6118
rect 24768 6054 24820 6060
rect 24676 5772 24728 5778
rect 24780 5760 24808 6054
rect 24872 5914 24900 6190
rect 24860 5908 24912 5914
rect 24860 5850 24912 5856
rect 24952 5772 25004 5778
rect 24780 5732 24952 5760
rect 24676 5714 24728 5720
rect 24952 5714 25004 5720
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24780 4486 24808 5306
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24216 4072 24268 4078
rect 24216 4014 24268 4020
rect 24584 4072 24636 4078
rect 24584 4014 24636 4020
rect 24032 3936 24084 3942
rect 24032 3878 24084 3884
rect 24124 3936 24176 3942
rect 24124 3878 24176 3884
rect 24400 3936 24452 3942
rect 24400 3878 24452 3884
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 23848 3392 23900 3398
rect 23848 3334 23900 3340
rect 23860 2990 23888 3334
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 23860 2650 23888 2926
rect 24044 2836 24072 3878
rect 24136 3482 24164 3878
rect 24412 3482 24440 3878
rect 24136 3454 24348 3482
rect 24412 3454 24624 3482
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24124 2848 24176 2854
rect 24044 2808 24124 2836
rect 24124 2790 24176 2796
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 23756 2032 23808 2038
rect 23756 1974 23808 1980
rect 23664 1964 23716 1970
rect 23664 1906 23716 1912
rect 23570 1864 23626 1873
rect 23570 1799 23626 1808
rect 23112 1760 23164 1766
rect 23112 1702 23164 1708
rect 23676 1714 23704 1906
rect 23768 1873 23796 1974
rect 23860 1902 23888 2586
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 23940 2304 23992 2310
rect 23940 2246 23992 2252
rect 23848 1896 23900 1902
rect 23754 1864 23810 1873
rect 23848 1838 23900 1844
rect 23754 1799 23810 1808
rect 23754 1728 23810 1737
rect 23676 1686 23754 1714
rect 23168 1660 23476 1669
rect 23754 1663 23810 1672
rect 23168 1658 23174 1660
rect 23230 1658 23254 1660
rect 23310 1658 23334 1660
rect 23390 1658 23414 1660
rect 23470 1658 23476 1660
rect 23230 1606 23232 1658
rect 23412 1606 23414 1658
rect 23168 1604 23174 1606
rect 23230 1604 23254 1606
rect 23310 1604 23334 1606
rect 23390 1604 23414 1606
rect 23470 1604 23476 1606
rect 23168 1595 23476 1604
rect 23572 1488 23624 1494
rect 23572 1430 23624 1436
rect 23020 1216 23072 1222
rect 23020 1158 23072 1164
rect 23388 1216 23440 1222
rect 23478 1184 23534 1193
rect 23440 1164 23478 1170
rect 23388 1158 23478 1164
rect 23400 1142 23478 1158
rect 23478 1119 23534 1128
rect 23584 882 23612 1430
rect 23664 1352 23716 1358
rect 23860 1306 23888 1838
rect 23952 1358 23980 2246
rect 23716 1300 23888 1306
rect 23664 1294 23888 1300
rect 23940 1352 23992 1358
rect 23940 1294 23992 1300
rect 23676 1278 23888 1294
rect 23662 912 23718 921
rect 23572 876 23624 882
rect 23662 847 23718 856
rect 23572 818 23624 824
rect 23676 814 23704 847
rect 23860 814 23888 1278
rect 24044 1222 24072 2450
rect 24136 1766 24164 2790
rect 24228 2650 24256 3334
rect 24320 2774 24348 3454
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24504 3058 24532 3334
rect 24492 3052 24544 3058
rect 24492 2994 24544 3000
rect 24320 2746 24532 2774
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 24400 2440 24452 2446
rect 24398 2408 24400 2417
rect 24452 2408 24454 2417
rect 24398 2343 24454 2352
rect 24504 1970 24532 2746
rect 24596 2394 24624 3454
rect 24688 2553 24716 3878
rect 24780 3602 24808 4422
rect 24860 4072 24912 4078
rect 24860 4014 24912 4020
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 24872 3233 24900 4014
rect 24964 3534 24992 5714
rect 25424 5370 25452 12242
rect 25688 11688 25740 11694
rect 25688 11630 25740 11636
rect 25700 11354 25728 11630
rect 25688 11348 25740 11354
rect 25688 11290 25740 11296
rect 25884 11257 25912 16594
rect 25976 16046 26004 17070
rect 26068 16980 26096 19246
rect 26160 18698 26188 21354
rect 26252 20074 26280 21422
rect 26424 21344 26476 21350
rect 26424 21286 26476 21292
rect 26332 20936 26384 20942
rect 26332 20878 26384 20884
rect 26344 20534 26372 20878
rect 26332 20528 26384 20534
rect 26332 20470 26384 20476
rect 26252 20046 26372 20074
rect 26240 19236 26292 19242
rect 26240 19178 26292 19184
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 26252 17338 26280 19178
rect 26344 18766 26372 20046
rect 26436 19514 26464 21286
rect 26424 19508 26476 19514
rect 26424 19450 26476 19456
rect 26516 19168 26568 19174
rect 26516 19110 26568 19116
rect 26700 19168 26752 19174
rect 26700 19110 26752 19116
rect 26332 18760 26384 18766
rect 26332 18702 26384 18708
rect 26344 17678 26372 18702
rect 26528 18465 26556 19110
rect 26514 18456 26570 18465
rect 26514 18391 26570 18400
rect 26608 18216 26660 18222
rect 26608 18158 26660 18164
rect 26424 18080 26476 18086
rect 26424 18022 26476 18028
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26240 17332 26292 17338
rect 26240 17274 26292 17280
rect 26148 16992 26200 16998
rect 26068 16952 26148 16980
rect 26148 16934 26200 16940
rect 26238 16960 26294 16969
rect 26056 16448 26108 16454
rect 26056 16390 26108 16396
rect 25964 16040 26016 16046
rect 25964 15982 26016 15988
rect 26068 15570 26096 16390
rect 26056 15564 26108 15570
rect 26056 15506 26108 15512
rect 25964 15360 26016 15366
rect 25964 15302 26016 15308
rect 25976 14482 26004 15302
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 25976 12306 26004 14418
rect 26068 13977 26096 15506
rect 26160 15484 26188 16934
rect 26238 16895 26294 16904
rect 26252 15638 26280 16895
rect 26344 16561 26372 17478
rect 26436 16794 26464 18022
rect 26516 17876 26568 17882
rect 26516 17818 26568 17824
rect 26424 16788 26476 16794
rect 26424 16730 26476 16736
rect 26330 16552 26386 16561
rect 26330 16487 26386 16496
rect 26332 16448 26384 16454
rect 26332 16390 26384 16396
rect 26344 15910 26372 16390
rect 26332 15904 26384 15910
rect 26332 15846 26384 15852
rect 26240 15632 26292 15638
rect 26240 15574 26292 15580
rect 26240 15496 26292 15502
rect 26160 15456 26240 15484
rect 26240 15438 26292 15444
rect 26528 15162 26556 17818
rect 26620 16250 26648 18158
rect 26712 17377 26740 19110
rect 26804 18970 26832 21422
rect 26963 20700 27271 20709
rect 26963 20698 26969 20700
rect 27025 20698 27049 20700
rect 27105 20698 27129 20700
rect 27185 20698 27209 20700
rect 27265 20698 27271 20700
rect 27025 20646 27027 20698
rect 27207 20646 27209 20698
rect 26963 20644 26969 20646
rect 27025 20644 27049 20646
rect 27105 20644 27129 20646
rect 27185 20644 27209 20646
rect 27265 20644 27271 20646
rect 26963 20635 27271 20644
rect 27344 20392 27396 20398
rect 27344 20334 27396 20340
rect 27356 19922 27384 20334
rect 27344 19916 27396 19922
rect 27344 19858 27396 19864
rect 26884 19848 26936 19854
rect 26884 19790 26936 19796
rect 26896 19310 26924 19790
rect 26963 19612 27271 19621
rect 26963 19610 26969 19612
rect 27025 19610 27049 19612
rect 27105 19610 27129 19612
rect 27185 19610 27209 19612
rect 27265 19610 27271 19612
rect 27025 19558 27027 19610
rect 27207 19558 27209 19610
rect 26963 19556 26969 19558
rect 27025 19556 27049 19558
rect 27105 19556 27129 19558
rect 27185 19556 27209 19558
rect 27265 19556 27271 19558
rect 26963 19547 27271 19556
rect 27356 19334 27384 19858
rect 27540 19854 27568 21490
rect 27896 21480 27948 21486
rect 27896 21422 27948 21428
rect 27528 19848 27580 19854
rect 27528 19790 27580 19796
rect 26884 19304 26936 19310
rect 27356 19306 27476 19334
rect 26884 19246 26936 19252
rect 26792 18964 26844 18970
rect 26792 18906 26844 18912
rect 26804 17746 26832 18906
rect 26896 18290 26924 19246
rect 27068 18760 27120 18766
rect 27068 18702 27120 18708
rect 27080 18630 27108 18702
rect 27068 18624 27120 18630
rect 27068 18566 27120 18572
rect 26963 18524 27271 18533
rect 26963 18522 26969 18524
rect 27025 18522 27049 18524
rect 27105 18522 27129 18524
rect 27185 18522 27209 18524
rect 27265 18522 27271 18524
rect 27025 18470 27027 18522
rect 27207 18470 27209 18522
rect 26963 18468 26969 18470
rect 27025 18468 27049 18470
rect 27105 18468 27129 18470
rect 27185 18468 27209 18470
rect 27265 18468 27271 18470
rect 26963 18459 27271 18468
rect 26884 18284 26936 18290
rect 26884 18226 26936 18232
rect 27160 17876 27212 17882
rect 27160 17818 27212 17824
rect 27172 17746 27200 17818
rect 26792 17740 26844 17746
rect 26792 17682 26844 17688
rect 27160 17740 27212 17746
rect 27160 17682 27212 17688
rect 26698 17368 26754 17377
rect 26698 17303 26754 17312
rect 26700 16992 26752 16998
rect 26804 16980 26832 17682
rect 26884 17672 26936 17678
rect 26884 17614 26936 17620
rect 26752 16952 26832 16980
rect 26700 16934 26752 16940
rect 26608 16244 26660 16250
rect 26608 16186 26660 16192
rect 26712 16046 26740 16934
rect 26792 16448 26844 16454
rect 26792 16390 26844 16396
rect 26804 16250 26832 16390
rect 26792 16244 26844 16250
rect 26792 16186 26844 16192
rect 26700 16040 26752 16046
rect 26620 16000 26700 16028
rect 26620 15638 26648 16000
rect 26700 15982 26752 15988
rect 26792 16040 26844 16046
rect 26792 15982 26844 15988
rect 26700 15904 26752 15910
rect 26700 15846 26752 15852
rect 26608 15632 26660 15638
rect 26608 15574 26660 15580
rect 26712 15201 26740 15846
rect 26804 15706 26832 15982
rect 26792 15700 26844 15706
rect 26792 15642 26844 15648
rect 26792 15428 26844 15434
rect 26792 15370 26844 15376
rect 26698 15192 26754 15201
rect 26516 15156 26568 15162
rect 26698 15127 26754 15136
rect 26516 15098 26568 15104
rect 26424 15088 26476 15094
rect 26424 15030 26476 15036
rect 26148 14816 26200 14822
rect 26148 14758 26200 14764
rect 26054 13968 26110 13977
rect 26054 13903 26110 13912
rect 26160 13870 26188 14758
rect 26436 14482 26464 15030
rect 26804 14958 26832 15370
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26792 14952 26844 14958
rect 26792 14894 26844 14900
rect 26424 14476 26476 14482
rect 26424 14418 26476 14424
rect 26436 13870 26464 14418
rect 26148 13864 26200 13870
rect 26148 13806 26200 13812
rect 26424 13864 26476 13870
rect 26424 13806 26476 13812
rect 26056 13728 26108 13734
rect 26056 13670 26108 13676
rect 26068 13433 26096 13670
rect 26436 13530 26464 13806
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 26054 13424 26110 13433
rect 26054 13359 26110 13368
rect 26344 13376 26372 13466
rect 26516 13388 26568 13394
rect 25964 12300 26016 12306
rect 25964 12242 26016 12248
rect 26068 11762 26096 13359
rect 26344 13348 26516 13376
rect 26516 13330 26568 13336
rect 26620 12986 26648 14894
rect 26700 14476 26752 14482
rect 26700 14418 26752 14424
rect 26712 13512 26740 14418
rect 26792 14272 26844 14278
rect 26792 14214 26844 14220
rect 26804 13954 26832 14214
rect 26896 14074 26924 17614
rect 26963 17436 27271 17445
rect 26963 17434 26969 17436
rect 27025 17434 27049 17436
rect 27105 17434 27129 17436
rect 27185 17434 27209 17436
rect 27265 17434 27271 17436
rect 27025 17382 27027 17434
rect 27207 17382 27209 17434
rect 26963 17380 26969 17382
rect 27025 17380 27049 17382
rect 27105 17380 27129 17382
rect 27185 17380 27209 17382
rect 27265 17380 27271 17382
rect 26963 17371 27271 17380
rect 27252 17332 27304 17338
rect 27252 17274 27304 17280
rect 27264 17241 27292 17274
rect 27250 17232 27306 17241
rect 27250 17167 27306 17176
rect 27344 17128 27396 17134
rect 27344 17070 27396 17076
rect 27252 16992 27304 16998
rect 27158 16960 27214 16969
rect 27214 16940 27252 16946
rect 27214 16934 27304 16940
rect 27214 16918 27292 16934
rect 27158 16895 27214 16904
rect 27172 16454 27200 16895
rect 27160 16448 27212 16454
rect 27160 16390 27212 16396
rect 26963 16348 27271 16357
rect 26963 16346 26969 16348
rect 27025 16346 27049 16348
rect 27105 16346 27129 16348
rect 27185 16346 27209 16348
rect 27265 16346 27271 16348
rect 27025 16294 27027 16346
rect 27207 16294 27209 16346
rect 26963 16292 26969 16294
rect 27025 16292 27049 16294
rect 27105 16292 27129 16294
rect 27185 16292 27209 16294
rect 27265 16292 27271 16294
rect 26963 16283 27271 16292
rect 27252 16040 27304 16046
rect 27252 15982 27304 15988
rect 27264 15348 27292 15982
rect 27356 15706 27384 17070
rect 27448 16658 27476 19306
rect 27620 18624 27672 18630
rect 27620 18566 27672 18572
rect 27804 18624 27856 18630
rect 27804 18566 27856 18572
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27436 16652 27488 16658
rect 27436 16594 27488 16600
rect 27448 16046 27476 16594
rect 27436 16040 27488 16046
rect 27436 15982 27488 15988
rect 27434 15736 27490 15745
rect 27344 15700 27396 15706
rect 27434 15671 27490 15680
rect 27344 15642 27396 15648
rect 27264 15320 27384 15348
rect 26963 15260 27271 15269
rect 26963 15258 26969 15260
rect 27025 15258 27049 15260
rect 27105 15258 27129 15260
rect 27185 15258 27209 15260
rect 27265 15258 27271 15260
rect 27025 15206 27027 15258
rect 27207 15206 27209 15258
rect 26963 15204 26969 15206
rect 27025 15204 27049 15206
rect 27105 15204 27129 15206
rect 27185 15204 27209 15206
rect 27265 15204 27271 15206
rect 26963 15195 27271 15204
rect 27356 15162 27384 15320
rect 27344 15156 27396 15162
rect 27344 15098 27396 15104
rect 27068 15020 27120 15026
rect 27252 15020 27304 15026
rect 27120 14980 27252 15008
rect 27068 14962 27120 14968
rect 27252 14962 27304 14968
rect 27344 14952 27396 14958
rect 27344 14894 27396 14900
rect 26976 14612 27028 14618
rect 26976 14554 27028 14560
rect 26988 14278 27016 14554
rect 27066 14512 27122 14521
rect 27066 14447 27122 14456
rect 27080 14414 27108 14447
rect 27068 14408 27120 14414
rect 27068 14350 27120 14356
rect 26976 14272 27028 14278
rect 26976 14214 27028 14220
rect 26963 14172 27271 14181
rect 26963 14170 26969 14172
rect 27025 14170 27049 14172
rect 27105 14170 27129 14172
rect 27185 14170 27209 14172
rect 27265 14170 27271 14172
rect 27025 14118 27027 14170
rect 27207 14118 27209 14170
rect 26963 14116 26969 14118
rect 27025 14116 27049 14118
rect 27105 14116 27129 14118
rect 27185 14116 27209 14118
rect 27265 14116 27271 14118
rect 26963 14107 27271 14116
rect 26884 14068 26936 14074
rect 26884 14010 26936 14016
rect 26804 13938 26924 13954
rect 26804 13932 26936 13938
rect 26804 13926 26884 13932
rect 26884 13874 26936 13880
rect 27068 13728 27120 13734
rect 27068 13670 27120 13676
rect 27080 13530 27108 13670
rect 26884 13524 26936 13530
rect 26712 13484 26884 13512
rect 26884 13466 26936 13472
rect 27068 13524 27120 13530
rect 27068 13466 27120 13472
rect 26963 13084 27271 13093
rect 26963 13082 26969 13084
rect 27025 13082 27049 13084
rect 27105 13082 27129 13084
rect 27185 13082 27209 13084
rect 27265 13082 27271 13084
rect 27025 13030 27027 13082
rect 27207 13030 27209 13082
rect 26963 13028 26969 13030
rect 27025 13028 27049 13030
rect 27105 13028 27129 13030
rect 27185 13028 27209 13030
rect 27265 13028 27271 13030
rect 26963 13019 27271 13028
rect 26608 12980 26660 12986
rect 26608 12922 26660 12928
rect 26424 12776 26476 12782
rect 26424 12718 26476 12724
rect 26148 12640 26200 12646
rect 26148 12582 26200 12588
rect 26160 12442 26188 12582
rect 26148 12436 26200 12442
rect 26148 12378 26200 12384
rect 26160 12306 26188 12378
rect 26436 12306 26464 12718
rect 26516 12640 26568 12646
rect 26516 12582 26568 12588
rect 26148 12300 26200 12306
rect 26148 12242 26200 12248
rect 26424 12300 26476 12306
rect 26424 12242 26476 12248
rect 26528 11898 26556 12582
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 26516 11892 26568 11898
rect 26516 11834 26568 11840
rect 26792 11892 26844 11898
rect 26896 11880 26924 12174
rect 26963 11996 27271 12005
rect 26963 11994 26969 11996
rect 27025 11994 27049 11996
rect 27105 11994 27129 11996
rect 27185 11994 27209 11996
rect 27265 11994 27271 11996
rect 27025 11942 27027 11994
rect 27207 11942 27209 11994
rect 26963 11940 26969 11942
rect 27025 11940 27049 11942
rect 27105 11940 27129 11942
rect 27185 11940 27209 11942
rect 27265 11940 27271 11942
rect 26963 11931 27271 11940
rect 26844 11852 26924 11880
rect 26792 11834 26844 11840
rect 26056 11756 26108 11762
rect 26056 11698 26108 11704
rect 26054 11656 26110 11665
rect 26054 11591 26110 11600
rect 25870 11248 25926 11257
rect 25870 11183 25926 11192
rect 25688 10804 25740 10810
rect 25608 10764 25688 10792
rect 25412 5364 25464 5370
rect 25412 5306 25464 5312
rect 25228 4616 25280 4622
rect 25134 4584 25190 4593
rect 25228 4558 25280 4564
rect 25134 4519 25190 4528
rect 25044 4480 25096 4486
rect 25044 4422 25096 4428
rect 24952 3528 25004 3534
rect 24952 3470 25004 3476
rect 24858 3224 24914 3233
rect 24858 3159 24914 3168
rect 24964 3108 24992 3470
rect 24872 3080 24992 3108
rect 24674 2544 24730 2553
rect 24674 2479 24730 2488
rect 24872 2417 24900 3080
rect 25056 2774 25084 4422
rect 24964 2746 25084 2774
rect 24964 2689 24992 2746
rect 24950 2680 25006 2689
rect 24950 2615 25006 2624
rect 24964 2446 24992 2615
rect 24952 2440 25004 2446
rect 24858 2408 24914 2417
rect 24596 2366 24716 2394
rect 24584 2304 24636 2310
rect 24584 2246 24636 2252
rect 24492 1964 24544 1970
rect 24492 1906 24544 1912
rect 24124 1760 24176 1766
rect 24124 1702 24176 1708
rect 24492 1760 24544 1766
rect 24492 1702 24544 1708
rect 24136 1358 24164 1702
rect 24124 1352 24176 1358
rect 24124 1294 24176 1300
rect 24032 1216 24084 1222
rect 24032 1158 24084 1164
rect 23020 808 23072 814
rect 23020 750 23072 756
rect 23664 808 23716 814
rect 23664 750 23716 756
rect 23848 808 23900 814
rect 23848 750 23900 756
rect 23032 406 23060 750
rect 23756 740 23808 746
rect 23756 682 23808 688
rect 23168 572 23476 581
rect 23168 570 23174 572
rect 23230 570 23254 572
rect 23310 570 23334 572
rect 23390 570 23414 572
rect 23470 570 23476 572
rect 23230 518 23232 570
rect 23412 518 23414 570
rect 23168 516 23174 518
rect 23230 516 23254 518
rect 23310 516 23334 518
rect 23390 516 23414 518
rect 23470 516 23476 518
rect 23168 507 23476 516
rect 23768 474 23796 682
rect 24136 678 24164 1294
rect 24504 814 24532 1702
rect 24596 882 24624 2246
rect 24688 1601 24716 2366
rect 24952 2382 25004 2388
rect 24858 2343 24914 2352
rect 24674 1592 24730 1601
rect 24674 1527 24730 1536
rect 24872 1426 24900 2343
rect 24952 1488 25004 1494
rect 24952 1430 25004 1436
rect 24860 1420 24912 1426
rect 24860 1362 24912 1368
rect 24964 1057 24992 1430
rect 24950 1048 25006 1057
rect 24950 983 25006 992
rect 24584 876 24636 882
rect 25148 864 25176 4519
rect 25240 3670 25268 4558
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 25228 3664 25280 3670
rect 25516 3641 25544 3878
rect 25228 3606 25280 3612
rect 25502 3632 25558 3641
rect 25608 3602 25636 10764
rect 25688 10746 25740 10752
rect 25688 10600 25740 10606
rect 25688 10542 25740 10548
rect 25700 9722 25728 10542
rect 26068 10538 26096 11591
rect 26332 11212 26384 11218
rect 26332 11154 26384 11160
rect 26056 10532 26108 10538
rect 26056 10474 26108 10480
rect 26240 10464 26292 10470
rect 26240 10406 26292 10412
rect 25688 9716 25740 9722
rect 25688 9658 25740 9664
rect 26252 9586 26280 10406
rect 26240 9580 26292 9586
rect 26240 9522 26292 9528
rect 25688 9512 25740 9518
rect 25688 9454 25740 9460
rect 25700 9178 25728 9454
rect 25872 9444 25924 9450
rect 25872 9386 25924 9392
rect 25688 9172 25740 9178
rect 25688 9114 25740 9120
rect 25780 9036 25832 9042
rect 25780 8978 25832 8984
rect 25686 5944 25742 5953
rect 25686 5879 25742 5888
rect 25700 5778 25728 5879
rect 25688 5772 25740 5778
rect 25688 5714 25740 5720
rect 25502 3567 25558 3576
rect 25596 3596 25648 3602
rect 25596 3538 25648 3544
rect 25608 3466 25636 3538
rect 25596 3460 25648 3466
rect 25596 3402 25648 3408
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 25504 3392 25556 3398
rect 25504 3334 25556 3340
rect 25240 2514 25268 3334
rect 25228 2508 25280 2514
rect 25228 2450 25280 2456
rect 25412 1352 25464 1358
rect 25412 1294 25464 1300
rect 25320 1216 25372 1222
rect 25320 1158 25372 1164
rect 25332 1018 25360 1158
rect 25424 1018 25452 1294
rect 25320 1012 25372 1018
rect 25320 954 25372 960
rect 25412 1012 25464 1018
rect 25412 954 25464 960
rect 25516 950 25544 3334
rect 25596 2304 25648 2310
rect 25596 2246 25648 2252
rect 25504 944 25556 950
rect 25504 886 25556 892
rect 25228 876 25280 882
rect 25148 836 25228 864
rect 24584 818 24636 824
rect 25228 818 25280 824
rect 24492 808 24544 814
rect 24492 750 24544 756
rect 24124 672 24176 678
rect 24124 614 24176 620
rect 25608 474 25636 2246
rect 25700 1290 25728 5714
rect 25792 4554 25820 8978
rect 25884 8566 25912 9386
rect 26146 9072 26202 9081
rect 25964 9036 26016 9042
rect 26146 9007 26148 9016
rect 25964 8978 26016 8984
rect 26200 9007 26202 9016
rect 26148 8978 26200 8984
rect 25872 8560 25924 8566
rect 25872 8502 25924 8508
rect 25976 8430 26004 8978
rect 26344 8634 26372 11154
rect 26424 11144 26476 11150
rect 26424 11086 26476 11092
rect 26436 10062 26464 11086
rect 26424 10056 26476 10062
rect 26424 9998 26476 10004
rect 26436 9042 26464 9998
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 26528 8634 26556 11834
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 26332 8628 26384 8634
rect 26332 8570 26384 8576
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 25964 8424 26016 8430
rect 25964 8366 26016 8372
rect 26424 8356 26476 8362
rect 26424 8298 26476 8304
rect 25872 8288 25924 8294
rect 25872 8230 25924 8236
rect 25884 7478 25912 8230
rect 25872 7472 25924 7478
rect 25872 7414 25924 7420
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 26252 7002 26280 7278
rect 26240 6996 26292 7002
rect 26240 6938 26292 6944
rect 25964 6792 26016 6798
rect 25964 6734 26016 6740
rect 25872 6656 25924 6662
rect 25872 6598 25924 6604
rect 25884 5137 25912 6598
rect 25976 5914 26004 6734
rect 26056 6656 26108 6662
rect 26056 6598 26108 6604
rect 25964 5908 26016 5914
rect 25964 5850 26016 5856
rect 25964 5704 26016 5710
rect 25964 5646 26016 5652
rect 25976 5166 26004 5646
rect 25964 5160 26016 5166
rect 25870 5128 25926 5137
rect 25964 5102 26016 5108
rect 25870 5063 25926 5072
rect 25884 4808 25912 5063
rect 25884 4780 26004 4808
rect 25870 4720 25926 4729
rect 25870 4655 25926 4664
rect 25780 4548 25832 4554
rect 25780 4490 25832 4496
rect 25778 4040 25834 4049
rect 25778 3975 25834 3984
rect 25792 3466 25820 3975
rect 25884 3602 25912 4655
rect 25976 4486 26004 4780
rect 25964 4480 26016 4486
rect 25964 4422 26016 4428
rect 25964 4072 26016 4078
rect 25964 4014 26016 4020
rect 25872 3596 25924 3602
rect 25872 3538 25924 3544
rect 25780 3460 25832 3466
rect 25780 3402 25832 3408
rect 25872 3392 25924 3398
rect 25872 3334 25924 3340
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 25792 2650 25820 2926
rect 25780 2644 25832 2650
rect 25780 2586 25832 2592
rect 25792 1902 25820 2586
rect 25780 1896 25832 1902
rect 25780 1838 25832 1844
rect 25792 1494 25820 1838
rect 25780 1488 25832 1494
rect 25780 1430 25832 1436
rect 25688 1284 25740 1290
rect 25688 1226 25740 1232
rect 25688 672 25740 678
rect 25688 614 25740 620
rect 23756 468 23808 474
rect 23756 410 23808 416
rect 25596 468 25648 474
rect 25596 410 25648 416
rect 23020 400 23072 406
rect 23020 342 23072 348
rect 22836 332 22888 338
rect 22836 274 22888 280
rect 25700 241 25728 614
rect 25884 406 25912 3334
rect 25976 3058 26004 4014
rect 25964 3052 26016 3058
rect 25964 2994 26016 3000
rect 25964 2916 26016 2922
rect 25964 2858 26016 2864
rect 25976 1426 26004 2858
rect 26068 2825 26096 6598
rect 26332 6316 26384 6322
rect 26332 6258 26384 6264
rect 26148 6180 26200 6186
rect 26148 6122 26200 6128
rect 26160 4146 26188 6122
rect 26344 5817 26372 6258
rect 26330 5808 26386 5817
rect 26240 5772 26292 5778
rect 26330 5743 26386 5752
rect 26240 5714 26292 5720
rect 26252 4826 26280 5714
rect 26436 5234 26464 8298
rect 26620 7954 26648 11494
rect 26700 11348 26752 11354
rect 26700 11290 26752 11296
rect 26712 10266 26740 11290
rect 26884 11144 26936 11150
rect 26884 11086 26936 11092
rect 26896 10538 26924 11086
rect 26963 10908 27271 10917
rect 26963 10906 26969 10908
rect 27025 10906 27049 10908
rect 27105 10906 27129 10908
rect 27185 10906 27209 10908
rect 27265 10906 27271 10908
rect 27025 10854 27027 10906
rect 27207 10854 27209 10906
rect 26963 10852 26969 10854
rect 27025 10852 27049 10854
rect 27105 10852 27129 10854
rect 27185 10852 27209 10854
rect 27265 10852 27271 10854
rect 26963 10843 27271 10852
rect 26884 10532 26936 10538
rect 26884 10474 26936 10480
rect 26700 10260 26752 10266
rect 26700 10202 26752 10208
rect 26884 10260 26936 10266
rect 26884 10202 26936 10208
rect 26700 9580 26752 9586
rect 26700 9522 26752 9528
rect 26712 9042 26740 9522
rect 26792 9512 26844 9518
rect 26792 9454 26844 9460
rect 26804 9178 26832 9454
rect 26896 9178 26924 10202
rect 26963 9820 27271 9829
rect 26963 9818 26969 9820
rect 27025 9818 27049 9820
rect 27105 9818 27129 9820
rect 27185 9818 27209 9820
rect 27265 9818 27271 9820
rect 27025 9766 27027 9818
rect 27207 9766 27209 9818
rect 26963 9764 26969 9766
rect 27025 9764 27049 9766
rect 27105 9764 27129 9766
rect 27185 9764 27209 9766
rect 27265 9764 27271 9766
rect 26963 9755 27271 9764
rect 26792 9172 26844 9178
rect 26792 9114 26844 9120
rect 26884 9172 26936 9178
rect 26884 9114 26936 9120
rect 26700 9036 26752 9042
rect 26700 8978 26752 8984
rect 26884 8832 26936 8838
rect 26884 8774 26936 8780
rect 26896 8498 26924 8774
rect 26963 8732 27271 8741
rect 26963 8730 26969 8732
rect 27025 8730 27049 8732
rect 27105 8730 27129 8732
rect 27185 8730 27209 8732
rect 27265 8730 27271 8732
rect 27025 8678 27027 8730
rect 27207 8678 27209 8730
rect 26963 8676 26969 8678
rect 27025 8676 27049 8678
rect 27105 8676 27129 8678
rect 27185 8676 27209 8678
rect 27265 8676 27271 8678
rect 26963 8667 27271 8676
rect 26884 8492 26936 8498
rect 26884 8434 26936 8440
rect 26608 7948 26660 7954
rect 26608 7890 26660 7896
rect 26516 6180 26568 6186
rect 26516 6122 26568 6128
rect 26528 5846 26556 6122
rect 26516 5840 26568 5846
rect 26516 5782 26568 5788
rect 26424 5228 26476 5234
rect 26424 5170 26476 5176
rect 26620 5114 26648 7890
rect 26792 7880 26844 7886
rect 26792 7822 26844 7828
rect 26804 7342 26832 7822
rect 26963 7644 27271 7653
rect 26963 7642 26969 7644
rect 27025 7642 27049 7644
rect 27105 7642 27129 7644
rect 27185 7642 27209 7644
rect 27265 7642 27271 7644
rect 27025 7590 27027 7642
rect 27207 7590 27209 7642
rect 26963 7588 26969 7590
rect 27025 7588 27049 7590
rect 27105 7588 27129 7590
rect 27185 7588 27209 7590
rect 27265 7588 27271 7590
rect 26963 7579 27271 7588
rect 26792 7336 26844 7342
rect 26792 7278 26844 7284
rect 26976 7336 27028 7342
rect 26976 7278 27028 7284
rect 26700 6928 26752 6934
rect 26700 6870 26752 6876
rect 26712 6254 26740 6870
rect 26804 6254 26832 7278
rect 26988 7002 27016 7278
rect 26976 6996 27028 7002
rect 26976 6938 27028 6944
rect 27356 6730 27384 14894
rect 27448 14822 27476 15671
rect 27436 14816 27488 14822
rect 27436 14758 27488 14764
rect 27448 12646 27476 14758
rect 27540 14498 27568 17138
rect 27632 14618 27660 18566
rect 27712 16992 27764 16998
rect 27712 16934 27764 16940
rect 27724 16697 27752 16934
rect 27710 16688 27766 16697
rect 27710 16623 27766 16632
rect 27712 16244 27764 16250
rect 27712 16186 27764 16192
rect 27724 14822 27752 16186
rect 27816 16153 27844 18566
rect 27908 18290 27936 21422
rect 28092 21078 28120 22102
rect 28172 22092 28224 22098
rect 28172 22034 28224 22040
rect 28080 21072 28132 21078
rect 28080 21014 28132 21020
rect 28184 20874 28212 22034
rect 28356 22024 28408 22030
rect 28356 21966 28408 21972
rect 28368 21010 28396 21966
rect 28540 21344 28592 21350
rect 28540 21286 28592 21292
rect 28552 21078 28580 21286
rect 28540 21072 28592 21078
rect 28540 21014 28592 21020
rect 28356 21004 28408 21010
rect 28356 20946 28408 20952
rect 28264 20936 28316 20942
rect 28264 20878 28316 20884
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 28172 20868 28224 20874
rect 28172 20810 28224 20816
rect 28172 20256 28224 20262
rect 28172 20198 28224 20204
rect 28078 20088 28134 20097
rect 28078 20023 28134 20032
rect 28092 19718 28120 20023
rect 27988 19712 28040 19718
rect 27988 19654 28040 19660
rect 28080 19712 28132 19718
rect 28080 19654 28132 19660
rect 27896 18284 27948 18290
rect 27896 18226 27948 18232
rect 27896 16584 27948 16590
rect 27896 16526 27948 16532
rect 27802 16144 27858 16153
rect 27802 16079 27858 16088
rect 27804 15972 27856 15978
rect 27804 15914 27856 15920
rect 27816 15706 27844 15914
rect 27804 15700 27856 15706
rect 27804 15642 27856 15648
rect 27816 14929 27844 15642
rect 27802 14920 27858 14929
rect 27802 14855 27858 14864
rect 27712 14816 27764 14822
rect 27712 14758 27764 14764
rect 27620 14612 27672 14618
rect 27620 14554 27672 14560
rect 27540 14470 27660 14498
rect 27528 14408 27580 14414
rect 27528 14350 27580 14356
rect 27540 13190 27568 14350
rect 27632 13938 27660 14470
rect 27620 13932 27672 13938
rect 27620 13874 27672 13880
rect 27618 13424 27674 13433
rect 27618 13359 27620 13368
rect 27672 13359 27674 13368
rect 27620 13330 27672 13336
rect 27528 13184 27580 13190
rect 27528 13126 27580 13132
rect 27804 12844 27856 12850
rect 27804 12786 27856 12792
rect 27436 12640 27488 12646
rect 27436 12582 27488 12588
rect 27448 12442 27476 12582
rect 27436 12436 27488 12442
rect 27436 12378 27488 12384
rect 27528 11892 27580 11898
rect 27528 11834 27580 11840
rect 27540 11694 27568 11834
rect 27618 11792 27674 11801
rect 27618 11727 27674 11736
rect 27632 11694 27660 11727
rect 27528 11688 27580 11694
rect 27528 11630 27580 11636
rect 27620 11688 27672 11694
rect 27620 11630 27672 11636
rect 27436 11348 27488 11354
rect 27436 11290 27488 11296
rect 27448 8430 27476 11290
rect 27540 8838 27568 11630
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 27816 8634 27844 12786
rect 27908 12442 27936 16526
rect 28000 14482 28028 19654
rect 28184 16658 28212 20198
rect 28276 18426 28304 20878
rect 28460 19922 28488 20878
rect 28540 20460 28592 20466
rect 28540 20402 28592 20408
rect 28448 19916 28500 19922
rect 28448 19858 28500 19864
rect 28264 18420 28316 18426
rect 28264 18362 28316 18368
rect 28354 17912 28410 17921
rect 28354 17847 28410 17856
rect 28368 17542 28396 17847
rect 28356 17536 28408 17542
rect 28356 17478 28408 17484
rect 28264 17060 28316 17066
rect 28316 17020 28488 17048
rect 28264 17002 28316 17008
rect 28080 16652 28132 16658
rect 28080 16594 28132 16600
rect 28172 16652 28224 16658
rect 28172 16594 28224 16600
rect 27988 14476 28040 14482
rect 27988 14418 28040 14424
rect 28092 14074 28120 16594
rect 28184 14550 28212 16594
rect 28264 16108 28316 16114
rect 28264 16050 28316 16056
rect 28172 14544 28224 14550
rect 28172 14486 28224 14492
rect 28080 14068 28132 14074
rect 28080 14010 28132 14016
rect 28184 13870 28212 14486
rect 28172 13864 28224 13870
rect 28172 13806 28224 13812
rect 28172 13728 28224 13734
rect 28000 13688 28172 13716
rect 28000 12617 28028 13688
rect 28172 13670 28224 13676
rect 28276 13530 28304 16050
rect 28354 15736 28410 15745
rect 28354 15671 28410 15680
rect 28368 15570 28396 15671
rect 28356 15564 28408 15570
rect 28356 15506 28408 15512
rect 28356 15360 28408 15366
rect 28356 15302 28408 15308
rect 28368 15162 28396 15302
rect 28356 15156 28408 15162
rect 28356 15098 28408 15104
rect 28356 14612 28408 14618
rect 28356 14554 28408 14560
rect 28368 14385 28396 14554
rect 28354 14376 28410 14385
rect 28354 14311 28410 14320
rect 28264 13524 28316 13530
rect 28264 13466 28316 13472
rect 28172 13456 28224 13462
rect 28172 13398 28224 13404
rect 28080 12640 28132 12646
rect 27986 12608 28042 12617
rect 28080 12582 28132 12588
rect 27986 12543 28042 12552
rect 27896 12436 27948 12442
rect 27896 12378 27948 12384
rect 27896 9376 27948 9382
rect 27896 9318 27948 9324
rect 27908 9178 27936 9318
rect 27896 9172 27948 9178
rect 27896 9114 27948 9120
rect 27896 8832 27948 8838
rect 27896 8774 27948 8780
rect 27620 8628 27672 8634
rect 27620 8570 27672 8576
rect 27804 8628 27856 8634
rect 27804 8570 27856 8576
rect 27436 8424 27488 8430
rect 27436 8366 27488 8372
rect 27632 7954 27660 8570
rect 27908 8022 27936 8774
rect 27896 8016 27948 8022
rect 27896 7958 27948 7964
rect 27620 7948 27672 7954
rect 27620 7890 27672 7896
rect 27804 7880 27856 7886
rect 27804 7822 27856 7828
rect 27436 7744 27488 7750
rect 27436 7686 27488 7692
rect 27528 7744 27580 7750
rect 27528 7686 27580 7692
rect 27448 7342 27476 7686
rect 27436 7336 27488 7342
rect 27436 7278 27488 7284
rect 27436 6928 27488 6934
rect 27436 6870 27488 6876
rect 27344 6724 27396 6730
rect 27344 6666 27396 6672
rect 26963 6556 27271 6565
rect 26963 6554 26969 6556
rect 27025 6554 27049 6556
rect 27105 6554 27129 6556
rect 27185 6554 27209 6556
rect 27265 6554 27271 6556
rect 27025 6502 27027 6554
rect 27207 6502 27209 6554
rect 26963 6500 26969 6502
rect 27025 6500 27049 6502
rect 27105 6500 27129 6502
rect 27185 6500 27209 6502
rect 27265 6500 27271 6502
rect 26963 6491 27271 6500
rect 26700 6248 26752 6254
rect 26700 6190 26752 6196
rect 26792 6248 26844 6254
rect 26792 6190 26844 6196
rect 27448 6202 27476 6870
rect 27540 6322 27568 7686
rect 27816 6798 27844 7822
rect 27908 7002 27936 7958
rect 27896 6996 27948 7002
rect 27896 6938 27948 6944
rect 28000 6798 28028 12543
rect 28092 12238 28120 12582
rect 28080 12232 28132 12238
rect 28080 12174 28132 12180
rect 28184 11762 28212 13398
rect 28172 11756 28224 11762
rect 28172 11698 28224 11704
rect 28264 11552 28316 11558
rect 28264 11494 28316 11500
rect 28080 11076 28132 11082
rect 28080 11018 28132 11024
rect 28092 8498 28120 11018
rect 28276 10674 28304 11494
rect 28264 10668 28316 10674
rect 28264 10610 28316 10616
rect 28368 10418 28396 14311
rect 28184 10390 28396 10418
rect 28184 8906 28212 10390
rect 28264 10056 28316 10062
rect 28460 10010 28488 17020
rect 28552 15366 28580 20402
rect 28736 19310 28764 22170
rect 30472 21888 30524 21894
rect 30472 21830 30524 21836
rect 30012 21344 30064 21350
rect 30012 21286 30064 21292
rect 30288 21344 30340 21350
rect 30288 21286 30340 21292
rect 28816 20936 28868 20942
rect 28816 20878 28868 20884
rect 29000 20936 29052 20942
rect 29000 20878 29052 20884
rect 29552 20936 29604 20942
rect 29552 20878 29604 20884
rect 28828 20262 28856 20878
rect 28816 20256 28868 20262
rect 28816 20198 28868 20204
rect 28828 20058 28856 20198
rect 28816 20052 28868 20058
rect 28816 19994 28868 20000
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 28724 19304 28776 19310
rect 28724 19246 28776 19252
rect 28632 19168 28684 19174
rect 28632 19110 28684 19116
rect 28644 18698 28672 19110
rect 28816 18828 28868 18834
rect 28816 18770 28868 18776
rect 28632 18692 28684 18698
rect 28632 18634 28684 18640
rect 28644 18154 28672 18634
rect 28724 18216 28776 18222
rect 28724 18158 28776 18164
rect 28632 18148 28684 18154
rect 28632 18090 28684 18096
rect 28736 17882 28764 18158
rect 28724 17876 28776 17882
rect 28724 17818 28776 17824
rect 28632 17808 28684 17814
rect 28632 17750 28684 17756
rect 28644 17270 28672 17750
rect 28736 17649 28764 17818
rect 28828 17814 28856 18770
rect 28816 17808 28868 17814
rect 28816 17750 28868 17756
rect 28722 17640 28778 17649
rect 28722 17575 28778 17584
rect 28724 17332 28776 17338
rect 28724 17274 28776 17280
rect 28632 17264 28684 17270
rect 28632 17206 28684 17212
rect 28644 17066 28672 17206
rect 28736 17134 28764 17274
rect 28724 17128 28776 17134
rect 28776 17076 28856 17082
rect 28724 17070 28856 17076
rect 28632 17060 28684 17066
rect 28736 17054 28856 17070
rect 28632 17002 28684 17008
rect 28644 15609 28672 17002
rect 28724 16992 28776 16998
rect 28724 16934 28776 16940
rect 28736 16289 28764 16934
rect 28828 16726 28856 17054
rect 28816 16720 28868 16726
rect 28816 16662 28868 16668
rect 28722 16280 28778 16289
rect 28722 16215 28778 16224
rect 28816 15904 28868 15910
rect 28816 15846 28868 15852
rect 28630 15600 28686 15609
rect 28630 15535 28686 15544
rect 28632 15496 28684 15502
rect 28684 15456 28764 15484
rect 28632 15438 28684 15444
rect 28540 15360 28592 15366
rect 28540 15302 28592 15308
rect 28540 15156 28592 15162
rect 28540 15098 28592 15104
rect 28552 13841 28580 15098
rect 28632 14272 28684 14278
rect 28632 14214 28684 14220
rect 28538 13832 28594 13841
rect 28538 13767 28594 13776
rect 28644 13462 28672 14214
rect 28632 13456 28684 13462
rect 28632 13398 28684 13404
rect 28632 12640 28684 12646
rect 28632 12582 28684 12588
rect 28540 12300 28592 12306
rect 28540 12242 28592 12248
rect 28552 11558 28580 12242
rect 28644 11898 28672 12582
rect 28632 11892 28684 11898
rect 28632 11834 28684 11840
rect 28540 11552 28592 11558
rect 28540 11494 28592 11500
rect 28540 11144 28592 11150
rect 28540 11086 28592 11092
rect 28552 10606 28580 11086
rect 28540 10600 28592 10606
rect 28540 10542 28592 10548
rect 28264 9998 28316 10004
rect 28276 9722 28304 9998
rect 28368 9982 28488 10010
rect 28264 9716 28316 9722
rect 28264 9658 28316 9664
rect 28172 8900 28224 8906
rect 28172 8842 28224 8848
rect 28264 8832 28316 8838
rect 28264 8774 28316 8780
rect 28080 8492 28132 8498
rect 28080 8434 28132 8440
rect 28172 8084 28224 8090
rect 28172 8026 28224 8032
rect 27804 6792 27856 6798
rect 27804 6734 27856 6740
rect 27988 6792 28040 6798
rect 27988 6734 28040 6740
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 27448 6174 27568 6202
rect 26700 6112 26752 6118
rect 26700 6054 26752 6060
rect 27252 6112 27304 6118
rect 27252 6054 27304 6060
rect 27344 6112 27396 6118
rect 27344 6054 27396 6060
rect 26528 5086 26648 5114
rect 26240 4820 26292 4826
rect 26240 4762 26292 4768
rect 26528 4146 26556 5086
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 26620 4146 26648 4966
rect 26148 4140 26200 4146
rect 26148 4082 26200 4088
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26608 4140 26660 4146
rect 26608 4082 26660 4088
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 26436 3058 26464 3878
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26424 3052 26476 3058
rect 26424 2994 26476 3000
rect 26439 2904 26467 2994
rect 26436 2876 26467 2904
rect 26054 2816 26110 2825
rect 26054 2751 26110 2760
rect 26240 2508 26292 2514
rect 26240 2450 26292 2456
rect 26056 2440 26108 2446
rect 26056 2382 26108 2388
rect 26068 2310 26096 2382
rect 26056 2304 26108 2310
rect 26252 2281 26280 2450
rect 26332 2440 26384 2446
rect 26332 2382 26384 2388
rect 26056 2246 26108 2252
rect 26238 2272 26294 2281
rect 26238 2207 26294 2216
rect 26344 1834 26372 2382
rect 26436 2145 26464 2876
rect 26422 2136 26478 2145
rect 26422 2071 26478 2080
rect 26436 1902 26464 2071
rect 26424 1896 26476 1902
rect 26424 1838 26476 1844
rect 26528 1850 26556 3470
rect 26620 2774 26648 3878
rect 26712 3058 26740 6054
rect 27264 5914 27292 6054
rect 27252 5908 27304 5914
rect 27252 5850 27304 5856
rect 26884 5704 26936 5710
rect 26884 5646 26936 5652
rect 26896 5370 26924 5646
rect 26963 5468 27271 5477
rect 26963 5466 26969 5468
rect 27025 5466 27049 5468
rect 27105 5466 27129 5468
rect 27185 5466 27209 5468
rect 27265 5466 27271 5468
rect 27025 5414 27027 5466
rect 27207 5414 27209 5466
rect 26963 5412 26969 5414
rect 27025 5412 27049 5414
rect 27105 5412 27129 5414
rect 27185 5412 27209 5414
rect 27265 5412 27271 5414
rect 26963 5403 27271 5412
rect 26884 5364 26936 5370
rect 26884 5306 26936 5312
rect 27068 5364 27120 5370
rect 27068 5306 27120 5312
rect 27080 5030 27108 5306
rect 27068 5024 27120 5030
rect 27068 4966 27120 4972
rect 26792 4480 26844 4486
rect 26792 4422 26844 4428
rect 26884 4480 26936 4486
rect 26884 4422 26936 4428
rect 26700 3052 26752 3058
rect 26700 2994 26752 3000
rect 26804 2961 26832 4422
rect 26790 2952 26846 2961
rect 26790 2887 26846 2896
rect 26792 2848 26844 2854
rect 26792 2790 26844 2796
rect 26620 2746 26740 2774
rect 26712 2009 26740 2746
rect 26804 2689 26832 2790
rect 26790 2680 26846 2689
rect 26790 2615 26846 2624
rect 26792 2440 26844 2446
rect 26792 2382 26844 2388
rect 26804 2145 26832 2382
rect 26790 2136 26846 2145
rect 26790 2071 26846 2080
rect 26698 2000 26754 2009
rect 26698 1935 26754 1944
rect 26896 1884 26924 4422
rect 26963 4380 27271 4389
rect 26963 4378 26969 4380
rect 27025 4378 27049 4380
rect 27105 4378 27129 4380
rect 27185 4378 27209 4380
rect 27265 4378 27271 4380
rect 27025 4326 27027 4378
rect 27207 4326 27209 4378
rect 26963 4324 26969 4326
rect 27025 4324 27049 4326
rect 27105 4324 27129 4326
rect 27185 4324 27209 4326
rect 27265 4324 27271 4326
rect 26963 4315 27271 4324
rect 26963 3292 27271 3301
rect 26963 3290 26969 3292
rect 27025 3290 27049 3292
rect 27105 3290 27129 3292
rect 27185 3290 27209 3292
rect 27265 3290 27271 3292
rect 27025 3238 27027 3290
rect 27207 3238 27209 3290
rect 26963 3236 26969 3238
rect 27025 3236 27049 3238
rect 27105 3236 27129 3238
rect 27185 3236 27209 3238
rect 27265 3236 27271 3238
rect 26963 3227 27271 3236
rect 26976 3052 27028 3058
rect 26976 2994 27028 3000
rect 26988 2825 27016 2994
rect 27250 2952 27306 2961
rect 27250 2887 27306 2896
rect 26974 2816 27030 2825
rect 26974 2751 27030 2760
rect 27264 2514 27292 2887
rect 27252 2508 27304 2514
rect 27252 2450 27304 2456
rect 26963 2204 27271 2213
rect 26963 2202 26969 2204
rect 27025 2202 27049 2204
rect 27105 2202 27129 2204
rect 27185 2202 27209 2204
rect 27265 2202 27271 2204
rect 27025 2150 27027 2202
rect 27207 2150 27209 2202
rect 26963 2148 26969 2150
rect 27025 2148 27049 2150
rect 27105 2148 27129 2150
rect 27185 2148 27209 2150
rect 27265 2148 27271 2150
rect 26963 2139 27271 2148
rect 26976 1896 27028 1902
rect 26896 1856 26976 1884
rect 26332 1828 26384 1834
rect 26528 1822 26832 1850
rect 26976 1838 27028 1844
rect 26332 1770 26384 1776
rect 26056 1760 26108 1766
rect 26424 1760 26476 1766
rect 26056 1702 26108 1708
rect 26422 1728 26424 1737
rect 26476 1728 26478 1737
rect 25964 1420 26016 1426
rect 25964 1362 26016 1368
rect 26068 1193 26096 1702
rect 26422 1663 26478 1672
rect 26148 1216 26200 1222
rect 26054 1184 26110 1193
rect 26148 1158 26200 1164
rect 26054 1119 26110 1128
rect 26160 950 26188 1158
rect 26148 944 26200 950
rect 26148 886 26200 892
rect 26436 882 26464 1663
rect 26516 1488 26568 1494
rect 26516 1430 26568 1436
rect 26698 1456 26754 1465
rect 26528 1340 26556 1430
rect 26698 1391 26754 1400
rect 26608 1352 26660 1358
rect 26528 1312 26608 1340
rect 26608 1294 26660 1300
rect 26424 876 26476 882
rect 26424 818 26476 824
rect 26608 808 26660 814
rect 26712 796 26740 1391
rect 26804 814 26832 1822
rect 26884 1556 26936 1562
rect 26884 1498 26936 1504
rect 26896 882 26924 1498
rect 26976 1352 27028 1358
rect 26976 1294 27028 1300
rect 26988 1222 27016 1294
rect 26976 1216 27028 1222
rect 26976 1158 27028 1164
rect 26963 1116 27271 1125
rect 26963 1114 26969 1116
rect 27025 1114 27049 1116
rect 27105 1114 27129 1116
rect 27185 1114 27209 1116
rect 27265 1114 27271 1116
rect 27025 1062 27027 1114
rect 27207 1062 27209 1114
rect 26963 1060 26969 1062
rect 27025 1060 27049 1062
rect 27105 1060 27129 1062
rect 27185 1060 27209 1062
rect 27265 1060 27271 1062
rect 26963 1051 27271 1060
rect 27356 882 27384 6054
rect 27540 5166 27568 6174
rect 28000 5778 28028 6734
rect 28080 6316 28132 6322
rect 28080 6258 28132 6264
rect 27988 5772 28040 5778
rect 27988 5714 28040 5720
rect 27896 5636 27948 5642
rect 27896 5578 27948 5584
rect 27804 5568 27856 5574
rect 27724 5528 27804 5556
rect 27528 5160 27580 5166
rect 27528 5102 27580 5108
rect 27540 4758 27568 5102
rect 27528 4752 27580 4758
rect 27528 4694 27580 4700
rect 27436 4072 27488 4078
rect 27436 4014 27488 4020
rect 27448 3602 27476 4014
rect 27528 3936 27580 3942
rect 27528 3878 27580 3884
rect 27436 3596 27488 3602
rect 27436 3538 27488 3544
rect 27448 2582 27476 3538
rect 27436 2576 27488 2582
rect 27436 2518 27488 2524
rect 27436 2440 27488 2446
rect 27436 2382 27488 2388
rect 27448 1562 27476 2382
rect 27436 1556 27488 1562
rect 27436 1498 27488 1504
rect 26884 876 26936 882
rect 26884 818 26936 824
rect 27344 876 27396 882
rect 27344 818 27396 824
rect 27540 814 27568 3878
rect 27618 3088 27674 3097
rect 27618 3023 27674 3032
rect 27632 2446 27660 3023
rect 27620 2440 27672 2446
rect 27620 2382 27672 2388
rect 27724 1970 27752 5528
rect 27804 5510 27856 5516
rect 27908 4690 27936 5578
rect 28092 5370 28120 6258
rect 28080 5364 28132 5370
rect 28080 5306 28132 5312
rect 27896 4684 27948 4690
rect 27896 4626 27948 4632
rect 27988 4684 28040 4690
rect 27988 4626 28040 4632
rect 28000 3602 28028 4626
rect 28184 4078 28212 8026
rect 28276 6798 28304 8774
rect 28368 8430 28396 9982
rect 28448 9920 28500 9926
rect 28448 9862 28500 9868
rect 28736 9874 28764 15456
rect 28828 13734 28856 15846
rect 28816 13728 28868 13734
rect 28816 13670 28868 13676
rect 28816 13184 28868 13190
rect 28816 13126 28868 13132
rect 28828 12434 28856 13126
rect 28920 12986 28948 19790
rect 29012 15162 29040 20878
rect 29184 20460 29236 20466
rect 29184 20402 29236 20408
rect 29092 19848 29144 19854
rect 29092 19790 29144 19796
rect 29000 15156 29052 15162
rect 29000 15098 29052 15104
rect 29000 14952 29052 14958
rect 29000 14894 29052 14900
rect 28908 12980 28960 12986
rect 28908 12922 28960 12928
rect 29012 12442 29040 14894
rect 29104 14074 29132 19790
rect 29196 19310 29224 20402
rect 29276 20392 29328 20398
rect 29276 20334 29328 20340
rect 29460 20392 29512 20398
rect 29460 20334 29512 20340
rect 29184 19304 29236 19310
rect 29184 19246 29236 19252
rect 29196 18834 29224 19246
rect 29184 18828 29236 18834
rect 29184 18770 29236 18776
rect 29196 18222 29224 18770
rect 29184 18216 29236 18222
rect 29184 18158 29236 18164
rect 29182 18048 29238 18057
rect 29182 17983 29238 17992
rect 29196 16794 29224 17983
rect 29184 16788 29236 16794
rect 29184 16730 29236 16736
rect 29184 16040 29236 16046
rect 29182 16008 29184 16017
rect 29236 16008 29238 16017
rect 29182 15943 29238 15952
rect 29182 15464 29238 15473
rect 29182 15399 29238 15408
rect 29196 14958 29224 15399
rect 29184 14952 29236 14958
rect 29184 14894 29236 14900
rect 29288 14618 29316 20334
rect 29472 19242 29500 20334
rect 29460 19236 29512 19242
rect 29460 19178 29512 19184
rect 29366 18320 29422 18329
rect 29422 18278 29500 18306
rect 29366 18255 29422 18264
rect 29368 18216 29420 18222
rect 29368 18158 29420 18164
rect 29380 17814 29408 18158
rect 29368 17808 29420 17814
rect 29368 17750 29420 17756
rect 29380 17338 29408 17750
rect 29368 17332 29420 17338
rect 29368 17274 29420 17280
rect 29366 17096 29422 17105
rect 29366 17031 29422 17040
rect 29380 16998 29408 17031
rect 29368 16992 29420 16998
rect 29368 16934 29420 16940
rect 29366 16280 29422 16289
rect 29366 16215 29422 16224
rect 29380 15570 29408 16215
rect 29368 15564 29420 15570
rect 29368 15506 29420 15512
rect 29472 15162 29500 18278
rect 29564 15434 29592 20878
rect 29644 20800 29696 20806
rect 29696 20760 29776 20788
rect 29644 20742 29696 20748
rect 29748 20466 29776 20760
rect 29736 20460 29788 20466
rect 29736 20402 29788 20408
rect 29644 20256 29696 20262
rect 29644 20198 29696 20204
rect 29656 19242 29684 20198
rect 29644 19236 29696 19242
rect 29644 19178 29696 19184
rect 29644 18080 29696 18086
rect 29644 18022 29696 18028
rect 29656 17678 29684 18022
rect 29644 17672 29696 17678
rect 29644 17614 29696 17620
rect 29656 17134 29684 17614
rect 29644 17128 29696 17134
rect 29644 17070 29696 17076
rect 29656 16726 29684 17070
rect 29644 16720 29696 16726
rect 29644 16662 29696 16668
rect 29748 16572 29776 20402
rect 30024 20330 30052 21286
rect 30300 21146 30328 21286
rect 30484 21146 30512 21830
rect 31300 21344 31352 21350
rect 31300 21286 31352 21292
rect 30758 21244 31066 21253
rect 30758 21242 30764 21244
rect 30820 21242 30844 21244
rect 30900 21242 30924 21244
rect 30980 21242 31004 21244
rect 31060 21242 31066 21244
rect 30820 21190 30822 21242
rect 31002 21190 31004 21242
rect 30758 21188 30764 21190
rect 30820 21188 30844 21190
rect 30900 21188 30924 21190
rect 30980 21188 31004 21190
rect 31060 21188 31066 21190
rect 30758 21179 31066 21188
rect 30288 21140 30340 21146
rect 30288 21082 30340 21088
rect 30472 21140 30524 21146
rect 30472 21082 30524 21088
rect 30012 20324 30064 20330
rect 30012 20266 30064 20272
rect 29828 20256 29880 20262
rect 29828 20198 29880 20204
rect 29656 16544 29776 16572
rect 29552 15428 29604 15434
rect 29552 15370 29604 15376
rect 29460 15156 29512 15162
rect 29460 15098 29512 15104
rect 29368 15088 29420 15094
rect 29368 15030 29420 15036
rect 29184 14612 29236 14618
rect 29184 14554 29236 14560
rect 29276 14612 29328 14618
rect 29276 14554 29328 14560
rect 29196 14482 29224 14554
rect 29184 14476 29236 14482
rect 29184 14418 29236 14424
rect 29092 14068 29144 14074
rect 29092 14010 29144 14016
rect 29090 13832 29146 13841
rect 29090 13767 29146 13776
rect 29000 12436 29052 12442
rect 28828 12406 28948 12434
rect 28816 12096 28868 12102
rect 28816 12038 28868 12044
rect 28828 10062 28856 12038
rect 28920 11218 28948 12406
rect 29000 12378 29052 12384
rect 28908 11212 28960 11218
rect 28908 11154 28960 11160
rect 29000 10464 29052 10470
rect 29000 10406 29052 10412
rect 28816 10056 28868 10062
rect 28816 9998 28868 10004
rect 28356 8424 28408 8430
rect 28356 8366 28408 8372
rect 28460 7954 28488 9862
rect 28736 9846 28948 9874
rect 28816 9648 28868 9654
rect 28816 9590 28868 9596
rect 28540 9376 28592 9382
rect 28540 9318 28592 9324
rect 28552 9178 28580 9318
rect 28540 9172 28592 9178
rect 28540 9114 28592 9120
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28644 8090 28672 8570
rect 28632 8084 28684 8090
rect 28632 8026 28684 8032
rect 28448 7948 28500 7954
rect 28448 7890 28500 7896
rect 28448 7744 28500 7750
rect 28448 7686 28500 7692
rect 28632 7744 28684 7750
rect 28632 7686 28684 7692
rect 28460 7546 28488 7686
rect 28448 7540 28500 7546
rect 28448 7482 28500 7488
rect 28264 6792 28316 6798
rect 28264 6734 28316 6740
rect 28538 6352 28594 6361
rect 28538 6287 28594 6296
rect 28356 6180 28408 6186
rect 28356 6122 28408 6128
rect 28368 5030 28396 6122
rect 28552 5370 28580 6287
rect 28540 5364 28592 5370
rect 28540 5306 28592 5312
rect 28356 5024 28408 5030
rect 28356 4966 28408 4972
rect 28368 4622 28396 4966
rect 28356 4616 28408 4622
rect 28540 4616 28592 4622
rect 28408 4564 28488 4570
rect 28356 4558 28488 4564
rect 28540 4558 28592 4564
rect 28368 4542 28488 4558
rect 28172 4072 28224 4078
rect 28172 4014 28224 4020
rect 28184 3738 28212 4014
rect 28356 3936 28408 3942
rect 28356 3878 28408 3884
rect 28368 3777 28396 3878
rect 28354 3768 28410 3777
rect 28172 3732 28224 3738
rect 28354 3703 28410 3712
rect 28172 3674 28224 3680
rect 27988 3596 28040 3602
rect 27988 3538 28040 3544
rect 27802 3496 27858 3505
rect 27802 3431 27858 3440
rect 27816 1986 27844 3431
rect 28000 2514 28028 3538
rect 28460 3534 28488 4542
rect 28356 3528 28408 3534
rect 28356 3470 28408 3476
rect 28448 3528 28500 3534
rect 28448 3470 28500 3476
rect 28368 3210 28396 3470
rect 28092 3182 28396 3210
rect 27988 2508 28040 2514
rect 27988 2450 28040 2456
rect 27712 1964 27764 1970
rect 27816 1958 28028 1986
rect 27712 1906 27764 1912
rect 28000 1562 28028 1958
rect 27988 1556 28040 1562
rect 27988 1498 28040 1504
rect 26660 768 26740 796
rect 26792 808 26844 814
rect 26608 750 26660 756
rect 26792 750 26844 756
rect 27528 808 27580 814
rect 27528 750 27580 756
rect 26056 672 26108 678
rect 26056 614 26108 620
rect 25872 400 25924 406
rect 25872 342 25924 348
rect 26068 338 26096 614
rect 26056 332 26108 338
rect 26056 274 26108 280
rect 25686 232 25742 241
rect 25686 167 25742 176
rect 22744 128 22796 134
rect 22744 70 22796 76
rect 26804 66 26832 750
rect 28092 105 28120 3182
rect 28172 3120 28224 3126
rect 28172 3062 28224 3068
rect 28184 2106 28212 3062
rect 28460 2650 28488 3470
rect 28448 2644 28500 2650
rect 28448 2586 28500 2592
rect 28172 2100 28224 2106
rect 28172 2042 28224 2048
rect 28356 1556 28408 1562
rect 28356 1498 28408 1504
rect 28368 202 28396 1498
rect 28552 1018 28580 4558
rect 28644 3602 28672 7686
rect 28724 7472 28776 7478
rect 28724 7414 28776 7420
rect 28632 3596 28684 3602
rect 28632 3538 28684 3544
rect 28736 2514 28764 7414
rect 28724 2508 28776 2514
rect 28724 2450 28776 2456
rect 28828 1970 28856 9590
rect 28920 8090 28948 9846
rect 29012 9586 29040 10406
rect 29000 9580 29052 9586
rect 29000 9522 29052 9528
rect 28908 8084 28960 8090
rect 28908 8026 28960 8032
rect 29012 7886 29040 9522
rect 29104 8430 29132 13767
rect 29182 13288 29238 13297
rect 29182 13223 29238 13232
rect 29196 10130 29224 13223
rect 29380 12714 29408 15030
rect 29656 14906 29684 16544
rect 29736 16040 29788 16046
rect 29840 16028 29868 20198
rect 30758 20156 31066 20165
rect 30758 20154 30764 20156
rect 30820 20154 30844 20156
rect 30900 20154 30924 20156
rect 30980 20154 31004 20156
rect 31060 20154 31066 20156
rect 30820 20102 30822 20154
rect 31002 20102 31004 20154
rect 30758 20100 30764 20102
rect 30820 20100 30844 20102
rect 30900 20100 30924 20102
rect 30980 20100 31004 20102
rect 31060 20100 31066 20102
rect 30758 20091 31066 20100
rect 30472 19712 30524 19718
rect 30472 19654 30524 19660
rect 30104 19168 30156 19174
rect 30104 19110 30156 19116
rect 30196 19168 30248 19174
rect 30196 19110 30248 19116
rect 30380 19168 30432 19174
rect 30380 19110 30432 19116
rect 29920 18080 29972 18086
rect 29920 18022 29972 18028
rect 29932 17542 29960 18022
rect 29920 17536 29972 17542
rect 29920 17478 29972 17484
rect 30012 17536 30064 17542
rect 30012 17478 30064 17484
rect 29932 17105 29960 17478
rect 29918 17096 29974 17105
rect 29918 17031 29974 17040
rect 29920 16992 29972 16998
rect 29920 16934 29972 16940
rect 29932 16794 29960 16934
rect 29920 16788 29972 16794
rect 29920 16730 29972 16736
rect 29788 16000 29868 16028
rect 29736 15982 29788 15988
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29736 15428 29788 15434
rect 29736 15370 29788 15376
rect 29472 14878 29684 14906
rect 29368 12708 29420 12714
rect 29368 12650 29420 12656
rect 29472 12594 29500 14878
rect 29748 14074 29776 15370
rect 29736 14068 29788 14074
rect 29736 14010 29788 14016
rect 29644 14000 29696 14006
rect 29644 13942 29696 13948
rect 29552 13796 29604 13802
rect 29552 13738 29604 13744
rect 29564 12850 29592 13738
rect 29552 12844 29604 12850
rect 29656 12832 29684 13942
rect 29840 12986 29868 15438
rect 29920 15088 29972 15094
rect 29920 15030 29972 15036
rect 29932 13938 29960 15030
rect 30024 14958 30052 17478
rect 30116 17066 30144 19110
rect 30208 18698 30236 19110
rect 30392 18970 30420 19110
rect 30484 18970 30512 19654
rect 30564 19304 30616 19310
rect 30564 19246 30616 19252
rect 30380 18964 30432 18970
rect 30380 18906 30432 18912
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 30196 18692 30248 18698
rect 30196 18634 30248 18640
rect 30208 18222 30236 18634
rect 30380 18624 30432 18630
rect 30380 18566 30432 18572
rect 30196 18216 30248 18222
rect 30196 18158 30248 18164
rect 30288 18080 30340 18086
rect 30288 18022 30340 18028
rect 30300 17785 30328 18022
rect 30286 17776 30342 17785
rect 30208 17734 30286 17762
rect 30104 17060 30156 17066
rect 30104 17002 30156 17008
rect 30102 16960 30158 16969
rect 30102 16895 30158 16904
rect 30116 16114 30144 16895
rect 30104 16108 30156 16114
rect 30104 16050 30156 16056
rect 30012 14952 30064 14958
rect 30012 14894 30064 14900
rect 30012 14476 30064 14482
rect 30012 14418 30064 14424
rect 29920 13932 29972 13938
rect 29920 13874 29972 13880
rect 29828 12980 29880 12986
rect 29828 12922 29880 12928
rect 29656 12804 29868 12832
rect 29552 12786 29604 12792
rect 29380 12566 29500 12594
rect 29380 12238 29408 12566
rect 29368 12232 29420 12238
rect 29368 12174 29420 12180
rect 29380 11218 29408 12174
rect 29368 11212 29420 11218
rect 29368 11154 29420 11160
rect 29276 11008 29328 11014
rect 29276 10950 29328 10956
rect 29184 10124 29236 10130
rect 29184 10066 29236 10072
rect 29184 9512 29236 9518
rect 29184 9454 29236 9460
rect 29092 8424 29144 8430
rect 29092 8366 29144 8372
rect 29092 8288 29144 8294
rect 29092 8230 29144 8236
rect 29000 7880 29052 7886
rect 28906 7848 28962 7857
rect 29000 7822 29052 7828
rect 28906 7783 28962 7792
rect 28920 5114 28948 7783
rect 29104 7342 29132 8230
rect 29196 7342 29224 9454
rect 29288 8634 29316 10950
rect 29368 10668 29420 10674
rect 29368 10610 29420 10616
rect 29276 8628 29328 8634
rect 29276 8570 29328 8576
rect 29092 7336 29144 7342
rect 29092 7278 29144 7284
rect 29184 7336 29236 7342
rect 29184 7278 29236 7284
rect 29000 7200 29052 7206
rect 29000 7142 29052 7148
rect 29012 5234 29040 7142
rect 29000 5228 29052 5234
rect 29000 5170 29052 5176
rect 28920 5086 29040 5114
rect 29012 3738 29040 5086
rect 29000 3732 29052 3738
rect 29000 3674 29052 3680
rect 29104 3058 29132 7278
rect 29288 6254 29316 8570
rect 29380 8498 29408 10610
rect 29460 10600 29512 10606
rect 29564 10588 29592 12786
rect 29840 12458 29868 12804
rect 30024 12782 30052 14418
rect 30116 13802 30144 16050
rect 30208 16046 30236 17734
rect 30286 17711 30342 17720
rect 30288 17196 30340 17202
rect 30288 17138 30340 17144
rect 30300 16658 30328 17138
rect 30392 16794 30420 18566
rect 30380 16788 30432 16794
rect 30380 16730 30432 16736
rect 30288 16652 30340 16658
rect 30288 16594 30340 16600
rect 30380 16652 30432 16658
rect 30380 16594 30432 16600
rect 30392 16250 30420 16594
rect 30484 16250 30512 18906
rect 30576 17338 30604 19246
rect 30758 19068 31066 19077
rect 30758 19066 30764 19068
rect 30820 19066 30844 19068
rect 30900 19066 30924 19068
rect 30980 19066 31004 19068
rect 31060 19066 31066 19068
rect 30820 19014 30822 19066
rect 31002 19014 31004 19066
rect 30758 19012 30764 19014
rect 30820 19012 30844 19014
rect 30900 19012 30924 19014
rect 30980 19012 31004 19014
rect 31060 19012 31066 19014
rect 30758 19003 31066 19012
rect 30758 17980 31066 17989
rect 30758 17978 30764 17980
rect 30820 17978 30844 17980
rect 30900 17978 30924 17980
rect 30980 17978 31004 17980
rect 31060 17978 31066 17980
rect 30820 17926 30822 17978
rect 31002 17926 31004 17978
rect 30758 17924 30764 17926
rect 30820 17924 30844 17926
rect 30900 17924 30924 17926
rect 30980 17924 31004 17926
rect 31060 17924 31066 17926
rect 30758 17915 31066 17924
rect 30656 17876 30708 17882
rect 30656 17818 30708 17824
rect 30564 17332 30616 17338
rect 30564 17274 30616 17280
rect 30380 16244 30432 16250
rect 30380 16186 30432 16192
rect 30472 16244 30524 16250
rect 30472 16186 30524 16192
rect 30196 16040 30248 16046
rect 30196 15982 30248 15988
rect 30196 15904 30248 15910
rect 30196 15846 30248 15852
rect 30472 15904 30524 15910
rect 30472 15846 30524 15852
rect 30208 14958 30236 15846
rect 30484 14958 30512 15846
rect 30196 14952 30248 14958
rect 30196 14894 30248 14900
rect 30472 14952 30524 14958
rect 30472 14894 30524 14900
rect 30208 14482 30236 14894
rect 30196 14476 30248 14482
rect 30196 14418 30248 14424
rect 30576 14074 30604 17274
rect 30668 15162 30696 17818
rect 30758 16892 31066 16901
rect 30758 16890 30764 16892
rect 30820 16890 30844 16892
rect 30900 16890 30924 16892
rect 30980 16890 31004 16892
rect 31060 16890 31066 16892
rect 30820 16838 30822 16890
rect 31002 16838 31004 16890
rect 30758 16836 30764 16838
rect 30820 16836 30844 16838
rect 30900 16836 30924 16838
rect 30980 16836 31004 16838
rect 31060 16836 31066 16838
rect 30758 16827 31066 16836
rect 31116 16652 31168 16658
rect 31116 16594 31168 16600
rect 30758 15804 31066 15813
rect 30758 15802 30764 15804
rect 30820 15802 30844 15804
rect 30900 15802 30924 15804
rect 30980 15802 31004 15804
rect 31060 15802 31066 15804
rect 30820 15750 30822 15802
rect 31002 15750 31004 15802
rect 30758 15748 30764 15750
rect 30820 15748 30844 15750
rect 30900 15748 30924 15750
rect 30980 15748 31004 15750
rect 31060 15748 31066 15750
rect 30758 15739 31066 15748
rect 30656 15156 30708 15162
rect 30656 15098 30708 15104
rect 30758 14716 31066 14725
rect 30758 14714 30764 14716
rect 30820 14714 30844 14716
rect 30900 14714 30924 14716
rect 30980 14714 31004 14716
rect 31060 14714 31066 14716
rect 30820 14662 30822 14714
rect 31002 14662 31004 14714
rect 30758 14660 30764 14662
rect 30820 14660 30844 14662
rect 30900 14660 30924 14662
rect 30980 14660 31004 14662
rect 31060 14660 31066 14662
rect 30758 14651 31066 14660
rect 30564 14068 30616 14074
rect 30564 14010 30616 14016
rect 30472 13932 30524 13938
rect 30472 13874 30524 13880
rect 30104 13796 30156 13802
rect 30104 13738 30156 13744
rect 30012 12776 30064 12782
rect 29656 12430 29868 12458
rect 29932 12736 30012 12764
rect 29656 11830 29684 12430
rect 29644 11824 29696 11830
rect 29644 11766 29696 11772
rect 29512 10560 29592 10588
rect 29460 10542 29512 10548
rect 29368 8492 29420 8498
rect 29368 8434 29420 8440
rect 29380 7342 29408 8434
rect 29368 7336 29420 7342
rect 29368 7278 29420 7284
rect 29276 6248 29328 6254
rect 29276 6190 29328 6196
rect 29366 6216 29422 6225
rect 29366 6151 29422 6160
rect 29184 5568 29236 5574
rect 29184 5510 29236 5516
rect 29196 4826 29224 5510
rect 29184 4820 29236 4826
rect 29184 4762 29236 4768
rect 29182 4176 29238 4185
rect 29182 4111 29238 4120
rect 29092 3052 29144 3058
rect 29092 2994 29144 3000
rect 29104 2446 29132 2994
rect 29092 2440 29144 2446
rect 29092 2382 29144 2388
rect 29196 2106 29224 4111
rect 29276 2984 29328 2990
rect 29276 2926 29328 2932
rect 29184 2100 29236 2106
rect 29184 2042 29236 2048
rect 28816 1964 28868 1970
rect 28816 1906 28868 1912
rect 29000 1896 29052 1902
rect 28998 1864 29000 1873
rect 29052 1864 29054 1873
rect 28998 1799 29054 1808
rect 28724 1760 28776 1766
rect 28724 1702 28776 1708
rect 28630 1456 28686 1465
rect 28630 1391 28632 1400
rect 28684 1391 28686 1400
rect 28632 1362 28684 1368
rect 28736 1329 28764 1702
rect 29012 1426 29040 1799
rect 29000 1420 29052 1426
rect 29000 1362 29052 1368
rect 28722 1320 28778 1329
rect 28722 1255 28778 1264
rect 28632 1216 28684 1222
rect 28632 1158 28684 1164
rect 28540 1012 28592 1018
rect 28540 954 28592 960
rect 28644 270 28672 1158
rect 29288 785 29316 2926
rect 29380 2650 29408 6151
rect 29472 5914 29500 10542
rect 29656 8566 29684 11766
rect 29932 10810 29960 12736
rect 30012 12718 30064 12724
rect 30484 12306 30512 13874
rect 30758 13628 31066 13637
rect 30758 13626 30764 13628
rect 30820 13626 30844 13628
rect 30900 13626 30924 13628
rect 30980 13626 31004 13628
rect 31060 13626 31066 13628
rect 30820 13574 30822 13626
rect 31002 13574 31004 13626
rect 30758 13572 30764 13574
rect 30820 13572 30844 13574
rect 30900 13572 30924 13574
rect 30980 13572 31004 13574
rect 31060 13572 31066 13574
rect 30758 13563 31066 13572
rect 30758 12540 31066 12549
rect 30758 12538 30764 12540
rect 30820 12538 30844 12540
rect 30900 12538 30924 12540
rect 30980 12538 31004 12540
rect 31060 12538 31066 12540
rect 30820 12486 30822 12538
rect 31002 12486 31004 12538
rect 30758 12484 30764 12486
rect 30820 12484 30844 12486
rect 30900 12484 30924 12486
rect 30980 12484 31004 12486
rect 31060 12484 31066 12486
rect 30758 12475 31066 12484
rect 30472 12300 30524 12306
rect 30472 12242 30524 12248
rect 30288 11212 30340 11218
rect 30288 11154 30340 11160
rect 30010 11112 30066 11121
rect 30010 11047 30012 11056
rect 30064 11047 30066 11056
rect 30012 11018 30064 11024
rect 29920 10804 29972 10810
rect 29920 10746 29972 10752
rect 29736 10464 29788 10470
rect 29736 10406 29788 10412
rect 29748 9654 29776 10406
rect 29932 10266 29960 10746
rect 30300 10742 30328 11154
rect 30288 10736 30340 10742
rect 30288 10678 30340 10684
rect 30484 10538 30512 12242
rect 30758 11452 31066 11461
rect 30758 11450 30764 11452
rect 30820 11450 30844 11452
rect 30900 11450 30924 11452
rect 30980 11450 31004 11452
rect 31060 11450 31066 11452
rect 30820 11398 30822 11450
rect 31002 11398 31004 11450
rect 30758 11396 30764 11398
rect 30820 11396 30844 11398
rect 30900 11396 30924 11398
rect 30980 11396 31004 11398
rect 31060 11396 31066 11398
rect 30758 11387 31066 11396
rect 30472 10532 30524 10538
rect 30472 10474 30524 10480
rect 29920 10260 29972 10266
rect 29920 10202 29972 10208
rect 30012 9920 30064 9926
rect 30012 9862 30064 9868
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 29736 9648 29788 9654
rect 29736 9590 29788 9596
rect 30024 9042 30052 9862
rect 30012 9036 30064 9042
rect 30012 8978 30064 8984
rect 29644 8560 29696 8566
rect 29644 8502 29696 8508
rect 29552 7880 29604 7886
rect 29552 7822 29604 7828
rect 29460 5908 29512 5914
rect 29460 5850 29512 5856
rect 29458 5672 29514 5681
rect 29458 5607 29514 5616
rect 29472 5574 29500 5607
rect 29460 5568 29512 5574
rect 29460 5510 29512 5516
rect 29564 4146 29592 7822
rect 29656 6458 29684 8502
rect 30116 7954 30144 9862
rect 30484 9518 30512 10474
rect 30758 10364 31066 10373
rect 30758 10362 30764 10364
rect 30820 10362 30844 10364
rect 30900 10362 30924 10364
rect 30980 10362 31004 10364
rect 31060 10362 31066 10364
rect 30820 10310 30822 10362
rect 31002 10310 31004 10362
rect 30758 10308 30764 10310
rect 30820 10308 30844 10310
rect 30900 10308 30924 10310
rect 30980 10308 31004 10310
rect 31060 10308 31066 10310
rect 30758 10299 31066 10308
rect 30472 9512 30524 9518
rect 30472 9454 30524 9460
rect 30288 9376 30340 9382
rect 30288 9318 30340 9324
rect 30196 8628 30248 8634
rect 30196 8570 30248 8576
rect 30208 8090 30236 8570
rect 30196 8084 30248 8090
rect 30196 8026 30248 8032
rect 30104 7948 30156 7954
rect 30104 7890 30156 7896
rect 30104 7744 30156 7750
rect 30104 7686 30156 7692
rect 29736 7200 29788 7206
rect 29736 7142 29788 7148
rect 29644 6452 29696 6458
rect 29644 6394 29696 6400
rect 29552 4140 29604 4146
rect 29552 4082 29604 4088
rect 29564 3466 29592 4082
rect 29552 3460 29604 3466
rect 29552 3402 29604 3408
rect 29748 2774 29776 7142
rect 30116 4690 30144 7686
rect 30300 6866 30328 9318
rect 30288 6860 30340 6866
rect 30288 6802 30340 6808
rect 30104 4684 30156 4690
rect 30104 4626 30156 4632
rect 29656 2746 29776 2774
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 29460 2440 29512 2446
rect 29460 2382 29512 2388
rect 29368 2304 29420 2310
rect 29368 2246 29420 2252
rect 29380 1562 29408 2246
rect 29368 1556 29420 1562
rect 29368 1498 29420 1504
rect 29368 1420 29420 1426
rect 29472 1408 29500 2382
rect 29656 2106 29684 2746
rect 29644 2100 29696 2106
rect 29644 2042 29696 2048
rect 30484 1465 30512 9454
rect 30758 9276 31066 9285
rect 30758 9274 30764 9276
rect 30820 9274 30844 9276
rect 30900 9274 30924 9276
rect 30980 9274 31004 9276
rect 31060 9274 31066 9276
rect 30820 9222 30822 9274
rect 31002 9222 31004 9274
rect 30758 9220 30764 9222
rect 30820 9220 30844 9222
rect 30900 9220 30924 9222
rect 30980 9220 31004 9222
rect 31060 9220 31066 9222
rect 30758 9211 31066 9220
rect 31128 9178 31156 16594
rect 31312 14550 31340 21286
rect 31392 20324 31444 20330
rect 31392 20266 31444 20272
rect 31300 14544 31352 14550
rect 31300 14486 31352 14492
rect 31404 13297 31432 20266
rect 31390 13288 31446 13297
rect 31390 13223 31446 13232
rect 31116 9172 31168 9178
rect 31116 9114 31168 9120
rect 30758 8188 31066 8197
rect 30758 8186 30764 8188
rect 30820 8186 30844 8188
rect 30900 8186 30924 8188
rect 30980 8186 31004 8188
rect 31060 8186 31066 8188
rect 30820 8134 30822 8186
rect 31002 8134 31004 8186
rect 30758 8132 30764 8134
rect 30820 8132 30844 8134
rect 30900 8132 30924 8134
rect 30980 8132 31004 8134
rect 31060 8132 31066 8134
rect 30758 8123 31066 8132
rect 30758 7100 31066 7109
rect 30758 7098 30764 7100
rect 30820 7098 30844 7100
rect 30900 7098 30924 7100
rect 30980 7098 31004 7100
rect 31060 7098 31066 7100
rect 30820 7046 30822 7098
rect 31002 7046 31004 7098
rect 30758 7044 30764 7046
rect 30820 7044 30844 7046
rect 30900 7044 30924 7046
rect 30980 7044 31004 7046
rect 31060 7044 31066 7046
rect 30758 7035 31066 7044
rect 30758 6012 31066 6021
rect 30758 6010 30764 6012
rect 30820 6010 30844 6012
rect 30900 6010 30924 6012
rect 30980 6010 31004 6012
rect 31060 6010 31066 6012
rect 30820 5958 30822 6010
rect 31002 5958 31004 6010
rect 30758 5956 30764 5958
rect 30820 5956 30844 5958
rect 30900 5956 30924 5958
rect 30980 5956 31004 5958
rect 31060 5956 31066 5958
rect 30758 5947 31066 5956
rect 30758 4924 31066 4933
rect 30758 4922 30764 4924
rect 30820 4922 30844 4924
rect 30900 4922 30924 4924
rect 30980 4922 31004 4924
rect 31060 4922 31066 4924
rect 30820 4870 30822 4922
rect 31002 4870 31004 4922
rect 30758 4868 30764 4870
rect 30820 4868 30844 4870
rect 30900 4868 30924 4870
rect 30980 4868 31004 4870
rect 31060 4868 31066 4870
rect 30758 4859 31066 4868
rect 30758 3836 31066 3845
rect 30758 3834 30764 3836
rect 30820 3834 30844 3836
rect 30900 3834 30924 3836
rect 30980 3834 31004 3836
rect 31060 3834 31066 3836
rect 30820 3782 30822 3834
rect 31002 3782 31004 3834
rect 30758 3780 30764 3782
rect 30820 3780 30844 3782
rect 30900 3780 30924 3782
rect 30980 3780 31004 3782
rect 31060 3780 31066 3782
rect 30758 3771 31066 3780
rect 30758 2748 31066 2757
rect 30758 2746 30764 2748
rect 30820 2746 30844 2748
rect 30900 2746 30924 2748
rect 30980 2746 31004 2748
rect 31060 2746 31066 2748
rect 30820 2694 30822 2746
rect 31002 2694 31004 2746
rect 30758 2692 30764 2694
rect 30820 2692 30844 2694
rect 30900 2692 30924 2694
rect 30980 2692 31004 2694
rect 31060 2692 31066 2694
rect 30758 2683 31066 2692
rect 30758 1660 31066 1669
rect 30758 1658 30764 1660
rect 30820 1658 30844 1660
rect 30900 1658 30924 1660
rect 30980 1658 31004 1660
rect 31060 1658 31066 1660
rect 30820 1606 30822 1658
rect 31002 1606 31004 1658
rect 30758 1604 30764 1606
rect 30820 1604 30844 1606
rect 30900 1604 30924 1606
rect 30980 1604 31004 1606
rect 31060 1604 31066 1606
rect 30758 1595 31066 1604
rect 29420 1380 29500 1408
rect 30470 1456 30526 1465
rect 30470 1391 30526 1400
rect 29368 1362 29420 1368
rect 29368 1216 29420 1222
rect 29368 1158 29420 1164
rect 29274 776 29330 785
rect 29274 711 29330 720
rect 29380 377 29408 1158
rect 29472 814 29500 1380
rect 29460 808 29512 814
rect 29460 750 29512 756
rect 30758 572 31066 581
rect 30758 570 30764 572
rect 30820 570 30844 572
rect 30900 570 30924 572
rect 30980 570 31004 572
rect 31060 570 31066 572
rect 30820 518 30822 570
rect 31002 518 31004 570
rect 30758 516 30764 518
rect 30820 516 30844 518
rect 30900 516 30924 518
rect 30980 516 31004 518
rect 31060 516 31066 518
rect 30758 507 31066 516
rect 29366 368 29422 377
rect 29366 303 29422 312
rect 28632 264 28684 270
rect 28632 206 28684 212
rect 28356 196 28408 202
rect 28356 138 28408 144
rect 28078 96 28134 105
rect 18878 31 18934 40
rect 19708 60 19760 66
rect 18604 2 18656 8
rect 19708 2 19760 8
rect 26792 60 26844 66
rect 28078 31 28134 40
rect 26792 2 26844 8
<< via2 >>
rect 8850 22244 8852 22264
rect 8852 22244 8904 22264
rect 8904 22244 8906 22264
rect 1674 21528 1730 21584
rect 8850 22208 8906 22244
rect 9678 22244 9680 22264
rect 9680 22244 9732 22264
rect 9732 22244 9734 22264
rect 9678 22208 9734 22244
rect 1030 18828 1086 18864
rect 1582 20340 1584 20360
rect 1584 20340 1636 20360
rect 1636 20340 1638 20360
rect 1582 20304 1638 20340
rect 1582 19352 1638 19408
rect 1030 18808 1032 18828
rect 1032 18808 1084 18828
rect 1084 18808 1086 18828
rect 1582 18708 1584 18728
rect 1584 18708 1636 18728
rect 1636 18708 1638 18728
rect 1582 18672 1638 18708
rect 1674 17584 1730 17640
rect 2042 16088 2098 16144
rect 1950 15000 2006 15056
rect 1398 14476 1454 14512
rect 1398 14456 1400 14476
rect 1400 14456 1452 14476
rect 1452 14456 1454 14476
rect 2134 15408 2190 15464
rect 1030 9424 1086 9480
rect 1030 3848 1086 3904
rect 1398 11092 1400 11112
rect 1400 11092 1452 11112
rect 1452 11092 1454 11112
rect 1398 11056 1454 11092
rect 1674 11328 1730 11384
rect 1674 10104 1730 10160
rect 2134 13640 2190 13696
rect 2226 12552 2282 12608
rect 2134 10668 2190 10704
rect 2134 10648 2136 10668
rect 2136 10648 2188 10668
rect 2188 10648 2190 10668
rect 1766 7792 1822 7848
rect 1674 7248 1730 7304
rect 1766 6976 1822 7032
rect 1950 7384 2006 7440
rect 1582 4664 1638 4720
rect 2042 5752 2098 5808
rect 2042 3576 2098 3632
rect 1766 3440 1822 3496
rect 1674 3032 1730 3088
rect 1398 2760 1454 2816
rect 1858 2624 1914 2680
rect 2042 1944 2098 2000
rect 2410 11872 2466 11928
rect 3974 21528 4030 21584
rect 7194 22072 7250 22128
rect 4199 21786 4255 21788
rect 4279 21786 4335 21788
rect 4359 21786 4415 21788
rect 4439 21786 4495 21788
rect 4199 21734 4245 21786
rect 4245 21734 4255 21786
rect 4279 21734 4309 21786
rect 4309 21734 4321 21786
rect 4321 21734 4335 21786
rect 4359 21734 4373 21786
rect 4373 21734 4385 21786
rect 4385 21734 4415 21786
rect 4439 21734 4449 21786
rect 4449 21734 4495 21786
rect 4199 21732 4255 21734
rect 4279 21732 4335 21734
rect 4359 21732 4415 21734
rect 4439 21732 4495 21734
rect 4199 20698 4255 20700
rect 4279 20698 4335 20700
rect 4359 20698 4415 20700
rect 4439 20698 4495 20700
rect 4199 20646 4245 20698
rect 4245 20646 4255 20698
rect 4279 20646 4309 20698
rect 4309 20646 4321 20698
rect 4321 20646 4335 20698
rect 4359 20646 4373 20698
rect 4373 20646 4385 20698
rect 4385 20646 4415 20698
rect 4439 20646 4449 20698
rect 4449 20646 4495 20698
rect 4199 20644 4255 20646
rect 4279 20644 4335 20646
rect 4359 20644 4415 20646
rect 4439 20644 4495 20646
rect 4199 19610 4255 19612
rect 4279 19610 4335 19612
rect 4359 19610 4415 19612
rect 4439 19610 4495 19612
rect 4199 19558 4245 19610
rect 4245 19558 4255 19610
rect 4279 19558 4309 19610
rect 4309 19558 4321 19610
rect 4321 19558 4335 19610
rect 4359 19558 4373 19610
rect 4373 19558 4385 19610
rect 4385 19558 4415 19610
rect 4439 19558 4449 19610
rect 4449 19558 4495 19610
rect 4199 19556 4255 19558
rect 4279 19556 4335 19558
rect 4359 19556 4415 19558
rect 4439 19556 4495 19558
rect 3882 19080 3938 19136
rect 3698 18672 3754 18728
rect 3606 17856 3662 17912
rect 3330 14592 3386 14648
rect 3146 13388 3202 13424
rect 3146 13368 3148 13388
rect 3148 13368 3200 13388
rect 3200 13368 3202 13388
rect 3054 12688 3110 12744
rect 2686 12144 2742 12200
rect 3514 15544 3570 15600
rect 4618 18944 4674 19000
rect 5814 21664 5870 21720
rect 4199 18522 4255 18524
rect 4279 18522 4335 18524
rect 4359 18522 4415 18524
rect 4439 18522 4495 18524
rect 4199 18470 4245 18522
rect 4245 18470 4255 18522
rect 4279 18470 4309 18522
rect 4309 18470 4321 18522
rect 4321 18470 4335 18522
rect 4359 18470 4373 18522
rect 4373 18470 4385 18522
rect 4385 18470 4415 18522
rect 4439 18470 4449 18522
rect 4449 18470 4495 18522
rect 4199 18468 4255 18470
rect 4279 18468 4335 18470
rect 4359 18468 4415 18470
rect 4439 18468 4495 18470
rect 4199 17434 4255 17436
rect 4279 17434 4335 17436
rect 4359 17434 4415 17436
rect 4439 17434 4495 17436
rect 4199 17382 4245 17434
rect 4245 17382 4255 17434
rect 4279 17382 4309 17434
rect 4309 17382 4321 17434
rect 4321 17382 4335 17434
rect 4359 17382 4373 17434
rect 4373 17382 4385 17434
rect 4385 17382 4415 17434
rect 4439 17382 4449 17434
rect 4449 17382 4495 17434
rect 4199 17380 4255 17382
rect 4279 17380 4335 17382
rect 4359 17380 4415 17382
rect 4439 17380 4495 17382
rect 4199 16346 4255 16348
rect 4279 16346 4335 16348
rect 4359 16346 4415 16348
rect 4439 16346 4495 16348
rect 4199 16294 4245 16346
rect 4245 16294 4255 16346
rect 4279 16294 4309 16346
rect 4309 16294 4321 16346
rect 4321 16294 4335 16346
rect 4359 16294 4373 16346
rect 4373 16294 4385 16346
rect 4385 16294 4415 16346
rect 4439 16294 4449 16346
rect 4449 16294 4495 16346
rect 4199 16292 4255 16294
rect 4279 16292 4335 16294
rect 4359 16292 4415 16294
rect 4439 16292 4495 16294
rect 4802 18808 4858 18864
rect 5170 19488 5226 19544
rect 5078 18400 5134 18456
rect 4986 18128 5042 18184
rect 4710 16904 4766 16960
rect 4434 15988 4436 16008
rect 4436 15988 4488 16008
rect 4488 15988 4490 16008
rect 4434 15952 4490 15988
rect 4199 15258 4255 15260
rect 4279 15258 4335 15260
rect 4359 15258 4415 15260
rect 4439 15258 4495 15260
rect 4199 15206 4245 15258
rect 4245 15206 4255 15258
rect 4279 15206 4309 15258
rect 4309 15206 4321 15258
rect 4321 15206 4335 15258
rect 4359 15206 4373 15258
rect 4373 15206 4385 15258
rect 4385 15206 4415 15258
rect 4439 15206 4449 15258
rect 4449 15206 4495 15258
rect 4199 15204 4255 15206
rect 4279 15204 4335 15206
rect 4359 15204 4415 15206
rect 4439 15204 4495 15206
rect 3974 15000 4030 15056
rect 4434 14476 4490 14512
rect 4434 14456 4436 14476
rect 4436 14456 4488 14476
rect 4488 14456 4490 14476
rect 3330 13268 3332 13288
rect 3332 13268 3384 13288
rect 3384 13268 3386 13288
rect 3330 13232 3386 13268
rect 3514 12824 3570 12880
rect 3238 11076 3294 11112
rect 3238 11056 3240 11076
rect 3240 11056 3292 11076
rect 3292 11056 3294 11076
rect 3238 10376 3294 10432
rect 3146 10240 3202 10296
rect 2870 9016 2926 9072
rect 3146 8916 3148 8936
rect 3148 8916 3200 8936
rect 3200 8916 3202 8936
rect 3146 8880 3202 8916
rect 2594 6704 2650 6760
rect 2594 5208 2650 5264
rect 2686 4936 2742 4992
rect 2870 4936 2926 4992
rect 3146 7112 3202 7168
rect 3514 11464 3570 11520
rect 3698 11056 3754 11112
rect 4199 14170 4255 14172
rect 4279 14170 4335 14172
rect 4359 14170 4415 14172
rect 4439 14170 4495 14172
rect 4199 14118 4245 14170
rect 4245 14118 4255 14170
rect 4279 14118 4309 14170
rect 4309 14118 4321 14170
rect 4321 14118 4335 14170
rect 4359 14118 4373 14170
rect 4373 14118 4385 14170
rect 4385 14118 4415 14170
rect 4439 14118 4449 14170
rect 4449 14118 4495 14170
rect 4199 14116 4255 14118
rect 4279 14116 4335 14118
rect 4359 14116 4415 14118
rect 4439 14116 4495 14118
rect 4199 13082 4255 13084
rect 4279 13082 4335 13084
rect 4359 13082 4415 13084
rect 4439 13082 4495 13084
rect 4199 13030 4245 13082
rect 4245 13030 4255 13082
rect 4279 13030 4309 13082
rect 4309 13030 4321 13082
rect 4321 13030 4335 13082
rect 4359 13030 4373 13082
rect 4373 13030 4385 13082
rect 4385 13030 4415 13082
rect 4439 13030 4449 13082
rect 4449 13030 4495 13082
rect 4199 13028 4255 13030
rect 4279 13028 4335 13030
rect 4359 13028 4415 13030
rect 4439 13028 4495 13030
rect 4250 12688 4306 12744
rect 4199 11994 4255 11996
rect 4279 11994 4335 11996
rect 4359 11994 4415 11996
rect 4439 11994 4495 11996
rect 4199 11942 4245 11994
rect 4245 11942 4255 11994
rect 4279 11942 4309 11994
rect 4309 11942 4321 11994
rect 4321 11942 4335 11994
rect 4359 11942 4373 11994
rect 4373 11942 4385 11994
rect 4385 11942 4415 11994
rect 4439 11942 4449 11994
rect 4449 11942 4495 11994
rect 4199 11940 4255 11942
rect 4279 11940 4335 11942
rect 4359 11940 4415 11942
rect 4439 11940 4495 11942
rect 3882 11228 3884 11248
rect 3884 11228 3936 11248
rect 3936 11228 3938 11248
rect 3882 11192 3938 11228
rect 4199 10906 4255 10908
rect 4279 10906 4335 10908
rect 4359 10906 4415 10908
rect 4439 10906 4495 10908
rect 4199 10854 4245 10906
rect 4245 10854 4255 10906
rect 4279 10854 4309 10906
rect 4309 10854 4321 10906
rect 4321 10854 4335 10906
rect 4359 10854 4373 10906
rect 4373 10854 4385 10906
rect 4385 10854 4415 10906
rect 4439 10854 4449 10906
rect 4449 10854 4495 10906
rect 4199 10852 4255 10854
rect 4279 10852 4335 10854
rect 4359 10852 4415 10854
rect 4439 10852 4495 10854
rect 3974 10376 4030 10432
rect 4066 9968 4122 10024
rect 4066 9832 4122 9888
rect 3974 8492 4030 8528
rect 3974 8472 3976 8492
rect 3976 8472 4028 8492
rect 4028 8472 4030 8492
rect 4199 9818 4255 9820
rect 4279 9818 4335 9820
rect 4359 9818 4415 9820
rect 4439 9818 4495 9820
rect 4199 9766 4245 9818
rect 4245 9766 4255 9818
rect 4279 9766 4309 9818
rect 4309 9766 4321 9818
rect 4321 9766 4335 9818
rect 4359 9766 4373 9818
rect 4373 9766 4385 9818
rect 4385 9766 4415 9818
rect 4439 9766 4449 9818
rect 4449 9766 4495 9818
rect 4199 9764 4255 9766
rect 4279 9764 4335 9766
rect 4359 9764 4415 9766
rect 4439 9764 4495 9766
rect 4894 17992 4950 18048
rect 4894 16632 4950 16688
rect 5354 18536 5410 18592
rect 5354 18284 5410 18320
rect 5354 18264 5356 18284
rect 5356 18264 5408 18284
rect 5408 18264 5410 18284
rect 5078 15136 5134 15192
rect 5354 17720 5410 17776
rect 5722 20848 5778 20904
rect 5630 18400 5686 18456
rect 5814 20748 5816 20768
rect 5816 20748 5868 20768
rect 5868 20748 5870 20768
rect 5814 20712 5870 20748
rect 6182 21120 6238 21176
rect 5998 20032 6054 20088
rect 5998 19932 6000 19952
rect 6000 19932 6052 19952
rect 6052 19932 6054 19952
rect 5998 19896 6054 19932
rect 6182 20340 6184 20360
rect 6184 20340 6236 20360
rect 6236 20340 6238 20360
rect 6182 20304 6238 20340
rect 6826 21392 6882 21448
rect 7194 21120 7250 21176
rect 7286 20596 7342 20632
rect 7286 20576 7288 20596
rect 7288 20576 7340 20596
rect 7340 20576 7342 20596
rect 6826 19760 6882 19816
rect 6642 19352 6698 19408
rect 5262 16904 5318 16960
rect 5170 14728 5226 14784
rect 5354 15000 5410 15056
rect 4894 13504 4950 13560
rect 5446 13368 5502 13424
rect 5814 15000 5870 15056
rect 5998 15272 6054 15328
rect 5630 14184 5686 14240
rect 5722 14068 5778 14104
rect 5722 14048 5724 14068
rect 5724 14048 5776 14068
rect 5776 14048 5778 14068
rect 6550 17992 6606 18048
rect 6458 16224 6514 16280
rect 6182 14592 6238 14648
rect 6366 14456 6422 14512
rect 7378 18536 7434 18592
rect 6826 18128 6882 18184
rect 6826 17076 6828 17096
rect 6828 17076 6880 17096
rect 6880 17076 6882 17096
rect 6826 17040 6882 17076
rect 7562 19216 7618 19272
rect 7194 15000 7250 15056
rect 7470 16360 7526 16416
rect 7746 17856 7802 17912
rect 7994 21242 8050 21244
rect 8074 21242 8130 21244
rect 8154 21242 8210 21244
rect 8234 21242 8290 21244
rect 7994 21190 8040 21242
rect 8040 21190 8050 21242
rect 8074 21190 8104 21242
rect 8104 21190 8116 21242
rect 8116 21190 8130 21242
rect 8154 21190 8168 21242
rect 8168 21190 8180 21242
rect 8180 21190 8210 21242
rect 8234 21190 8244 21242
rect 8244 21190 8290 21242
rect 7994 21188 8050 21190
rect 8074 21188 8130 21190
rect 8154 21188 8210 21190
rect 8234 21188 8290 21190
rect 8022 21004 8078 21040
rect 8022 20984 8024 21004
rect 8024 20984 8076 21004
rect 8076 20984 8078 21004
rect 8574 21256 8630 21312
rect 8850 21664 8906 21720
rect 8850 20884 8852 20904
rect 8852 20884 8904 20904
rect 8904 20884 8906 20904
rect 8482 20712 8538 20768
rect 8390 20324 8446 20360
rect 8390 20304 8392 20324
rect 8392 20304 8444 20324
rect 8444 20304 8446 20324
rect 7994 20154 8050 20156
rect 8074 20154 8130 20156
rect 8154 20154 8210 20156
rect 8234 20154 8290 20156
rect 7994 20102 8040 20154
rect 8040 20102 8050 20154
rect 8074 20102 8104 20154
rect 8104 20102 8116 20154
rect 8116 20102 8130 20154
rect 8154 20102 8168 20154
rect 8168 20102 8180 20154
rect 8180 20102 8210 20154
rect 8234 20102 8244 20154
rect 8244 20102 8290 20154
rect 7994 20100 8050 20102
rect 8074 20100 8130 20102
rect 8154 20100 8210 20102
rect 8234 20100 8290 20102
rect 8482 20032 8538 20088
rect 8850 20848 8906 20884
rect 8850 20576 8906 20632
rect 8850 19896 8906 19952
rect 7994 19066 8050 19068
rect 8074 19066 8130 19068
rect 8154 19066 8210 19068
rect 8234 19066 8290 19068
rect 7994 19014 8040 19066
rect 8040 19014 8050 19066
rect 8074 19014 8104 19066
rect 8104 19014 8116 19066
rect 8116 19014 8130 19066
rect 8154 19014 8168 19066
rect 8168 19014 8180 19066
rect 8180 19014 8210 19066
rect 8234 19014 8244 19066
rect 8244 19014 8290 19066
rect 7994 19012 8050 19014
rect 8074 19012 8130 19014
rect 8154 19012 8210 19014
rect 8234 19012 8290 19014
rect 8850 19116 8852 19136
rect 8852 19116 8904 19136
rect 8904 19116 8906 19136
rect 8850 19080 8906 19116
rect 8114 18536 8170 18592
rect 8298 18536 8354 18592
rect 7994 17978 8050 17980
rect 8074 17978 8130 17980
rect 8154 17978 8210 17980
rect 8234 17978 8290 17980
rect 7994 17926 8040 17978
rect 8040 17926 8050 17978
rect 8074 17926 8104 17978
rect 8104 17926 8116 17978
rect 8116 17926 8130 17978
rect 8154 17926 8168 17978
rect 8168 17926 8180 17978
rect 8180 17926 8210 17978
rect 8234 17926 8244 17978
rect 8244 17926 8290 17978
rect 7994 17924 8050 17926
rect 8074 17924 8130 17926
rect 8154 17924 8210 17926
rect 8234 17924 8290 17926
rect 8666 17992 8722 18048
rect 7838 17584 7894 17640
rect 7746 17448 7802 17504
rect 7994 16890 8050 16892
rect 8074 16890 8130 16892
rect 8154 16890 8210 16892
rect 8234 16890 8290 16892
rect 7994 16838 8040 16890
rect 8040 16838 8050 16890
rect 8074 16838 8104 16890
rect 8104 16838 8116 16890
rect 8116 16838 8130 16890
rect 8154 16838 8168 16890
rect 8168 16838 8180 16890
rect 8180 16838 8210 16890
rect 8234 16838 8244 16890
rect 8244 16838 8290 16890
rect 7994 16836 8050 16838
rect 8074 16836 8130 16838
rect 8154 16836 8210 16838
rect 8234 16836 8290 16838
rect 8390 16768 8446 16824
rect 7994 15802 8050 15804
rect 8074 15802 8130 15804
rect 8154 15802 8210 15804
rect 8234 15802 8290 15804
rect 7994 15750 8040 15802
rect 8040 15750 8050 15802
rect 8074 15750 8104 15802
rect 8104 15750 8116 15802
rect 8116 15750 8130 15802
rect 8154 15750 8168 15802
rect 8168 15750 8180 15802
rect 8180 15750 8210 15802
rect 8234 15750 8244 15802
rect 8244 15750 8290 15802
rect 7994 15748 8050 15750
rect 8074 15748 8130 15750
rect 8154 15748 8210 15750
rect 8234 15748 8290 15750
rect 7746 15272 7802 15328
rect 7654 15136 7710 15192
rect 7102 14728 7158 14784
rect 6734 14456 6790 14512
rect 5262 12688 5318 12744
rect 4199 8730 4255 8732
rect 4279 8730 4335 8732
rect 4359 8730 4415 8732
rect 4439 8730 4495 8732
rect 4199 8678 4245 8730
rect 4245 8678 4255 8730
rect 4279 8678 4309 8730
rect 4309 8678 4321 8730
rect 4321 8678 4335 8730
rect 4359 8678 4373 8730
rect 4373 8678 4385 8730
rect 4385 8678 4415 8730
rect 4439 8678 4449 8730
rect 4449 8678 4495 8730
rect 4199 8676 4255 8678
rect 4279 8676 4335 8678
rect 4359 8676 4415 8678
rect 4439 8676 4495 8678
rect 3514 5888 3570 5944
rect 3054 3712 3110 3768
rect 3054 1536 3110 1592
rect 3238 4564 3240 4584
rect 3240 4564 3292 4584
rect 3292 4564 3294 4584
rect 3238 4528 3294 4564
rect 4066 7928 4122 7984
rect 4199 7642 4255 7644
rect 4279 7642 4335 7644
rect 4359 7642 4415 7644
rect 4439 7642 4495 7644
rect 4199 7590 4245 7642
rect 4245 7590 4255 7642
rect 4279 7590 4309 7642
rect 4309 7590 4321 7642
rect 4321 7590 4335 7642
rect 4359 7590 4373 7642
rect 4373 7590 4385 7642
rect 4385 7590 4415 7642
rect 4439 7590 4449 7642
rect 4449 7590 4495 7642
rect 4199 7588 4255 7590
rect 4279 7588 4335 7590
rect 4359 7588 4415 7590
rect 4439 7588 4495 7590
rect 5446 11600 5502 11656
rect 5078 11328 5134 11384
rect 4199 6554 4255 6556
rect 4279 6554 4335 6556
rect 4359 6554 4415 6556
rect 4439 6554 4495 6556
rect 4199 6502 4245 6554
rect 4245 6502 4255 6554
rect 4279 6502 4309 6554
rect 4309 6502 4321 6554
rect 4321 6502 4335 6554
rect 4359 6502 4373 6554
rect 4373 6502 4385 6554
rect 4385 6502 4415 6554
rect 4439 6502 4449 6554
rect 4449 6502 4495 6554
rect 4199 6500 4255 6502
rect 4279 6500 4335 6502
rect 4359 6500 4415 6502
rect 4439 6500 4495 6502
rect 4802 5480 4858 5536
rect 4199 5466 4255 5468
rect 4279 5466 4335 5468
rect 4359 5466 4415 5468
rect 4439 5466 4495 5468
rect 4199 5414 4245 5466
rect 4245 5414 4255 5466
rect 4279 5414 4309 5466
rect 4309 5414 4321 5466
rect 4321 5414 4335 5466
rect 4359 5414 4373 5466
rect 4373 5414 4385 5466
rect 4385 5414 4415 5466
rect 4439 5414 4449 5466
rect 4449 5414 4495 5466
rect 4199 5412 4255 5414
rect 4279 5412 4335 5414
rect 4359 5412 4415 5414
rect 4439 5412 4495 5414
rect 4066 4564 4068 4584
rect 4068 4564 4120 4584
rect 4120 4564 4122 4584
rect 4066 4528 4122 4564
rect 4199 4378 4255 4380
rect 4279 4378 4335 4380
rect 4359 4378 4415 4380
rect 4439 4378 4495 4380
rect 4199 4326 4245 4378
rect 4245 4326 4255 4378
rect 4279 4326 4309 4378
rect 4309 4326 4321 4378
rect 4321 4326 4335 4378
rect 4359 4326 4373 4378
rect 4373 4326 4385 4378
rect 4385 4326 4415 4378
rect 4439 4326 4449 4378
rect 4449 4326 4495 4378
rect 4199 4324 4255 4326
rect 4279 4324 4335 4326
rect 4359 4324 4415 4326
rect 4439 4324 4495 4326
rect 4526 4140 4582 4176
rect 4526 4120 4528 4140
rect 4528 4120 4580 4140
rect 4580 4120 4582 4140
rect 4158 3712 4214 3768
rect 3790 2624 3846 2680
rect 3238 2352 3294 2408
rect 4199 3290 4255 3292
rect 4279 3290 4335 3292
rect 4359 3290 4415 3292
rect 4439 3290 4495 3292
rect 4199 3238 4245 3290
rect 4245 3238 4255 3290
rect 4279 3238 4309 3290
rect 4309 3238 4321 3290
rect 4321 3238 4335 3290
rect 4359 3238 4373 3290
rect 4373 3238 4385 3290
rect 4385 3238 4415 3290
rect 4439 3238 4449 3290
rect 4449 3238 4495 3290
rect 4199 3236 4255 3238
rect 4279 3236 4335 3238
rect 4359 3236 4415 3238
rect 4439 3236 4495 3238
rect 4158 2796 4160 2816
rect 4160 2796 4212 2816
rect 4212 2796 4214 2816
rect 4158 2760 4214 2796
rect 3974 2388 3976 2408
rect 3976 2388 4028 2408
rect 4028 2388 4030 2408
rect 3974 2352 4030 2388
rect 4199 2202 4255 2204
rect 4279 2202 4335 2204
rect 4359 2202 4415 2204
rect 4439 2202 4495 2204
rect 4199 2150 4245 2202
rect 4245 2150 4255 2202
rect 4279 2150 4309 2202
rect 4309 2150 4321 2202
rect 4321 2150 4335 2202
rect 4359 2150 4373 2202
rect 4373 2150 4385 2202
rect 4385 2150 4415 2202
rect 4439 2150 4449 2202
rect 4449 2150 4495 2202
rect 4199 2148 4255 2150
rect 4279 2148 4335 2150
rect 4359 2148 4415 2150
rect 4439 2148 4495 2150
rect 4526 1944 4582 2000
rect 6458 12416 6514 12472
rect 5906 11872 5962 11928
rect 5262 9424 5318 9480
rect 5262 9052 5264 9072
rect 5264 9052 5316 9072
rect 5316 9052 5318 9072
rect 5262 9016 5318 9052
rect 5446 8780 5448 8800
rect 5448 8780 5500 8800
rect 5500 8780 5502 8800
rect 5446 8744 5502 8780
rect 5630 9632 5686 9688
rect 5078 2624 5134 2680
rect 4526 1400 4582 1456
rect 4250 1300 4252 1320
rect 4252 1300 4304 1320
rect 4304 1300 4306 1320
rect 4250 1264 4306 1300
rect 4199 1114 4255 1116
rect 4279 1114 4335 1116
rect 4359 1114 4415 1116
rect 4439 1114 4495 1116
rect 4199 1062 4245 1114
rect 4245 1062 4255 1114
rect 4279 1062 4309 1114
rect 4309 1062 4321 1114
rect 4321 1062 4335 1114
rect 4359 1062 4373 1114
rect 4373 1062 4385 1114
rect 4385 1062 4415 1114
rect 4439 1062 4449 1114
rect 4449 1062 4495 1114
rect 4199 1060 4255 1062
rect 4279 1060 4335 1062
rect 4359 1060 4415 1062
rect 4439 1060 4495 1062
rect 4986 756 4988 776
rect 4988 756 5040 776
rect 5040 756 5042 776
rect 4986 720 5042 756
rect 5262 6160 5318 6216
rect 5446 4528 5502 4584
rect 5354 3984 5410 4040
rect 5814 9424 5870 9480
rect 5722 8336 5778 8392
rect 6182 11464 6238 11520
rect 5906 8064 5962 8120
rect 5906 6840 5962 6896
rect 7010 14068 7066 14104
rect 7010 14048 7012 14068
rect 7012 14048 7064 14068
rect 7064 14048 7066 14068
rect 7286 14184 7342 14240
rect 7102 13232 7158 13288
rect 7378 12416 7434 12472
rect 5722 5888 5778 5944
rect 5906 2896 5962 2952
rect 6090 6316 6146 6352
rect 6366 10104 6422 10160
rect 9218 20052 9274 20088
rect 9218 20032 9220 20052
rect 9220 20032 9272 20052
rect 9272 20032 9274 20052
rect 9494 19488 9550 19544
rect 8574 15000 8630 15056
rect 7994 14714 8050 14716
rect 8074 14714 8130 14716
rect 8154 14714 8210 14716
rect 8234 14714 8290 14716
rect 7994 14662 8040 14714
rect 8040 14662 8050 14714
rect 8074 14662 8104 14714
rect 8104 14662 8116 14714
rect 8116 14662 8130 14714
rect 8154 14662 8168 14714
rect 8168 14662 8180 14714
rect 8180 14662 8210 14714
rect 8234 14662 8244 14714
rect 8244 14662 8290 14714
rect 7994 14660 8050 14662
rect 8074 14660 8130 14662
rect 8154 14660 8210 14662
rect 8234 14660 8290 14662
rect 7994 13626 8050 13628
rect 8074 13626 8130 13628
rect 8154 13626 8210 13628
rect 8234 13626 8290 13628
rect 7994 13574 8040 13626
rect 8040 13574 8050 13626
rect 8074 13574 8104 13626
rect 8104 13574 8116 13626
rect 8116 13574 8130 13626
rect 8154 13574 8168 13626
rect 8168 13574 8180 13626
rect 8180 13574 8210 13626
rect 8234 13574 8244 13626
rect 8244 13574 8290 13626
rect 7994 13572 8050 13574
rect 8074 13572 8130 13574
rect 8154 13572 8210 13574
rect 8234 13572 8290 13574
rect 7654 13504 7710 13560
rect 9402 17584 9458 17640
rect 8850 16224 8906 16280
rect 9034 16224 9090 16280
rect 9218 17176 9274 17232
rect 9310 16768 9366 16824
rect 9126 15408 9182 15464
rect 9218 15020 9274 15056
rect 9218 15000 9220 15020
rect 9220 15000 9272 15020
rect 9272 15000 9274 15020
rect 9218 14864 9274 14920
rect 10322 21936 10378 21992
rect 9770 19896 9826 19952
rect 9678 18536 9734 18592
rect 9678 18400 9734 18456
rect 9862 17720 9918 17776
rect 9770 17584 9826 17640
rect 9494 15544 9550 15600
rect 9862 16224 9918 16280
rect 9678 14048 9734 14104
rect 7994 12538 8050 12540
rect 8074 12538 8130 12540
rect 8154 12538 8210 12540
rect 8234 12538 8290 12540
rect 7994 12486 8040 12538
rect 8040 12486 8050 12538
rect 8074 12486 8104 12538
rect 8104 12486 8116 12538
rect 8116 12486 8130 12538
rect 8154 12486 8168 12538
rect 8168 12486 8180 12538
rect 8180 12486 8210 12538
rect 8234 12486 8244 12538
rect 8244 12486 8290 12538
rect 7994 12484 8050 12486
rect 8074 12484 8130 12486
rect 8154 12484 8210 12486
rect 8234 12484 8290 12486
rect 6550 9832 6606 9888
rect 7378 11464 7434 11520
rect 7994 11450 8050 11452
rect 8074 11450 8130 11452
rect 8154 11450 8210 11452
rect 8234 11450 8290 11452
rect 7994 11398 8040 11450
rect 8040 11398 8050 11450
rect 8074 11398 8104 11450
rect 8104 11398 8116 11450
rect 8116 11398 8130 11450
rect 8154 11398 8168 11450
rect 8168 11398 8180 11450
rect 8180 11398 8210 11450
rect 8234 11398 8244 11450
rect 8244 11398 8290 11450
rect 7994 11396 8050 11398
rect 8074 11396 8130 11398
rect 8154 11396 8210 11398
rect 8234 11396 8290 11398
rect 7010 9832 7066 9888
rect 6274 8336 6330 8392
rect 6550 7928 6606 7984
rect 6090 6296 6092 6316
rect 6092 6296 6144 6316
rect 6144 6296 6146 6316
rect 6366 5616 6422 5672
rect 6734 7928 6790 7984
rect 6918 8064 6974 8120
rect 7470 9036 7526 9072
rect 7470 9016 7472 9036
rect 7472 9016 7524 9036
rect 7524 9016 7526 9036
rect 7994 10362 8050 10364
rect 8074 10362 8130 10364
rect 8154 10362 8210 10364
rect 8234 10362 8290 10364
rect 7994 10310 8040 10362
rect 8040 10310 8050 10362
rect 8074 10310 8104 10362
rect 8104 10310 8116 10362
rect 8116 10310 8130 10362
rect 8154 10310 8168 10362
rect 8168 10310 8180 10362
rect 8180 10310 8210 10362
rect 8234 10310 8244 10362
rect 8244 10310 8290 10362
rect 7994 10308 8050 10310
rect 8074 10308 8130 10310
rect 8154 10308 8210 10310
rect 8234 10308 8290 10310
rect 8850 11328 8906 11384
rect 9126 12724 9128 12744
rect 9128 12724 9180 12744
rect 9180 12724 9182 12744
rect 9126 12688 9182 12724
rect 9862 14320 9918 14376
rect 10322 20596 10378 20632
rect 10322 20576 10324 20596
rect 10324 20576 10376 20596
rect 10376 20576 10378 20596
rect 10322 18944 10378 19000
rect 9126 11872 9182 11928
rect 7994 9274 8050 9276
rect 8074 9274 8130 9276
rect 8154 9274 8210 9276
rect 8234 9274 8290 9276
rect 7994 9222 8040 9274
rect 8040 9222 8050 9274
rect 8074 9222 8104 9274
rect 8104 9222 8116 9274
rect 8116 9222 8130 9274
rect 8154 9222 8168 9274
rect 8168 9222 8180 9274
rect 8180 9222 8210 9274
rect 8234 9222 8244 9274
rect 8244 9222 8290 9274
rect 7994 9220 8050 9222
rect 8074 9220 8130 9222
rect 8154 9220 8210 9222
rect 8234 9220 8290 9222
rect 7194 6840 7250 6896
rect 7378 6976 7434 7032
rect 7654 7112 7710 7168
rect 7994 8186 8050 8188
rect 8074 8186 8130 8188
rect 8154 8186 8210 8188
rect 8234 8186 8290 8188
rect 7994 8134 8040 8186
rect 8040 8134 8050 8186
rect 8074 8134 8104 8186
rect 8104 8134 8116 8186
rect 8116 8134 8130 8186
rect 8154 8134 8168 8186
rect 8168 8134 8180 8186
rect 8180 8134 8210 8186
rect 8234 8134 8244 8186
rect 8244 8134 8290 8186
rect 7994 8132 8050 8134
rect 8074 8132 8130 8134
rect 8154 8132 8210 8134
rect 8234 8132 8290 8134
rect 8114 7520 8170 7576
rect 8666 7656 8722 7712
rect 7994 7098 8050 7100
rect 8074 7098 8130 7100
rect 8154 7098 8210 7100
rect 8234 7098 8290 7100
rect 7994 7046 8040 7098
rect 8040 7046 8050 7098
rect 8074 7046 8104 7098
rect 8104 7046 8116 7098
rect 8116 7046 8130 7098
rect 8154 7046 8168 7098
rect 8168 7046 8180 7098
rect 8180 7046 8210 7098
rect 8234 7046 8244 7098
rect 8244 7046 8290 7098
rect 7994 7044 8050 7046
rect 8074 7044 8130 7046
rect 8154 7044 8210 7046
rect 8234 7044 8290 7046
rect 10230 16632 10286 16688
rect 10322 14592 10378 14648
rect 10138 14048 10194 14104
rect 12438 21936 12494 21992
rect 11789 21786 11845 21788
rect 11869 21786 11925 21788
rect 11949 21786 12005 21788
rect 12029 21786 12085 21788
rect 11789 21734 11835 21786
rect 11835 21734 11845 21786
rect 11869 21734 11899 21786
rect 11899 21734 11911 21786
rect 11911 21734 11925 21786
rect 11949 21734 11963 21786
rect 11963 21734 11975 21786
rect 11975 21734 12005 21786
rect 12029 21734 12039 21786
rect 12039 21734 12085 21786
rect 11789 21732 11845 21734
rect 11869 21732 11925 21734
rect 11949 21732 12005 21734
rect 12029 21732 12085 21734
rect 11058 21428 11060 21448
rect 11060 21428 11112 21448
rect 11112 21428 11114 21448
rect 10874 21256 10930 21312
rect 11058 21392 11114 21428
rect 10782 20848 10838 20904
rect 10874 20304 10930 20360
rect 10874 18944 10930 19000
rect 10506 15952 10562 16008
rect 10690 16360 10746 16416
rect 10690 15952 10746 16008
rect 11058 19624 11114 19680
rect 11058 19252 11060 19272
rect 11060 19252 11112 19272
rect 11112 19252 11114 19272
rect 11058 19216 11114 19252
rect 11242 17720 11298 17776
rect 11058 17448 11114 17504
rect 9862 12688 9918 12744
rect 9770 11328 9826 11384
rect 9770 11056 9826 11112
rect 10414 13640 10470 13696
rect 10046 12980 10102 13016
rect 10046 12960 10048 12980
rect 10048 12960 10100 12980
rect 10100 12960 10102 12980
rect 10874 13776 10930 13832
rect 10782 13640 10838 13696
rect 11426 16668 11428 16688
rect 11428 16668 11480 16688
rect 11480 16668 11482 16688
rect 11426 16632 11482 16668
rect 11426 15544 11482 15600
rect 11518 15136 11574 15192
rect 11334 14764 11336 14784
rect 11336 14764 11388 14784
rect 11388 14764 11390 14784
rect 11334 14728 11390 14764
rect 11242 14320 11298 14376
rect 11242 14184 11298 14240
rect 10966 12688 11022 12744
rect 11058 12552 11114 12608
rect 9954 10648 10010 10704
rect 9126 9016 9182 9072
rect 10046 9560 10102 9616
rect 10322 9016 10378 9072
rect 11426 14320 11482 14376
rect 11518 13676 11520 13696
rect 11520 13676 11572 13696
rect 11572 13676 11574 13696
rect 11518 13640 11574 13676
rect 12714 21256 12770 21312
rect 11702 20848 11758 20904
rect 11789 20698 11845 20700
rect 11869 20698 11925 20700
rect 11949 20698 12005 20700
rect 12029 20698 12085 20700
rect 11789 20646 11835 20698
rect 11835 20646 11845 20698
rect 11869 20646 11899 20698
rect 11899 20646 11911 20698
rect 11911 20646 11925 20698
rect 11949 20646 11963 20698
rect 11963 20646 11975 20698
rect 11975 20646 12005 20698
rect 12029 20646 12039 20698
rect 12039 20646 12085 20698
rect 11789 20644 11845 20646
rect 11869 20644 11925 20646
rect 11949 20644 12005 20646
rect 12029 20644 12085 20646
rect 11978 20304 12034 20360
rect 11789 19610 11845 19612
rect 11869 19610 11925 19612
rect 11949 19610 12005 19612
rect 12029 19610 12085 19612
rect 11789 19558 11835 19610
rect 11835 19558 11845 19610
rect 11869 19558 11899 19610
rect 11899 19558 11911 19610
rect 11911 19558 11925 19610
rect 11949 19558 11963 19610
rect 11963 19558 11975 19610
rect 11975 19558 12005 19610
rect 12029 19558 12039 19610
rect 12039 19558 12085 19610
rect 11789 19556 11845 19558
rect 11869 19556 11925 19558
rect 11949 19556 12005 19558
rect 12029 19556 12085 19558
rect 12530 20440 12586 20496
rect 11789 18522 11845 18524
rect 11869 18522 11925 18524
rect 11949 18522 12005 18524
rect 12029 18522 12085 18524
rect 11789 18470 11835 18522
rect 11835 18470 11845 18522
rect 11869 18470 11899 18522
rect 11899 18470 11911 18522
rect 11911 18470 11925 18522
rect 11949 18470 11963 18522
rect 11963 18470 11975 18522
rect 11975 18470 12005 18522
rect 12029 18470 12039 18522
rect 12039 18470 12085 18522
rect 11789 18468 11845 18470
rect 11869 18468 11925 18470
rect 11949 18468 12005 18470
rect 12029 18468 12085 18470
rect 11789 17434 11845 17436
rect 11869 17434 11925 17436
rect 11949 17434 12005 17436
rect 12029 17434 12085 17436
rect 11789 17382 11835 17434
rect 11835 17382 11845 17434
rect 11869 17382 11899 17434
rect 11899 17382 11911 17434
rect 11911 17382 11925 17434
rect 11949 17382 11963 17434
rect 11963 17382 11975 17434
rect 11975 17382 12005 17434
rect 12029 17382 12039 17434
rect 12039 17382 12085 17434
rect 11789 17380 11845 17382
rect 11869 17380 11925 17382
rect 11949 17380 12005 17382
rect 12029 17380 12085 17382
rect 11789 16346 11845 16348
rect 11869 16346 11925 16348
rect 11949 16346 12005 16348
rect 12029 16346 12085 16348
rect 11789 16294 11835 16346
rect 11835 16294 11845 16346
rect 11869 16294 11899 16346
rect 11899 16294 11911 16346
rect 11911 16294 11925 16346
rect 11949 16294 11963 16346
rect 11963 16294 11975 16346
rect 11975 16294 12005 16346
rect 12029 16294 12039 16346
rect 12039 16294 12085 16346
rect 11789 16292 11845 16294
rect 11869 16292 11925 16294
rect 11949 16292 12005 16294
rect 12029 16292 12085 16294
rect 11794 15680 11850 15736
rect 12346 18128 12402 18184
rect 11789 15258 11845 15260
rect 11869 15258 11925 15260
rect 11949 15258 12005 15260
rect 12029 15258 12085 15260
rect 11789 15206 11835 15258
rect 11835 15206 11845 15258
rect 11869 15206 11899 15258
rect 11899 15206 11911 15258
rect 11911 15206 11925 15258
rect 11949 15206 11963 15258
rect 11963 15206 11975 15258
rect 11975 15206 12005 15258
rect 12029 15206 12039 15258
rect 12039 15206 12085 15258
rect 11789 15204 11845 15206
rect 11869 15204 11925 15206
rect 11949 15204 12005 15206
rect 12029 15204 12085 15206
rect 11789 14170 11845 14172
rect 11869 14170 11925 14172
rect 11949 14170 12005 14172
rect 12029 14170 12085 14172
rect 11789 14118 11835 14170
rect 11835 14118 11845 14170
rect 11869 14118 11899 14170
rect 11899 14118 11911 14170
rect 11911 14118 11925 14170
rect 11949 14118 11963 14170
rect 11963 14118 11975 14170
rect 11975 14118 12005 14170
rect 12029 14118 12039 14170
rect 12039 14118 12085 14170
rect 11789 14116 11845 14118
rect 11869 14116 11925 14118
rect 11949 14116 12005 14118
rect 12029 14116 12085 14118
rect 11518 13252 11574 13288
rect 11518 13232 11520 13252
rect 11520 13232 11572 13252
rect 11572 13232 11574 13252
rect 11886 13776 11942 13832
rect 12714 19488 12770 19544
rect 12898 19216 12954 19272
rect 12806 16632 12862 16688
rect 12622 14728 12678 14784
rect 12070 13504 12126 13560
rect 11886 13232 11942 13288
rect 12070 13232 12126 13288
rect 11789 13082 11845 13084
rect 11869 13082 11925 13084
rect 11949 13082 12005 13084
rect 12029 13082 12085 13084
rect 11789 13030 11835 13082
rect 11835 13030 11845 13082
rect 11869 13030 11899 13082
rect 11899 13030 11911 13082
rect 11911 13030 11925 13082
rect 11949 13030 11963 13082
rect 11963 13030 11975 13082
rect 11975 13030 12005 13082
rect 12029 13030 12039 13082
rect 12039 13030 12085 13082
rect 11789 13028 11845 13030
rect 11869 13028 11925 13030
rect 11949 13028 12005 13030
rect 12029 13028 12085 13030
rect 11978 12724 11980 12744
rect 11980 12724 12032 12744
rect 12032 12724 12034 12744
rect 11978 12688 12034 12724
rect 11978 12436 12034 12472
rect 11978 12416 11980 12436
rect 11980 12416 12032 12436
rect 12032 12416 12034 12436
rect 11789 11994 11845 11996
rect 11869 11994 11925 11996
rect 11949 11994 12005 11996
rect 12029 11994 12085 11996
rect 11789 11942 11835 11994
rect 11835 11942 11845 11994
rect 11869 11942 11899 11994
rect 11899 11942 11911 11994
rect 11911 11942 11925 11994
rect 11949 11942 11963 11994
rect 11963 11942 11975 11994
rect 11975 11942 12005 11994
rect 12029 11942 12039 11994
rect 12039 11942 12085 11994
rect 11789 11940 11845 11942
rect 11869 11940 11925 11942
rect 11949 11940 12005 11942
rect 12029 11940 12085 11942
rect 11426 11600 11482 11656
rect 11610 11636 11612 11656
rect 11612 11636 11664 11656
rect 11664 11636 11666 11656
rect 11610 11600 11666 11636
rect 11518 10956 11520 10976
rect 11520 10956 11572 10976
rect 11572 10956 11574 10976
rect 11518 10920 11574 10956
rect 12070 11348 12126 11384
rect 12070 11328 12072 11348
rect 12072 11328 12124 11348
rect 12124 11328 12126 11348
rect 12990 15000 13046 15056
rect 12622 12552 12678 12608
rect 13358 20304 13414 20360
rect 13818 20476 13820 20496
rect 13820 20476 13872 20496
rect 13872 20476 13874 20496
rect 13818 20440 13874 20476
rect 13266 14592 13322 14648
rect 11789 10906 11845 10908
rect 11869 10906 11925 10908
rect 11949 10906 12005 10908
rect 12029 10906 12085 10908
rect 11789 10854 11835 10906
rect 11835 10854 11845 10906
rect 11869 10854 11899 10906
rect 11899 10854 11911 10906
rect 11911 10854 11925 10906
rect 11949 10854 11963 10906
rect 11963 10854 11975 10906
rect 11975 10854 12005 10906
rect 12029 10854 12039 10906
rect 12039 10854 12085 10906
rect 11789 10852 11845 10854
rect 11869 10852 11925 10854
rect 11949 10852 12005 10854
rect 12029 10852 12085 10854
rect 11334 10512 11390 10568
rect 10782 9424 10838 9480
rect 9862 8744 9918 8800
rect 7994 6010 8050 6012
rect 8074 6010 8130 6012
rect 8154 6010 8210 6012
rect 8234 6010 8290 6012
rect 7994 5958 8040 6010
rect 8040 5958 8050 6010
rect 8074 5958 8104 6010
rect 8104 5958 8116 6010
rect 8116 5958 8130 6010
rect 8154 5958 8168 6010
rect 8168 5958 8180 6010
rect 8180 5958 8210 6010
rect 8234 5958 8244 6010
rect 8244 5958 8290 6010
rect 7994 5956 8050 5958
rect 8074 5956 8130 5958
rect 8154 5956 8210 5958
rect 8234 5956 8290 5958
rect 7194 3848 7250 3904
rect 7994 4922 8050 4924
rect 8074 4922 8130 4924
rect 8154 4922 8210 4924
rect 8234 4922 8290 4924
rect 7994 4870 8040 4922
rect 8040 4870 8050 4922
rect 8074 4870 8104 4922
rect 8104 4870 8116 4922
rect 8116 4870 8130 4922
rect 8154 4870 8168 4922
rect 8168 4870 8180 4922
rect 8180 4870 8210 4922
rect 8234 4870 8244 4922
rect 8244 4870 8290 4922
rect 7994 4868 8050 4870
rect 8074 4868 8130 4870
rect 8154 4868 8210 4870
rect 8234 4868 8290 4870
rect 8758 4936 8814 4992
rect 9126 6024 9182 6080
rect 8942 5516 8944 5536
rect 8944 5516 8996 5536
rect 8996 5516 8998 5536
rect 8942 5480 8998 5516
rect 7994 3834 8050 3836
rect 8074 3834 8130 3836
rect 8154 3834 8210 3836
rect 8234 3834 8290 3836
rect 7994 3782 8040 3834
rect 8040 3782 8050 3834
rect 8074 3782 8104 3834
rect 8104 3782 8116 3834
rect 8116 3782 8130 3834
rect 8154 3782 8168 3834
rect 8168 3782 8180 3834
rect 8180 3782 8210 3834
rect 8234 3782 8244 3834
rect 8244 3782 8290 3834
rect 7994 3780 8050 3782
rect 8074 3780 8130 3782
rect 8154 3780 8210 3782
rect 8234 3780 8290 3782
rect 8298 3476 8300 3496
rect 8300 3476 8352 3496
rect 8352 3476 8354 3496
rect 6550 2388 6552 2408
rect 6552 2388 6604 2408
rect 6604 2388 6606 2408
rect 6550 2352 6606 2388
rect 6274 1808 6330 1864
rect 5630 1128 5686 1184
rect 3790 40 3846 96
rect 8298 3440 8354 3476
rect 7654 3168 7710 3224
rect 7994 2746 8050 2748
rect 8074 2746 8130 2748
rect 8154 2746 8210 2748
rect 8234 2746 8290 2748
rect 7994 2694 8040 2746
rect 8040 2694 8050 2746
rect 8074 2694 8104 2746
rect 8104 2694 8116 2746
rect 8116 2694 8130 2746
rect 8154 2694 8168 2746
rect 8168 2694 8180 2746
rect 8180 2694 8210 2746
rect 8234 2694 8244 2746
rect 8244 2694 8290 2746
rect 7994 2692 8050 2694
rect 8074 2692 8130 2694
rect 8154 2692 8210 2694
rect 8234 2692 8290 2694
rect 6642 1536 6698 1592
rect 7994 1658 8050 1660
rect 8074 1658 8130 1660
rect 8154 1658 8210 1660
rect 8234 1658 8290 1660
rect 7994 1606 8040 1658
rect 8040 1606 8050 1658
rect 8074 1606 8104 1658
rect 8104 1606 8116 1658
rect 8116 1606 8130 1658
rect 8154 1606 8168 1658
rect 8168 1606 8180 1658
rect 8180 1606 8210 1658
rect 8234 1606 8244 1658
rect 8244 1606 8290 1658
rect 7994 1604 8050 1606
rect 8074 1604 8130 1606
rect 8154 1604 8210 1606
rect 8234 1604 8290 1606
rect 8666 3304 8722 3360
rect 9586 7656 9642 7712
rect 9402 7112 9458 7168
rect 9402 6840 9458 6896
rect 9402 6704 9458 6760
rect 9770 6704 9826 6760
rect 9218 4936 9274 4992
rect 9402 4664 9458 4720
rect 8666 2760 8722 2816
rect 9770 3032 9826 3088
rect 10690 8336 10746 8392
rect 10598 7812 10654 7848
rect 10598 7792 10600 7812
rect 10600 7792 10652 7812
rect 10652 7792 10654 7812
rect 10506 7520 10562 7576
rect 10506 6976 10562 7032
rect 9494 2488 9550 2544
rect 9494 2216 9550 2272
rect 9494 2080 9550 2136
rect 9402 1128 9458 1184
rect 10598 6160 10654 6216
rect 11789 9818 11845 9820
rect 11869 9818 11925 9820
rect 11949 9818 12005 9820
rect 12029 9818 12085 9820
rect 11789 9766 11835 9818
rect 11835 9766 11845 9818
rect 11869 9766 11899 9818
rect 11899 9766 11911 9818
rect 11911 9766 11925 9818
rect 11949 9766 11963 9818
rect 11963 9766 11975 9818
rect 11975 9766 12005 9818
rect 12029 9766 12039 9818
rect 12039 9766 12085 9818
rect 11789 9764 11845 9766
rect 11869 9764 11925 9766
rect 11949 9764 12005 9766
rect 12029 9764 12085 9766
rect 11886 9560 11942 9616
rect 11426 9016 11482 9072
rect 11789 8730 11845 8732
rect 11869 8730 11925 8732
rect 11949 8730 12005 8732
rect 12029 8730 12085 8732
rect 11789 8678 11835 8730
rect 11835 8678 11845 8730
rect 11869 8678 11899 8730
rect 11899 8678 11911 8730
rect 11911 8678 11925 8730
rect 11949 8678 11963 8730
rect 11963 8678 11975 8730
rect 11975 8678 12005 8730
rect 12029 8678 12039 8730
rect 12039 8678 12085 8730
rect 11789 8676 11845 8678
rect 11869 8676 11925 8678
rect 11949 8676 12005 8678
rect 12029 8676 12085 8678
rect 12254 9424 12310 9480
rect 11610 7384 11666 7440
rect 11789 7642 11845 7644
rect 11869 7642 11925 7644
rect 11949 7642 12005 7644
rect 12029 7642 12085 7644
rect 11789 7590 11835 7642
rect 11835 7590 11845 7642
rect 11869 7590 11899 7642
rect 11899 7590 11911 7642
rect 11911 7590 11925 7642
rect 11949 7590 11963 7642
rect 11963 7590 11975 7642
rect 11975 7590 12005 7642
rect 12029 7590 12039 7642
rect 12039 7590 12085 7642
rect 11789 7588 11845 7590
rect 11869 7588 11925 7590
rect 11949 7588 12005 7590
rect 12029 7588 12085 7590
rect 10874 6196 10876 6216
rect 10876 6196 10928 6216
rect 10928 6196 10930 6216
rect 10874 6160 10930 6196
rect 11150 5072 11206 5128
rect 11789 6554 11845 6556
rect 11869 6554 11925 6556
rect 11949 6554 12005 6556
rect 12029 6554 12085 6556
rect 11789 6502 11835 6554
rect 11835 6502 11845 6554
rect 11869 6502 11899 6554
rect 11899 6502 11911 6554
rect 11911 6502 11925 6554
rect 11949 6502 11963 6554
rect 11963 6502 11975 6554
rect 11975 6502 12005 6554
rect 12029 6502 12039 6554
rect 12039 6502 12085 6554
rect 11789 6500 11845 6502
rect 11869 6500 11925 6502
rect 11949 6500 12005 6502
rect 12029 6500 12085 6502
rect 13082 12416 13138 12472
rect 13174 12008 13230 12064
rect 12898 10512 12954 10568
rect 13358 12960 13414 13016
rect 13450 12008 13506 12064
rect 13634 17040 13690 17096
rect 13726 16768 13782 16824
rect 15198 21528 15254 21584
rect 17958 21528 18014 21584
rect 14002 17992 14058 18048
rect 13910 17060 13966 17096
rect 13910 17040 13912 17060
rect 13912 17040 13964 17060
rect 13964 17040 13966 17060
rect 13910 16496 13966 16552
rect 13818 16224 13874 16280
rect 15584 21242 15640 21244
rect 15664 21242 15720 21244
rect 15744 21242 15800 21244
rect 15824 21242 15880 21244
rect 15584 21190 15630 21242
rect 15630 21190 15640 21242
rect 15664 21190 15694 21242
rect 15694 21190 15706 21242
rect 15706 21190 15720 21242
rect 15744 21190 15758 21242
rect 15758 21190 15770 21242
rect 15770 21190 15800 21242
rect 15824 21190 15834 21242
rect 15834 21190 15880 21242
rect 15584 21188 15640 21190
rect 15664 21188 15720 21190
rect 15744 21188 15800 21190
rect 15824 21188 15880 21190
rect 14554 20304 14610 20360
rect 14370 18944 14426 19000
rect 21638 22208 21694 22264
rect 19246 22072 19302 22128
rect 19379 21786 19435 21788
rect 19459 21786 19515 21788
rect 19539 21786 19595 21788
rect 19619 21786 19675 21788
rect 19379 21734 19425 21786
rect 19425 21734 19435 21786
rect 19459 21734 19489 21786
rect 19489 21734 19501 21786
rect 19501 21734 19515 21786
rect 19539 21734 19553 21786
rect 19553 21734 19565 21786
rect 19565 21734 19595 21786
rect 19619 21734 19629 21786
rect 19629 21734 19675 21786
rect 19379 21732 19435 21734
rect 19459 21732 19515 21734
rect 19539 21732 19595 21734
rect 19619 21732 19675 21734
rect 18510 20984 18566 21040
rect 16118 20440 16174 20496
rect 15584 20154 15640 20156
rect 15664 20154 15720 20156
rect 15744 20154 15800 20156
rect 15824 20154 15880 20156
rect 15584 20102 15630 20154
rect 15630 20102 15640 20154
rect 15664 20102 15694 20154
rect 15694 20102 15706 20154
rect 15706 20102 15720 20154
rect 15744 20102 15758 20154
rect 15758 20102 15770 20154
rect 15770 20102 15800 20154
rect 15824 20102 15834 20154
rect 15834 20102 15880 20154
rect 15584 20100 15640 20102
rect 15664 20100 15720 20102
rect 15744 20100 15800 20102
rect 15824 20100 15880 20102
rect 14370 18672 14426 18728
rect 14278 18264 14334 18320
rect 14278 17448 14334 17504
rect 14002 14592 14058 14648
rect 13818 12960 13874 13016
rect 14370 13912 14426 13968
rect 14278 13640 14334 13696
rect 13818 12552 13874 12608
rect 13450 11600 13506 11656
rect 12622 7792 12678 7848
rect 12530 7112 12586 7168
rect 11789 5466 11845 5468
rect 11869 5466 11925 5468
rect 11949 5466 12005 5468
rect 12029 5466 12085 5468
rect 11789 5414 11835 5466
rect 11835 5414 11845 5466
rect 11869 5414 11899 5466
rect 11899 5414 11911 5466
rect 11911 5414 11925 5466
rect 11949 5414 11963 5466
rect 11963 5414 11975 5466
rect 11975 5414 12005 5466
rect 12029 5414 12039 5466
rect 12039 5414 12085 5466
rect 11789 5412 11845 5414
rect 11869 5412 11925 5414
rect 11949 5412 12005 5414
rect 12029 5412 12085 5414
rect 11789 4378 11845 4380
rect 11869 4378 11925 4380
rect 11949 4378 12005 4380
rect 12029 4378 12085 4380
rect 11789 4326 11835 4378
rect 11835 4326 11845 4378
rect 11869 4326 11899 4378
rect 11899 4326 11911 4378
rect 11911 4326 11925 4378
rect 11949 4326 11963 4378
rect 11963 4326 11975 4378
rect 11975 4326 12005 4378
rect 12029 4326 12039 4378
rect 12039 4326 12085 4378
rect 11789 4324 11845 4326
rect 11869 4324 11925 4326
rect 11949 4324 12005 4326
rect 12029 4324 12085 4326
rect 11150 3168 11206 3224
rect 10690 1808 10746 1864
rect 10598 1536 10654 1592
rect 11789 3290 11845 3292
rect 11869 3290 11925 3292
rect 11949 3290 12005 3292
rect 12029 3290 12085 3292
rect 11789 3238 11835 3290
rect 11835 3238 11845 3290
rect 11869 3238 11899 3290
rect 11899 3238 11911 3290
rect 11911 3238 11925 3290
rect 11949 3238 11963 3290
rect 11963 3238 11975 3290
rect 11975 3238 12005 3290
rect 12029 3238 12039 3290
rect 12039 3238 12085 3290
rect 11789 3236 11845 3238
rect 11869 3236 11925 3238
rect 11949 3236 12005 3238
rect 12029 3236 12085 3238
rect 12162 3032 12218 3088
rect 11242 1980 11244 2000
rect 11244 1980 11296 2000
rect 11296 1980 11298 2000
rect 11242 1944 11298 1980
rect 11334 1400 11390 1456
rect 11789 2202 11845 2204
rect 11869 2202 11925 2204
rect 11949 2202 12005 2204
rect 12029 2202 12085 2204
rect 11789 2150 11835 2202
rect 11835 2150 11845 2202
rect 11869 2150 11899 2202
rect 11899 2150 11911 2202
rect 11911 2150 11925 2202
rect 11949 2150 11963 2202
rect 11963 2150 11975 2202
rect 11975 2150 12005 2202
rect 12029 2150 12039 2202
rect 12039 2150 12085 2202
rect 11789 2148 11845 2150
rect 11869 2148 11925 2150
rect 11949 2148 12005 2150
rect 12029 2148 12085 2150
rect 11978 1944 12034 2000
rect 13726 9968 13782 10024
rect 14462 12824 14518 12880
rect 14830 17740 14886 17776
rect 14830 17720 14832 17740
rect 14832 17720 14884 17740
rect 14884 17720 14886 17740
rect 14922 16632 14978 16688
rect 15106 19352 15162 19408
rect 15290 19216 15346 19272
rect 15382 19080 15438 19136
rect 15014 16224 15070 16280
rect 14738 15680 14794 15736
rect 14830 14864 14886 14920
rect 14922 14592 14978 14648
rect 15584 19066 15640 19068
rect 15664 19066 15720 19068
rect 15744 19066 15800 19068
rect 15824 19066 15880 19068
rect 15584 19014 15630 19066
rect 15630 19014 15640 19066
rect 15664 19014 15694 19066
rect 15694 19014 15706 19066
rect 15706 19014 15720 19066
rect 15744 19014 15758 19066
rect 15758 19014 15770 19066
rect 15770 19014 15800 19066
rect 15824 19014 15834 19066
rect 15834 19014 15880 19066
rect 15584 19012 15640 19014
rect 15664 19012 15720 19014
rect 15744 19012 15800 19014
rect 15824 19012 15880 19014
rect 16394 19216 16450 19272
rect 15584 17978 15640 17980
rect 15664 17978 15720 17980
rect 15744 17978 15800 17980
rect 15824 17978 15880 17980
rect 15584 17926 15630 17978
rect 15630 17926 15640 17978
rect 15664 17926 15694 17978
rect 15694 17926 15706 17978
rect 15706 17926 15720 17978
rect 15744 17926 15758 17978
rect 15758 17926 15770 17978
rect 15770 17926 15800 17978
rect 15824 17926 15834 17978
rect 15834 17926 15880 17978
rect 15584 17924 15640 17926
rect 15664 17924 15720 17926
rect 15744 17924 15800 17926
rect 15824 17924 15880 17926
rect 15584 16890 15640 16892
rect 15664 16890 15720 16892
rect 15744 16890 15800 16892
rect 15824 16890 15880 16892
rect 15584 16838 15630 16890
rect 15630 16838 15640 16890
rect 15664 16838 15694 16890
rect 15694 16838 15706 16890
rect 15706 16838 15720 16890
rect 15744 16838 15758 16890
rect 15758 16838 15770 16890
rect 15770 16838 15800 16890
rect 15824 16838 15834 16890
rect 15834 16838 15880 16890
rect 15584 16836 15640 16838
rect 15664 16836 15720 16838
rect 15744 16836 15800 16838
rect 15824 16836 15880 16838
rect 15584 15802 15640 15804
rect 15664 15802 15720 15804
rect 15744 15802 15800 15804
rect 15824 15802 15880 15804
rect 15584 15750 15630 15802
rect 15630 15750 15640 15802
rect 15664 15750 15694 15802
rect 15694 15750 15706 15802
rect 15706 15750 15720 15802
rect 15744 15750 15758 15802
rect 15758 15750 15770 15802
rect 15770 15750 15800 15802
rect 15824 15750 15834 15802
rect 15834 15750 15880 15802
rect 15584 15748 15640 15750
rect 15664 15748 15720 15750
rect 15744 15748 15800 15750
rect 15824 15748 15880 15750
rect 18050 19896 18106 19952
rect 18326 19488 18382 19544
rect 16578 16904 16634 16960
rect 16210 15952 16266 16008
rect 16118 15428 16174 15464
rect 16118 15408 16120 15428
rect 16120 15408 16172 15428
rect 16172 15408 16174 15428
rect 16118 14864 16174 14920
rect 15584 14714 15640 14716
rect 15664 14714 15720 14716
rect 15744 14714 15800 14716
rect 15824 14714 15880 14716
rect 15584 14662 15630 14714
rect 15630 14662 15640 14714
rect 15664 14662 15694 14714
rect 15694 14662 15706 14714
rect 15706 14662 15720 14714
rect 15744 14662 15758 14714
rect 15758 14662 15770 14714
rect 15770 14662 15800 14714
rect 15824 14662 15834 14714
rect 15834 14662 15880 14714
rect 15584 14660 15640 14662
rect 15664 14660 15720 14662
rect 15744 14660 15800 14662
rect 15824 14660 15880 14662
rect 15584 13626 15640 13628
rect 15664 13626 15720 13628
rect 15744 13626 15800 13628
rect 15824 13626 15880 13628
rect 15584 13574 15630 13626
rect 15630 13574 15640 13626
rect 15664 13574 15694 13626
rect 15694 13574 15706 13626
rect 15706 13574 15720 13626
rect 15744 13574 15758 13626
rect 15758 13574 15770 13626
rect 15770 13574 15800 13626
rect 15824 13574 15834 13626
rect 15834 13574 15880 13626
rect 15584 13572 15640 13574
rect 15664 13572 15720 13574
rect 15744 13572 15800 13574
rect 15824 13572 15880 13574
rect 15290 12280 15346 12336
rect 13450 7928 13506 7984
rect 13726 6860 13782 6896
rect 13726 6840 13728 6860
rect 13728 6840 13780 6860
rect 13780 6840 13782 6860
rect 13542 6160 13598 6216
rect 13358 5888 13414 5944
rect 12346 1808 12402 1864
rect 11978 1536 12034 1592
rect 7994 570 8050 572
rect 8074 570 8130 572
rect 8154 570 8210 572
rect 8234 570 8290 572
rect 7994 518 8040 570
rect 8040 518 8050 570
rect 8074 518 8104 570
rect 8104 518 8116 570
rect 8116 518 8130 570
rect 8154 518 8168 570
rect 8168 518 8180 570
rect 8180 518 8210 570
rect 8234 518 8244 570
rect 8244 518 8290 570
rect 7994 516 8050 518
rect 8074 516 8130 518
rect 8154 516 8210 518
rect 8234 516 8290 518
rect 6918 312 6974 368
rect 11789 1114 11845 1116
rect 11869 1114 11925 1116
rect 11949 1114 12005 1116
rect 12029 1114 12085 1116
rect 11789 1062 11835 1114
rect 11835 1062 11845 1114
rect 11869 1062 11899 1114
rect 11899 1062 11911 1114
rect 11911 1062 11925 1114
rect 11949 1062 11963 1114
rect 11963 1062 11975 1114
rect 11975 1062 12005 1114
rect 12029 1062 12039 1114
rect 12039 1062 12085 1114
rect 11789 1060 11845 1062
rect 11869 1060 11925 1062
rect 11949 1060 12005 1062
rect 12029 1060 12085 1062
rect 6274 176 6330 232
rect 12070 876 12126 912
rect 12070 856 12072 876
rect 12072 856 12124 876
rect 12124 856 12126 876
rect 14462 7520 14518 7576
rect 14278 7112 14334 7168
rect 14646 6996 14702 7032
rect 14646 6976 14648 6996
rect 14648 6976 14700 6996
rect 14700 6976 14702 6996
rect 13726 5752 13782 5808
rect 13634 5208 13690 5264
rect 13910 4256 13966 4312
rect 13726 3984 13782 4040
rect 12162 584 12218 640
rect 15014 11872 15070 11928
rect 16578 15952 16634 16008
rect 15584 12538 15640 12540
rect 15664 12538 15720 12540
rect 15744 12538 15800 12540
rect 15824 12538 15880 12540
rect 15584 12486 15630 12538
rect 15630 12486 15640 12538
rect 15664 12486 15694 12538
rect 15694 12486 15706 12538
rect 15706 12486 15720 12538
rect 15744 12486 15758 12538
rect 15758 12486 15770 12538
rect 15770 12486 15800 12538
rect 15824 12486 15834 12538
rect 15834 12486 15880 12538
rect 15584 12484 15640 12486
rect 15664 12484 15720 12486
rect 15744 12484 15800 12486
rect 15824 12484 15880 12486
rect 15566 12164 15622 12200
rect 15566 12144 15568 12164
rect 15568 12144 15620 12164
rect 15620 12144 15622 12164
rect 15584 11450 15640 11452
rect 15664 11450 15720 11452
rect 15744 11450 15800 11452
rect 15824 11450 15880 11452
rect 15584 11398 15630 11450
rect 15630 11398 15640 11450
rect 15664 11398 15694 11450
rect 15694 11398 15706 11450
rect 15706 11398 15720 11450
rect 15744 11398 15758 11450
rect 15758 11398 15770 11450
rect 15770 11398 15800 11450
rect 15824 11398 15834 11450
rect 15834 11398 15880 11450
rect 15584 11396 15640 11398
rect 15664 11396 15720 11398
rect 15744 11396 15800 11398
rect 15824 11396 15880 11398
rect 15474 11212 15530 11248
rect 15474 11192 15476 11212
rect 15476 11192 15528 11212
rect 15528 11192 15530 11212
rect 15584 10362 15640 10364
rect 15664 10362 15720 10364
rect 15744 10362 15800 10364
rect 15824 10362 15880 10364
rect 15584 10310 15630 10362
rect 15630 10310 15640 10362
rect 15664 10310 15694 10362
rect 15694 10310 15706 10362
rect 15706 10310 15720 10362
rect 15744 10310 15758 10362
rect 15758 10310 15770 10362
rect 15770 10310 15800 10362
rect 15824 10310 15834 10362
rect 15834 10310 15880 10362
rect 15584 10308 15640 10310
rect 15664 10308 15720 10310
rect 15744 10308 15800 10310
rect 15824 10308 15880 10310
rect 15584 9274 15640 9276
rect 15664 9274 15720 9276
rect 15744 9274 15800 9276
rect 15824 9274 15880 9276
rect 15584 9222 15630 9274
rect 15630 9222 15640 9274
rect 15664 9222 15694 9274
rect 15694 9222 15706 9274
rect 15706 9222 15720 9274
rect 15744 9222 15758 9274
rect 15758 9222 15770 9274
rect 15770 9222 15800 9274
rect 15824 9222 15834 9274
rect 15834 9222 15880 9274
rect 15584 9220 15640 9222
rect 15664 9220 15720 9222
rect 15744 9220 15800 9222
rect 15824 9220 15880 9222
rect 16946 16768 17002 16824
rect 18326 18536 18382 18592
rect 17866 17196 17922 17232
rect 17866 17176 17868 17196
rect 17868 17176 17920 17196
rect 17920 17176 17922 17196
rect 17866 16768 17922 16824
rect 17866 16496 17922 16552
rect 17222 15988 17224 16008
rect 17224 15988 17276 16008
rect 17276 15988 17278 16008
rect 17222 15952 17278 15988
rect 16854 15428 16910 15464
rect 16854 15408 16856 15428
rect 16856 15408 16908 15428
rect 16908 15408 16910 15428
rect 16302 12724 16304 12744
rect 16304 12724 16356 12744
rect 16356 12724 16358 12744
rect 16302 12688 16358 12724
rect 16210 12008 16266 12064
rect 15934 8472 15990 8528
rect 15584 8186 15640 8188
rect 15664 8186 15720 8188
rect 15744 8186 15800 8188
rect 15824 8186 15880 8188
rect 15584 8134 15630 8186
rect 15630 8134 15640 8186
rect 15664 8134 15694 8186
rect 15694 8134 15706 8186
rect 15706 8134 15720 8186
rect 15744 8134 15758 8186
rect 15758 8134 15770 8186
rect 15770 8134 15800 8186
rect 15824 8134 15834 8186
rect 15834 8134 15880 8186
rect 15584 8132 15640 8134
rect 15664 8132 15720 8134
rect 15744 8132 15800 8134
rect 15824 8132 15880 8134
rect 16118 9152 16174 9208
rect 16762 13368 16818 13424
rect 16946 14048 17002 14104
rect 18142 14048 18198 14104
rect 17682 13912 17738 13968
rect 16946 13232 17002 13288
rect 17958 13232 18014 13288
rect 18694 17584 18750 17640
rect 19062 20848 19118 20904
rect 19246 21020 19248 21040
rect 19248 21020 19300 21040
rect 19300 21020 19302 21040
rect 19246 20984 19302 21020
rect 19379 20698 19435 20700
rect 19459 20698 19515 20700
rect 19539 20698 19595 20700
rect 19619 20698 19675 20700
rect 19379 20646 19425 20698
rect 19425 20646 19435 20698
rect 19459 20646 19489 20698
rect 19489 20646 19501 20698
rect 19501 20646 19515 20698
rect 19539 20646 19553 20698
rect 19553 20646 19565 20698
rect 19565 20646 19595 20698
rect 19619 20646 19629 20698
rect 19629 20646 19675 20698
rect 19379 20644 19435 20646
rect 19459 20644 19515 20646
rect 19539 20644 19595 20646
rect 19619 20644 19675 20646
rect 19379 19610 19435 19612
rect 19459 19610 19515 19612
rect 19539 19610 19595 19612
rect 19619 19610 19675 19612
rect 19379 19558 19425 19610
rect 19425 19558 19435 19610
rect 19459 19558 19489 19610
rect 19489 19558 19501 19610
rect 19501 19558 19515 19610
rect 19539 19558 19553 19610
rect 19553 19558 19565 19610
rect 19565 19558 19595 19610
rect 19619 19558 19629 19610
rect 19629 19558 19675 19610
rect 19379 19556 19435 19558
rect 19459 19556 19515 19558
rect 19539 19556 19595 19558
rect 19619 19556 19675 19558
rect 19379 18522 19435 18524
rect 19459 18522 19515 18524
rect 19539 18522 19595 18524
rect 19619 18522 19675 18524
rect 19379 18470 19425 18522
rect 19425 18470 19435 18522
rect 19459 18470 19489 18522
rect 19489 18470 19501 18522
rect 19501 18470 19515 18522
rect 19539 18470 19553 18522
rect 19553 18470 19565 18522
rect 19565 18470 19595 18522
rect 19619 18470 19629 18522
rect 19629 18470 19675 18522
rect 19379 18468 19435 18470
rect 19459 18468 19515 18470
rect 19539 18468 19595 18470
rect 19619 18468 19675 18470
rect 19379 17434 19435 17436
rect 19459 17434 19515 17436
rect 19539 17434 19595 17436
rect 19619 17434 19675 17436
rect 19379 17382 19425 17434
rect 19425 17382 19435 17434
rect 19459 17382 19489 17434
rect 19489 17382 19501 17434
rect 19501 17382 19515 17434
rect 19539 17382 19553 17434
rect 19553 17382 19565 17434
rect 19565 17382 19595 17434
rect 19619 17382 19629 17434
rect 19629 17382 19675 17434
rect 19379 17380 19435 17382
rect 19459 17380 19515 17382
rect 19539 17380 19595 17382
rect 19619 17380 19675 17382
rect 19522 16632 19578 16688
rect 20902 20712 20958 20768
rect 19890 17448 19946 17504
rect 22466 22228 22522 22264
rect 22466 22208 22468 22228
rect 22468 22208 22520 22228
rect 22520 22208 22522 22228
rect 22282 21936 22338 21992
rect 22006 21564 22008 21584
rect 22008 21564 22060 21584
rect 22060 21564 22062 21584
rect 22006 21528 22062 21564
rect 21454 19488 21510 19544
rect 20810 18808 20866 18864
rect 21086 18672 21142 18728
rect 19890 16904 19946 16960
rect 19379 16346 19435 16348
rect 19459 16346 19515 16348
rect 19539 16346 19595 16348
rect 19619 16346 19675 16348
rect 19379 16294 19425 16346
rect 19425 16294 19435 16346
rect 19459 16294 19489 16346
rect 19489 16294 19501 16346
rect 19501 16294 19515 16346
rect 19539 16294 19553 16346
rect 19553 16294 19565 16346
rect 19565 16294 19595 16346
rect 19619 16294 19629 16346
rect 19629 16294 19675 16346
rect 19379 16292 19435 16294
rect 19459 16292 19515 16294
rect 19539 16292 19595 16294
rect 19619 16292 19675 16294
rect 18878 13912 18934 13968
rect 19379 15258 19435 15260
rect 19459 15258 19515 15260
rect 19539 15258 19595 15260
rect 19619 15258 19675 15260
rect 19379 15206 19425 15258
rect 19425 15206 19435 15258
rect 19459 15206 19489 15258
rect 19489 15206 19501 15258
rect 19501 15206 19515 15258
rect 19539 15206 19553 15258
rect 19553 15206 19565 15258
rect 19565 15206 19595 15258
rect 19619 15206 19629 15258
rect 19629 15206 19675 15258
rect 19379 15204 19435 15206
rect 19459 15204 19515 15206
rect 19539 15204 19595 15206
rect 19619 15204 19675 15206
rect 19246 14456 19302 14512
rect 19522 14320 19578 14376
rect 20442 17584 20498 17640
rect 20626 17584 20682 17640
rect 20258 16904 20314 16960
rect 19379 14170 19435 14172
rect 19459 14170 19515 14172
rect 19539 14170 19595 14172
rect 19619 14170 19675 14172
rect 19379 14118 19425 14170
rect 19425 14118 19435 14170
rect 19459 14118 19489 14170
rect 19489 14118 19501 14170
rect 19501 14118 19515 14170
rect 19539 14118 19553 14170
rect 19553 14118 19565 14170
rect 19565 14118 19595 14170
rect 19619 14118 19629 14170
rect 19629 14118 19675 14170
rect 19379 14116 19435 14118
rect 19459 14116 19515 14118
rect 19539 14116 19595 14118
rect 19619 14116 19675 14118
rect 16394 9832 16450 9888
rect 16302 9016 16358 9072
rect 15934 7928 15990 7984
rect 15584 7098 15640 7100
rect 15664 7098 15720 7100
rect 15744 7098 15800 7100
rect 15824 7098 15880 7100
rect 15584 7046 15630 7098
rect 15630 7046 15640 7098
rect 15664 7046 15694 7098
rect 15694 7046 15706 7098
rect 15706 7046 15720 7098
rect 15744 7046 15758 7098
rect 15758 7046 15770 7098
rect 15770 7046 15800 7098
rect 15824 7046 15834 7098
rect 15834 7046 15880 7098
rect 15584 7044 15640 7046
rect 15664 7044 15720 7046
rect 15744 7044 15800 7046
rect 15824 7044 15880 7046
rect 15290 6296 15346 6352
rect 15584 6010 15640 6012
rect 15664 6010 15720 6012
rect 15744 6010 15800 6012
rect 15824 6010 15880 6012
rect 15584 5958 15630 6010
rect 15630 5958 15640 6010
rect 15664 5958 15694 6010
rect 15694 5958 15706 6010
rect 15706 5958 15720 6010
rect 15744 5958 15758 6010
rect 15758 5958 15770 6010
rect 15770 5958 15800 6010
rect 15824 5958 15834 6010
rect 15834 5958 15880 6010
rect 15584 5956 15640 5958
rect 15664 5956 15720 5958
rect 15744 5956 15800 5958
rect 15824 5956 15880 5958
rect 15198 5616 15254 5672
rect 14738 2760 14794 2816
rect 15014 1944 15070 2000
rect 14462 584 14518 640
rect 15584 4922 15640 4924
rect 15664 4922 15720 4924
rect 15744 4922 15800 4924
rect 15824 4922 15880 4924
rect 15584 4870 15630 4922
rect 15630 4870 15640 4922
rect 15664 4870 15694 4922
rect 15694 4870 15706 4922
rect 15706 4870 15720 4922
rect 15744 4870 15758 4922
rect 15758 4870 15770 4922
rect 15770 4870 15800 4922
rect 15824 4870 15834 4922
rect 15834 4870 15880 4922
rect 15584 4868 15640 4870
rect 15664 4868 15720 4870
rect 15744 4868 15800 4870
rect 15824 4868 15880 4870
rect 15474 4004 15530 4040
rect 15474 3984 15476 4004
rect 15476 3984 15528 4004
rect 15528 3984 15530 4004
rect 15584 3834 15640 3836
rect 15664 3834 15720 3836
rect 15744 3834 15800 3836
rect 15824 3834 15880 3836
rect 15584 3782 15630 3834
rect 15630 3782 15640 3834
rect 15664 3782 15694 3834
rect 15694 3782 15706 3834
rect 15706 3782 15720 3834
rect 15744 3782 15758 3834
rect 15758 3782 15770 3834
rect 15770 3782 15800 3834
rect 15824 3782 15834 3834
rect 15834 3782 15880 3834
rect 15584 3780 15640 3782
rect 15664 3780 15720 3782
rect 15744 3780 15800 3782
rect 15824 3780 15880 3782
rect 16762 9288 16818 9344
rect 16762 9036 16818 9072
rect 16762 9016 16764 9036
rect 16764 9016 16816 9036
rect 16816 9016 16818 9036
rect 17038 9016 17094 9072
rect 16578 8336 16634 8392
rect 16210 6704 16266 6760
rect 16394 7112 16450 7168
rect 15934 3440 15990 3496
rect 16578 7404 16634 7440
rect 16578 7384 16580 7404
rect 16580 7384 16632 7404
rect 16632 7384 16634 7404
rect 16578 6860 16634 6896
rect 16578 6840 16580 6860
rect 16580 6840 16632 6860
rect 16632 6840 16634 6860
rect 17222 9288 17278 9344
rect 16946 7520 17002 7576
rect 17038 7248 17094 7304
rect 17038 6840 17094 6896
rect 16486 5888 16542 5944
rect 17130 6704 17186 6760
rect 17498 9424 17554 9480
rect 17406 8916 17408 8936
rect 17408 8916 17460 8936
rect 17460 8916 17462 8936
rect 17406 8880 17462 8916
rect 16394 2896 16450 2952
rect 15584 2746 15640 2748
rect 15664 2746 15720 2748
rect 15744 2746 15800 2748
rect 15824 2746 15880 2748
rect 15584 2694 15630 2746
rect 15630 2694 15640 2746
rect 15664 2694 15694 2746
rect 15694 2694 15706 2746
rect 15706 2694 15720 2746
rect 15744 2694 15758 2746
rect 15758 2694 15770 2746
rect 15770 2694 15800 2746
rect 15824 2694 15834 2746
rect 15834 2694 15880 2746
rect 15584 2692 15640 2694
rect 15664 2692 15720 2694
rect 15744 2692 15800 2694
rect 15824 2692 15880 2694
rect 17222 3476 17224 3496
rect 17224 3476 17276 3496
rect 17276 3476 17278 3496
rect 15584 1658 15640 1660
rect 15664 1658 15720 1660
rect 15744 1658 15800 1660
rect 15824 1658 15880 1660
rect 15584 1606 15630 1658
rect 15630 1606 15640 1658
rect 15664 1606 15694 1658
rect 15694 1606 15706 1658
rect 15706 1606 15720 1658
rect 15744 1606 15758 1658
rect 15758 1606 15770 1658
rect 15770 1606 15800 1658
rect 15824 1606 15834 1658
rect 15834 1606 15880 1658
rect 15584 1604 15640 1606
rect 15664 1604 15720 1606
rect 15744 1604 15800 1606
rect 15824 1604 15880 1606
rect 17222 3440 17278 3476
rect 16762 2216 16818 2272
rect 16302 1536 16358 1592
rect 16210 1400 16266 1456
rect 17774 9324 17776 9344
rect 17776 9324 17828 9344
rect 17828 9324 17830 9344
rect 17774 9288 17830 9324
rect 17774 9152 17830 9208
rect 20902 16632 20958 16688
rect 21086 16652 21142 16688
rect 21086 16632 21088 16652
rect 21088 16632 21140 16652
rect 21140 16632 21142 16652
rect 21178 15000 21234 15056
rect 19379 13082 19435 13084
rect 19459 13082 19515 13084
rect 19539 13082 19595 13084
rect 19619 13082 19675 13084
rect 19379 13030 19425 13082
rect 19425 13030 19435 13082
rect 19459 13030 19489 13082
rect 19489 13030 19501 13082
rect 19501 13030 19515 13082
rect 19539 13030 19553 13082
rect 19553 13030 19565 13082
rect 19565 13030 19595 13082
rect 19619 13030 19629 13082
rect 19629 13030 19675 13082
rect 19379 13028 19435 13030
rect 19459 13028 19515 13030
rect 19539 13028 19595 13030
rect 19619 13028 19675 13030
rect 20074 13252 20130 13288
rect 20074 13232 20076 13252
rect 20076 13232 20128 13252
rect 20128 13232 20130 13252
rect 19379 11994 19435 11996
rect 19459 11994 19515 11996
rect 19539 11994 19595 11996
rect 19619 11994 19675 11996
rect 19379 11942 19425 11994
rect 19425 11942 19435 11994
rect 19459 11942 19489 11994
rect 19489 11942 19501 11994
rect 19501 11942 19515 11994
rect 19539 11942 19553 11994
rect 19553 11942 19565 11994
rect 19565 11942 19595 11994
rect 19619 11942 19629 11994
rect 19629 11942 19675 11994
rect 19379 11940 19435 11942
rect 19459 11940 19515 11942
rect 19539 11940 19595 11942
rect 19619 11940 19675 11942
rect 18878 10668 18934 10704
rect 18878 10648 18880 10668
rect 18880 10648 18932 10668
rect 18932 10648 18934 10668
rect 18234 9016 18290 9072
rect 17774 5072 17830 5128
rect 17774 4276 17830 4312
rect 17774 4256 17776 4276
rect 17776 4256 17828 4276
rect 17828 4256 17830 4276
rect 17590 3032 17646 3088
rect 17406 1536 17462 1592
rect 18418 8916 18420 8936
rect 18420 8916 18472 8936
rect 18472 8916 18474 8936
rect 18418 8880 18474 8916
rect 20442 11056 20498 11112
rect 19379 10906 19435 10908
rect 19459 10906 19515 10908
rect 19539 10906 19595 10908
rect 19619 10906 19675 10908
rect 19379 10854 19425 10906
rect 19425 10854 19435 10906
rect 19459 10854 19489 10906
rect 19489 10854 19501 10906
rect 19501 10854 19515 10906
rect 19539 10854 19553 10906
rect 19553 10854 19565 10906
rect 19565 10854 19595 10906
rect 19619 10854 19629 10906
rect 19629 10854 19675 10906
rect 19379 10852 19435 10854
rect 19459 10852 19515 10854
rect 19539 10852 19595 10854
rect 19619 10852 19675 10854
rect 19338 10668 19394 10704
rect 19338 10648 19340 10668
rect 19340 10648 19392 10668
rect 19392 10648 19394 10668
rect 23570 21936 23626 21992
rect 22742 21528 22798 21584
rect 21914 18400 21970 18456
rect 22098 17584 22154 17640
rect 22190 16496 22246 16552
rect 21730 13388 21786 13424
rect 21730 13368 21732 13388
rect 21732 13368 21784 13388
rect 21784 13368 21786 13388
rect 24490 21548 24546 21584
rect 24490 21528 24492 21548
rect 24492 21528 24544 21548
rect 24544 21528 24546 21548
rect 23174 21242 23230 21244
rect 23254 21242 23310 21244
rect 23334 21242 23390 21244
rect 23414 21242 23470 21244
rect 23174 21190 23220 21242
rect 23220 21190 23230 21242
rect 23254 21190 23284 21242
rect 23284 21190 23296 21242
rect 23296 21190 23310 21242
rect 23334 21190 23348 21242
rect 23348 21190 23360 21242
rect 23360 21190 23390 21242
rect 23414 21190 23424 21242
rect 23424 21190 23470 21242
rect 23174 21188 23230 21190
rect 23254 21188 23310 21190
rect 23334 21188 23390 21190
rect 23414 21188 23470 21190
rect 22834 21020 22836 21040
rect 22836 21020 22888 21040
rect 22888 21020 22890 21040
rect 22834 20984 22890 21020
rect 22926 20848 22982 20904
rect 22650 18264 22706 18320
rect 23662 20712 23718 20768
rect 23174 20154 23230 20156
rect 23254 20154 23310 20156
rect 23334 20154 23390 20156
rect 23414 20154 23470 20156
rect 23174 20102 23220 20154
rect 23220 20102 23230 20154
rect 23254 20102 23284 20154
rect 23284 20102 23296 20154
rect 23296 20102 23310 20154
rect 23334 20102 23348 20154
rect 23348 20102 23360 20154
rect 23360 20102 23390 20154
rect 23414 20102 23424 20154
rect 23424 20102 23470 20154
rect 23174 20100 23230 20102
rect 23254 20100 23310 20102
rect 23334 20100 23390 20102
rect 23414 20100 23470 20102
rect 23570 20032 23626 20088
rect 23174 19066 23230 19068
rect 23254 19066 23310 19068
rect 23334 19066 23390 19068
rect 23414 19066 23470 19068
rect 23174 19014 23220 19066
rect 23220 19014 23230 19066
rect 23254 19014 23284 19066
rect 23284 19014 23296 19066
rect 23296 19014 23310 19066
rect 23334 19014 23348 19066
rect 23348 19014 23360 19066
rect 23360 19014 23390 19066
rect 23414 19014 23424 19066
rect 23424 19014 23470 19066
rect 23174 19012 23230 19014
rect 23254 19012 23310 19014
rect 23334 19012 23390 19014
rect 23414 19012 23470 19014
rect 23570 18672 23626 18728
rect 23386 18128 23442 18184
rect 23174 17978 23230 17980
rect 23254 17978 23310 17980
rect 23334 17978 23390 17980
rect 23414 17978 23470 17980
rect 23174 17926 23220 17978
rect 23220 17926 23230 17978
rect 23254 17926 23284 17978
rect 23284 17926 23296 17978
rect 23296 17926 23310 17978
rect 23334 17926 23348 17978
rect 23348 17926 23360 17978
rect 23360 17926 23390 17978
rect 23414 17926 23424 17978
rect 23424 17926 23470 17978
rect 23174 17924 23230 17926
rect 23254 17924 23310 17926
rect 23334 17924 23390 17926
rect 23414 17924 23470 17926
rect 22926 17312 22982 17368
rect 23110 17176 23166 17232
rect 23754 17856 23810 17912
rect 23662 17176 23718 17232
rect 23018 16904 23074 16960
rect 23174 16890 23230 16892
rect 23254 16890 23310 16892
rect 23334 16890 23390 16892
rect 23414 16890 23470 16892
rect 23174 16838 23220 16890
rect 23220 16838 23230 16890
rect 23254 16838 23284 16890
rect 23284 16838 23296 16890
rect 23296 16838 23310 16890
rect 23334 16838 23348 16890
rect 23348 16838 23360 16890
rect 23360 16838 23390 16890
rect 23414 16838 23424 16890
rect 23424 16838 23470 16890
rect 23174 16836 23230 16838
rect 23254 16836 23310 16838
rect 23334 16836 23390 16838
rect 23414 16836 23470 16838
rect 23938 18536 23994 18592
rect 24030 17992 24086 18048
rect 24674 19488 24730 19544
rect 25134 21120 25190 21176
rect 24306 17856 24362 17912
rect 24214 17448 24270 17504
rect 23846 16496 23902 16552
rect 23174 15802 23230 15804
rect 23254 15802 23310 15804
rect 23334 15802 23390 15804
rect 23414 15802 23470 15804
rect 23174 15750 23220 15802
rect 23220 15750 23230 15802
rect 23254 15750 23284 15802
rect 23284 15750 23296 15802
rect 23296 15750 23310 15802
rect 23334 15750 23348 15802
rect 23348 15750 23360 15802
rect 23360 15750 23390 15802
rect 23414 15750 23424 15802
rect 23424 15750 23470 15802
rect 23174 15748 23230 15750
rect 23254 15748 23310 15750
rect 23334 15748 23390 15750
rect 23414 15748 23470 15750
rect 23386 15544 23442 15600
rect 23570 14728 23626 14784
rect 23174 14714 23230 14716
rect 23254 14714 23310 14716
rect 23334 14714 23390 14716
rect 23414 14714 23470 14716
rect 23174 14662 23220 14714
rect 23220 14662 23230 14714
rect 23254 14662 23284 14714
rect 23284 14662 23296 14714
rect 23296 14662 23310 14714
rect 23334 14662 23348 14714
rect 23348 14662 23360 14714
rect 23360 14662 23390 14714
rect 23414 14662 23424 14714
rect 23424 14662 23470 14714
rect 23174 14660 23230 14662
rect 23254 14660 23310 14662
rect 23334 14660 23390 14662
rect 23414 14660 23470 14662
rect 22742 13368 22798 13424
rect 22926 12860 22928 12880
rect 22928 12860 22980 12880
rect 22980 12860 22982 12880
rect 22926 12824 22982 12860
rect 23174 13626 23230 13628
rect 23254 13626 23310 13628
rect 23334 13626 23390 13628
rect 23414 13626 23470 13628
rect 23174 13574 23220 13626
rect 23220 13574 23230 13626
rect 23254 13574 23284 13626
rect 23284 13574 23296 13626
rect 23296 13574 23310 13626
rect 23334 13574 23348 13626
rect 23348 13574 23360 13626
rect 23360 13574 23390 13626
rect 23414 13574 23424 13626
rect 23424 13574 23470 13626
rect 23174 13572 23230 13574
rect 23254 13572 23310 13574
rect 23334 13572 23390 13574
rect 23414 13572 23470 13574
rect 24858 18672 24914 18728
rect 24674 17992 24730 18048
rect 26969 21786 27025 21788
rect 27049 21786 27105 21788
rect 27129 21786 27185 21788
rect 27209 21786 27265 21788
rect 26969 21734 27015 21786
rect 27015 21734 27025 21786
rect 27049 21734 27079 21786
rect 27079 21734 27091 21786
rect 27091 21734 27105 21786
rect 27129 21734 27143 21786
rect 27143 21734 27155 21786
rect 27155 21734 27185 21786
rect 27209 21734 27219 21786
rect 27219 21734 27265 21786
rect 26969 21732 27025 21734
rect 27049 21732 27105 21734
rect 27129 21732 27185 21734
rect 27209 21732 27265 21734
rect 25318 18536 25374 18592
rect 24490 16496 24546 16552
rect 24766 16632 24822 16688
rect 24766 16088 24822 16144
rect 24490 15136 24546 15192
rect 24950 15020 25006 15056
rect 24950 15000 24952 15020
rect 24952 15000 25004 15020
rect 25004 15000 25006 15020
rect 24398 13812 24400 13832
rect 24400 13812 24452 13832
rect 24452 13812 24454 13832
rect 24398 13776 24454 13812
rect 19379 9818 19435 9820
rect 19459 9818 19515 9820
rect 19539 9818 19595 9820
rect 19619 9818 19675 9820
rect 19379 9766 19425 9818
rect 19425 9766 19435 9818
rect 19459 9766 19489 9818
rect 19489 9766 19501 9818
rect 19501 9766 19515 9818
rect 19539 9766 19553 9818
rect 19553 9766 19565 9818
rect 19565 9766 19595 9818
rect 19619 9766 19629 9818
rect 19629 9766 19675 9818
rect 19379 9764 19435 9766
rect 19459 9764 19515 9766
rect 19539 9764 19595 9766
rect 19619 9764 19675 9766
rect 18326 7384 18382 7440
rect 18694 7384 18750 7440
rect 19379 8730 19435 8732
rect 19459 8730 19515 8732
rect 19539 8730 19595 8732
rect 19619 8730 19675 8732
rect 19379 8678 19425 8730
rect 19425 8678 19435 8730
rect 19459 8678 19489 8730
rect 19489 8678 19501 8730
rect 19501 8678 19515 8730
rect 19539 8678 19553 8730
rect 19553 8678 19565 8730
rect 19565 8678 19595 8730
rect 19619 8678 19629 8730
rect 19629 8678 19675 8730
rect 19379 8676 19435 8678
rect 19459 8676 19515 8678
rect 19539 8676 19595 8678
rect 19619 8676 19675 8678
rect 19379 7642 19435 7644
rect 19459 7642 19515 7644
rect 19539 7642 19595 7644
rect 19619 7642 19675 7644
rect 19379 7590 19425 7642
rect 19425 7590 19435 7642
rect 19459 7590 19489 7642
rect 19489 7590 19501 7642
rect 19501 7590 19515 7642
rect 19539 7590 19553 7642
rect 19553 7590 19565 7642
rect 19565 7590 19595 7642
rect 19619 7590 19629 7642
rect 19629 7590 19675 7642
rect 19379 7588 19435 7590
rect 19459 7588 19515 7590
rect 19539 7588 19595 7590
rect 19619 7588 19675 7590
rect 19379 6554 19435 6556
rect 19459 6554 19515 6556
rect 19539 6554 19595 6556
rect 19619 6554 19675 6556
rect 19379 6502 19425 6554
rect 19425 6502 19435 6554
rect 19459 6502 19489 6554
rect 19489 6502 19501 6554
rect 19501 6502 19515 6554
rect 19539 6502 19553 6554
rect 19553 6502 19565 6554
rect 19565 6502 19595 6554
rect 19619 6502 19629 6554
rect 19629 6502 19675 6554
rect 19379 6500 19435 6502
rect 19459 6500 19515 6502
rect 19539 6500 19595 6502
rect 19619 6500 19675 6502
rect 18878 4936 18934 4992
rect 19379 5466 19435 5468
rect 19459 5466 19515 5468
rect 19539 5466 19595 5468
rect 19619 5466 19675 5468
rect 19379 5414 19425 5466
rect 19425 5414 19435 5466
rect 19459 5414 19489 5466
rect 19489 5414 19501 5466
rect 19501 5414 19515 5466
rect 19539 5414 19553 5466
rect 19553 5414 19565 5466
rect 19565 5414 19595 5466
rect 19619 5414 19629 5466
rect 19629 5414 19675 5466
rect 19379 5412 19435 5414
rect 19459 5412 19515 5414
rect 19539 5412 19595 5414
rect 19619 5412 19675 5414
rect 23174 12538 23230 12540
rect 23254 12538 23310 12540
rect 23334 12538 23390 12540
rect 23414 12538 23470 12540
rect 23174 12486 23220 12538
rect 23220 12486 23230 12538
rect 23254 12486 23284 12538
rect 23284 12486 23296 12538
rect 23296 12486 23310 12538
rect 23334 12486 23348 12538
rect 23348 12486 23360 12538
rect 23360 12486 23390 12538
rect 23414 12486 23424 12538
rect 23424 12486 23470 12538
rect 23174 12484 23230 12486
rect 23254 12484 23310 12486
rect 23334 12484 23390 12486
rect 23414 12484 23470 12486
rect 23754 12552 23810 12608
rect 24306 13368 24362 13424
rect 24122 11756 24178 11792
rect 24122 11736 24124 11756
rect 24124 11736 24176 11756
rect 24176 11736 24178 11756
rect 23174 11450 23230 11452
rect 23254 11450 23310 11452
rect 23334 11450 23390 11452
rect 23414 11450 23470 11452
rect 23174 11398 23220 11450
rect 23220 11398 23230 11450
rect 23254 11398 23284 11450
rect 23284 11398 23296 11450
rect 23296 11398 23310 11450
rect 23334 11398 23348 11450
rect 23348 11398 23360 11450
rect 23360 11398 23390 11450
rect 23414 11398 23424 11450
rect 23424 11398 23470 11450
rect 23174 11396 23230 11398
rect 23254 11396 23310 11398
rect 23334 11396 23390 11398
rect 23414 11396 23470 11398
rect 23174 10362 23230 10364
rect 23254 10362 23310 10364
rect 23334 10362 23390 10364
rect 23414 10362 23470 10364
rect 23174 10310 23220 10362
rect 23220 10310 23230 10362
rect 23254 10310 23284 10362
rect 23284 10310 23296 10362
rect 23296 10310 23310 10362
rect 23334 10310 23348 10362
rect 23348 10310 23360 10362
rect 23360 10310 23390 10362
rect 23414 10310 23424 10362
rect 23424 10310 23470 10362
rect 23174 10308 23230 10310
rect 23254 10308 23310 10310
rect 23334 10308 23390 10310
rect 23414 10308 23470 10310
rect 23174 9274 23230 9276
rect 23254 9274 23310 9276
rect 23334 9274 23390 9276
rect 23414 9274 23470 9276
rect 23174 9222 23220 9274
rect 23220 9222 23230 9274
rect 23254 9222 23284 9274
rect 23284 9222 23296 9274
rect 23296 9222 23310 9274
rect 23334 9222 23348 9274
rect 23348 9222 23360 9274
rect 23360 9222 23390 9274
rect 23414 9222 23424 9274
rect 23424 9222 23470 9274
rect 23174 9220 23230 9222
rect 23254 9220 23310 9222
rect 23334 9220 23390 9222
rect 23414 9220 23470 9222
rect 22926 9016 22982 9072
rect 20166 6704 20222 6760
rect 18510 3576 18566 3632
rect 15584 570 15640 572
rect 15664 570 15720 572
rect 15744 570 15800 572
rect 15824 570 15880 572
rect 15584 518 15630 570
rect 15630 518 15640 570
rect 15664 518 15694 570
rect 15694 518 15706 570
rect 15706 518 15720 570
rect 15744 518 15758 570
rect 15758 518 15770 570
rect 15770 518 15800 570
rect 15824 518 15834 570
rect 15834 518 15880 570
rect 15584 516 15640 518
rect 15664 516 15720 518
rect 15744 516 15800 518
rect 15824 516 15880 518
rect 16486 584 16542 640
rect 18234 40 18290 96
rect 19379 4378 19435 4380
rect 19459 4378 19515 4380
rect 19539 4378 19595 4380
rect 19619 4378 19675 4380
rect 19379 4326 19425 4378
rect 19425 4326 19435 4378
rect 19459 4326 19489 4378
rect 19489 4326 19501 4378
rect 19501 4326 19515 4378
rect 19539 4326 19553 4378
rect 19553 4326 19565 4378
rect 19565 4326 19595 4378
rect 19619 4326 19629 4378
rect 19629 4326 19675 4378
rect 19379 4324 19435 4326
rect 19459 4324 19515 4326
rect 19539 4324 19595 4326
rect 19619 4324 19675 4326
rect 19379 3290 19435 3292
rect 19459 3290 19515 3292
rect 19539 3290 19595 3292
rect 19619 3290 19675 3292
rect 19379 3238 19425 3290
rect 19425 3238 19435 3290
rect 19459 3238 19489 3290
rect 19489 3238 19501 3290
rect 19501 3238 19515 3290
rect 19539 3238 19553 3290
rect 19553 3238 19565 3290
rect 19565 3238 19595 3290
rect 19619 3238 19629 3290
rect 19629 3238 19675 3290
rect 19379 3236 19435 3238
rect 19459 3236 19515 3238
rect 19539 3236 19595 3238
rect 19619 3236 19675 3238
rect 19246 2216 19302 2272
rect 19379 2202 19435 2204
rect 19459 2202 19515 2204
rect 19539 2202 19595 2204
rect 19619 2202 19675 2204
rect 19379 2150 19425 2202
rect 19425 2150 19435 2202
rect 19459 2150 19489 2202
rect 19489 2150 19501 2202
rect 19501 2150 19515 2202
rect 19539 2150 19553 2202
rect 19553 2150 19565 2202
rect 19565 2150 19595 2202
rect 19619 2150 19629 2202
rect 19629 2150 19675 2202
rect 19379 2148 19435 2150
rect 19459 2148 19515 2150
rect 19539 2148 19595 2150
rect 19619 2148 19675 2150
rect 19379 1114 19435 1116
rect 19459 1114 19515 1116
rect 19539 1114 19595 1116
rect 19619 1114 19675 1116
rect 19379 1062 19425 1114
rect 19425 1062 19435 1114
rect 19459 1062 19489 1114
rect 19489 1062 19501 1114
rect 19501 1062 19515 1114
rect 19539 1062 19553 1114
rect 19553 1062 19565 1114
rect 19565 1062 19595 1114
rect 19619 1062 19629 1114
rect 19629 1062 19675 1114
rect 19379 1060 19435 1062
rect 19459 1060 19515 1062
rect 19539 1060 19595 1062
rect 19619 1060 19675 1062
rect 18878 584 18934 640
rect 18878 40 18934 96
rect 22006 7828 22008 7848
rect 22008 7828 22060 7848
rect 22060 7828 22062 7848
rect 20718 3984 20774 4040
rect 20994 3032 21050 3088
rect 22006 7792 22062 7828
rect 23174 8186 23230 8188
rect 23254 8186 23310 8188
rect 23334 8186 23390 8188
rect 23414 8186 23470 8188
rect 23174 8134 23220 8186
rect 23220 8134 23230 8186
rect 23254 8134 23284 8186
rect 23284 8134 23296 8186
rect 23296 8134 23310 8186
rect 23334 8134 23348 8186
rect 23348 8134 23360 8186
rect 23360 8134 23390 8186
rect 23414 8134 23424 8186
rect 23424 8134 23470 8186
rect 23174 8132 23230 8134
rect 23254 8132 23310 8134
rect 23334 8132 23390 8134
rect 23414 8132 23470 8134
rect 22558 7948 22614 7984
rect 22558 7928 22560 7948
rect 22560 7928 22612 7948
rect 22612 7928 22614 7948
rect 23478 7284 23480 7304
rect 23480 7284 23532 7304
rect 23532 7284 23534 7304
rect 23478 7248 23534 7284
rect 23174 7098 23230 7100
rect 23254 7098 23310 7100
rect 23334 7098 23390 7100
rect 23414 7098 23470 7100
rect 23174 7046 23220 7098
rect 23220 7046 23230 7098
rect 23254 7046 23284 7098
rect 23284 7046 23296 7098
rect 23296 7046 23310 7098
rect 23334 7046 23348 7098
rect 23348 7046 23360 7098
rect 23360 7046 23390 7098
rect 23414 7046 23424 7098
rect 23424 7046 23470 7098
rect 23174 7044 23230 7046
rect 23254 7044 23310 7046
rect 23334 7044 23390 7046
rect 23414 7044 23470 7046
rect 22190 6296 22246 6352
rect 23386 6160 23442 6216
rect 22650 5888 22706 5944
rect 22650 4664 22706 4720
rect 23174 6010 23230 6012
rect 23254 6010 23310 6012
rect 23334 6010 23390 6012
rect 23414 6010 23470 6012
rect 23174 5958 23220 6010
rect 23220 5958 23230 6010
rect 23254 5958 23284 6010
rect 23284 5958 23296 6010
rect 23296 5958 23310 6010
rect 23334 5958 23348 6010
rect 23348 5958 23360 6010
rect 23360 5958 23390 6010
rect 23414 5958 23424 6010
rect 23424 5958 23470 6010
rect 23174 5956 23230 5958
rect 23254 5956 23310 5958
rect 23334 5956 23390 5958
rect 23414 5956 23470 5958
rect 23110 5616 23166 5672
rect 23174 4922 23230 4924
rect 23254 4922 23310 4924
rect 23334 4922 23390 4924
rect 23414 4922 23470 4924
rect 23174 4870 23220 4922
rect 23220 4870 23230 4922
rect 23254 4870 23284 4922
rect 23284 4870 23296 4922
rect 23296 4870 23310 4922
rect 23334 4870 23348 4922
rect 23348 4870 23360 4922
rect 23360 4870 23390 4922
rect 23414 4870 23424 4922
rect 23424 4870 23470 4922
rect 23174 4868 23230 4870
rect 23254 4868 23310 4870
rect 23334 4868 23390 4870
rect 23414 4868 23470 4870
rect 24030 5888 24086 5944
rect 23174 3834 23230 3836
rect 23254 3834 23310 3836
rect 23334 3834 23390 3836
rect 23414 3834 23470 3836
rect 23174 3782 23220 3834
rect 23220 3782 23230 3834
rect 23254 3782 23284 3834
rect 23284 3782 23296 3834
rect 23296 3782 23310 3834
rect 23334 3782 23348 3834
rect 23348 3782 23360 3834
rect 23360 3782 23390 3834
rect 23414 3782 23424 3834
rect 23424 3782 23470 3834
rect 23174 3780 23230 3782
rect 23254 3780 23310 3782
rect 23334 3780 23390 3782
rect 23414 3780 23470 3782
rect 23570 3712 23626 3768
rect 20442 2896 20498 2952
rect 20534 2624 20590 2680
rect 20534 1672 20590 1728
rect 21822 2624 21878 2680
rect 21086 2216 21142 2272
rect 21638 2080 21694 2136
rect 20994 1536 21050 1592
rect 21546 992 21602 1048
rect 23174 2746 23230 2748
rect 23254 2746 23310 2748
rect 23334 2746 23390 2748
rect 23414 2746 23470 2748
rect 23174 2694 23220 2746
rect 23220 2694 23230 2746
rect 23254 2694 23284 2746
rect 23284 2694 23296 2746
rect 23296 2694 23310 2746
rect 23334 2694 23348 2746
rect 23348 2694 23360 2746
rect 23360 2694 23390 2746
rect 23414 2694 23424 2746
rect 23424 2694 23470 2746
rect 23174 2692 23230 2694
rect 23254 2692 23310 2694
rect 23334 2692 23390 2694
rect 23414 2692 23470 2694
rect 22650 1536 22706 1592
rect 20810 448 20866 504
rect 20718 312 20774 368
rect 22926 1672 22982 1728
rect 24490 12844 24546 12880
rect 24490 12824 24492 12844
rect 24492 12824 24544 12844
rect 24544 12824 24546 12844
rect 25410 14728 25466 14784
rect 25778 17584 25834 17640
rect 25778 14456 25834 14512
rect 24858 9424 24914 9480
rect 25134 7384 25190 7440
rect 24582 6840 24638 6896
rect 23570 1808 23626 1864
rect 23754 1808 23810 1864
rect 23754 1672 23810 1728
rect 23174 1658 23230 1660
rect 23254 1658 23310 1660
rect 23334 1658 23390 1660
rect 23414 1658 23470 1660
rect 23174 1606 23220 1658
rect 23220 1606 23230 1658
rect 23254 1606 23284 1658
rect 23284 1606 23296 1658
rect 23296 1606 23310 1658
rect 23334 1606 23348 1658
rect 23348 1606 23360 1658
rect 23360 1606 23390 1658
rect 23414 1606 23424 1658
rect 23424 1606 23470 1658
rect 23174 1604 23230 1606
rect 23254 1604 23310 1606
rect 23334 1604 23390 1606
rect 23414 1604 23470 1606
rect 23478 1128 23534 1184
rect 23662 856 23718 912
rect 24398 2388 24400 2408
rect 24400 2388 24452 2408
rect 24452 2388 24454 2408
rect 24398 2352 24454 2388
rect 26514 18400 26570 18456
rect 26238 16904 26294 16960
rect 26330 16496 26386 16552
rect 26969 20698 27025 20700
rect 27049 20698 27105 20700
rect 27129 20698 27185 20700
rect 27209 20698 27265 20700
rect 26969 20646 27015 20698
rect 27015 20646 27025 20698
rect 27049 20646 27079 20698
rect 27079 20646 27091 20698
rect 27091 20646 27105 20698
rect 27129 20646 27143 20698
rect 27143 20646 27155 20698
rect 27155 20646 27185 20698
rect 27209 20646 27219 20698
rect 27219 20646 27265 20698
rect 26969 20644 27025 20646
rect 27049 20644 27105 20646
rect 27129 20644 27185 20646
rect 27209 20644 27265 20646
rect 26969 19610 27025 19612
rect 27049 19610 27105 19612
rect 27129 19610 27185 19612
rect 27209 19610 27265 19612
rect 26969 19558 27015 19610
rect 27015 19558 27025 19610
rect 27049 19558 27079 19610
rect 27079 19558 27091 19610
rect 27091 19558 27105 19610
rect 27129 19558 27143 19610
rect 27143 19558 27155 19610
rect 27155 19558 27185 19610
rect 27209 19558 27219 19610
rect 27219 19558 27265 19610
rect 26969 19556 27025 19558
rect 27049 19556 27105 19558
rect 27129 19556 27185 19558
rect 27209 19556 27265 19558
rect 26969 18522 27025 18524
rect 27049 18522 27105 18524
rect 27129 18522 27185 18524
rect 27209 18522 27265 18524
rect 26969 18470 27015 18522
rect 27015 18470 27025 18522
rect 27049 18470 27079 18522
rect 27079 18470 27091 18522
rect 27091 18470 27105 18522
rect 27129 18470 27143 18522
rect 27143 18470 27155 18522
rect 27155 18470 27185 18522
rect 27209 18470 27219 18522
rect 27219 18470 27265 18522
rect 26969 18468 27025 18470
rect 27049 18468 27105 18470
rect 27129 18468 27185 18470
rect 27209 18468 27265 18470
rect 26698 17312 26754 17368
rect 26698 15136 26754 15192
rect 26054 13912 26110 13968
rect 26054 13368 26110 13424
rect 26969 17434 27025 17436
rect 27049 17434 27105 17436
rect 27129 17434 27185 17436
rect 27209 17434 27265 17436
rect 26969 17382 27015 17434
rect 27015 17382 27025 17434
rect 27049 17382 27079 17434
rect 27079 17382 27091 17434
rect 27091 17382 27105 17434
rect 27129 17382 27143 17434
rect 27143 17382 27155 17434
rect 27155 17382 27185 17434
rect 27209 17382 27219 17434
rect 27219 17382 27265 17434
rect 26969 17380 27025 17382
rect 27049 17380 27105 17382
rect 27129 17380 27185 17382
rect 27209 17380 27265 17382
rect 27250 17176 27306 17232
rect 27158 16904 27214 16960
rect 26969 16346 27025 16348
rect 27049 16346 27105 16348
rect 27129 16346 27185 16348
rect 27209 16346 27265 16348
rect 26969 16294 27015 16346
rect 27015 16294 27025 16346
rect 27049 16294 27079 16346
rect 27079 16294 27091 16346
rect 27091 16294 27105 16346
rect 27129 16294 27143 16346
rect 27143 16294 27155 16346
rect 27155 16294 27185 16346
rect 27209 16294 27219 16346
rect 27219 16294 27265 16346
rect 26969 16292 27025 16294
rect 27049 16292 27105 16294
rect 27129 16292 27185 16294
rect 27209 16292 27265 16294
rect 27434 15680 27490 15736
rect 26969 15258 27025 15260
rect 27049 15258 27105 15260
rect 27129 15258 27185 15260
rect 27209 15258 27265 15260
rect 26969 15206 27015 15258
rect 27015 15206 27025 15258
rect 27049 15206 27079 15258
rect 27079 15206 27091 15258
rect 27091 15206 27105 15258
rect 27129 15206 27143 15258
rect 27143 15206 27155 15258
rect 27155 15206 27185 15258
rect 27209 15206 27219 15258
rect 27219 15206 27265 15258
rect 26969 15204 27025 15206
rect 27049 15204 27105 15206
rect 27129 15204 27185 15206
rect 27209 15204 27265 15206
rect 27066 14456 27122 14512
rect 26969 14170 27025 14172
rect 27049 14170 27105 14172
rect 27129 14170 27185 14172
rect 27209 14170 27265 14172
rect 26969 14118 27015 14170
rect 27015 14118 27025 14170
rect 27049 14118 27079 14170
rect 27079 14118 27091 14170
rect 27091 14118 27105 14170
rect 27129 14118 27143 14170
rect 27143 14118 27155 14170
rect 27155 14118 27185 14170
rect 27209 14118 27219 14170
rect 27219 14118 27265 14170
rect 26969 14116 27025 14118
rect 27049 14116 27105 14118
rect 27129 14116 27185 14118
rect 27209 14116 27265 14118
rect 26969 13082 27025 13084
rect 27049 13082 27105 13084
rect 27129 13082 27185 13084
rect 27209 13082 27265 13084
rect 26969 13030 27015 13082
rect 27015 13030 27025 13082
rect 27049 13030 27079 13082
rect 27079 13030 27091 13082
rect 27091 13030 27105 13082
rect 27129 13030 27143 13082
rect 27143 13030 27155 13082
rect 27155 13030 27185 13082
rect 27209 13030 27219 13082
rect 27219 13030 27265 13082
rect 26969 13028 27025 13030
rect 27049 13028 27105 13030
rect 27129 13028 27185 13030
rect 27209 13028 27265 13030
rect 26969 11994 27025 11996
rect 27049 11994 27105 11996
rect 27129 11994 27185 11996
rect 27209 11994 27265 11996
rect 26969 11942 27015 11994
rect 27015 11942 27025 11994
rect 27049 11942 27079 11994
rect 27079 11942 27091 11994
rect 27091 11942 27105 11994
rect 27129 11942 27143 11994
rect 27143 11942 27155 11994
rect 27155 11942 27185 11994
rect 27209 11942 27219 11994
rect 27219 11942 27265 11994
rect 26969 11940 27025 11942
rect 27049 11940 27105 11942
rect 27129 11940 27185 11942
rect 27209 11940 27265 11942
rect 26054 11600 26110 11656
rect 25870 11192 25926 11248
rect 25134 4528 25190 4584
rect 24858 3168 24914 3224
rect 24674 2488 24730 2544
rect 24950 2624 25006 2680
rect 23174 570 23230 572
rect 23254 570 23310 572
rect 23334 570 23390 572
rect 23414 570 23470 572
rect 23174 518 23220 570
rect 23220 518 23230 570
rect 23254 518 23284 570
rect 23284 518 23296 570
rect 23296 518 23310 570
rect 23334 518 23348 570
rect 23348 518 23360 570
rect 23360 518 23390 570
rect 23414 518 23424 570
rect 23424 518 23470 570
rect 23174 516 23230 518
rect 23254 516 23310 518
rect 23334 516 23390 518
rect 23414 516 23470 518
rect 24858 2352 24914 2408
rect 24674 1536 24730 1592
rect 24950 992 25006 1048
rect 25502 3576 25558 3632
rect 25686 5888 25742 5944
rect 26146 9036 26202 9072
rect 26146 9016 26148 9036
rect 26148 9016 26200 9036
rect 26200 9016 26202 9036
rect 25870 5072 25926 5128
rect 25870 4664 25926 4720
rect 25778 3984 25834 4040
rect 26330 5752 26386 5808
rect 26969 10906 27025 10908
rect 27049 10906 27105 10908
rect 27129 10906 27185 10908
rect 27209 10906 27265 10908
rect 26969 10854 27015 10906
rect 27015 10854 27025 10906
rect 27049 10854 27079 10906
rect 27079 10854 27091 10906
rect 27091 10854 27105 10906
rect 27129 10854 27143 10906
rect 27143 10854 27155 10906
rect 27155 10854 27185 10906
rect 27209 10854 27219 10906
rect 27219 10854 27265 10906
rect 26969 10852 27025 10854
rect 27049 10852 27105 10854
rect 27129 10852 27185 10854
rect 27209 10852 27265 10854
rect 26969 9818 27025 9820
rect 27049 9818 27105 9820
rect 27129 9818 27185 9820
rect 27209 9818 27265 9820
rect 26969 9766 27015 9818
rect 27015 9766 27025 9818
rect 27049 9766 27079 9818
rect 27079 9766 27091 9818
rect 27091 9766 27105 9818
rect 27129 9766 27143 9818
rect 27143 9766 27155 9818
rect 27155 9766 27185 9818
rect 27209 9766 27219 9818
rect 27219 9766 27265 9818
rect 26969 9764 27025 9766
rect 27049 9764 27105 9766
rect 27129 9764 27185 9766
rect 27209 9764 27265 9766
rect 26969 8730 27025 8732
rect 27049 8730 27105 8732
rect 27129 8730 27185 8732
rect 27209 8730 27265 8732
rect 26969 8678 27015 8730
rect 27015 8678 27025 8730
rect 27049 8678 27079 8730
rect 27079 8678 27091 8730
rect 27091 8678 27105 8730
rect 27129 8678 27143 8730
rect 27143 8678 27155 8730
rect 27155 8678 27185 8730
rect 27209 8678 27219 8730
rect 27219 8678 27265 8730
rect 26969 8676 27025 8678
rect 27049 8676 27105 8678
rect 27129 8676 27185 8678
rect 27209 8676 27265 8678
rect 26969 7642 27025 7644
rect 27049 7642 27105 7644
rect 27129 7642 27185 7644
rect 27209 7642 27265 7644
rect 26969 7590 27015 7642
rect 27015 7590 27025 7642
rect 27049 7590 27079 7642
rect 27079 7590 27091 7642
rect 27091 7590 27105 7642
rect 27129 7590 27143 7642
rect 27143 7590 27155 7642
rect 27155 7590 27185 7642
rect 27209 7590 27219 7642
rect 27219 7590 27265 7642
rect 26969 7588 27025 7590
rect 27049 7588 27105 7590
rect 27129 7588 27185 7590
rect 27209 7588 27265 7590
rect 27710 16632 27766 16688
rect 28078 20032 28134 20088
rect 27802 16088 27858 16144
rect 27802 14864 27858 14920
rect 27618 13388 27674 13424
rect 27618 13368 27620 13388
rect 27620 13368 27672 13388
rect 27672 13368 27674 13388
rect 27618 11736 27674 11792
rect 28354 17856 28410 17912
rect 28354 15680 28410 15736
rect 28354 14320 28410 14376
rect 27986 12552 28042 12608
rect 26969 6554 27025 6556
rect 27049 6554 27105 6556
rect 27129 6554 27185 6556
rect 27209 6554 27265 6556
rect 26969 6502 27015 6554
rect 27015 6502 27025 6554
rect 27049 6502 27079 6554
rect 27079 6502 27091 6554
rect 27091 6502 27105 6554
rect 27129 6502 27143 6554
rect 27143 6502 27155 6554
rect 27155 6502 27185 6554
rect 27209 6502 27219 6554
rect 27219 6502 27265 6554
rect 26969 6500 27025 6502
rect 27049 6500 27105 6502
rect 27129 6500 27185 6502
rect 27209 6500 27265 6502
rect 28722 17584 28778 17640
rect 28722 16224 28778 16280
rect 28630 15544 28686 15600
rect 28538 13776 28594 13832
rect 26054 2760 26110 2816
rect 26238 2216 26294 2272
rect 26422 2080 26478 2136
rect 26969 5466 27025 5468
rect 27049 5466 27105 5468
rect 27129 5466 27185 5468
rect 27209 5466 27265 5468
rect 26969 5414 27015 5466
rect 27015 5414 27025 5466
rect 27049 5414 27079 5466
rect 27079 5414 27091 5466
rect 27091 5414 27105 5466
rect 27129 5414 27143 5466
rect 27143 5414 27155 5466
rect 27155 5414 27185 5466
rect 27209 5414 27219 5466
rect 27219 5414 27265 5466
rect 26969 5412 27025 5414
rect 27049 5412 27105 5414
rect 27129 5412 27185 5414
rect 27209 5412 27265 5414
rect 26790 2896 26846 2952
rect 26790 2624 26846 2680
rect 26790 2080 26846 2136
rect 26698 1944 26754 2000
rect 26969 4378 27025 4380
rect 27049 4378 27105 4380
rect 27129 4378 27185 4380
rect 27209 4378 27265 4380
rect 26969 4326 27015 4378
rect 27015 4326 27025 4378
rect 27049 4326 27079 4378
rect 27079 4326 27091 4378
rect 27091 4326 27105 4378
rect 27129 4326 27143 4378
rect 27143 4326 27155 4378
rect 27155 4326 27185 4378
rect 27209 4326 27219 4378
rect 27219 4326 27265 4378
rect 26969 4324 27025 4326
rect 27049 4324 27105 4326
rect 27129 4324 27185 4326
rect 27209 4324 27265 4326
rect 26969 3290 27025 3292
rect 27049 3290 27105 3292
rect 27129 3290 27185 3292
rect 27209 3290 27265 3292
rect 26969 3238 27015 3290
rect 27015 3238 27025 3290
rect 27049 3238 27079 3290
rect 27079 3238 27091 3290
rect 27091 3238 27105 3290
rect 27129 3238 27143 3290
rect 27143 3238 27155 3290
rect 27155 3238 27185 3290
rect 27209 3238 27219 3290
rect 27219 3238 27265 3290
rect 26969 3236 27025 3238
rect 27049 3236 27105 3238
rect 27129 3236 27185 3238
rect 27209 3236 27265 3238
rect 27250 2896 27306 2952
rect 26974 2760 27030 2816
rect 26969 2202 27025 2204
rect 27049 2202 27105 2204
rect 27129 2202 27185 2204
rect 27209 2202 27265 2204
rect 26969 2150 27015 2202
rect 27015 2150 27025 2202
rect 27049 2150 27079 2202
rect 27079 2150 27091 2202
rect 27091 2150 27105 2202
rect 27129 2150 27143 2202
rect 27143 2150 27155 2202
rect 27155 2150 27185 2202
rect 27209 2150 27219 2202
rect 27219 2150 27265 2202
rect 26969 2148 27025 2150
rect 27049 2148 27105 2150
rect 27129 2148 27185 2150
rect 27209 2148 27265 2150
rect 26422 1708 26424 1728
rect 26424 1708 26476 1728
rect 26476 1708 26478 1728
rect 26422 1672 26478 1708
rect 26054 1128 26110 1184
rect 26698 1400 26754 1456
rect 26969 1114 27025 1116
rect 27049 1114 27105 1116
rect 27129 1114 27185 1116
rect 27209 1114 27265 1116
rect 26969 1062 27015 1114
rect 27015 1062 27025 1114
rect 27049 1062 27079 1114
rect 27079 1062 27091 1114
rect 27091 1062 27105 1114
rect 27129 1062 27143 1114
rect 27143 1062 27155 1114
rect 27155 1062 27185 1114
rect 27209 1062 27219 1114
rect 27219 1062 27265 1114
rect 26969 1060 27025 1062
rect 27049 1060 27105 1062
rect 27129 1060 27185 1062
rect 27209 1060 27265 1062
rect 27618 3032 27674 3088
rect 29182 17992 29238 18048
rect 29182 15988 29184 16008
rect 29184 15988 29236 16008
rect 29236 15988 29238 16008
rect 29182 15952 29238 15988
rect 29182 15408 29238 15464
rect 29366 18264 29422 18320
rect 29366 17040 29422 17096
rect 29366 16224 29422 16280
rect 30764 21242 30820 21244
rect 30844 21242 30900 21244
rect 30924 21242 30980 21244
rect 31004 21242 31060 21244
rect 30764 21190 30810 21242
rect 30810 21190 30820 21242
rect 30844 21190 30874 21242
rect 30874 21190 30886 21242
rect 30886 21190 30900 21242
rect 30924 21190 30938 21242
rect 30938 21190 30950 21242
rect 30950 21190 30980 21242
rect 31004 21190 31014 21242
rect 31014 21190 31060 21242
rect 30764 21188 30820 21190
rect 30844 21188 30900 21190
rect 30924 21188 30980 21190
rect 31004 21188 31060 21190
rect 29090 13776 29146 13832
rect 28538 6296 28594 6352
rect 28354 3712 28410 3768
rect 27802 3440 27858 3496
rect 25686 176 25742 232
rect 29182 13232 29238 13288
rect 30764 20154 30820 20156
rect 30844 20154 30900 20156
rect 30924 20154 30980 20156
rect 31004 20154 31060 20156
rect 30764 20102 30810 20154
rect 30810 20102 30820 20154
rect 30844 20102 30874 20154
rect 30874 20102 30886 20154
rect 30886 20102 30900 20154
rect 30924 20102 30938 20154
rect 30938 20102 30950 20154
rect 30950 20102 30980 20154
rect 31004 20102 31014 20154
rect 31014 20102 31060 20154
rect 30764 20100 30820 20102
rect 30844 20100 30900 20102
rect 30924 20100 30980 20102
rect 31004 20100 31060 20102
rect 29918 17040 29974 17096
rect 30102 16904 30158 16960
rect 28906 7792 28962 7848
rect 30286 17720 30342 17776
rect 30764 19066 30820 19068
rect 30844 19066 30900 19068
rect 30924 19066 30980 19068
rect 31004 19066 31060 19068
rect 30764 19014 30810 19066
rect 30810 19014 30820 19066
rect 30844 19014 30874 19066
rect 30874 19014 30886 19066
rect 30886 19014 30900 19066
rect 30924 19014 30938 19066
rect 30938 19014 30950 19066
rect 30950 19014 30980 19066
rect 31004 19014 31014 19066
rect 31014 19014 31060 19066
rect 30764 19012 30820 19014
rect 30844 19012 30900 19014
rect 30924 19012 30980 19014
rect 31004 19012 31060 19014
rect 30764 17978 30820 17980
rect 30844 17978 30900 17980
rect 30924 17978 30980 17980
rect 31004 17978 31060 17980
rect 30764 17926 30810 17978
rect 30810 17926 30820 17978
rect 30844 17926 30874 17978
rect 30874 17926 30886 17978
rect 30886 17926 30900 17978
rect 30924 17926 30938 17978
rect 30938 17926 30950 17978
rect 30950 17926 30980 17978
rect 31004 17926 31014 17978
rect 31014 17926 31060 17978
rect 30764 17924 30820 17926
rect 30844 17924 30900 17926
rect 30924 17924 30980 17926
rect 31004 17924 31060 17926
rect 30764 16890 30820 16892
rect 30844 16890 30900 16892
rect 30924 16890 30980 16892
rect 31004 16890 31060 16892
rect 30764 16838 30810 16890
rect 30810 16838 30820 16890
rect 30844 16838 30874 16890
rect 30874 16838 30886 16890
rect 30886 16838 30900 16890
rect 30924 16838 30938 16890
rect 30938 16838 30950 16890
rect 30950 16838 30980 16890
rect 31004 16838 31014 16890
rect 31014 16838 31060 16890
rect 30764 16836 30820 16838
rect 30844 16836 30900 16838
rect 30924 16836 30980 16838
rect 31004 16836 31060 16838
rect 30764 15802 30820 15804
rect 30844 15802 30900 15804
rect 30924 15802 30980 15804
rect 31004 15802 31060 15804
rect 30764 15750 30810 15802
rect 30810 15750 30820 15802
rect 30844 15750 30874 15802
rect 30874 15750 30886 15802
rect 30886 15750 30900 15802
rect 30924 15750 30938 15802
rect 30938 15750 30950 15802
rect 30950 15750 30980 15802
rect 31004 15750 31014 15802
rect 31014 15750 31060 15802
rect 30764 15748 30820 15750
rect 30844 15748 30900 15750
rect 30924 15748 30980 15750
rect 31004 15748 31060 15750
rect 30764 14714 30820 14716
rect 30844 14714 30900 14716
rect 30924 14714 30980 14716
rect 31004 14714 31060 14716
rect 30764 14662 30810 14714
rect 30810 14662 30820 14714
rect 30844 14662 30874 14714
rect 30874 14662 30886 14714
rect 30886 14662 30900 14714
rect 30924 14662 30938 14714
rect 30938 14662 30950 14714
rect 30950 14662 30980 14714
rect 31004 14662 31014 14714
rect 31014 14662 31060 14714
rect 30764 14660 30820 14662
rect 30844 14660 30900 14662
rect 30924 14660 30980 14662
rect 31004 14660 31060 14662
rect 29366 6160 29422 6216
rect 29182 4120 29238 4176
rect 28998 1844 29000 1864
rect 29000 1844 29052 1864
rect 29052 1844 29054 1864
rect 28998 1808 29054 1844
rect 28630 1420 28686 1456
rect 28630 1400 28632 1420
rect 28632 1400 28684 1420
rect 28684 1400 28686 1420
rect 28722 1264 28778 1320
rect 30764 13626 30820 13628
rect 30844 13626 30900 13628
rect 30924 13626 30980 13628
rect 31004 13626 31060 13628
rect 30764 13574 30810 13626
rect 30810 13574 30820 13626
rect 30844 13574 30874 13626
rect 30874 13574 30886 13626
rect 30886 13574 30900 13626
rect 30924 13574 30938 13626
rect 30938 13574 30950 13626
rect 30950 13574 30980 13626
rect 31004 13574 31014 13626
rect 31014 13574 31060 13626
rect 30764 13572 30820 13574
rect 30844 13572 30900 13574
rect 30924 13572 30980 13574
rect 31004 13572 31060 13574
rect 30764 12538 30820 12540
rect 30844 12538 30900 12540
rect 30924 12538 30980 12540
rect 31004 12538 31060 12540
rect 30764 12486 30810 12538
rect 30810 12486 30820 12538
rect 30844 12486 30874 12538
rect 30874 12486 30886 12538
rect 30886 12486 30900 12538
rect 30924 12486 30938 12538
rect 30938 12486 30950 12538
rect 30950 12486 30980 12538
rect 31004 12486 31014 12538
rect 31014 12486 31060 12538
rect 30764 12484 30820 12486
rect 30844 12484 30900 12486
rect 30924 12484 30980 12486
rect 31004 12484 31060 12486
rect 30010 11076 30066 11112
rect 30010 11056 30012 11076
rect 30012 11056 30064 11076
rect 30064 11056 30066 11076
rect 30764 11450 30820 11452
rect 30844 11450 30900 11452
rect 30924 11450 30980 11452
rect 31004 11450 31060 11452
rect 30764 11398 30810 11450
rect 30810 11398 30820 11450
rect 30844 11398 30874 11450
rect 30874 11398 30886 11450
rect 30886 11398 30900 11450
rect 30924 11398 30938 11450
rect 30938 11398 30950 11450
rect 30950 11398 30980 11450
rect 31004 11398 31014 11450
rect 31014 11398 31060 11450
rect 30764 11396 30820 11398
rect 30844 11396 30900 11398
rect 30924 11396 30980 11398
rect 31004 11396 31060 11398
rect 29458 5616 29514 5672
rect 30764 10362 30820 10364
rect 30844 10362 30900 10364
rect 30924 10362 30980 10364
rect 31004 10362 31060 10364
rect 30764 10310 30810 10362
rect 30810 10310 30820 10362
rect 30844 10310 30874 10362
rect 30874 10310 30886 10362
rect 30886 10310 30900 10362
rect 30924 10310 30938 10362
rect 30938 10310 30950 10362
rect 30950 10310 30980 10362
rect 31004 10310 31014 10362
rect 31014 10310 31060 10362
rect 30764 10308 30820 10310
rect 30844 10308 30900 10310
rect 30924 10308 30980 10310
rect 31004 10308 31060 10310
rect 30764 9274 30820 9276
rect 30844 9274 30900 9276
rect 30924 9274 30980 9276
rect 31004 9274 31060 9276
rect 30764 9222 30810 9274
rect 30810 9222 30820 9274
rect 30844 9222 30874 9274
rect 30874 9222 30886 9274
rect 30886 9222 30900 9274
rect 30924 9222 30938 9274
rect 30938 9222 30950 9274
rect 30950 9222 30980 9274
rect 31004 9222 31014 9274
rect 31014 9222 31060 9274
rect 30764 9220 30820 9222
rect 30844 9220 30900 9222
rect 30924 9220 30980 9222
rect 31004 9220 31060 9222
rect 31390 13232 31446 13288
rect 30764 8186 30820 8188
rect 30844 8186 30900 8188
rect 30924 8186 30980 8188
rect 31004 8186 31060 8188
rect 30764 8134 30810 8186
rect 30810 8134 30820 8186
rect 30844 8134 30874 8186
rect 30874 8134 30886 8186
rect 30886 8134 30900 8186
rect 30924 8134 30938 8186
rect 30938 8134 30950 8186
rect 30950 8134 30980 8186
rect 31004 8134 31014 8186
rect 31014 8134 31060 8186
rect 30764 8132 30820 8134
rect 30844 8132 30900 8134
rect 30924 8132 30980 8134
rect 31004 8132 31060 8134
rect 30764 7098 30820 7100
rect 30844 7098 30900 7100
rect 30924 7098 30980 7100
rect 31004 7098 31060 7100
rect 30764 7046 30810 7098
rect 30810 7046 30820 7098
rect 30844 7046 30874 7098
rect 30874 7046 30886 7098
rect 30886 7046 30900 7098
rect 30924 7046 30938 7098
rect 30938 7046 30950 7098
rect 30950 7046 30980 7098
rect 31004 7046 31014 7098
rect 31014 7046 31060 7098
rect 30764 7044 30820 7046
rect 30844 7044 30900 7046
rect 30924 7044 30980 7046
rect 31004 7044 31060 7046
rect 30764 6010 30820 6012
rect 30844 6010 30900 6012
rect 30924 6010 30980 6012
rect 31004 6010 31060 6012
rect 30764 5958 30810 6010
rect 30810 5958 30820 6010
rect 30844 5958 30874 6010
rect 30874 5958 30886 6010
rect 30886 5958 30900 6010
rect 30924 5958 30938 6010
rect 30938 5958 30950 6010
rect 30950 5958 30980 6010
rect 31004 5958 31014 6010
rect 31014 5958 31060 6010
rect 30764 5956 30820 5958
rect 30844 5956 30900 5958
rect 30924 5956 30980 5958
rect 31004 5956 31060 5958
rect 30764 4922 30820 4924
rect 30844 4922 30900 4924
rect 30924 4922 30980 4924
rect 31004 4922 31060 4924
rect 30764 4870 30810 4922
rect 30810 4870 30820 4922
rect 30844 4870 30874 4922
rect 30874 4870 30886 4922
rect 30886 4870 30900 4922
rect 30924 4870 30938 4922
rect 30938 4870 30950 4922
rect 30950 4870 30980 4922
rect 31004 4870 31014 4922
rect 31014 4870 31060 4922
rect 30764 4868 30820 4870
rect 30844 4868 30900 4870
rect 30924 4868 30980 4870
rect 31004 4868 31060 4870
rect 30764 3834 30820 3836
rect 30844 3834 30900 3836
rect 30924 3834 30980 3836
rect 31004 3834 31060 3836
rect 30764 3782 30810 3834
rect 30810 3782 30820 3834
rect 30844 3782 30874 3834
rect 30874 3782 30886 3834
rect 30886 3782 30900 3834
rect 30924 3782 30938 3834
rect 30938 3782 30950 3834
rect 30950 3782 30980 3834
rect 31004 3782 31014 3834
rect 31014 3782 31060 3834
rect 30764 3780 30820 3782
rect 30844 3780 30900 3782
rect 30924 3780 30980 3782
rect 31004 3780 31060 3782
rect 30764 2746 30820 2748
rect 30844 2746 30900 2748
rect 30924 2746 30980 2748
rect 31004 2746 31060 2748
rect 30764 2694 30810 2746
rect 30810 2694 30820 2746
rect 30844 2694 30874 2746
rect 30874 2694 30886 2746
rect 30886 2694 30900 2746
rect 30924 2694 30938 2746
rect 30938 2694 30950 2746
rect 30950 2694 30980 2746
rect 31004 2694 31014 2746
rect 31014 2694 31060 2746
rect 30764 2692 30820 2694
rect 30844 2692 30900 2694
rect 30924 2692 30980 2694
rect 31004 2692 31060 2694
rect 30764 1658 30820 1660
rect 30844 1658 30900 1660
rect 30924 1658 30980 1660
rect 31004 1658 31060 1660
rect 30764 1606 30810 1658
rect 30810 1606 30820 1658
rect 30844 1606 30874 1658
rect 30874 1606 30886 1658
rect 30886 1606 30900 1658
rect 30924 1606 30938 1658
rect 30938 1606 30950 1658
rect 30950 1606 30980 1658
rect 31004 1606 31014 1658
rect 31014 1606 31060 1658
rect 30764 1604 30820 1606
rect 30844 1604 30900 1606
rect 30924 1604 30980 1606
rect 31004 1604 31060 1606
rect 30470 1400 30526 1456
rect 29274 720 29330 776
rect 30764 570 30820 572
rect 30844 570 30900 572
rect 30924 570 30980 572
rect 31004 570 31060 572
rect 30764 518 30810 570
rect 30810 518 30820 570
rect 30844 518 30874 570
rect 30874 518 30886 570
rect 30886 518 30900 570
rect 30924 518 30938 570
rect 30938 518 30950 570
rect 30950 518 30980 570
rect 31004 518 31014 570
rect 31014 518 31060 570
rect 30764 516 30820 518
rect 30844 516 30900 518
rect 30924 516 30980 518
rect 31004 516 31060 518
rect 29366 312 29422 368
rect 28078 40 28134 96
<< metal3 >>
rect 8845 22268 8911 22269
rect 9673 22268 9739 22269
rect 8845 22264 8892 22268
rect 8956 22266 8962 22268
rect 9622 22266 9628 22268
rect 8845 22208 8850 22264
rect 8845 22204 8892 22208
rect 8956 22206 9002 22266
rect 9582 22206 9628 22266
rect 9692 22264 9739 22268
rect 9734 22208 9739 22264
rect 8956 22204 8962 22206
rect 9622 22204 9628 22206
rect 9692 22204 9739 22208
rect 8845 22203 8911 22204
rect 9673 22203 9739 22204
rect 21633 22266 21699 22269
rect 22461 22266 22527 22269
rect 21633 22264 22527 22266
rect 21633 22208 21638 22264
rect 21694 22208 22466 22264
rect 22522 22208 22527 22264
rect 21633 22206 22527 22208
rect 21633 22203 21699 22206
rect 22461 22203 22527 22206
rect 6862 22068 6868 22132
rect 6932 22130 6938 22132
rect 7189 22130 7255 22133
rect 6932 22128 7255 22130
rect 6932 22072 7194 22128
rect 7250 22072 7255 22128
rect 6932 22070 7255 22072
rect 6932 22068 6938 22070
rect 7189 22067 7255 22070
rect 19241 22130 19307 22133
rect 25446 22130 25452 22132
rect 19241 22128 25452 22130
rect 19241 22072 19246 22128
rect 19302 22072 25452 22128
rect 19241 22070 25452 22072
rect 19241 22067 19307 22070
rect 25446 22068 25452 22070
rect 25516 22068 25522 22132
rect 10317 21994 10383 21997
rect 12433 21996 12499 21997
rect 12382 21994 12388 21996
rect 2730 21992 10383 21994
rect 2730 21936 10322 21992
rect 10378 21936 10383 21992
rect 2730 21934 10383 21936
rect 12346 21934 12388 21994
rect 12452 21994 12499 21996
rect 12452 21992 12544 21994
rect 12494 21936 12544 21992
rect 1669 21586 1735 21589
rect 2730 21586 2790 21934
rect 10317 21931 10383 21934
rect 12382 21932 12388 21934
rect 12452 21934 12544 21936
rect 12452 21932 12499 21934
rect 21950 21932 21956 21996
rect 22020 21994 22026 21996
rect 22277 21994 22343 21997
rect 23565 21996 23631 21997
rect 23565 21994 23612 21996
rect 22020 21992 22343 21994
rect 22020 21936 22282 21992
rect 22338 21936 22343 21992
rect 22020 21934 22343 21936
rect 23520 21992 23612 21994
rect 23520 21936 23570 21992
rect 23520 21934 23612 21936
rect 22020 21932 22026 21934
rect 12433 21931 12499 21932
rect 22277 21931 22343 21934
rect 23565 21932 23612 21934
rect 23676 21932 23682 21996
rect 23565 21931 23631 21932
rect 4189 21792 4505 21793
rect 4189 21728 4195 21792
rect 4259 21728 4275 21792
rect 4339 21728 4355 21792
rect 4419 21728 4435 21792
rect 4499 21728 4505 21792
rect 4189 21727 4505 21728
rect 11779 21792 12095 21793
rect 11779 21728 11785 21792
rect 11849 21728 11865 21792
rect 11929 21728 11945 21792
rect 12009 21728 12025 21792
rect 12089 21728 12095 21792
rect 11779 21727 12095 21728
rect 19369 21792 19685 21793
rect 19369 21728 19375 21792
rect 19439 21728 19455 21792
rect 19519 21728 19535 21792
rect 19599 21728 19615 21792
rect 19679 21728 19685 21792
rect 19369 21727 19685 21728
rect 26959 21792 27275 21793
rect 26959 21728 26965 21792
rect 27029 21728 27045 21792
rect 27109 21728 27125 21792
rect 27189 21728 27205 21792
rect 27269 21728 27275 21792
rect 26959 21727 27275 21728
rect 5809 21722 5875 21725
rect 8845 21722 8911 21725
rect 5809 21720 8911 21722
rect 5809 21664 5814 21720
rect 5870 21664 8850 21720
rect 8906 21664 8911 21720
rect 5809 21662 8911 21664
rect 5809 21659 5875 21662
rect 8845 21659 8911 21662
rect 1669 21584 2790 21586
rect 1669 21528 1674 21584
rect 1730 21528 2790 21584
rect 1669 21526 2790 21528
rect 3969 21586 4035 21589
rect 11094 21586 11100 21588
rect 3969 21584 11100 21586
rect 3969 21528 3974 21584
rect 4030 21528 11100 21584
rect 3969 21526 11100 21528
rect 1669 21523 1735 21526
rect 3969 21523 4035 21526
rect 11094 21524 11100 21526
rect 11164 21524 11170 21588
rect 13118 21524 13124 21588
rect 13188 21586 13194 21588
rect 15193 21586 15259 21589
rect 13188 21584 15259 21586
rect 13188 21528 15198 21584
rect 15254 21528 15259 21584
rect 13188 21526 15259 21528
rect 13188 21524 13194 21526
rect 15193 21523 15259 21526
rect 16982 21524 16988 21588
rect 17052 21586 17058 21588
rect 17953 21586 18019 21589
rect 17052 21584 18019 21586
rect 17052 21528 17958 21584
rect 18014 21528 18019 21584
rect 17052 21526 18019 21528
rect 17052 21524 17058 21526
rect 17953 21523 18019 21526
rect 22001 21586 22067 21589
rect 22737 21586 22803 21589
rect 24485 21586 24551 21589
rect 22001 21584 24551 21586
rect 22001 21528 22006 21584
rect 22062 21528 22742 21584
rect 22798 21528 24490 21584
rect 24546 21528 24551 21584
rect 22001 21526 24551 21528
rect 22001 21523 22067 21526
rect 22737 21523 22803 21526
rect 24485 21523 24551 21526
rect 6821 21450 6887 21453
rect 11053 21450 11119 21453
rect 24894 21450 24900 21452
rect 6821 21448 11119 21450
rect 6821 21392 6826 21448
rect 6882 21392 11058 21448
rect 11114 21392 11119 21448
rect 6821 21390 11119 21392
rect 6821 21387 6887 21390
rect 11053 21387 11119 21390
rect 22694 21390 24900 21450
rect 8569 21314 8635 21317
rect 10869 21314 10935 21317
rect 12709 21314 12775 21317
rect 22694 21314 22754 21390
rect 24894 21388 24900 21390
rect 24964 21388 24970 21452
rect 8569 21312 12775 21314
rect 8569 21256 8574 21312
rect 8630 21256 10874 21312
rect 10930 21256 12714 21312
rect 12770 21256 12775 21312
rect 8569 21254 12775 21256
rect 8569 21251 8635 21254
rect 10869 21251 10935 21254
rect 12709 21251 12775 21254
rect 22050 21254 22754 21314
rect 7984 21248 8300 21249
rect 7984 21184 7990 21248
rect 8054 21184 8070 21248
rect 8134 21184 8150 21248
rect 8214 21184 8230 21248
rect 8294 21184 8300 21248
rect 7984 21183 8300 21184
rect 15574 21248 15890 21249
rect 15574 21184 15580 21248
rect 15644 21184 15660 21248
rect 15724 21184 15740 21248
rect 15804 21184 15820 21248
rect 15884 21184 15890 21248
rect 15574 21183 15890 21184
rect 6177 21178 6243 21181
rect 7189 21178 7255 21181
rect 6177 21176 7255 21178
rect 6177 21120 6182 21176
rect 6238 21120 7194 21176
rect 7250 21120 7255 21176
rect 6177 21118 7255 21120
rect 6177 21115 6243 21118
rect 7189 21115 7255 21118
rect 8017 21042 8083 21045
rect 18505 21042 18571 21045
rect 8017 21040 18571 21042
rect 8017 20984 8022 21040
rect 8078 20984 18510 21040
rect 18566 20984 18571 21040
rect 8017 20982 18571 20984
rect 8017 20979 8083 20982
rect 18505 20979 18571 20982
rect 19241 21042 19307 21045
rect 22050 21042 22110 21254
rect 23164 21248 23480 21249
rect 23164 21184 23170 21248
rect 23234 21184 23250 21248
rect 23314 21184 23330 21248
rect 23394 21184 23410 21248
rect 23474 21184 23480 21248
rect 23164 21183 23480 21184
rect 30754 21248 31070 21249
rect 30754 21184 30760 21248
rect 30824 21184 30840 21248
rect 30904 21184 30920 21248
rect 30984 21184 31000 21248
rect 31064 21184 31070 21248
rect 30754 21183 31070 21184
rect 25129 21178 25195 21181
rect 26366 21178 26372 21180
rect 25129 21176 26372 21178
rect 25129 21120 25134 21176
rect 25190 21120 26372 21176
rect 25129 21118 26372 21120
rect 25129 21115 25195 21118
rect 26366 21116 26372 21118
rect 26436 21116 26442 21180
rect 22829 21042 22895 21045
rect 19241 21040 22110 21042
rect 19241 20984 19246 21040
rect 19302 20984 22110 21040
rect 19241 20982 22110 20984
rect 22326 21040 22895 21042
rect 22326 20984 22834 21040
rect 22890 20984 22895 21040
rect 22326 20982 22895 20984
rect 19241 20979 19307 20982
rect 5717 20906 5783 20909
rect 8845 20906 8911 20909
rect 5717 20904 8911 20906
rect 5717 20848 5722 20904
rect 5778 20848 8850 20904
rect 8906 20848 8911 20904
rect 5717 20846 8911 20848
rect 5717 20843 5783 20846
rect 8845 20843 8911 20846
rect 10777 20906 10843 20909
rect 11697 20906 11763 20909
rect 10777 20904 11763 20906
rect 10777 20848 10782 20904
rect 10838 20848 11702 20904
rect 11758 20848 11763 20904
rect 10777 20846 11763 20848
rect 10777 20843 10843 20846
rect 11697 20843 11763 20846
rect 19057 20906 19123 20909
rect 22326 20906 22386 20982
rect 22829 20979 22895 20982
rect 22921 20908 22987 20909
rect 22870 20906 22876 20908
rect 19057 20904 22386 20906
rect 19057 20848 19062 20904
rect 19118 20848 22386 20904
rect 19057 20846 22386 20848
rect 22830 20846 22876 20906
rect 22940 20904 22987 20908
rect 22982 20848 22987 20904
rect 19057 20843 19123 20846
rect 22870 20844 22876 20846
rect 22940 20844 22987 20848
rect 22921 20843 22987 20844
rect 5809 20770 5875 20773
rect 8477 20770 8543 20773
rect 5809 20768 8543 20770
rect 5809 20712 5814 20768
rect 5870 20712 8482 20768
rect 8538 20712 8543 20768
rect 5809 20710 8543 20712
rect 5809 20707 5875 20710
rect 8477 20707 8543 20710
rect 20897 20770 20963 20773
rect 22502 20770 22508 20772
rect 20897 20768 22508 20770
rect 20897 20712 20902 20768
rect 20958 20712 22508 20768
rect 20897 20710 22508 20712
rect 20897 20707 20963 20710
rect 22502 20708 22508 20710
rect 22572 20708 22578 20772
rect 23657 20770 23723 20773
rect 24158 20770 24164 20772
rect 23657 20768 24164 20770
rect 23657 20712 23662 20768
rect 23718 20712 24164 20768
rect 23657 20710 24164 20712
rect 23657 20707 23723 20710
rect 24158 20708 24164 20710
rect 24228 20708 24234 20772
rect 4189 20704 4505 20705
rect 4189 20640 4195 20704
rect 4259 20640 4275 20704
rect 4339 20640 4355 20704
rect 4419 20640 4435 20704
rect 4499 20640 4505 20704
rect 4189 20639 4505 20640
rect 11779 20704 12095 20705
rect 11779 20640 11785 20704
rect 11849 20640 11865 20704
rect 11929 20640 11945 20704
rect 12009 20640 12025 20704
rect 12089 20640 12095 20704
rect 11779 20639 12095 20640
rect 19369 20704 19685 20705
rect 19369 20640 19375 20704
rect 19439 20640 19455 20704
rect 19519 20640 19535 20704
rect 19599 20640 19615 20704
rect 19679 20640 19685 20704
rect 19369 20639 19685 20640
rect 26959 20704 27275 20705
rect 26959 20640 26965 20704
rect 27029 20640 27045 20704
rect 27109 20640 27125 20704
rect 27189 20640 27205 20704
rect 27269 20640 27275 20704
rect 26959 20639 27275 20640
rect 7281 20634 7347 20637
rect 8845 20634 8911 20637
rect 10317 20636 10383 20637
rect 10317 20634 10364 20636
rect 7281 20632 8911 20634
rect 7281 20576 7286 20632
rect 7342 20576 8850 20632
rect 8906 20576 8911 20632
rect 7281 20574 8911 20576
rect 10272 20632 10364 20634
rect 10272 20576 10322 20632
rect 10272 20574 10364 20576
rect 7281 20571 7347 20574
rect 8845 20571 8911 20574
rect 10317 20572 10364 20574
rect 10428 20572 10434 20636
rect 10317 20571 10383 20572
rect 8886 20498 8892 20500
rect 2730 20438 8892 20498
rect 1577 20362 1643 20365
rect 2730 20362 2790 20438
rect 8886 20436 8892 20438
rect 8956 20436 8962 20500
rect 10910 20436 10916 20500
rect 10980 20498 10986 20500
rect 12525 20498 12591 20501
rect 10980 20496 12591 20498
rect 10980 20440 12530 20496
rect 12586 20440 12591 20496
rect 10980 20438 12591 20440
rect 10980 20436 10986 20438
rect 12525 20435 12591 20438
rect 13670 20436 13676 20500
rect 13740 20498 13746 20500
rect 13813 20498 13879 20501
rect 16113 20500 16179 20501
rect 13740 20496 13879 20498
rect 13740 20440 13818 20496
rect 13874 20440 13879 20496
rect 13740 20438 13879 20440
rect 13740 20436 13746 20438
rect 13813 20435 13879 20438
rect 16062 20436 16068 20500
rect 16132 20498 16179 20500
rect 16132 20496 16224 20498
rect 16174 20440 16224 20496
rect 16132 20438 16224 20440
rect 16132 20436 16179 20438
rect 16113 20435 16179 20436
rect 1577 20360 2790 20362
rect 1577 20304 1582 20360
rect 1638 20304 2790 20360
rect 1577 20302 2790 20304
rect 6177 20362 6243 20365
rect 8385 20362 8451 20365
rect 6177 20360 8451 20362
rect 6177 20304 6182 20360
rect 6238 20304 8390 20360
rect 8446 20304 8451 20360
rect 6177 20302 8451 20304
rect 1577 20299 1643 20302
rect 6177 20299 6243 20302
rect 8385 20299 8451 20302
rect 10869 20362 10935 20365
rect 11973 20362 12039 20365
rect 13353 20362 13419 20365
rect 10869 20360 13419 20362
rect 10869 20304 10874 20360
rect 10930 20304 11978 20360
rect 12034 20304 13358 20360
rect 13414 20304 13419 20360
rect 10869 20302 13419 20304
rect 10869 20299 10935 20302
rect 11973 20299 12039 20302
rect 13353 20299 13419 20302
rect 14549 20364 14615 20365
rect 14549 20360 14596 20364
rect 14660 20362 14666 20364
rect 14549 20304 14554 20360
rect 14549 20300 14596 20304
rect 14660 20302 14706 20362
rect 14660 20300 14666 20302
rect 14549 20299 14615 20300
rect 7984 20160 8300 20161
rect 7984 20096 7990 20160
rect 8054 20096 8070 20160
rect 8134 20096 8150 20160
rect 8214 20096 8230 20160
rect 8294 20096 8300 20160
rect 7984 20095 8300 20096
rect 15574 20160 15890 20161
rect 15574 20096 15580 20160
rect 15644 20096 15660 20160
rect 15724 20096 15740 20160
rect 15804 20096 15820 20160
rect 15884 20096 15890 20160
rect 15574 20095 15890 20096
rect 23164 20160 23480 20161
rect 23164 20096 23170 20160
rect 23234 20096 23250 20160
rect 23314 20096 23330 20160
rect 23394 20096 23410 20160
rect 23474 20096 23480 20160
rect 23164 20095 23480 20096
rect 30754 20160 31070 20161
rect 30754 20096 30760 20160
rect 30824 20096 30840 20160
rect 30904 20096 30920 20160
rect 30984 20096 31000 20160
rect 31064 20096 31070 20160
rect 30754 20095 31070 20096
rect 5993 20090 6059 20093
rect 5812 20088 6059 20090
rect 5812 20032 5998 20088
rect 6054 20032 6059 20088
rect 5812 20030 6059 20032
rect 5812 19682 5872 20030
rect 5993 20027 6059 20030
rect 8477 20090 8543 20093
rect 9213 20090 9279 20093
rect 8477 20088 9279 20090
rect 8477 20032 8482 20088
rect 8538 20032 9218 20088
rect 9274 20032 9279 20088
rect 8477 20030 9279 20032
rect 8477 20027 8543 20030
rect 9213 20027 9279 20030
rect 23565 20090 23631 20093
rect 28073 20090 28139 20093
rect 23565 20088 28139 20090
rect 23565 20032 23570 20088
rect 23626 20032 28078 20088
rect 28134 20032 28139 20088
rect 23565 20030 28139 20032
rect 23565 20027 23631 20030
rect 28073 20027 28139 20030
rect 5993 19954 6059 19957
rect 8845 19954 8911 19957
rect 5993 19952 8911 19954
rect 5993 19896 5998 19952
rect 6054 19896 8850 19952
rect 8906 19896 8911 19952
rect 5993 19894 8911 19896
rect 5993 19891 6059 19894
rect 8845 19891 8911 19894
rect 9765 19954 9831 19957
rect 18045 19954 18111 19957
rect 9765 19952 18111 19954
rect 9765 19896 9770 19952
rect 9826 19896 18050 19952
rect 18106 19896 18111 19952
rect 9765 19894 18111 19896
rect 9765 19891 9831 19894
rect 18045 19891 18111 19894
rect 6821 19818 6887 19821
rect 9438 19818 9444 19820
rect 6821 19816 9444 19818
rect 6821 19760 6826 19816
rect 6882 19760 9444 19816
rect 6821 19758 9444 19760
rect 6821 19755 6887 19758
rect 9438 19756 9444 19758
rect 9508 19756 9514 19820
rect 11053 19682 11119 19685
rect 5812 19680 11162 19682
rect 5812 19624 11058 19680
rect 11114 19624 11162 19680
rect 5812 19622 11162 19624
rect 11053 19619 11162 19622
rect 4189 19616 4505 19617
rect 4189 19552 4195 19616
rect 4259 19552 4275 19616
rect 4339 19552 4355 19616
rect 4419 19552 4435 19616
rect 4499 19552 4505 19616
rect 4189 19551 4505 19552
rect 5165 19546 5231 19549
rect 9489 19546 9555 19549
rect 5165 19544 9555 19546
rect 5165 19488 5170 19544
rect 5226 19488 9494 19544
rect 9550 19488 9555 19544
rect 5165 19486 9555 19488
rect 5165 19483 5231 19486
rect 9489 19483 9555 19486
rect 1577 19410 1643 19413
rect 2078 19410 2084 19412
rect 1577 19408 2084 19410
rect 1577 19352 1582 19408
rect 1638 19352 2084 19408
rect 1577 19350 2084 19352
rect 1577 19347 1643 19350
rect 2078 19348 2084 19350
rect 2148 19348 2154 19412
rect 6637 19410 6703 19413
rect 6862 19410 6868 19412
rect 6637 19408 6868 19410
rect 6637 19352 6642 19408
rect 6698 19352 6868 19408
rect 6637 19350 6868 19352
rect 6637 19347 6703 19350
rect 6862 19348 6868 19350
rect 6932 19348 6938 19412
rect 11102 19410 11162 19619
rect 11779 19616 12095 19617
rect 11779 19552 11785 19616
rect 11849 19552 11865 19616
rect 11929 19552 11945 19616
rect 12009 19552 12025 19616
rect 12089 19552 12095 19616
rect 11779 19551 12095 19552
rect 19369 19616 19685 19617
rect 19369 19552 19375 19616
rect 19439 19552 19455 19616
rect 19519 19552 19535 19616
rect 19599 19552 19615 19616
rect 19679 19552 19685 19616
rect 19369 19551 19685 19552
rect 26959 19616 27275 19617
rect 26959 19552 26965 19616
rect 27029 19552 27045 19616
rect 27109 19552 27125 19616
rect 27189 19552 27205 19616
rect 27269 19552 27275 19616
rect 26959 19551 27275 19552
rect 12709 19546 12775 19549
rect 18321 19546 18387 19549
rect 12709 19544 18387 19546
rect 12709 19488 12714 19544
rect 12770 19488 18326 19544
rect 18382 19488 18387 19544
rect 12709 19486 18387 19488
rect 12709 19483 12775 19486
rect 18321 19483 18387 19486
rect 21449 19546 21515 19549
rect 24669 19546 24735 19549
rect 21449 19544 24735 19546
rect 21449 19488 21454 19544
rect 21510 19488 24674 19544
rect 24730 19488 24735 19544
rect 21449 19486 24735 19488
rect 21449 19483 21515 19486
rect 24669 19483 24735 19486
rect 15101 19410 15167 19413
rect 11102 19408 15167 19410
rect 11102 19352 15106 19408
rect 15162 19352 15167 19408
rect 11102 19350 15167 19352
rect 12942 19277 13002 19350
rect 15101 19347 15167 19350
rect 7046 19212 7052 19276
rect 7116 19274 7122 19276
rect 7557 19274 7623 19277
rect 11053 19274 11119 19277
rect 11462 19274 11468 19276
rect 7116 19272 7623 19274
rect 7116 19216 7562 19272
rect 7618 19216 7623 19272
rect 7116 19214 7623 19216
rect 7116 19212 7122 19214
rect 7557 19211 7623 19214
rect 7744 19214 8908 19274
rect 3877 19138 3943 19141
rect 7744 19138 7804 19214
rect 8848 19141 8908 19214
rect 11053 19272 11468 19274
rect 11053 19216 11058 19272
rect 11114 19216 11468 19272
rect 11053 19214 11468 19216
rect 11053 19211 11119 19214
rect 11462 19212 11468 19214
rect 11532 19212 11538 19276
rect 12893 19272 13002 19277
rect 12893 19216 12898 19272
rect 12954 19216 13002 19272
rect 12893 19214 13002 19216
rect 12893 19211 12959 19214
rect 14222 19212 14228 19276
rect 14292 19274 14298 19276
rect 15285 19274 15351 19277
rect 16389 19276 16455 19277
rect 16389 19274 16436 19276
rect 14292 19272 15351 19274
rect 14292 19216 15290 19272
rect 15346 19216 15351 19272
rect 14292 19214 15351 19216
rect 16344 19272 16436 19274
rect 16344 19216 16394 19272
rect 16344 19214 16436 19216
rect 14292 19212 14298 19214
rect 15285 19211 15351 19214
rect 16389 19212 16436 19214
rect 16500 19212 16506 19276
rect 16389 19211 16455 19212
rect 3877 19136 7804 19138
rect 3877 19080 3882 19136
rect 3938 19080 7804 19136
rect 3877 19078 7804 19080
rect 8845 19136 8911 19141
rect 15377 19140 15443 19141
rect 8845 19080 8850 19136
rect 8906 19080 8911 19136
rect 3877 19075 3943 19078
rect 8845 19075 8911 19080
rect 15326 19076 15332 19140
rect 15396 19138 15443 19140
rect 15396 19136 15488 19138
rect 15438 19080 15488 19136
rect 15396 19078 15488 19080
rect 15396 19076 15443 19078
rect 15377 19075 15443 19076
rect 7984 19072 8300 19073
rect 7984 19008 7990 19072
rect 8054 19008 8070 19072
rect 8134 19008 8150 19072
rect 8214 19008 8230 19072
rect 8294 19008 8300 19072
rect 7984 19007 8300 19008
rect 15574 19072 15890 19073
rect 15574 19008 15580 19072
rect 15644 19008 15660 19072
rect 15724 19008 15740 19072
rect 15804 19008 15820 19072
rect 15884 19008 15890 19072
rect 15574 19007 15890 19008
rect 23164 19072 23480 19073
rect 23164 19008 23170 19072
rect 23234 19008 23250 19072
rect 23314 19008 23330 19072
rect 23394 19008 23410 19072
rect 23474 19008 23480 19072
rect 23164 19007 23480 19008
rect 30754 19072 31070 19073
rect 30754 19008 30760 19072
rect 30824 19008 30840 19072
rect 30904 19008 30920 19072
rect 30984 19008 31000 19072
rect 31064 19008 31070 19072
rect 30754 19007 31070 19008
rect 4613 19002 4679 19005
rect 5022 19002 5028 19004
rect 4613 19000 5028 19002
rect 4613 18944 4618 19000
rect 4674 18944 5028 19000
rect 4613 18942 5028 18944
rect 4613 18939 4679 18942
rect 5022 18940 5028 18942
rect 5092 18940 5098 19004
rect 10317 19002 10383 19005
rect 10869 19002 10935 19005
rect 14365 19002 14431 19005
rect 10317 19000 10935 19002
rect 10317 18944 10322 19000
rect 10378 18944 10874 19000
rect 10930 18944 10935 19000
rect 10317 18942 10935 18944
rect 10317 18939 10383 18942
rect 10869 18939 10935 18942
rect 12804 19000 14431 19002
rect 12804 18944 14370 19000
rect 14426 18944 14431 19000
rect 12804 18942 14431 18944
rect 1025 18866 1091 18869
rect 4797 18866 4863 18869
rect 1025 18864 4863 18866
rect 1025 18808 1030 18864
rect 1086 18808 4802 18864
rect 4858 18808 4863 18864
rect 1025 18806 4863 18808
rect 1025 18803 1091 18806
rect 4797 18803 4863 18806
rect 7598 18804 7604 18868
rect 7668 18866 7674 18868
rect 12804 18866 12864 18942
rect 14365 18939 14431 18942
rect 20805 18866 20871 18869
rect 7668 18806 12864 18866
rect 14230 18864 20871 18866
rect 14230 18808 20810 18864
rect 20866 18808 20871 18864
rect 14230 18806 20871 18808
rect 7668 18804 7674 18806
rect 1577 18730 1643 18733
rect 3693 18730 3759 18733
rect 1577 18728 3759 18730
rect 1577 18672 1582 18728
rect 1638 18672 3698 18728
rect 3754 18672 3759 18728
rect 1577 18670 3759 18672
rect 1577 18667 1643 18670
rect 3693 18667 3759 18670
rect 7782 18668 7788 18732
rect 7852 18730 7858 18732
rect 14230 18730 14290 18806
rect 20805 18803 20871 18806
rect 7852 18670 14290 18730
rect 14365 18730 14431 18733
rect 21081 18730 21147 18733
rect 14365 18728 21147 18730
rect 14365 18672 14370 18728
rect 14426 18672 21086 18728
rect 21142 18672 21147 18728
rect 14365 18670 21147 18672
rect 7852 18668 7858 18670
rect 14365 18667 14431 18670
rect 21081 18667 21147 18670
rect 23565 18730 23631 18733
rect 24853 18730 24919 18733
rect 23565 18728 24919 18730
rect 23565 18672 23570 18728
rect 23626 18672 24858 18728
rect 24914 18672 24919 18728
rect 23565 18670 24919 18672
rect 23565 18667 23631 18670
rect 24853 18667 24919 18670
rect 5349 18594 5415 18597
rect 7373 18594 7439 18597
rect 8109 18594 8175 18597
rect 5349 18592 8175 18594
rect 5349 18536 5354 18592
rect 5410 18536 7378 18592
rect 7434 18536 8114 18592
rect 8170 18536 8175 18592
rect 5349 18534 8175 18536
rect 5349 18531 5415 18534
rect 7373 18531 7439 18534
rect 8109 18531 8175 18534
rect 8293 18594 8359 18597
rect 9673 18594 9739 18597
rect 18321 18594 18387 18597
rect 8293 18592 9739 18594
rect 8293 18536 8298 18592
rect 8354 18536 9678 18592
rect 9734 18536 9739 18592
rect 8293 18534 9739 18536
rect 8293 18531 8359 18534
rect 9673 18531 9739 18534
rect 13126 18592 18387 18594
rect 13126 18536 18326 18592
rect 18382 18536 18387 18592
rect 13126 18534 18387 18536
rect 4189 18528 4505 18529
rect 4189 18464 4195 18528
rect 4259 18464 4275 18528
rect 4339 18464 4355 18528
rect 4419 18464 4435 18528
rect 4499 18464 4505 18528
rect 4189 18463 4505 18464
rect 11779 18528 12095 18529
rect 11779 18464 11785 18528
rect 11849 18464 11865 18528
rect 11929 18464 11945 18528
rect 12009 18464 12025 18528
rect 12089 18464 12095 18528
rect 11779 18463 12095 18464
rect 5073 18458 5139 18461
rect 5390 18458 5396 18460
rect 5073 18456 5396 18458
rect 5073 18400 5078 18456
rect 5134 18400 5396 18456
rect 5073 18398 5396 18400
rect 5073 18395 5139 18398
rect 5390 18396 5396 18398
rect 5460 18396 5466 18460
rect 5625 18458 5691 18461
rect 9673 18458 9739 18461
rect 5625 18456 9739 18458
rect 5625 18400 5630 18456
rect 5686 18400 9678 18456
rect 9734 18400 9739 18456
rect 5625 18398 9739 18400
rect 5625 18395 5691 18398
rect 9673 18395 9739 18398
rect 5349 18322 5415 18325
rect 13126 18322 13186 18534
rect 18321 18531 18387 18534
rect 23933 18594 23999 18597
rect 25313 18594 25379 18597
rect 23933 18592 25379 18594
rect 23933 18536 23938 18592
rect 23994 18536 25318 18592
rect 25374 18536 25379 18592
rect 23933 18534 25379 18536
rect 23933 18531 23999 18534
rect 25313 18531 25379 18534
rect 19369 18528 19685 18529
rect 19369 18464 19375 18528
rect 19439 18464 19455 18528
rect 19519 18464 19535 18528
rect 19599 18464 19615 18528
rect 19679 18464 19685 18528
rect 19369 18463 19685 18464
rect 26959 18528 27275 18529
rect 26959 18464 26965 18528
rect 27029 18464 27045 18528
rect 27109 18464 27125 18528
rect 27189 18464 27205 18528
rect 27269 18464 27275 18528
rect 26959 18463 27275 18464
rect 21909 18458 21975 18461
rect 26509 18458 26575 18461
rect 21909 18456 26575 18458
rect 21909 18400 21914 18456
rect 21970 18400 26514 18456
rect 26570 18400 26575 18456
rect 21909 18398 26575 18400
rect 21909 18395 21975 18398
rect 26509 18395 26575 18398
rect 14273 18322 14339 18325
rect 5349 18320 13186 18322
rect 5349 18264 5354 18320
rect 5410 18264 13186 18320
rect 5349 18262 13186 18264
rect 13310 18320 14339 18322
rect 13310 18264 14278 18320
rect 14334 18264 14339 18320
rect 13310 18262 14339 18264
rect 5349 18259 5415 18262
rect 4654 18124 4660 18188
rect 4724 18186 4730 18188
rect 4981 18186 5047 18189
rect 4724 18184 5047 18186
rect 4724 18128 4986 18184
rect 5042 18128 5047 18184
rect 4724 18126 5047 18128
rect 4724 18124 4730 18126
rect 4981 18123 5047 18126
rect 6821 18186 6887 18189
rect 12341 18186 12407 18189
rect 12566 18186 12572 18188
rect 6821 18184 8954 18186
rect 6821 18128 6826 18184
rect 6882 18128 8954 18184
rect 6821 18126 8954 18128
rect 6821 18123 6887 18126
rect 4889 18052 4955 18053
rect 4838 17988 4844 18052
rect 4908 18050 4955 18052
rect 4908 18048 5000 18050
rect 4950 17992 5000 18048
rect 4908 17990 5000 17992
rect 4908 17988 4955 17990
rect 5942 17988 5948 18052
rect 6012 18050 6018 18052
rect 6545 18050 6611 18053
rect 8661 18052 8727 18053
rect 8661 18050 8708 18052
rect 6012 18048 6611 18050
rect 6012 17992 6550 18048
rect 6606 17992 6611 18048
rect 6012 17990 6611 17992
rect 8616 18048 8708 18050
rect 8616 17992 8666 18048
rect 8616 17990 8708 17992
rect 6012 17988 6018 17990
rect 4889 17987 4955 17988
rect 6545 17987 6611 17990
rect 8661 17988 8708 17990
rect 8772 17988 8778 18052
rect 8894 18050 8954 18126
rect 12341 18184 12572 18186
rect 12341 18128 12346 18184
rect 12402 18128 12572 18184
rect 12341 18126 12572 18128
rect 12341 18123 12407 18126
rect 12566 18124 12572 18126
rect 12636 18124 12642 18188
rect 13310 18050 13370 18262
rect 14273 18259 14339 18262
rect 22645 18322 22711 18325
rect 29361 18322 29427 18325
rect 22645 18320 29427 18322
rect 22645 18264 22650 18320
rect 22706 18264 29366 18320
rect 29422 18264 29427 18320
rect 22645 18262 29427 18264
rect 22645 18259 22711 18262
rect 29361 18259 29427 18262
rect 23381 18186 23447 18189
rect 24710 18186 24716 18188
rect 23381 18184 24716 18186
rect 23381 18128 23386 18184
rect 23442 18128 24716 18184
rect 23381 18126 24716 18128
rect 23381 18123 23447 18126
rect 24710 18124 24716 18126
rect 24780 18124 24786 18188
rect 8894 17990 13370 18050
rect 13997 18052 14063 18053
rect 13997 18048 14044 18052
rect 14108 18050 14114 18052
rect 24025 18050 24091 18053
rect 24669 18050 24735 18053
rect 29177 18050 29243 18053
rect 13997 17992 14002 18048
rect 13997 17988 14044 17992
rect 14108 17990 14154 18050
rect 24025 18048 24548 18050
rect 24025 17992 24030 18048
rect 24086 17992 24548 18048
rect 24025 17990 24548 17992
rect 14108 17988 14114 17990
rect 8661 17987 8727 17988
rect 13997 17987 14063 17988
rect 24025 17987 24091 17990
rect 7984 17984 8300 17985
rect 7984 17920 7990 17984
rect 8054 17920 8070 17984
rect 8134 17920 8150 17984
rect 8214 17920 8230 17984
rect 8294 17920 8300 17984
rect 7984 17919 8300 17920
rect 15574 17984 15890 17985
rect 15574 17920 15580 17984
rect 15644 17920 15660 17984
rect 15724 17920 15740 17984
rect 15804 17920 15820 17984
rect 15884 17920 15890 17984
rect 15574 17919 15890 17920
rect 23164 17984 23480 17985
rect 23164 17920 23170 17984
rect 23234 17920 23250 17984
rect 23314 17920 23330 17984
rect 23394 17920 23410 17984
rect 23474 17920 23480 17984
rect 23164 17919 23480 17920
rect 3601 17914 3667 17917
rect 7741 17914 7807 17917
rect 3601 17912 7807 17914
rect 3601 17856 3606 17912
rect 3662 17856 7746 17912
rect 7802 17856 7807 17912
rect 3601 17854 7807 17856
rect 3601 17851 3667 17854
rect 7741 17851 7807 17854
rect 23749 17914 23815 17917
rect 24301 17914 24367 17917
rect 23749 17912 24367 17914
rect 23749 17856 23754 17912
rect 23810 17856 24306 17912
rect 24362 17856 24367 17912
rect 23749 17854 24367 17856
rect 24488 17914 24548 17990
rect 24669 18048 29243 18050
rect 24669 17992 24674 18048
rect 24730 17992 29182 18048
rect 29238 17992 29243 18048
rect 24669 17990 29243 17992
rect 24669 17987 24735 17990
rect 29177 17987 29243 17990
rect 30754 17984 31070 17985
rect 30754 17920 30760 17984
rect 30824 17920 30840 17984
rect 30904 17920 30920 17984
rect 30984 17920 31000 17984
rect 31064 17920 31070 17984
rect 30754 17919 31070 17920
rect 28349 17914 28415 17917
rect 24488 17912 28415 17914
rect 24488 17856 28354 17912
rect 28410 17856 28415 17912
rect 24488 17854 28415 17856
rect 23749 17851 23815 17854
rect 24301 17851 24367 17854
rect 28349 17851 28415 17854
rect 5349 17778 5415 17781
rect 9857 17778 9923 17781
rect 5349 17776 9923 17778
rect 5349 17720 5354 17776
rect 5410 17720 9862 17776
rect 9918 17720 9923 17776
rect 5349 17718 9923 17720
rect 5349 17715 5415 17718
rect 9857 17715 9923 17718
rect 11237 17778 11303 17781
rect 14825 17778 14891 17781
rect 30281 17778 30347 17781
rect 11237 17776 30347 17778
rect 11237 17720 11242 17776
rect 11298 17720 14830 17776
rect 14886 17720 30286 17776
rect 30342 17720 30347 17776
rect 11237 17718 30347 17720
rect 11237 17715 11303 17718
rect 14825 17715 14891 17718
rect 30281 17715 30347 17718
rect 1669 17642 1735 17645
rect 7833 17642 7899 17645
rect 9397 17642 9463 17645
rect 1669 17640 6930 17642
rect 1669 17584 1674 17640
rect 1730 17584 6930 17640
rect 1669 17582 6930 17584
rect 1669 17579 1735 17582
rect 4189 17440 4505 17441
rect 4189 17376 4195 17440
rect 4259 17376 4275 17440
rect 4339 17376 4355 17440
rect 4419 17376 4435 17440
rect 4499 17376 4505 17440
rect 4189 17375 4505 17376
rect 6870 17370 6930 17582
rect 7833 17640 9463 17642
rect 7833 17584 7838 17640
rect 7894 17584 9402 17640
rect 9458 17584 9463 17640
rect 7833 17582 9463 17584
rect 7833 17579 7899 17582
rect 9397 17579 9463 17582
rect 9765 17642 9831 17645
rect 18689 17642 18755 17645
rect 20437 17642 20503 17645
rect 9765 17640 18755 17642
rect 9765 17584 9770 17640
rect 9826 17584 18694 17640
rect 18750 17584 18755 17640
rect 9765 17582 18755 17584
rect 9765 17579 9831 17582
rect 18689 17579 18755 17582
rect 19198 17640 20503 17642
rect 19198 17584 20442 17640
rect 20498 17584 20503 17640
rect 19198 17582 20503 17584
rect 7741 17506 7807 17509
rect 11053 17506 11119 17509
rect 7741 17504 11119 17506
rect 7741 17448 7746 17504
rect 7802 17448 11058 17504
rect 11114 17448 11119 17504
rect 7741 17446 11119 17448
rect 7741 17443 7807 17446
rect 11053 17443 11119 17446
rect 14273 17506 14339 17509
rect 19198 17506 19258 17582
rect 20437 17579 20503 17582
rect 20621 17642 20687 17645
rect 22093 17642 22159 17645
rect 20621 17640 22159 17642
rect 20621 17584 20626 17640
rect 20682 17584 22098 17640
rect 22154 17584 22159 17640
rect 20621 17582 22159 17584
rect 20621 17579 20687 17582
rect 22093 17579 22159 17582
rect 25773 17642 25839 17645
rect 28717 17642 28783 17645
rect 25773 17640 28783 17642
rect 25773 17584 25778 17640
rect 25834 17584 28722 17640
rect 28778 17584 28783 17640
rect 25773 17582 28783 17584
rect 25773 17579 25839 17582
rect 28717 17579 28783 17582
rect 14273 17504 19258 17506
rect 14273 17448 14278 17504
rect 14334 17448 19258 17504
rect 14273 17446 19258 17448
rect 19885 17506 19951 17509
rect 24209 17506 24275 17509
rect 19885 17504 24275 17506
rect 19885 17448 19890 17504
rect 19946 17448 24214 17504
rect 24270 17448 24275 17504
rect 19885 17446 24275 17448
rect 14273 17443 14339 17446
rect 19885 17443 19951 17446
rect 24209 17443 24275 17446
rect 11779 17440 12095 17441
rect 11779 17376 11785 17440
rect 11849 17376 11865 17440
rect 11929 17376 11945 17440
rect 12009 17376 12025 17440
rect 12089 17376 12095 17440
rect 11779 17375 12095 17376
rect 19369 17440 19685 17441
rect 19369 17376 19375 17440
rect 19439 17376 19455 17440
rect 19519 17376 19535 17440
rect 19599 17376 19615 17440
rect 19679 17376 19685 17440
rect 19369 17375 19685 17376
rect 26959 17440 27275 17441
rect 26959 17376 26965 17440
rect 27029 17376 27045 17440
rect 27109 17376 27125 17440
rect 27189 17376 27205 17440
rect 27269 17376 27275 17440
rect 26959 17375 27275 17376
rect 10358 17370 10364 17372
rect 6870 17310 10364 17370
rect 10358 17308 10364 17310
rect 10428 17308 10434 17372
rect 22921 17370 22987 17373
rect 26693 17370 26759 17373
rect 22921 17368 26759 17370
rect 22921 17312 22926 17368
rect 22982 17312 26698 17368
rect 26754 17312 26759 17368
rect 22921 17310 26759 17312
rect 22921 17307 22987 17310
rect 26693 17307 26759 17310
rect 9213 17234 9279 17237
rect 17861 17234 17927 17237
rect 23105 17234 23171 17237
rect 9213 17232 12450 17234
rect 9213 17176 9218 17232
rect 9274 17176 12450 17232
rect 9213 17174 12450 17176
rect 9213 17171 9279 17174
rect 6821 17098 6887 17101
rect 12390 17098 12450 17174
rect 17861 17232 23171 17234
rect 17861 17176 17866 17232
rect 17922 17176 23110 17232
rect 23166 17176 23171 17232
rect 17861 17174 23171 17176
rect 17861 17171 17927 17174
rect 23105 17171 23171 17174
rect 23657 17234 23723 17237
rect 27245 17234 27311 17237
rect 23657 17232 27311 17234
rect 23657 17176 23662 17232
rect 23718 17176 27250 17232
rect 27306 17176 27311 17232
rect 23657 17174 27311 17176
rect 23657 17171 23723 17174
rect 27245 17171 27311 17174
rect 13629 17098 13695 17101
rect 6821 17096 9690 17098
rect 6821 17040 6826 17096
rect 6882 17040 9690 17096
rect 6821 17038 9690 17040
rect 12390 17096 13695 17098
rect 12390 17040 13634 17096
rect 13690 17040 13695 17096
rect 12390 17038 13695 17040
rect 6821 17035 6887 17038
rect 4705 16962 4771 16965
rect 5257 16962 5323 16965
rect 4705 16960 5323 16962
rect 4705 16904 4710 16960
rect 4766 16904 5262 16960
rect 5318 16904 5323 16960
rect 4705 16902 5323 16904
rect 4705 16899 4771 16902
rect 5257 16899 5323 16902
rect 7984 16896 8300 16897
rect 7984 16832 7990 16896
rect 8054 16832 8070 16896
rect 8134 16832 8150 16896
rect 8214 16832 8230 16896
rect 8294 16832 8300 16896
rect 7984 16831 8300 16832
rect 8385 16826 8451 16829
rect 9305 16826 9371 16829
rect 8385 16824 9371 16826
rect 8385 16768 8390 16824
rect 8446 16768 9310 16824
rect 9366 16768 9371 16824
rect 8385 16766 9371 16768
rect 9630 16826 9690 17038
rect 13629 17035 13695 17038
rect 13905 17098 13971 17101
rect 29361 17098 29427 17101
rect 13905 17096 29427 17098
rect 13905 17040 13910 17096
rect 13966 17040 29366 17096
rect 29422 17040 29427 17096
rect 13905 17038 29427 17040
rect 13905 17035 13971 17038
rect 29361 17035 29427 17038
rect 29913 17098 29979 17101
rect 29913 17096 30114 17098
rect 29913 17040 29918 17096
rect 29974 17040 30114 17096
rect 29913 17038 30114 17040
rect 29913 17035 29979 17038
rect 30054 16965 30114 17038
rect 16573 16962 16639 16965
rect 19885 16962 19951 16965
rect 16573 16960 19951 16962
rect 16573 16904 16578 16960
rect 16634 16904 19890 16960
rect 19946 16904 19951 16960
rect 16573 16902 19951 16904
rect 16573 16899 16639 16902
rect 19885 16899 19951 16902
rect 20253 16962 20319 16965
rect 23013 16962 23079 16965
rect 26233 16962 26299 16965
rect 27153 16962 27219 16965
rect 20253 16960 23079 16962
rect 20253 16904 20258 16960
rect 20314 16904 23018 16960
rect 23074 16904 23079 16960
rect 20253 16902 23079 16904
rect 20253 16899 20319 16902
rect 23013 16899 23079 16902
rect 23982 16960 27219 16962
rect 23982 16904 26238 16960
rect 26294 16904 27158 16960
rect 27214 16904 27219 16960
rect 23982 16902 27219 16904
rect 30054 16960 30163 16965
rect 30054 16904 30102 16960
rect 30158 16904 30163 16960
rect 30054 16902 30163 16904
rect 15574 16896 15890 16897
rect 15574 16832 15580 16896
rect 15644 16832 15660 16896
rect 15724 16832 15740 16896
rect 15804 16832 15820 16896
rect 15884 16832 15890 16896
rect 15574 16831 15890 16832
rect 23164 16896 23480 16897
rect 23164 16832 23170 16896
rect 23234 16832 23250 16896
rect 23314 16832 23330 16896
rect 23394 16832 23410 16896
rect 23474 16832 23480 16896
rect 23164 16831 23480 16832
rect 13721 16826 13787 16829
rect 9630 16824 13787 16826
rect 9630 16768 13726 16824
rect 13782 16768 13787 16824
rect 9630 16766 13787 16768
rect 8385 16763 8451 16766
rect 9305 16763 9371 16766
rect 13721 16763 13787 16766
rect 16941 16826 17007 16829
rect 17861 16826 17927 16829
rect 16941 16824 22938 16826
rect 16941 16768 16946 16824
rect 17002 16768 17866 16824
rect 17922 16768 22938 16824
rect 16941 16766 22938 16768
rect 16941 16763 17007 16766
rect 17861 16763 17927 16766
rect 4889 16690 4955 16693
rect 10225 16690 10291 16693
rect 4889 16688 10291 16690
rect 4889 16632 4894 16688
rect 4950 16632 10230 16688
rect 10286 16632 10291 16688
rect 4889 16630 10291 16632
rect 4889 16627 4955 16630
rect 10225 16627 10291 16630
rect 11421 16690 11487 16693
rect 12801 16690 12867 16693
rect 11421 16688 12867 16690
rect 11421 16632 11426 16688
rect 11482 16632 12806 16688
rect 12862 16632 12867 16688
rect 11421 16630 12867 16632
rect 11421 16627 11487 16630
rect 12801 16627 12867 16630
rect 14917 16690 14983 16693
rect 15142 16690 15148 16692
rect 14917 16688 15148 16690
rect 14917 16632 14922 16688
rect 14978 16632 15148 16688
rect 14917 16630 15148 16632
rect 14917 16627 14983 16630
rect 15142 16628 15148 16630
rect 15212 16628 15218 16692
rect 19517 16690 19583 16693
rect 20897 16690 20963 16693
rect 19517 16688 20963 16690
rect 19517 16632 19522 16688
rect 19578 16632 20902 16688
rect 20958 16632 20963 16688
rect 19517 16630 20963 16632
rect 19517 16627 19583 16630
rect 20897 16627 20963 16630
rect 21081 16690 21147 16693
rect 22878 16690 22938 16766
rect 23982 16690 24042 16902
rect 26233 16899 26299 16902
rect 27153 16899 27219 16902
rect 30097 16899 30163 16902
rect 30754 16896 31070 16897
rect 30754 16832 30760 16896
rect 30824 16832 30840 16896
rect 30904 16832 30920 16896
rect 30984 16832 31000 16896
rect 31064 16832 31070 16896
rect 30754 16831 31070 16832
rect 21081 16688 22386 16690
rect 21081 16632 21086 16688
rect 21142 16632 22386 16688
rect 21081 16630 22386 16632
rect 22878 16630 24042 16690
rect 24761 16690 24827 16693
rect 27705 16690 27771 16693
rect 24761 16688 27771 16690
rect 24761 16632 24766 16688
rect 24822 16632 27710 16688
rect 27766 16632 27771 16688
rect 24761 16630 27771 16632
rect 21081 16627 21147 16630
rect 6862 16492 6868 16556
rect 6932 16554 6938 16556
rect 13905 16554 13971 16557
rect 6932 16552 13971 16554
rect 6932 16496 13910 16552
rect 13966 16496 13971 16552
rect 6932 16494 13971 16496
rect 6932 16492 6938 16494
rect 13905 16491 13971 16494
rect 17861 16554 17927 16557
rect 22185 16554 22251 16557
rect 17861 16552 22251 16554
rect 17861 16496 17866 16552
rect 17922 16496 22190 16552
rect 22246 16496 22251 16552
rect 17861 16494 22251 16496
rect 22326 16554 22386 16630
rect 24761 16627 24827 16630
rect 27705 16627 27771 16630
rect 23841 16554 23907 16557
rect 23974 16554 23980 16556
rect 22326 16552 23980 16554
rect 22326 16496 23846 16552
rect 23902 16496 23980 16552
rect 22326 16494 23980 16496
rect 17861 16491 17927 16494
rect 22185 16491 22251 16494
rect 23841 16491 23907 16494
rect 23974 16492 23980 16494
rect 24044 16492 24050 16556
rect 24485 16554 24551 16557
rect 26325 16554 26391 16557
rect 24485 16552 26391 16554
rect 24485 16496 24490 16552
rect 24546 16496 26330 16552
rect 26386 16496 26391 16552
rect 24485 16494 26391 16496
rect 24485 16491 24551 16494
rect 26325 16491 26391 16494
rect 7465 16418 7531 16421
rect 10685 16418 10751 16421
rect 7465 16416 10751 16418
rect 7465 16360 7470 16416
rect 7526 16360 10690 16416
rect 10746 16360 10751 16416
rect 7465 16358 10751 16360
rect 7465 16355 7531 16358
rect 10685 16355 10751 16358
rect 4189 16352 4505 16353
rect 4189 16288 4195 16352
rect 4259 16288 4275 16352
rect 4339 16288 4355 16352
rect 4419 16288 4435 16352
rect 4499 16288 4505 16352
rect 4189 16287 4505 16288
rect 11779 16352 12095 16353
rect 11779 16288 11785 16352
rect 11849 16288 11865 16352
rect 11929 16288 11945 16352
rect 12009 16288 12025 16352
rect 12089 16288 12095 16352
rect 11779 16287 12095 16288
rect 19369 16352 19685 16353
rect 19369 16288 19375 16352
rect 19439 16288 19455 16352
rect 19519 16288 19535 16352
rect 19599 16288 19615 16352
rect 19679 16288 19685 16352
rect 19369 16287 19685 16288
rect 26959 16352 27275 16353
rect 26959 16288 26965 16352
rect 27029 16288 27045 16352
rect 27109 16288 27125 16352
rect 27189 16288 27205 16352
rect 27269 16288 27275 16352
rect 26959 16287 27275 16288
rect 6453 16282 6519 16285
rect 8845 16282 8911 16285
rect 6453 16280 8911 16282
rect 6453 16224 6458 16280
rect 6514 16224 8850 16280
rect 8906 16224 8911 16280
rect 6453 16222 8911 16224
rect 6453 16219 6519 16222
rect 8845 16219 8911 16222
rect 9029 16282 9095 16285
rect 9857 16282 9923 16285
rect 9029 16280 9923 16282
rect 9029 16224 9034 16280
rect 9090 16224 9862 16280
rect 9918 16224 9923 16280
rect 9029 16222 9923 16224
rect 9029 16219 9095 16222
rect 9857 16219 9923 16222
rect 13813 16282 13879 16285
rect 15009 16282 15075 16285
rect 13813 16280 15075 16282
rect 13813 16224 13818 16280
rect 13874 16224 15014 16280
rect 15070 16224 15075 16280
rect 13813 16222 15075 16224
rect 13813 16219 13879 16222
rect 15009 16219 15075 16222
rect 27654 16220 27660 16284
rect 27724 16282 27730 16284
rect 28717 16282 28783 16285
rect 29361 16282 29427 16285
rect 27724 16280 29427 16282
rect 27724 16224 28722 16280
rect 28778 16224 29366 16280
rect 29422 16224 29427 16280
rect 27724 16222 29427 16224
rect 27724 16220 27730 16222
rect 28717 16219 28783 16222
rect 29361 16219 29427 16222
rect 2037 16146 2103 16149
rect 24761 16146 24827 16149
rect 27797 16146 27863 16149
rect 2037 16144 22110 16146
rect 2037 16088 2042 16144
rect 2098 16088 22110 16144
rect 2037 16086 22110 16088
rect 2037 16083 2103 16086
rect 4429 16010 4495 16013
rect 10501 16010 10567 16013
rect 4429 16008 10567 16010
rect 4429 15952 4434 16008
rect 4490 15952 10506 16008
rect 10562 15952 10567 16008
rect 4429 15950 10567 15952
rect 4429 15947 4495 15950
rect 10501 15947 10567 15950
rect 10685 16010 10751 16013
rect 16205 16010 16271 16013
rect 10685 16008 16271 16010
rect 10685 15952 10690 16008
rect 10746 15952 16210 16008
rect 16266 15952 16271 16008
rect 10685 15950 16271 15952
rect 10685 15947 10751 15950
rect 16205 15947 16271 15950
rect 16573 16010 16639 16013
rect 17217 16010 17283 16013
rect 16573 16008 17283 16010
rect 16573 15952 16578 16008
rect 16634 15952 17222 16008
rect 17278 15952 17283 16008
rect 16573 15950 17283 15952
rect 22050 16010 22110 16086
rect 24761 16144 27863 16146
rect 24761 16088 24766 16144
rect 24822 16088 27802 16144
rect 27858 16088 27863 16144
rect 24761 16086 27863 16088
rect 24761 16083 24827 16086
rect 27797 16083 27863 16086
rect 29177 16010 29243 16013
rect 22050 16008 29243 16010
rect 22050 15952 29182 16008
rect 29238 15952 29243 16008
rect 22050 15950 29243 15952
rect 16573 15947 16639 15950
rect 17217 15947 17283 15950
rect 29177 15947 29243 15950
rect 7984 15808 8300 15809
rect 7984 15744 7990 15808
rect 8054 15744 8070 15808
rect 8134 15744 8150 15808
rect 8214 15744 8230 15808
rect 8294 15744 8300 15808
rect 7984 15743 8300 15744
rect 15574 15808 15890 15809
rect 15574 15744 15580 15808
rect 15644 15744 15660 15808
rect 15724 15744 15740 15808
rect 15804 15744 15820 15808
rect 15884 15744 15890 15808
rect 15574 15743 15890 15744
rect 23164 15808 23480 15809
rect 23164 15744 23170 15808
rect 23234 15744 23250 15808
rect 23314 15744 23330 15808
rect 23394 15744 23410 15808
rect 23474 15744 23480 15808
rect 23164 15743 23480 15744
rect 30754 15808 31070 15809
rect 30754 15744 30760 15808
rect 30824 15744 30840 15808
rect 30904 15744 30920 15808
rect 30984 15744 31000 15808
rect 31064 15744 31070 15808
rect 30754 15743 31070 15744
rect 11789 15738 11855 15741
rect 14733 15738 14799 15741
rect 11789 15736 14799 15738
rect 11789 15680 11794 15736
rect 11850 15680 14738 15736
rect 14794 15680 14799 15736
rect 11789 15678 14799 15680
rect 11789 15675 11855 15678
rect 14733 15675 14799 15678
rect 27429 15738 27495 15741
rect 28349 15738 28415 15741
rect 27429 15736 28415 15738
rect 27429 15680 27434 15736
rect 27490 15680 28354 15736
rect 28410 15680 28415 15736
rect 27429 15678 28415 15680
rect 27429 15675 27495 15678
rect 28349 15675 28415 15678
rect 3509 15602 3575 15605
rect 9489 15602 9555 15605
rect 3509 15600 9555 15602
rect 3509 15544 3514 15600
rect 3570 15544 9494 15600
rect 9550 15544 9555 15600
rect 3509 15542 9555 15544
rect 3509 15539 3575 15542
rect 9489 15539 9555 15542
rect 11421 15602 11487 15605
rect 23381 15602 23447 15605
rect 28625 15602 28691 15605
rect 11421 15600 16590 15602
rect 11421 15544 11426 15600
rect 11482 15544 16590 15600
rect 11421 15542 16590 15544
rect 11421 15539 11487 15542
rect 2129 15466 2195 15469
rect 8518 15466 8524 15468
rect 2129 15464 8524 15466
rect 2129 15408 2134 15464
rect 2190 15408 8524 15464
rect 2129 15406 8524 15408
rect 2129 15403 2195 15406
rect 8518 15404 8524 15406
rect 8588 15404 8594 15468
rect 9121 15466 9187 15469
rect 16113 15466 16179 15469
rect 9121 15464 16179 15466
rect 9121 15408 9126 15464
rect 9182 15408 16118 15464
rect 16174 15408 16179 15464
rect 9121 15406 16179 15408
rect 16530 15466 16590 15542
rect 23381 15600 28691 15602
rect 23381 15544 23386 15600
rect 23442 15544 28630 15600
rect 28686 15544 28691 15600
rect 23381 15542 28691 15544
rect 23381 15539 23447 15542
rect 28625 15539 28691 15542
rect 16849 15466 16915 15469
rect 29177 15466 29243 15469
rect 16530 15464 29243 15466
rect 16530 15408 16854 15464
rect 16910 15408 29182 15464
rect 29238 15408 29243 15464
rect 16530 15406 29243 15408
rect 9121 15403 9187 15406
rect 16113 15403 16179 15406
rect 16849 15403 16915 15406
rect 29177 15403 29243 15406
rect 5993 15330 6059 15333
rect 7741 15330 7807 15333
rect 5993 15328 7807 15330
rect 5993 15272 5998 15328
rect 6054 15272 7746 15328
rect 7802 15272 7807 15328
rect 5993 15270 7807 15272
rect 5993 15267 6059 15270
rect 7741 15267 7807 15270
rect 4189 15264 4505 15265
rect 4189 15200 4195 15264
rect 4259 15200 4275 15264
rect 4339 15200 4355 15264
rect 4419 15200 4435 15264
rect 4499 15200 4505 15264
rect 4189 15199 4505 15200
rect 11779 15264 12095 15265
rect 11779 15200 11785 15264
rect 11849 15200 11865 15264
rect 11929 15200 11945 15264
rect 12009 15200 12025 15264
rect 12089 15200 12095 15264
rect 11779 15199 12095 15200
rect 19369 15264 19685 15265
rect 19369 15200 19375 15264
rect 19439 15200 19455 15264
rect 19519 15200 19535 15264
rect 19599 15200 19615 15264
rect 19679 15200 19685 15264
rect 19369 15199 19685 15200
rect 26959 15264 27275 15265
rect 26959 15200 26965 15264
rect 27029 15200 27045 15264
rect 27109 15200 27125 15264
rect 27189 15200 27205 15264
rect 27269 15200 27275 15264
rect 26959 15199 27275 15200
rect 5073 15194 5139 15197
rect 7649 15194 7715 15197
rect 11513 15194 11579 15197
rect 5073 15192 7482 15194
rect 5073 15136 5078 15192
rect 5134 15136 7482 15192
rect 5073 15134 7482 15136
rect 5073 15131 5139 15134
rect 1945 15058 2011 15061
rect 3969 15058 4035 15061
rect 5349 15058 5415 15061
rect 1945 15056 2790 15058
rect 1945 15000 1950 15056
rect 2006 15000 2790 15056
rect 1945 14998 2790 15000
rect 1945 14995 2011 14998
rect 2730 14922 2790 14998
rect 3969 15056 5415 15058
rect 3969 15000 3974 15056
rect 4030 15000 5354 15056
rect 5410 15000 5415 15056
rect 3969 14998 5415 15000
rect 3969 14995 4035 14998
rect 5349 14995 5415 14998
rect 5809 15058 5875 15061
rect 7189 15058 7255 15061
rect 5809 15056 7255 15058
rect 5809 15000 5814 15056
rect 5870 15000 7194 15056
rect 7250 15000 7255 15056
rect 5809 14998 7255 15000
rect 7422 15058 7482 15134
rect 7649 15192 11579 15194
rect 7649 15136 7654 15192
rect 7710 15136 11518 15192
rect 11574 15136 11579 15192
rect 7649 15134 11579 15136
rect 7649 15131 7715 15134
rect 11513 15131 11579 15134
rect 24485 15194 24551 15197
rect 26693 15194 26759 15197
rect 24485 15192 26759 15194
rect 24485 15136 24490 15192
rect 24546 15136 26698 15192
rect 26754 15136 26759 15192
rect 24485 15134 26759 15136
rect 24485 15131 24551 15134
rect 26693 15131 26759 15134
rect 8569 15058 8635 15061
rect 7422 15056 8635 15058
rect 7422 15000 8574 15056
rect 8630 15000 8635 15056
rect 7422 14998 8635 15000
rect 5809 14995 5875 14998
rect 7189 14995 7255 14998
rect 8569 14995 8635 14998
rect 9213 15058 9279 15061
rect 12985 15058 13051 15061
rect 9213 15056 13051 15058
rect 9213 15000 9218 15056
rect 9274 15000 12990 15056
rect 13046 15000 13051 15056
rect 9213 14998 13051 15000
rect 9213 14995 9279 14998
rect 12985 14995 13051 14998
rect 21173 15058 21239 15061
rect 24945 15058 25011 15061
rect 21173 15056 25011 15058
rect 21173 15000 21178 15056
rect 21234 15000 24950 15056
rect 25006 15000 25011 15056
rect 21173 14998 25011 15000
rect 21173 14995 21239 14998
rect 24945 14995 25011 14998
rect 9213 14922 9279 14925
rect 14825 14922 14891 14925
rect 2730 14920 9279 14922
rect 2730 14864 9218 14920
rect 9274 14864 9279 14920
rect 2730 14862 9279 14864
rect 9213 14859 9279 14862
rect 9630 14920 14891 14922
rect 9630 14864 14830 14920
rect 14886 14864 14891 14920
rect 9630 14862 14891 14864
rect 5165 14786 5231 14789
rect 7097 14786 7163 14789
rect 5165 14784 7163 14786
rect 5165 14728 5170 14784
rect 5226 14728 7102 14784
rect 7158 14728 7163 14784
rect 5165 14726 7163 14728
rect 5165 14723 5231 14726
rect 7097 14723 7163 14726
rect 7984 14720 8300 14721
rect 7984 14656 7990 14720
rect 8054 14656 8070 14720
rect 8134 14656 8150 14720
rect 8214 14656 8230 14720
rect 8294 14656 8300 14720
rect 7984 14655 8300 14656
rect 3325 14650 3391 14653
rect 6177 14650 6243 14653
rect 3325 14648 6243 14650
rect 3325 14592 3330 14648
rect 3386 14592 6182 14648
rect 6238 14592 6243 14648
rect 3325 14590 6243 14592
rect 3325 14587 3391 14590
rect 6177 14587 6243 14590
rect 1393 14514 1459 14517
rect 4429 14514 4495 14517
rect 6361 14514 6427 14517
rect 1393 14512 6427 14514
rect 1393 14456 1398 14512
rect 1454 14456 4434 14512
rect 4490 14456 6366 14512
rect 6422 14456 6427 14512
rect 1393 14454 6427 14456
rect 1393 14451 1459 14454
rect 4429 14451 4495 14454
rect 6361 14451 6427 14454
rect 6729 14514 6795 14517
rect 9630 14514 9690 14862
rect 14825 14859 14891 14862
rect 16113 14922 16179 14925
rect 27797 14922 27863 14925
rect 16113 14920 27863 14922
rect 16113 14864 16118 14920
rect 16174 14864 27802 14920
rect 27858 14864 27863 14920
rect 16113 14862 27863 14864
rect 16113 14859 16179 14862
rect 27797 14859 27863 14862
rect 11329 14786 11395 14789
rect 12617 14786 12683 14789
rect 11329 14784 12683 14786
rect 11329 14728 11334 14784
rect 11390 14728 12622 14784
rect 12678 14728 12683 14784
rect 11329 14726 12683 14728
rect 11329 14723 11395 14726
rect 12617 14723 12683 14726
rect 23565 14786 23631 14789
rect 25405 14786 25471 14789
rect 23565 14784 25471 14786
rect 23565 14728 23570 14784
rect 23626 14728 25410 14784
rect 25466 14728 25471 14784
rect 23565 14726 25471 14728
rect 23565 14723 23631 14726
rect 25405 14723 25471 14726
rect 15574 14720 15890 14721
rect 15574 14656 15580 14720
rect 15644 14656 15660 14720
rect 15724 14656 15740 14720
rect 15804 14656 15820 14720
rect 15884 14656 15890 14720
rect 15574 14655 15890 14656
rect 23164 14720 23480 14721
rect 23164 14656 23170 14720
rect 23234 14656 23250 14720
rect 23314 14656 23330 14720
rect 23394 14656 23410 14720
rect 23474 14656 23480 14720
rect 23164 14655 23480 14656
rect 30754 14720 31070 14721
rect 30754 14656 30760 14720
rect 30824 14656 30840 14720
rect 30904 14656 30920 14720
rect 30984 14656 31000 14720
rect 31064 14656 31070 14720
rect 30754 14655 31070 14656
rect 10317 14650 10383 14653
rect 13261 14650 13327 14653
rect 10317 14648 13327 14650
rect 10317 14592 10322 14648
rect 10378 14592 13266 14648
rect 13322 14592 13327 14648
rect 10317 14590 13327 14592
rect 10317 14587 10383 14590
rect 13261 14587 13327 14590
rect 13997 14650 14063 14653
rect 14917 14650 14983 14653
rect 13997 14648 14983 14650
rect 13997 14592 14002 14648
rect 14058 14592 14922 14648
rect 14978 14592 14983 14648
rect 13997 14590 14983 14592
rect 13997 14587 14063 14590
rect 14917 14587 14983 14590
rect 19241 14514 19307 14517
rect 6729 14512 9690 14514
rect 6729 14456 6734 14512
rect 6790 14456 9690 14512
rect 6729 14454 9690 14456
rect 12390 14512 19307 14514
rect 12390 14456 19246 14512
rect 19302 14456 19307 14512
rect 12390 14454 19307 14456
rect 6729 14451 6795 14454
rect 2078 14316 2084 14380
rect 2148 14378 2154 14380
rect 9857 14378 9923 14381
rect 2148 14376 9923 14378
rect 2148 14320 9862 14376
rect 9918 14320 9923 14376
rect 2148 14318 9923 14320
rect 2148 14316 2154 14318
rect 9857 14315 9923 14318
rect 11237 14378 11303 14381
rect 11421 14378 11487 14381
rect 11237 14376 11487 14378
rect 11237 14320 11242 14376
rect 11298 14320 11426 14376
rect 11482 14320 11487 14376
rect 11237 14318 11487 14320
rect 11237 14315 11303 14318
rect 11421 14315 11487 14318
rect 5625 14242 5691 14245
rect 7281 14242 7347 14245
rect 5625 14240 7347 14242
rect 5625 14184 5630 14240
rect 5686 14184 7286 14240
rect 7342 14184 7347 14240
rect 5625 14182 7347 14184
rect 5625 14179 5691 14182
rect 7281 14179 7347 14182
rect 9438 14180 9444 14244
rect 9508 14242 9514 14244
rect 11237 14242 11303 14245
rect 9508 14240 11303 14242
rect 9508 14184 11242 14240
rect 11298 14184 11303 14240
rect 9508 14182 11303 14184
rect 9508 14180 9514 14182
rect 11237 14179 11303 14182
rect 4189 14176 4505 14177
rect 4189 14112 4195 14176
rect 4259 14112 4275 14176
rect 4339 14112 4355 14176
rect 4419 14112 4435 14176
rect 4499 14112 4505 14176
rect 4189 14111 4505 14112
rect 11779 14176 12095 14177
rect 11779 14112 11785 14176
rect 11849 14112 11865 14176
rect 11929 14112 11945 14176
rect 12009 14112 12025 14176
rect 12089 14112 12095 14176
rect 11779 14111 12095 14112
rect 5717 14106 5783 14109
rect 7005 14106 7071 14109
rect 5717 14104 7071 14106
rect 5717 14048 5722 14104
rect 5778 14048 7010 14104
rect 7066 14048 7071 14104
rect 5717 14046 7071 14048
rect 5717 14043 5783 14046
rect 7005 14043 7071 14046
rect 9673 14106 9739 14109
rect 10133 14106 10199 14109
rect 9673 14104 10199 14106
rect 9673 14048 9678 14104
rect 9734 14048 10138 14104
rect 10194 14048 10199 14104
rect 9673 14046 10199 14048
rect 9673 14043 9739 14046
rect 10133 14043 10199 14046
rect 12390 13970 12450 14454
rect 19241 14451 19307 14454
rect 25773 14514 25839 14517
rect 27061 14514 27127 14517
rect 25773 14512 27127 14514
rect 25773 14456 25778 14512
rect 25834 14456 27066 14512
rect 27122 14456 27127 14512
rect 25773 14454 27127 14456
rect 25773 14451 25839 14454
rect 27061 14451 27127 14454
rect 19517 14378 19583 14381
rect 28349 14378 28415 14381
rect 19517 14376 28415 14378
rect 19517 14320 19522 14376
rect 19578 14320 28354 14376
rect 28410 14320 28415 14376
rect 19517 14318 28415 14320
rect 19517 14315 19583 14318
rect 28349 14315 28415 14318
rect 19369 14176 19685 14177
rect 19369 14112 19375 14176
rect 19439 14112 19455 14176
rect 19519 14112 19535 14176
rect 19599 14112 19615 14176
rect 19679 14112 19685 14176
rect 19369 14111 19685 14112
rect 26959 14176 27275 14177
rect 26959 14112 26965 14176
rect 27029 14112 27045 14176
rect 27109 14112 27125 14176
rect 27189 14112 27205 14176
rect 27269 14112 27275 14176
rect 26959 14111 27275 14112
rect 16941 14106 17007 14109
rect 18137 14106 18203 14109
rect 16941 14104 18203 14106
rect 16941 14048 16946 14104
rect 17002 14048 18142 14104
rect 18198 14048 18203 14104
rect 16941 14046 18203 14048
rect 16941 14043 17007 14046
rect 18137 14043 18203 14046
rect 6870 13910 12450 13970
rect 14365 13970 14431 13973
rect 17677 13970 17743 13973
rect 14365 13968 17743 13970
rect 14365 13912 14370 13968
rect 14426 13912 17682 13968
rect 17738 13912 17743 13968
rect 14365 13910 17743 13912
rect 2129 13698 2195 13701
rect 6870 13698 6930 13910
rect 14365 13907 14431 13910
rect 17677 13907 17743 13910
rect 18873 13970 18939 13973
rect 26049 13970 26115 13973
rect 18873 13968 26115 13970
rect 18873 13912 18878 13968
rect 18934 13912 26054 13968
rect 26110 13912 26115 13968
rect 18873 13910 26115 13912
rect 18873 13907 18939 13910
rect 26049 13907 26115 13910
rect 10869 13834 10935 13837
rect 11881 13834 11947 13837
rect 2129 13696 6930 13698
rect 2129 13640 2134 13696
rect 2190 13640 6930 13696
rect 2129 13638 6930 13640
rect 7790 13774 8586 13834
rect 2129 13635 2195 13638
rect 4889 13562 4955 13565
rect 7649 13562 7715 13565
rect 4889 13560 7715 13562
rect 4889 13504 4894 13560
rect 4950 13504 7654 13560
rect 7710 13504 7715 13560
rect 4889 13502 7715 13504
rect 4889 13499 4955 13502
rect 7649 13499 7715 13502
rect 3141 13426 3207 13429
rect 5441 13426 5507 13429
rect 7790 13426 7850 13774
rect 7984 13632 8300 13633
rect 7984 13568 7990 13632
rect 8054 13568 8070 13632
rect 8134 13568 8150 13632
rect 8214 13568 8230 13632
rect 8294 13568 8300 13632
rect 7984 13567 8300 13568
rect 8526 13562 8586 13774
rect 10869 13832 11947 13834
rect 10869 13776 10874 13832
rect 10930 13776 11886 13832
rect 11942 13776 11947 13832
rect 10869 13774 11947 13776
rect 10869 13771 10935 13774
rect 11881 13771 11947 13774
rect 24393 13834 24459 13837
rect 28533 13834 28599 13837
rect 29085 13834 29151 13837
rect 24393 13832 29151 13834
rect 24393 13776 24398 13832
rect 24454 13776 28538 13832
rect 28594 13776 29090 13832
rect 29146 13776 29151 13832
rect 24393 13774 29151 13776
rect 24393 13771 24459 13774
rect 28533 13771 28599 13774
rect 29085 13771 29151 13774
rect 8886 13636 8892 13700
rect 8956 13698 8962 13700
rect 10409 13698 10475 13701
rect 8956 13696 10475 13698
rect 8956 13640 10414 13696
rect 10470 13640 10475 13696
rect 8956 13638 10475 13640
rect 8956 13636 8962 13638
rect 10409 13635 10475 13638
rect 10777 13698 10843 13701
rect 11094 13698 11100 13700
rect 10777 13696 11100 13698
rect 10777 13640 10782 13696
rect 10838 13640 11100 13696
rect 10777 13638 11100 13640
rect 10777 13635 10843 13638
rect 11094 13636 11100 13638
rect 11164 13636 11170 13700
rect 11513 13698 11579 13701
rect 14273 13698 14339 13701
rect 11513 13696 14339 13698
rect 11513 13640 11518 13696
rect 11574 13640 14278 13696
rect 14334 13640 14339 13696
rect 11513 13638 14339 13640
rect 11513 13635 11579 13638
rect 14273 13635 14339 13638
rect 15574 13632 15890 13633
rect 15574 13568 15580 13632
rect 15644 13568 15660 13632
rect 15724 13568 15740 13632
rect 15804 13568 15820 13632
rect 15884 13568 15890 13632
rect 15574 13567 15890 13568
rect 23164 13632 23480 13633
rect 23164 13568 23170 13632
rect 23234 13568 23250 13632
rect 23314 13568 23330 13632
rect 23394 13568 23410 13632
rect 23474 13568 23480 13632
rect 23164 13567 23480 13568
rect 30754 13632 31070 13633
rect 30754 13568 30760 13632
rect 30824 13568 30840 13632
rect 30904 13568 30920 13632
rect 30984 13568 31000 13632
rect 31064 13568 31070 13632
rect 30754 13567 31070 13568
rect 12065 13562 12131 13565
rect 8526 13560 12131 13562
rect 8526 13504 12070 13560
rect 12126 13504 12131 13560
rect 8526 13502 12131 13504
rect 12065 13499 12131 13502
rect 3141 13424 7850 13426
rect 3141 13368 3146 13424
rect 3202 13368 5446 13424
rect 5502 13368 7850 13424
rect 3141 13366 7850 13368
rect 3141 13363 3207 13366
rect 5441 13363 5507 13366
rect 8518 13364 8524 13428
rect 8588 13426 8594 13428
rect 16757 13426 16823 13429
rect 8588 13424 16823 13426
rect 8588 13368 16762 13424
rect 16818 13368 16823 13424
rect 8588 13366 16823 13368
rect 8588 13364 8594 13366
rect 16757 13363 16823 13366
rect 21725 13426 21791 13429
rect 22737 13426 22803 13429
rect 24301 13426 24367 13429
rect 21725 13424 24367 13426
rect 21725 13368 21730 13424
rect 21786 13368 22742 13424
rect 22798 13368 24306 13424
rect 24362 13368 24367 13424
rect 21725 13366 24367 13368
rect 21725 13363 21791 13366
rect 22737 13363 22803 13366
rect 24301 13363 24367 13366
rect 26049 13426 26115 13429
rect 27613 13426 27679 13429
rect 26049 13424 27679 13426
rect 26049 13368 26054 13424
rect 26110 13368 27618 13424
rect 27674 13368 27679 13424
rect 26049 13366 27679 13368
rect 26049 13363 26115 13366
rect 27613 13363 27679 13366
rect 3325 13290 3391 13293
rect 3325 13288 4952 13290
rect 3325 13232 3330 13288
rect 3386 13232 4952 13288
rect 3325 13230 4952 13232
rect 3325 13227 3391 13230
rect 4189 13088 4505 13089
rect 4189 13024 4195 13088
rect 4259 13024 4275 13088
rect 4339 13024 4355 13088
rect 4419 13024 4435 13088
rect 4499 13024 4505 13088
rect 4189 13023 4505 13024
rect 4892 13018 4952 13230
rect 5022 13228 5028 13292
rect 5092 13228 5098 13292
rect 7097 13290 7163 13293
rect 11513 13290 11579 13293
rect 11881 13290 11947 13293
rect 7097 13288 11579 13290
rect 7097 13232 7102 13288
rect 7158 13232 11518 13288
rect 11574 13232 11579 13288
rect 7097 13230 11579 13232
rect 5030 13154 5090 13228
rect 7097 13227 7163 13230
rect 11513 13227 11579 13230
rect 11654 13288 11947 13290
rect 11654 13232 11886 13288
rect 11942 13232 11947 13288
rect 11654 13230 11947 13232
rect 11654 13154 11714 13230
rect 11881 13227 11947 13230
rect 12065 13290 12131 13293
rect 16941 13290 17007 13293
rect 17953 13290 18019 13293
rect 12065 13288 18019 13290
rect 12065 13232 12070 13288
rect 12126 13232 16946 13288
rect 17002 13232 17958 13288
rect 18014 13232 18019 13288
rect 12065 13230 18019 13232
rect 12065 13227 12131 13230
rect 16941 13227 17007 13230
rect 17953 13227 18019 13230
rect 20069 13290 20135 13293
rect 29177 13290 29243 13293
rect 31385 13290 31451 13293
rect 20069 13288 31451 13290
rect 20069 13232 20074 13288
rect 20130 13232 29182 13288
rect 29238 13232 31390 13288
rect 31446 13232 31451 13288
rect 20069 13230 31451 13232
rect 20069 13227 20135 13230
rect 29177 13227 29243 13230
rect 31385 13227 31451 13230
rect 5030 13094 11714 13154
rect 11779 13088 12095 13089
rect 11779 13024 11785 13088
rect 11849 13024 11865 13088
rect 11929 13024 11945 13088
rect 12009 13024 12025 13088
rect 12089 13024 12095 13088
rect 11779 13023 12095 13024
rect 19369 13088 19685 13089
rect 19369 13024 19375 13088
rect 19439 13024 19455 13088
rect 19519 13024 19535 13088
rect 19599 13024 19615 13088
rect 19679 13024 19685 13088
rect 19369 13023 19685 13024
rect 26959 13088 27275 13089
rect 26959 13024 26965 13088
rect 27029 13024 27045 13088
rect 27109 13024 27125 13088
rect 27189 13024 27205 13088
rect 27269 13024 27275 13088
rect 26959 13023 27275 13024
rect 10041 13018 10107 13021
rect 4892 13016 10107 13018
rect 4892 12960 10046 13016
rect 10102 12960 10107 13016
rect 4892 12958 10107 12960
rect 10041 12955 10107 12958
rect 13353 13018 13419 13021
rect 13813 13018 13879 13021
rect 13353 13016 13879 13018
rect 13353 12960 13358 13016
rect 13414 12960 13818 13016
rect 13874 12960 13879 13016
rect 13353 12958 13879 12960
rect 13353 12955 13419 12958
rect 13813 12955 13879 12958
rect 3509 12882 3575 12885
rect 14457 12882 14523 12885
rect 22921 12882 22987 12885
rect 24485 12882 24551 12885
rect 3509 12880 19350 12882
rect 3509 12824 3514 12880
rect 3570 12824 14462 12880
rect 14518 12824 19350 12880
rect 3509 12822 19350 12824
rect 3509 12819 3575 12822
rect 14457 12819 14523 12822
rect 3049 12746 3115 12749
rect 4245 12746 4311 12749
rect 3049 12744 4311 12746
rect 3049 12688 3054 12744
rect 3110 12688 4250 12744
rect 4306 12688 4311 12744
rect 3049 12686 4311 12688
rect 3049 12683 3115 12686
rect 4245 12683 4311 12686
rect 5257 12746 5323 12749
rect 9121 12746 9187 12749
rect 5257 12744 9187 12746
rect 5257 12688 5262 12744
rect 5318 12688 9126 12744
rect 9182 12688 9187 12744
rect 5257 12686 9187 12688
rect 5257 12683 5323 12686
rect 9121 12683 9187 12686
rect 9857 12746 9923 12749
rect 10961 12746 11027 12749
rect 9857 12744 11027 12746
rect 9857 12688 9862 12744
rect 9918 12688 10966 12744
rect 11022 12688 11027 12744
rect 9857 12686 11027 12688
rect 9857 12683 9923 12686
rect 10961 12683 11027 12686
rect 11973 12746 12039 12749
rect 16297 12746 16363 12749
rect 11973 12744 16363 12746
rect 11973 12688 11978 12744
rect 12034 12688 16302 12744
rect 16358 12688 16363 12744
rect 11973 12686 16363 12688
rect 19290 12746 19350 12822
rect 22921 12880 24551 12882
rect 22921 12824 22926 12880
rect 22982 12824 24490 12880
rect 24546 12824 24551 12880
rect 22921 12822 24551 12824
rect 22921 12819 22987 12822
rect 24485 12819 24551 12822
rect 27654 12746 27660 12748
rect 19290 12686 27660 12746
rect 11973 12683 12039 12686
rect 16297 12683 16363 12686
rect 27654 12684 27660 12686
rect 27724 12684 27730 12748
rect 2221 12610 2287 12613
rect 11053 12610 11119 12613
rect 12617 12610 12683 12613
rect 13813 12610 13879 12613
rect 2221 12608 3986 12610
rect 2221 12552 2226 12608
rect 2282 12552 3986 12608
rect 2221 12550 3986 12552
rect 2221 12547 2287 12550
rect 3926 12338 3986 12550
rect 11053 12608 13879 12610
rect 11053 12552 11058 12608
rect 11114 12552 12622 12608
rect 12678 12552 13818 12608
rect 13874 12552 13879 12608
rect 11053 12550 13879 12552
rect 11053 12547 11119 12550
rect 12617 12547 12683 12550
rect 13813 12547 13879 12550
rect 23749 12610 23815 12613
rect 27981 12610 28047 12613
rect 23749 12608 28047 12610
rect 23749 12552 23754 12608
rect 23810 12552 27986 12608
rect 28042 12552 28047 12608
rect 23749 12550 28047 12552
rect 23749 12547 23815 12550
rect 27981 12547 28047 12550
rect 7984 12544 8300 12545
rect 7984 12480 7990 12544
rect 8054 12480 8070 12544
rect 8134 12480 8150 12544
rect 8214 12480 8230 12544
rect 8294 12480 8300 12544
rect 7984 12479 8300 12480
rect 15574 12544 15890 12545
rect 15574 12480 15580 12544
rect 15644 12480 15660 12544
rect 15724 12480 15740 12544
rect 15804 12480 15820 12544
rect 15884 12480 15890 12544
rect 15574 12479 15890 12480
rect 23164 12544 23480 12545
rect 23164 12480 23170 12544
rect 23234 12480 23250 12544
rect 23314 12480 23330 12544
rect 23394 12480 23410 12544
rect 23474 12480 23480 12544
rect 23164 12479 23480 12480
rect 30754 12544 31070 12545
rect 30754 12480 30760 12544
rect 30824 12480 30840 12544
rect 30904 12480 30920 12544
rect 30984 12480 31000 12544
rect 31064 12480 31070 12544
rect 30754 12479 31070 12480
rect 6453 12474 6519 12477
rect 7373 12474 7439 12477
rect 6453 12472 7439 12474
rect 6453 12416 6458 12472
rect 6514 12416 7378 12472
rect 7434 12416 7439 12472
rect 6453 12414 7439 12416
rect 6453 12411 6519 12414
rect 7373 12411 7439 12414
rect 11973 12474 12039 12477
rect 13077 12474 13143 12477
rect 11973 12472 13143 12474
rect 11973 12416 11978 12472
rect 12034 12416 13082 12472
rect 13138 12416 13143 12472
rect 11973 12414 13143 12416
rect 11973 12411 12039 12414
rect 13077 12411 13143 12414
rect 15285 12338 15351 12341
rect 3926 12336 15351 12338
rect 3926 12280 15290 12336
rect 15346 12280 15351 12336
rect 3926 12278 15351 12280
rect 15285 12275 15351 12278
rect 2681 12202 2747 12205
rect 15561 12202 15627 12205
rect 2681 12200 15627 12202
rect 2681 12144 2686 12200
rect 2742 12144 15566 12200
rect 15622 12144 15627 12200
rect 2681 12142 15627 12144
rect 2681 12139 2747 12142
rect 15561 12139 15627 12142
rect 13169 12066 13235 12069
rect 13445 12066 13511 12069
rect 16205 12066 16271 12069
rect 13169 12064 16271 12066
rect 13169 12008 13174 12064
rect 13230 12008 13450 12064
rect 13506 12008 16210 12064
rect 16266 12008 16271 12064
rect 13169 12006 16271 12008
rect 13169 12003 13235 12006
rect 13445 12003 13511 12006
rect 16205 12003 16271 12006
rect 4189 12000 4505 12001
rect 4189 11936 4195 12000
rect 4259 11936 4275 12000
rect 4339 11936 4355 12000
rect 4419 11936 4435 12000
rect 4499 11936 4505 12000
rect 4189 11935 4505 11936
rect 11779 12000 12095 12001
rect 11779 11936 11785 12000
rect 11849 11936 11865 12000
rect 11929 11936 11945 12000
rect 12009 11936 12025 12000
rect 12089 11936 12095 12000
rect 11779 11935 12095 11936
rect 19369 12000 19685 12001
rect 19369 11936 19375 12000
rect 19439 11936 19455 12000
rect 19519 11936 19535 12000
rect 19599 11936 19615 12000
rect 19679 11936 19685 12000
rect 19369 11935 19685 11936
rect 26959 12000 27275 12001
rect 26959 11936 26965 12000
rect 27029 11936 27045 12000
rect 27109 11936 27125 12000
rect 27189 11936 27205 12000
rect 27269 11936 27275 12000
rect 26959 11935 27275 11936
rect 2405 11930 2471 11933
rect 5901 11930 5967 11933
rect 9121 11930 9187 11933
rect 15009 11930 15075 11933
rect 2405 11928 2790 11930
rect 2405 11872 2410 11928
rect 2466 11872 2790 11928
rect 2405 11870 2790 11872
rect 2405 11867 2471 11870
rect 2730 11794 2790 11870
rect 5901 11928 9187 11930
rect 5901 11872 5906 11928
rect 5962 11872 9126 11928
rect 9182 11872 9187 11928
rect 5901 11870 9187 11872
rect 5901 11867 5967 11870
rect 9121 11867 9187 11870
rect 12390 11928 15075 11930
rect 12390 11872 15014 11928
rect 15070 11872 15075 11928
rect 12390 11870 15075 11872
rect 12390 11794 12450 11870
rect 15009 11867 15075 11870
rect 2730 11734 12450 11794
rect 23974 11732 23980 11796
rect 24044 11794 24050 11796
rect 24117 11794 24183 11797
rect 27613 11794 27679 11797
rect 24044 11792 27679 11794
rect 24044 11736 24122 11792
rect 24178 11736 27618 11792
rect 27674 11736 27679 11792
rect 24044 11734 27679 11736
rect 24044 11732 24050 11734
rect 24117 11731 24183 11734
rect 27613 11731 27679 11734
rect 5441 11658 5507 11661
rect 11421 11658 11487 11661
rect 5441 11656 11487 11658
rect 5441 11600 5446 11656
rect 5502 11600 11426 11656
rect 11482 11600 11487 11656
rect 5441 11598 11487 11600
rect 5441 11595 5507 11598
rect 11421 11595 11487 11598
rect 11605 11658 11671 11661
rect 13445 11658 13511 11661
rect 11605 11656 13511 11658
rect 11605 11600 11610 11656
rect 11666 11600 13450 11656
rect 13506 11600 13511 11656
rect 11605 11598 13511 11600
rect 11605 11595 11671 11598
rect 13445 11595 13511 11598
rect 15142 11596 15148 11660
rect 15212 11658 15218 11660
rect 26049 11658 26115 11661
rect 15212 11656 26115 11658
rect 15212 11600 26054 11656
rect 26110 11600 26115 11656
rect 15212 11598 26115 11600
rect 15212 11596 15218 11598
rect 26049 11595 26115 11598
rect 3509 11522 3575 11525
rect 6177 11522 6243 11525
rect 7373 11522 7439 11525
rect 3509 11520 7439 11522
rect 3509 11464 3514 11520
rect 3570 11464 6182 11520
rect 6238 11464 7378 11520
rect 7434 11464 7439 11520
rect 3509 11462 7439 11464
rect 3509 11459 3575 11462
rect 6177 11459 6243 11462
rect 7373 11459 7439 11462
rect 7984 11456 8300 11457
rect 7984 11392 7990 11456
rect 8054 11392 8070 11456
rect 8134 11392 8150 11456
rect 8214 11392 8230 11456
rect 8294 11392 8300 11456
rect 7984 11391 8300 11392
rect 15574 11456 15890 11457
rect 15574 11392 15580 11456
rect 15644 11392 15660 11456
rect 15724 11392 15740 11456
rect 15804 11392 15820 11456
rect 15884 11392 15890 11456
rect 15574 11391 15890 11392
rect 23164 11456 23480 11457
rect 23164 11392 23170 11456
rect 23234 11392 23250 11456
rect 23314 11392 23330 11456
rect 23394 11392 23410 11456
rect 23474 11392 23480 11456
rect 23164 11391 23480 11392
rect 30754 11456 31070 11457
rect 30754 11392 30760 11456
rect 30824 11392 30840 11456
rect 30904 11392 30920 11456
rect 30984 11392 31000 11456
rect 31064 11392 31070 11456
rect 30754 11391 31070 11392
rect 1669 11386 1735 11389
rect 5073 11386 5139 11389
rect 1669 11384 5139 11386
rect 1669 11328 1674 11384
rect 1730 11328 5078 11384
rect 5134 11328 5139 11384
rect 1669 11326 5139 11328
rect 1669 11323 1735 11326
rect 5073 11323 5139 11326
rect 8518 11324 8524 11388
rect 8588 11386 8594 11388
rect 8845 11386 8911 11389
rect 8588 11384 8911 11386
rect 8588 11328 8850 11384
rect 8906 11328 8911 11384
rect 8588 11326 8911 11328
rect 8588 11324 8594 11326
rect 8845 11323 8911 11326
rect 9765 11386 9831 11389
rect 12065 11386 12131 11389
rect 9765 11384 12131 11386
rect 9765 11328 9770 11384
rect 9826 11328 12070 11384
rect 12126 11328 12131 11384
rect 9765 11326 12131 11328
rect 9765 11323 9831 11326
rect 12065 11323 12131 11326
rect 3877 11250 3943 11253
rect 15469 11250 15535 11253
rect 25865 11250 25931 11253
rect 3877 11248 25931 11250
rect 3877 11192 3882 11248
rect 3938 11192 15474 11248
rect 15530 11192 25870 11248
rect 25926 11192 25931 11248
rect 3877 11190 25931 11192
rect 3877 11187 3943 11190
rect 15469 11187 15535 11190
rect 25865 11187 25931 11190
rect 1393 11114 1459 11117
rect 3233 11114 3299 11117
rect 1393 11112 3299 11114
rect 1393 11056 1398 11112
rect 1454 11056 3238 11112
rect 3294 11056 3299 11112
rect 1393 11054 3299 11056
rect 1393 11051 1459 11054
rect 3233 11051 3299 11054
rect 3693 11114 3759 11117
rect 9765 11114 9831 11117
rect 3693 11112 9831 11114
rect 3693 11056 3698 11112
rect 3754 11056 9770 11112
rect 9826 11056 9831 11112
rect 3693 11054 9831 11056
rect 3693 11051 3759 11054
rect 9765 11051 9831 11054
rect 10358 11052 10364 11116
rect 10428 11052 10434 11116
rect 20437 11114 20503 11117
rect 30005 11114 30071 11117
rect 20437 11112 30071 11114
rect 20437 11056 20442 11112
rect 20498 11056 30010 11112
rect 30066 11056 30071 11112
rect 20437 11054 30071 11056
rect 10366 10978 10426 11052
rect 20437 11051 20503 11054
rect 30005 11051 30071 11054
rect 11513 10978 11579 10981
rect 10366 10976 11579 10978
rect 10366 10920 11518 10976
rect 11574 10920 11579 10976
rect 10366 10918 11579 10920
rect 11513 10915 11579 10918
rect 4189 10912 4505 10913
rect 4189 10848 4195 10912
rect 4259 10848 4275 10912
rect 4339 10848 4355 10912
rect 4419 10848 4435 10912
rect 4499 10848 4505 10912
rect 4189 10847 4505 10848
rect 11779 10912 12095 10913
rect 11779 10848 11785 10912
rect 11849 10848 11865 10912
rect 11929 10848 11945 10912
rect 12009 10848 12025 10912
rect 12089 10848 12095 10912
rect 11779 10847 12095 10848
rect 19369 10912 19685 10913
rect 19369 10848 19375 10912
rect 19439 10848 19455 10912
rect 19519 10848 19535 10912
rect 19599 10848 19615 10912
rect 19679 10848 19685 10912
rect 19369 10847 19685 10848
rect 26959 10912 27275 10913
rect 26959 10848 26965 10912
rect 27029 10848 27045 10912
rect 27109 10848 27125 10912
rect 27189 10848 27205 10912
rect 27269 10848 27275 10912
rect 26959 10847 27275 10848
rect 2129 10706 2195 10709
rect 9949 10706 10015 10709
rect 2129 10704 10015 10706
rect 2129 10648 2134 10704
rect 2190 10648 9954 10704
rect 10010 10648 10015 10704
rect 2129 10646 10015 10648
rect 2129 10643 2195 10646
rect 9949 10643 10015 10646
rect 18873 10706 18939 10709
rect 19333 10706 19399 10709
rect 18873 10704 19399 10706
rect 18873 10648 18878 10704
rect 18934 10648 19338 10704
rect 19394 10648 19399 10704
rect 18873 10646 19399 10648
rect 18873 10643 18939 10646
rect 19333 10643 19399 10646
rect 11329 10570 11395 10573
rect 12893 10570 12959 10573
rect 2730 10568 11395 10570
rect 2730 10512 11334 10568
rect 11390 10512 11395 10568
rect 2730 10510 11395 10512
rect 1669 10162 1735 10165
rect 2730 10162 2790 10510
rect 11329 10507 11395 10510
rect 12390 10568 12959 10570
rect 12390 10512 12898 10568
rect 12954 10512 12959 10568
rect 12390 10510 12959 10512
rect 3233 10434 3299 10437
rect 3969 10434 4035 10437
rect 3233 10432 4035 10434
rect 3233 10376 3238 10432
rect 3294 10376 3974 10432
rect 4030 10376 4035 10432
rect 3233 10374 4035 10376
rect 3233 10371 3299 10374
rect 3969 10371 4035 10374
rect 7984 10368 8300 10369
rect 7984 10304 7990 10368
rect 8054 10304 8070 10368
rect 8134 10304 8150 10368
rect 8214 10304 8230 10368
rect 8294 10304 8300 10368
rect 7984 10303 8300 10304
rect 3141 10298 3207 10301
rect 3141 10296 6562 10298
rect 3141 10240 3146 10296
rect 3202 10240 6562 10296
rect 3141 10238 6562 10240
rect 3141 10235 3207 10238
rect 6361 10162 6427 10165
rect 1669 10160 2790 10162
rect 1669 10104 1674 10160
rect 1730 10104 2790 10160
rect 1669 10102 2790 10104
rect 3926 10160 6427 10162
rect 3926 10104 6366 10160
rect 6422 10104 6427 10160
rect 3926 10102 6427 10104
rect 6502 10162 6562 10238
rect 12390 10162 12450 10510
rect 12893 10507 12959 10510
rect 15574 10368 15890 10369
rect 15574 10304 15580 10368
rect 15644 10304 15660 10368
rect 15724 10304 15740 10368
rect 15804 10304 15820 10368
rect 15884 10304 15890 10368
rect 15574 10303 15890 10304
rect 23164 10368 23480 10369
rect 23164 10304 23170 10368
rect 23234 10304 23250 10368
rect 23314 10304 23330 10368
rect 23394 10304 23410 10368
rect 23474 10304 23480 10368
rect 23164 10303 23480 10304
rect 30754 10368 31070 10369
rect 30754 10304 30760 10368
rect 30824 10304 30840 10368
rect 30904 10304 30920 10368
rect 30984 10304 31000 10368
rect 31064 10304 31070 10368
rect 30754 10303 31070 10304
rect 6502 10102 12450 10162
rect 1669 10099 1735 10102
rect 3926 9890 3986 10102
rect 6361 10099 6427 10102
rect 4061 10026 4127 10029
rect 13721 10026 13787 10029
rect 4061 10024 13787 10026
rect 4061 9968 4066 10024
rect 4122 9968 13726 10024
rect 13782 9968 13787 10024
rect 4061 9966 13787 9968
rect 4061 9963 4127 9966
rect 13721 9963 13787 9966
rect 4061 9890 4127 9893
rect 3926 9888 4127 9890
rect 3926 9832 4066 9888
rect 4122 9832 4127 9888
rect 3926 9830 4127 9832
rect 4061 9827 4127 9830
rect 6545 9890 6611 9893
rect 7005 9890 7071 9893
rect 6545 9888 7071 9890
rect 6545 9832 6550 9888
rect 6606 9832 7010 9888
rect 7066 9832 7071 9888
rect 6545 9830 7071 9832
rect 6545 9827 6611 9830
rect 7005 9827 7071 9830
rect 16389 9888 16455 9893
rect 16389 9832 16394 9888
rect 16450 9832 16455 9888
rect 16389 9827 16455 9832
rect 4189 9824 4505 9825
rect 4189 9760 4195 9824
rect 4259 9760 4275 9824
rect 4339 9760 4355 9824
rect 4419 9760 4435 9824
rect 4499 9760 4505 9824
rect 4189 9759 4505 9760
rect 11779 9824 12095 9825
rect 11779 9760 11785 9824
rect 11849 9760 11865 9824
rect 11929 9760 11945 9824
rect 12009 9760 12025 9824
rect 12089 9760 12095 9824
rect 11779 9759 12095 9760
rect 16392 9754 16452 9827
rect 19369 9824 19685 9825
rect 19369 9760 19375 9824
rect 19439 9760 19455 9824
rect 19519 9760 19535 9824
rect 19599 9760 19615 9824
rect 19679 9760 19685 9824
rect 19369 9759 19685 9760
rect 26959 9824 27275 9825
rect 26959 9760 26965 9824
rect 27029 9760 27045 9824
rect 27109 9760 27125 9824
rect 27189 9760 27205 9824
rect 27269 9760 27275 9824
rect 26959 9759 27275 9760
rect 16392 9694 17004 9754
rect 5625 9690 5691 9693
rect 5582 9688 5691 9690
rect 5582 9632 5630 9688
rect 5686 9632 5691 9688
rect 5582 9627 5691 9632
rect 1025 9482 1091 9485
rect 5257 9482 5323 9485
rect 1025 9480 5323 9482
rect 1025 9424 1030 9480
rect 1086 9424 5262 9480
rect 5318 9424 5323 9480
rect 1025 9422 5323 9424
rect 5582 9482 5642 9627
rect 10041 9618 10107 9621
rect 11881 9618 11947 9621
rect 10041 9616 11947 9618
rect 10041 9560 10046 9616
rect 10102 9560 11886 9616
rect 11942 9560 11947 9616
rect 10041 9558 11947 9560
rect 16944 9618 17004 9694
rect 16944 9558 17556 9618
rect 10041 9555 10107 9558
rect 11881 9555 11947 9558
rect 17496 9485 17556 9558
rect 5809 9482 5875 9485
rect 5582 9480 5875 9482
rect 5582 9424 5814 9480
rect 5870 9424 5875 9480
rect 5582 9422 5875 9424
rect 1025 9419 1091 9422
rect 5257 9419 5323 9422
rect 5809 9419 5875 9422
rect 10777 9482 10843 9485
rect 12249 9482 12315 9485
rect 10777 9480 12315 9482
rect 10777 9424 10782 9480
rect 10838 9424 12254 9480
rect 12310 9424 12315 9480
rect 10777 9422 12315 9424
rect 10777 9419 10843 9422
rect 12249 9419 12315 9422
rect 17493 9482 17559 9485
rect 24853 9482 24919 9485
rect 17493 9480 24919 9482
rect 17493 9424 17498 9480
rect 17554 9424 24858 9480
rect 24914 9424 24919 9480
rect 17493 9422 24919 9424
rect 17493 9419 17559 9422
rect 24853 9419 24919 9422
rect 16757 9346 16823 9349
rect 17217 9346 17283 9349
rect 17769 9346 17835 9349
rect 16757 9344 17835 9346
rect 16757 9288 16762 9344
rect 16818 9288 17222 9344
rect 17278 9288 17774 9344
rect 17830 9288 17835 9344
rect 16757 9286 17835 9288
rect 16757 9283 16823 9286
rect 17217 9283 17283 9286
rect 17769 9283 17835 9286
rect 7984 9280 8300 9281
rect 7984 9216 7990 9280
rect 8054 9216 8070 9280
rect 8134 9216 8150 9280
rect 8214 9216 8230 9280
rect 8294 9216 8300 9280
rect 7984 9215 8300 9216
rect 15574 9280 15890 9281
rect 15574 9216 15580 9280
rect 15644 9216 15660 9280
rect 15724 9216 15740 9280
rect 15804 9216 15820 9280
rect 15884 9216 15890 9280
rect 15574 9215 15890 9216
rect 23164 9280 23480 9281
rect 23164 9216 23170 9280
rect 23234 9216 23250 9280
rect 23314 9216 23330 9280
rect 23394 9216 23410 9280
rect 23474 9216 23480 9280
rect 23164 9215 23480 9216
rect 30754 9280 31070 9281
rect 30754 9216 30760 9280
rect 30824 9216 30840 9280
rect 30904 9216 30920 9280
rect 30984 9216 31000 9280
rect 31064 9216 31070 9280
rect 30754 9215 31070 9216
rect 16113 9210 16179 9213
rect 17769 9210 17835 9213
rect 16113 9208 17835 9210
rect 16113 9152 16118 9208
rect 16174 9152 17774 9208
rect 17830 9152 17835 9208
rect 16113 9150 17835 9152
rect 16113 9147 16179 9150
rect 17769 9147 17835 9150
rect 2865 9074 2931 9077
rect 5257 9074 5323 9077
rect 2865 9072 5323 9074
rect 2865 9016 2870 9072
rect 2926 9016 5262 9072
rect 5318 9016 5323 9072
rect 2865 9014 5323 9016
rect 2865 9011 2931 9014
rect 5257 9011 5323 9014
rect 7465 9074 7531 9077
rect 9121 9074 9187 9077
rect 7465 9072 9187 9074
rect 7465 9016 7470 9072
rect 7526 9016 9126 9072
rect 9182 9016 9187 9072
rect 7465 9014 9187 9016
rect 7465 9011 7531 9014
rect 9121 9011 9187 9014
rect 10317 9074 10383 9077
rect 11421 9074 11487 9077
rect 10317 9072 11487 9074
rect 10317 9016 10322 9072
rect 10378 9016 11426 9072
rect 11482 9016 11487 9072
rect 10317 9014 11487 9016
rect 10317 9011 10383 9014
rect 11421 9011 11487 9014
rect 16297 9074 16363 9077
rect 16757 9074 16823 9077
rect 16297 9072 16823 9074
rect 16297 9016 16302 9072
rect 16358 9016 16762 9072
rect 16818 9016 16823 9072
rect 16297 9014 16823 9016
rect 16297 9011 16363 9014
rect 16757 9011 16823 9014
rect 17033 9074 17099 9077
rect 18229 9074 18295 9077
rect 17033 9072 18295 9074
rect 17033 9016 17038 9072
rect 17094 9016 18234 9072
rect 18290 9016 18295 9072
rect 17033 9014 18295 9016
rect 17033 9011 17099 9014
rect 18229 9011 18295 9014
rect 22921 9074 22987 9077
rect 26141 9074 26207 9077
rect 22921 9072 26207 9074
rect 22921 9016 22926 9072
rect 22982 9016 26146 9072
rect 26202 9016 26207 9072
rect 22921 9014 26207 9016
rect 22921 9011 22987 9014
rect 26141 9011 26207 9014
rect 3141 8938 3207 8941
rect 14038 8938 14044 8940
rect 3141 8936 14044 8938
rect 3141 8880 3146 8936
rect 3202 8880 14044 8936
rect 3141 8878 14044 8880
rect 3141 8875 3207 8878
rect 14038 8876 14044 8878
rect 14108 8876 14114 8940
rect 17401 8938 17467 8941
rect 18413 8938 18479 8941
rect 17401 8936 18479 8938
rect 17401 8880 17406 8936
rect 17462 8880 18418 8936
rect 18474 8880 18479 8936
rect 17401 8878 18479 8880
rect 17401 8875 17467 8878
rect 18413 8875 18479 8878
rect 5441 8802 5507 8805
rect 9857 8802 9923 8805
rect 5441 8800 9923 8802
rect 5441 8744 5446 8800
rect 5502 8744 9862 8800
rect 9918 8744 9923 8800
rect 5441 8742 9923 8744
rect 5441 8739 5507 8742
rect 9857 8739 9923 8742
rect 4189 8736 4505 8737
rect 4189 8672 4195 8736
rect 4259 8672 4275 8736
rect 4339 8672 4355 8736
rect 4419 8672 4435 8736
rect 4499 8672 4505 8736
rect 4189 8671 4505 8672
rect 11779 8736 12095 8737
rect 11779 8672 11785 8736
rect 11849 8672 11865 8736
rect 11929 8672 11945 8736
rect 12009 8672 12025 8736
rect 12089 8672 12095 8736
rect 11779 8671 12095 8672
rect 19369 8736 19685 8737
rect 19369 8672 19375 8736
rect 19439 8672 19455 8736
rect 19519 8672 19535 8736
rect 19599 8672 19615 8736
rect 19679 8672 19685 8736
rect 19369 8671 19685 8672
rect 26959 8736 27275 8737
rect 26959 8672 26965 8736
rect 27029 8672 27045 8736
rect 27109 8672 27125 8736
rect 27189 8672 27205 8736
rect 27269 8672 27275 8736
rect 26959 8671 27275 8672
rect 3969 8530 4035 8533
rect 15929 8530 15995 8533
rect 3969 8528 15995 8530
rect 3969 8472 3974 8528
rect 4030 8472 15934 8528
rect 15990 8472 15995 8528
rect 3969 8470 15995 8472
rect 3969 8467 4035 8470
rect 15929 8467 15995 8470
rect 5717 8394 5783 8397
rect 6269 8394 6335 8397
rect 5717 8392 6335 8394
rect 5717 8336 5722 8392
rect 5778 8336 6274 8392
rect 6330 8336 6335 8392
rect 5717 8334 6335 8336
rect 5717 8331 5783 8334
rect 6269 8331 6335 8334
rect 10685 8394 10751 8397
rect 16573 8394 16639 8397
rect 10685 8392 16639 8394
rect 10685 8336 10690 8392
rect 10746 8336 16578 8392
rect 16634 8336 16639 8392
rect 10685 8334 16639 8336
rect 10685 8331 10751 8334
rect 16573 8331 16639 8334
rect 7984 8192 8300 8193
rect 7984 8128 7990 8192
rect 8054 8128 8070 8192
rect 8134 8128 8150 8192
rect 8214 8128 8230 8192
rect 8294 8128 8300 8192
rect 7984 8127 8300 8128
rect 15574 8192 15890 8193
rect 15574 8128 15580 8192
rect 15644 8128 15660 8192
rect 15724 8128 15740 8192
rect 15804 8128 15820 8192
rect 15884 8128 15890 8192
rect 15574 8127 15890 8128
rect 23164 8192 23480 8193
rect 23164 8128 23170 8192
rect 23234 8128 23250 8192
rect 23314 8128 23330 8192
rect 23394 8128 23410 8192
rect 23474 8128 23480 8192
rect 23164 8127 23480 8128
rect 30754 8192 31070 8193
rect 30754 8128 30760 8192
rect 30824 8128 30840 8192
rect 30904 8128 30920 8192
rect 30984 8128 31000 8192
rect 31064 8128 31070 8192
rect 30754 8127 31070 8128
rect 5901 8122 5967 8125
rect 6913 8122 6979 8125
rect 5901 8120 6979 8122
rect 5901 8064 5906 8120
rect 5962 8064 6918 8120
rect 6974 8064 6979 8120
rect 5901 8062 6979 8064
rect 5901 8059 5967 8062
rect 6913 8059 6979 8062
rect 4061 7986 4127 7989
rect 6545 7986 6611 7989
rect 4061 7984 6611 7986
rect 4061 7928 4066 7984
rect 4122 7928 6550 7984
rect 6606 7928 6611 7984
rect 4061 7926 6611 7928
rect 4061 7923 4127 7926
rect 6545 7923 6611 7926
rect 6729 7986 6795 7989
rect 13445 7986 13511 7989
rect 6729 7984 13511 7986
rect 6729 7928 6734 7984
rect 6790 7928 13450 7984
rect 13506 7928 13511 7984
rect 6729 7926 13511 7928
rect 6729 7923 6795 7926
rect 13445 7923 13511 7926
rect 15929 7986 15995 7989
rect 22553 7986 22619 7989
rect 15929 7984 22619 7986
rect 15929 7928 15934 7984
rect 15990 7928 22558 7984
rect 22614 7928 22619 7984
rect 15929 7926 22619 7928
rect 15929 7923 15995 7926
rect 22553 7923 22619 7926
rect 1761 7850 1827 7853
rect 10593 7850 10659 7853
rect 1761 7848 10659 7850
rect 1761 7792 1766 7848
rect 1822 7792 10598 7848
rect 10654 7792 10659 7848
rect 1761 7790 10659 7792
rect 1761 7787 1827 7790
rect 10593 7787 10659 7790
rect 11654 7790 12266 7850
rect 8661 7714 8727 7717
rect 9581 7714 9647 7717
rect 11654 7714 11714 7790
rect 8661 7712 11714 7714
rect 8661 7656 8666 7712
rect 8722 7656 9586 7712
rect 9642 7656 11714 7712
rect 8661 7654 11714 7656
rect 8661 7651 8727 7654
rect 9581 7651 9647 7654
rect 4189 7648 4505 7649
rect 4189 7584 4195 7648
rect 4259 7584 4275 7648
rect 4339 7584 4355 7648
rect 4419 7584 4435 7648
rect 4499 7584 4505 7648
rect 4189 7583 4505 7584
rect 11779 7648 12095 7649
rect 11779 7584 11785 7648
rect 11849 7584 11865 7648
rect 11929 7584 11945 7648
rect 12009 7584 12025 7648
rect 12089 7584 12095 7648
rect 11779 7583 12095 7584
rect 8109 7578 8175 7581
rect 10501 7578 10567 7581
rect 8109 7576 10567 7578
rect 8109 7520 8114 7576
rect 8170 7520 10506 7576
rect 10562 7520 10567 7576
rect 8109 7518 10567 7520
rect 8109 7515 8175 7518
rect 10501 7515 10567 7518
rect 1945 7442 2011 7445
rect 11605 7442 11671 7445
rect 1945 7440 11671 7442
rect 1945 7384 1950 7440
rect 2006 7384 11610 7440
rect 11666 7384 11671 7440
rect 1945 7382 11671 7384
rect 12206 7442 12266 7790
rect 12382 7788 12388 7852
rect 12452 7850 12458 7852
rect 12617 7850 12683 7853
rect 12452 7848 12683 7850
rect 12452 7792 12622 7848
rect 12678 7792 12683 7848
rect 12452 7790 12683 7792
rect 12452 7788 12458 7790
rect 12617 7787 12683 7790
rect 22001 7850 22067 7853
rect 28901 7850 28967 7853
rect 22001 7848 28967 7850
rect 22001 7792 22006 7848
rect 22062 7792 28906 7848
rect 28962 7792 28967 7848
rect 22001 7790 28967 7792
rect 22001 7787 22067 7790
rect 28901 7787 28967 7790
rect 19369 7648 19685 7649
rect 19369 7584 19375 7648
rect 19439 7584 19455 7648
rect 19519 7584 19535 7648
rect 19599 7584 19615 7648
rect 19679 7584 19685 7648
rect 19369 7583 19685 7584
rect 26959 7648 27275 7649
rect 26959 7584 26965 7648
rect 27029 7584 27045 7648
rect 27109 7584 27125 7648
rect 27189 7584 27205 7648
rect 27269 7584 27275 7648
rect 26959 7583 27275 7584
rect 14457 7578 14523 7581
rect 16941 7578 17007 7581
rect 14457 7576 17007 7578
rect 14457 7520 14462 7576
rect 14518 7520 16946 7576
rect 17002 7520 17007 7576
rect 14457 7518 17007 7520
rect 14457 7515 14523 7518
rect 16941 7515 17007 7518
rect 16573 7442 16639 7445
rect 18321 7442 18387 7445
rect 12206 7440 18387 7442
rect 12206 7384 16578 7440
rect 16634 7384 18326 7440
rect 18382 7384 18387 7440
rect 12206 7382 18387 7384
rect 1945 7379 2011 7382
rect 11605 7379 11671 7382
rect 16573 7379 16639 7382
rect 18321 7379 18387 7382
rect 18689 7442 18755 7445
rect 25129 7442 25195 7445
rect 18689 7440 25195 7442
rect 18689 7384 18694 7440
rect 18750 7384 25134 7440
rect 25190 7384 25195 7440
rect 18689 7382 25195 7384
rect 18689 7379 18755 7382
rect 25129 7379 25195 7382
rect 1669 7306 1735 7309
rect 17033 7306 17099 7309
rect 23473 7306 23539 7309
rect 1669 7304 17099 7306
rect 1669 7248 1674 7304
rect 1730 7248 17038 7304
rect 17094 7248 17099 7304
rect 1669 7246 17099 7248
rect 1669 7243 1735 7246
rect 17033 7243 17099 7246
rect 22050 7304 23539 7306
rect 22050 7248 23478 7304
rect 23534 7248 23539 7304
rect 22050 7246 23539 7248
rect 3141 7170 3207 7173
rect 7649 7170 7715 7173
rect 9397 7172 9463 7173
rect 9397 7170 9444 7172
rect 3141 7168 7715 7170
rect 3141 7112 3146 7168
rect 3202 7112 7654 7168
rect 7710 7112 7715 7168
rect 3141 7110 7715 7112
rect 9316 7168 9444 7170
rect 9508 7170 9514 7172
rect 12525 7170 12591 7173
rect 14273 7170 14339 7173
rect 9508 7168 14339 7170
rect 9316 7112 9402 7168
rect 9508 7112 12530 7168
rect 12586 7112 14278 7168
rect 14334 7112 14339 7168
rect 9316 7110 9444 7112
rect 3141 7107 3207 7110
rect 7649 7107 7715 7110
rect 9397 7108 9444 7110
rect 9508 7110 14339 7112
rect 9508 7108 9514 7110
rect 9397 7107 9463 7108
rect 12525 7107 12591 7110
rect 14273 7107 14339 7110
rect 16389 7170 16455 7173
rect 22050 7170 22110 7246
rect 23473 7243 23539 7246
rect 16389 7168 22110 7170
rect 16389 7112 16394 7168
rect 16450 7112 22110 7168
rect 16389 7110 22110 7112
rect 16389 7107 16455 7110
rect 7984 7104 8300 7105
rect 7984 7040 7990 7104
rect 8054 7040 8070 7104
rect 8134 7040 8150 7104
rect 8214 7040 8230 7104
rect 8294 7040 8300 7104
rect 7984 7039 8300 7040
rect 15574 7104 15890 7105
rect 15574 7040 15580 7104
rect 15644 7040 15660 7104
rect 15724 7040 15740 7104
rect 15804 7040 15820 7104
rect 15884 7040 15890 7104
rect 15574 7039 15890 7040
rect 23164 7104 23480 7105
rect 23164 7040 23170 7104
rect 23234 7040 23250 7104
rect 23314 7040 23330 7104
rect 23394 7040 23410 7104
rect 23474 7040 23480 7104
rect 23164 7039 23480 7040
rect 30754 7104 31070 7105
rect 30754 7040 30760 7104
rect 30824 7040 30840 7104
rect 30904 7040 30920 7104
rect 30984 7040 31000 7104
rect 31064 7040 31070 7104
rect 30754 7039 31070 7040
rect 1761 7034 1827 7037
rect 7373 7034 7439 7037
rect 1761 7032 7439 7034
rect 1761 6976 1766 7032
rect 1822 6976 7378 7032
rect 7434 6976 7439 7032
rect 1761 6974 7439 6976
rect 1761 6971 1827 6974
rect 7373 6971 7439 6974
rect 10501 7034 10567 7037
rect 14641 7034 14707 7037
rect 10501 7032 14707 7034
rect 10501 6976 10506 7032
rect 10562 6976 14646 7032
rect 14702 6976 14707 7032
rect 10501 6974 14707 6976
rect 10501 6971 10567 6974
rect 14641 6971 14707 6974
rect 5901 6898 5967 6901
rect 7189 6898 7255 6901
rect 5901 6896 7255 6898
rect 5901 6840 5906 6896
rect 5962 6840 7194 6896
rect 7250 6840 7255 6896
rect 5901 6838 7255 6840
rect 5901 6835 5967 6838
rect 7189 6835 7255 6838
rect 9397 6898 9463 6901
rect 13721 6898 13787 6901
rect 9397 6896 13787 6898
rect 9397 6840 9402 6896
rect 9458 6840 13726 6896
rect 13782 6840 13787 6896
rect 9397 6838 13787 6840
rect 9397 6835 9463 6838
rect 13721 6835 13787 6838
rect 16573 6898 16639 6901
rect 17033 6898 17099 6901
rect 24577 6898 24643 6901
rect 16573 6896 24643 6898
rect 16573 6840 16578 6896
rect 16634 6840 17038 6896
rect 17094 6840 24582 6896
rect 24638 6840 24643 6896
rect 16573 6838 24643 6840
rect 16573 6835 16639 6838
rect 17033 6835 17099 6838
rect 24577 6835 24643 6838
rect 2589 6762 2655 6765
rect 9397 6762 9463 6765
rect 2589 6760 9463 6762
rect 2589 6704 2594 6760
rect 2650 6704 9402 6760
rect 9458 6704 9463 6760
rect 2589 6702 9463 6704
rect 2589 6699 2655 6702
rect 9397 6699 9463 6702
rect 9765 6762 9831 6765
rect 16205 6762 16271 6765
rect 9765 6760 16271 6762
rect 9765 6704 9770 6760
rect 9826 6704 16210 6760
rect 16266 6704 16271 6760
rect 9765 6702 16271 6704
rect 9765 6699 9831 6702
rect 16205 6699 16271 6702
rect 17125 6762 17191 6765
rect 20161 6762 20227 6765
rect 17125 6760 20227 6762
rect 17125 6704 17130 6760
rect 17186 6704 20166 6760
rect 20222 6704 20227 6760
rect 17125 6702 20227 6704
rect 17125 6699 17191 6702
rect 20161 6699 20227 6702
rect 4189 6560 4505 6561
rect 4189 6496 4195 6560
rect 4259 6496 4275 6560
rect 4339 6496 4355 6560
rect 4419 6496 4435 6560
rect 4499 6496 4505 6560
rect 4189 6495 4505 6496
rect 11779 6560 12095 6561
rect 11779 6496 11785 6560
rect 11849 6496 11865 6560
rect 11929 6496 11945 6560
rect 12009 6496 12025 6560
rect 12089 6496 12095 6560
rect 11779 6495 12095 6496
rect 19369 6560 19685 6561
rect 19369 6496 19375 6560
rect 19439 6496 19455 6560
rect 19519 6496 19535 6560
rect 19599 6496 19615 6560
rect 19679 6496 19685 6560
rect 19369 6495 19685 6496
rect 26959 6560 27275 6561
rect 26959 6496 26965 6560
rect 27029 6496 27045 6560
rect 27109 6496 27125 6560
rect 27189 6496 27205 6560
rect 27269 6496 27275 6560
rect 26959 6495 27275 6496
rect 6085 6354 6151 6357
rect 15285 6354 15351 6357
rect 6085 6352 15351 6354
rect 6085 6296 6090 6352
rect 6146 6296 15290 6352
rect 15346 6296 15351 6352
rect 6085 6294 15351 6296
rect 6085 6291 6151 6294
rect 15285 6291 15351 6294
rect 22185 6354 22251 6357
rect 28533 6354 28599 6357
rect 22185 6352 28599 6354
rect 22185 6296 22190 6352
rect 22246 6296 28538 6352
rect 28594 6296 28599 6352
rect 22185 6294 28599 6296
rect 22185 6291 22251 6294
rect 28533 6291 28599 6294
rect 5257 6218 5323 6221
rect 10593 6218 10659 6221
rect 5257 6216 10659 6218
rect 5257 6160 5262 6216
rect 5318 6160 10598 6216
rect 10654 6160 10659 6216
rect 5257 6158 10659 6160
rect 5257 6155 5323 6158
rect 10593 6155 10659 6158
rect 10869 6218 10935 6221
rect 12198 6218 12204 6220
rect 10869 6216 12204 6218
rect 10869 6160 10874 6216
rect 10930 6160 12204 6216
rect 10869 6158 12204 6160
rect 10869 6155 10935 6158
rect 12198 6156 12204 6158
rect 12268 6156 12274 6220
rect 13537 6218 13603 6221
rect 12390 6216 13603 6218
rect 12390 6160 13542 6216
rect 13598 6160 13603 6216
rect 12390 6158 13603 6160
rect 9121 6082 9187 6085
rect 12390 6082 12450 6158
rect 13537 6155 13603 6158
rect 23381 6218 23447 6221
rect 29361 6218 29427 6221
rect 23381 6216 29427 6218
rect 23381 6160 23386 6216
rect 23442 6160 29366 6216
rect 29422 6160 29427 6216
rect 23381 6158 29427 6160
rect 23381 6155 23447 6158
rect 29361 6155 29427 6158
rect 9121 6080 12450 6082
rect 9121 6024 9126 6080
rect 9182 6024 12450 6080
rect 9121 6022 12450 6024
rect 9121 6019 9187 6022
rect 7984 6016 8300 6017
rect 7984 5952 7990 6016
rect 8054 5952 8070 6016
rect 8134 5952 8150 6016
rect 8214 5952 8230 6016
rect 8294 5952 8300 6016
rect 7984 5951 8300 5952
rect 15574 6016 15890 6017
rect 15574 5952 15580 6016
rect 15644 5952 15660 6016
rect 15724 5952 15740 6016
rect 15804 5952 15820 6016
rect 15884 5952 15890 6016
rect 15574 5951 15890 5952
rect 23164 6016 23480 6017
rect 23164 5952 23170 6016
rect 23234 5952 23250 6016
rect 23314 5952 23330 6016
rect 23394 5952 23410 6016
rect 23474 5952 23480 6016
rect 23164 5951 23480 5952
rect 30754 6016 31070 6017
rect 30754 5952 30760 6016
rect 30824 5952 30840 6016
rect 30904 5952 30920 6016
rect 30984 5952 31000 6016
rect 31064 5952 31070 6016
rect 30754 5951 31070 5952
rect 3509 5946 3575 5949
rect 5717 5946 5783 5949
rect 3509 5944 5783 5946
rect 3509 5888 3514 5944
rect 3570 5888 5722 5944
rect 5778 5888 5783 5944
rect 3509 5886 5783 5888
rect 3509 5883 3575 5886
rect 5717 5883 5783 5886
rect 13353 5946 13419 5949
rect 16481 5946 16547 5949
rect 22645 5946 22711 5949
rect 13353 5944 13922 5946
rect 13353 5888 13358 5944
rect 13414 5888 13922 5944
rect 13353 5886 13922 5888
rect 13353 5883 13419 5886
rect 2037 5810 2103 5813
rect 13721 5810 13787 5813
rect 2037 5808 13787 5810
rect 2037 5752 2042 5808
rect 2098 5752 13726 5808
rect 13782 5752 13787 5808
rect 2037 5750 13787 5752
rect 13862 5810 13922 5886
rect 16481 5944 22711 5946
rect 16481 5888 16486 5944
rect 16542 5888 22650 5944
rect 22706 5888 22711 5944
rect 16481 5886 22711 5888
rect 16481 5883 16547 5886
rect 22645 5883 22711 5886
rect 24025 5946 24091 5949
rect 25681 5946 25747 5949
rect 24025 5944 25747 5946
rect 24025 5888 24030 5944
rect 24086 5888 25686 5944
rect 25742 5888 25747 5944
rect 24025 5886 25747 5888
rect 24025 5883 24091 5886
rect 25681 5883 25747 5886
rect 26325 5810 26391 5813
rect 13862 5808 26391 5810
rect 13862 5752 26330 5808
rect 26386 5752 26391 5808
rect 13862 5750 26391 5752
rect 2037 5747 2103 5750
rect 13721 5747 13787 5750
rect 26325 5747 26391 5750
rect 6361 5674 6427 5677
rect 15193 5674 15259 5677
rect 6361 5672 15259 5674
rect 6361 5616 6366 5672
rect 6422 5616 15198 5672
rect 15254 5616 15259 5672
rect 6361 5614 15259 5616
rect 6361 5611 6427 5614
rect 15193 5611 15259 5614
rect 23105 5674 23171 5677
rect 29453 5674 29519 5677
rect 23105 5672 29519 5674
rect 23105 5616 23110 5672
rect 23166 5616 29458 5672
rect 29514 5616 29519 5672
rect 23105 5614 29519 5616
rect 23105 5611 23171 5614
rect 29453 5611 29519 5614
rect 4797 5538 4863 5541
rect 8937 5538 9003 5541
rect 4797 5536 9003 5538
rect 4797 5480 4802 5536
rect 4858 5480 8942 5536
rect 8998 5480 9003 5536
rect 4797 5478 9003 5480
rect 4797 5475 4863 5478
rect 8937 5475 9003 5478
rect 4189 5472 4505 5473
rect 4189 5408 4195 5472
rect 4259 5408 4275 5472
rect 4339 5408 4355 5472
rect 4419 5408 4435 5472
rect 4499 5408 4505 5472
rect 4189 5407 4505 5408
rect 11779 5472 12095 5473
rect 11779 5408 11785 5472
rect 11849 5408 11865 5472
rect 11929 5408 11945 5472
rect 12009 5408 12025 5472
rect 12089 5408 12095 5472
rect 11779 5407 12095 5408
rect 19369 5472 19685 5473
rect 19369 5408 19375 5472
rect 19439 5408 19455 5472
rect 19519 5408 19535 5472
rect 19599 5408 19615 5472
rect 19679 5408 19685 5472
rect 19369 5407 19685 5408
rect 26959 5472 27275 5473
rect 26959 5408 26965 5472
rect 27029 5408 27045 5472
rect 27109 5408 27125 5472
rect 27189 5408 27205 5472
rect 27269 5408 27275 5472
rect 26959 5407 27275 5408
rect 2589 5266 2655 5269
rect 13629 5266 13695 5269
rect 2589 5264 13695 5266
rect 2589 5208 2594 5264
rect 2650 5208 13634 5264
rect 13690 5208 13695 5264
rect 2589 5206 13695 5208
rect 2589 5203 2655 5206
rect 13629 5203 13695 5206
rect 11145 5130 11211 5133
rect 17769 5130 17835 5133
rect 25865 5130 25931 5133
rect 11145 5128 17835 5130
rect 11145 5072 11150 5128
rect 11206 5072 17774 5128
rect 17830 5072 17835 5128
rect 11145 5070 17835 5072
rect 11145 5067 11211 5070
rect 17769 5067 17835 5070
rect 19290 5128 25931 5130
rect 19290 5072 25870 5128
rect 25926 5072 25931 5128
rect 19290 5070 25931 5072
rect 2681 4994 2747 4997
rect 2865 4994 2931 4997
rect 2681 4992 2931 4994
rect 2681 4936 2686 4992
rect 2742 4936 2870 4992
rect 2926 4936 2931 4992
rect 2681 4934 2931 4936
rect 2681 4931 2747 4934
rect 2865 4931 2931 4934
rect 8753 4994 8819 4997
rect 9213 4994 9279 4997
rect 8753 4992 9279 4994
rect 8753 4936 8758 4992
rect 8814 4936 9218 4992
rect 9274 4936 9279 4992
rect 8753 4934 9279 4936
rect 8753 4931 8819 4934
rect 9213 4931 9279 4934
rect 18873 4994 18939 4997
rect 19290 4994 19350 5070
rect 25865 5067 25931 5070
rect 18873 4992 19350 4994
rect 18873 4936 18878 4992
rect 18934 4936 19350 4992
rect 18873 4934 19350 4936
rect 18873 4931 18939 4934
rect 7984 4928 8300 4929
rect 7984 4864 7990 4928
rect 8054 4864 8070 4928
rect 8134 4864 8150 4928
rect 8214 4864 8230 4928
rect 8294 4864 8300 4928
rect 7984 4863 8300 4864
rect 15574 4928 15890 4929
rect 15574 4864 15580 4928
rect 15644 4864 15660 4928
rect 15724 4864 15740 4928
rect 15804 4864 15820 4928
rect 15884 4864 15890 4928
rect 15574 4863 15890 4864
rect 23164 4928 23480 4929
rect 23164 4864 23170 4928
rect 23234 4864 23250 4928
rect 23314 4864 23330 4928
rect 23394 4864 23410 4928
rect 23474 4864 23480 4928
rect 23164 4863 23480 4864
rect 30754 4928 31070 4929
rect 30754 4864 30760 4928
rect 30824 4864 30840 4928
rect 30904 4864 30920 4928
rect 30984 4864 31000 4928
rect 31064 4864 31070 4928
rect 30754 4863 31070 4864
rect 1577 4722 1643 4725
rect 9397 4722 9463 4725
rect 1577 4720 9463 4722
rect 1577 4664 1582 4720
rect 1638 4664 9402 4720
rect 9458 4664 9463 4720
rect 1577 4662 9463 4664
rect 1577 4659 1643 4662
rect 9397 4659 9463 4662
rect 22645 4722 22711 4725
rect 25865 4722 25931 4725
rect 22645 4720 25931 4722
rect 22645 4664 22650 4720
rect 22706 4664 25870 4720
rect 25926 4664 25931 4720
rect 22645 4662 25931 4664
rect 22645 4659 22711 4662
rect 25865 4659 25931 4662
rect 3233 4586 3299 4589
rect 4061 4586 4127 4589
rect 3233 4584 4127 4586
rect 3233 4528 3238 4584
rect 3294 4528 4066 4584
rect 4122 4528 4127 4584
rect 3233 4526 4127 4528
rect 3233 4523 3299 4526
rect 4061 4523 4127 4526
rect 5441 4586 5507 4589
rect 25129 4586 25195 4589
rect 5441 4584 25195 4586
rect 5441 4528 5446 4584
rect 5502 4528 25134 4584
rect 25190 4528 25195 4584
rect 5441 4526 25195 4528
rect 5441 4523 5507 4526
rect 25129 4523 25195 4526
rect 4189 4384 4505 4385
rect 4189 4320 4195 4384
rect 4259 4320 4275 4384
rect 4339 4320 4355 4384
rect 4419 4320 4435 4384
rect 4499 4320 4505 4384
rect 4189 4319 4505 4320
rect 11779 4384 12095 4385
rect 11779 4320 11785 4384
rect 11849 4320 11865 4384
rect 11929 4320 11945 4384
rect 12009 4320 12025 4384
rect 12089 4320 12095 4384
rect 11779 4319 12095 4320
rect 19369 4384 19685 4385
rect 19369 4320 19375 4384
rect 19439 4320 19455 4384
rect 19519 4320 19535 4384
rect 19599 4320 19615 4384
rect 19679 4320 19685 4384
rect 19369 4319 19685 4320
rect 26959 4384 27275 4385
rect 26959 4320 26965 4384
rect 27029 4320 27045 4384
rect 27109 4320 27125 4384
rect 27189 4320 27205 4384
rect 27269 4320 27275 4384
rect 26959 4319 27275 4320
rect 13905 4314 13971 4317
rect 17769 4314 17835 4317
rect 13905 4312 17835 4314
rect 13905 4256 13910 4312
rect 13966 4256 17774 4312
rect 17830 4256 17835 4312
rect 13905 4254 17835 4256
rect 13905 4251 13971 4254
rect 17769 4251 17835 4254
rect 4521 4178 4587 4181
rect 29177 4178 29243 4181
rect 4521 4176 29243 4178
rect 4521 4120 4526 4176
rect 4582 4120 29182 4176
rect 29238 4120 29243 4176
rect 4521 4118 29243 4120
rect 4521 4115 4587 4118
rect 29177 4115 29243 4118
rect 5349 4042 5415 4045
rect 8518 4042 8524 4044
rect 5349 4040 8524 4042
rect 5349 3984 5354 4040
rect 5410 3984 8524 4040
rect 5349 3982 8524 3984
rect 5349 3979 5415 3982
rect 8518 3980 8524 3982
rect 8588 3980 8594 4044
rect 13721 4042 13787 4045
rect 15469 4042 15535 4045
rect 13721 4040 15535 4042
rect 13721 3984 13726 4040
rect 13782 3984 15474 4040
rect 15530 3984 15535 4040
rect 13721 3982 15535 3984
rect 13721 3979 13787 3982
rect 15469 3979 15535 3982
rect 20713 4042 20779 4045
rect 25773 4042 25839 4045
rect 20713 4040 25839 4042
rect 20713 3984 20718 4040
rect 20774 3984 25778 4040
rect 25834 3984 25839 4040
rect 20713 3982 25839 3984
rect 20713 3979 20779 3982
rect 25773 3979 25839 3982
rect 1025 3906 1091 3909
rect 7189 3906 7255 3909
rect 1025 3904 7255 3906
rect 1025 3848 1030 3904
rect 1086 3848 7194 3904
rect 7250 3848 7255 3904
rect 1025 3846 7255 3848
rect 1025 3843 1091 3846
rect 7189 3843 7255 3846
rect 7984 3840 8300 3841
rect 7984 3776 7990 3840
rect 8054 3776 8070 3840
rect 8134 3776 8150 3840
rect 8214 3776 8230 3840
rect 8294 3776 8300 3840
rect 7984 3775 8300 3776
rect 15574 3840 15890 3841
rect 15574 3776 15580 3840
rect 15644 3776 15660 3840
rect 15724 3776 15740 3840
rect 15804 3776 15820 3840
rect 15884 3776 15890 3840
rect 15574 3775 15890 3776
rect 23164 3840 23480 3841
rect 23164 3776 23170 3840
rect 23234 3776 23250 3840
rect 23314 3776 23330 3840
rect 23394 3776 23410 3840
rect 23474 3776 23480 3840
rect 23164 3775 23480 3776
rect 30754 3840 31070 3841
rect 30754 3776 30760 3840
rect 30824 3776 30840 3840
rect 30904 3776 30920 3840
rect 30984 3776 31000 3840
rect 31064 3776 31070 3840
rect 30754 3775 31070 3776
rect 3049 3770 3115 3773
rect 4153 3770 4219 3773
rect 3049 3768 4219 3770
rect 3049 3712 3054 3768
rect 3110 3712 4158 3768
rect 4214 3712 4219 3768
rect 3049 3710 4219 3712
rect 3049 3707 3115 3710
rect 4153 3707 4219 3710
rect 23565 3770 23631 3773
rect 28349 3770 28415 3773
rect 23565 3768 28415 3770
rect 23565 3712 23570 3768
rect 23626 3712 28354 3768
rect 28410 3712 28415 3768
rect 23565 3710 28415 3712
rect 23565 3707 23631 3710
rect 28349 3707 28415 3710
rect 2037 3634 2103 3637
rect 18505 3634 18571 3637
rect 25497 3634 25563 3637
rect 2037 3632 25563 3634
rect 2037 3576 2042 3632
rect 2098 3576 18510 3632
rect 18566 3576 25502 3632
rect 25558 3576 25563 3632
rect 2037 3574 25563 3576
rect 2037 3571 2103 3574
rect 18505 3571 18571 3574
rect 25497 3571 25563 3574
rect 1761 3498 1827 3501
rect 8293 3498 8359 3501
rect 15929 3498 15995 3501
rect 1761 3496 8218 3498
rect 1761 3440 1766 3496
rect 1822 3440 8218 3496
rect 1761 3438 8218 3440
rect 1761 3435 1827 3438
rect 8158 3362 8218 3438
rect 8293 3496 15995 3498
rect 8293 3440 8298 3496
rect 8354 3440 15934 3496
rect 15990 3440 15995 3496
rect 8293 3438 15995 3440
rect 8293 3435 8359 3438
rect 15929 3435 15995 3438
rect 17217 3498 17283 3501
rect 27797 3498 27863 3501
rect 17217 3496 27863 3498
rect 17217 3440 17222 3496
rect 17278 3440 27802 3496
rect 27858 3440 27863 3496
rect 17217 3438 27863 3440
rect 17217 3435 17283 3438
rect 27797 3435 27863 3438
rect 8661 3362 8727 3365
rect 8158 3360 8727 3362
rect 8158 3304 8666 3360
rect 8722 3304 8727 3360
rect 8158 3302 8727 3304
rect 8661 3299 8727 3302
rect 4189 3296 4505 3297
rect 4189 3232 4195 3296
rect 4259 3232 4275 3296
rect 4339 3232 4355 3296
rect 4419 3232 4435 3296
rect 4499 3232 4505 3296
rect 4189 3231 4505 3232
rect 11779 3296 12095 3297
rect 11779 3232 11785 3296
rect 11849 3232 11865 3296
rect 11929 3232 11945 3296
rect 12009 3232 12025 3296
rect 12089 3232 12095 3296
rect 11779 3231 12095 3232
rect 19369 3296 19685 3297
rect 19369 3232 19375 3296
rect 19439 3232 19455 3296
rect 19519 3232 19535 3296
rect 19599 3232 19615 3296
rect 19679 3232 19685 3296
rect 19369 3231 19685 3232
rect 26959 3296 27275 3297
rect 26959 3232 26965 3296
rect 27029 3232 27045 3296
rect 27109 3232 27125 3296
rect 27189 3232 27205 3296
rect 27269 3232 27275 3296
rect 26959 3231 27275 3232
rect 7649 3226 7715 3229
rect 11145 3226 11211 3229
rect 24853 3226 24919 3229
rect 7649 3224 11211 3226
rect 7649 3168 7654 3224
rect 7710 3168 11150 3224
rect 11206 3168 11211 3224
rect 7649 3166 11211 3168
rect 7649 3163 7715 3166
rect 11145 3163 11211 3166
rect 19750 3224 24919 3226
rect 19750 3168 24858 3224
rect 24914 3168 24919 3224
rect 19750 3166 24919 3168
rect 1669 3090 1735 3093
rect 9765 3090 9831 3093
rect 1669 3088 9831 3090
rect 1669 3032 1674 3088
rect 1730 3032 9770 3088
rect 9826 3032 9831 3088
rect 1669 3030 9831 3032
rect 1669 3027 1735 3030
rect 9765 3027 9831 3030
rect 12157 3090 12223 3093
rect 17585 3090 17651 3093
rect 19750 3090 19810 3166
rect 24853 3163 24919 3166
rect 12157 3088 19810 3090
rect 12157 3032 12162 3088
rect 12218 3032 17590 3088
rect 17646 3032 19810 3088
rect 12157 3030 19810 3032
rect 20989 3090 21055 3093
rect 27613 3090 27679 3093
rect 20989 3088 27679 3090
rect 20989 3032 20994 3088
rect 21050 3032 27618 3088
rect 27674 3032 27679 3088
rect 20989 3030 27679 3032
rect 12157 3027 12223 3030
rect 17585 3027 17651 3030
rect 20989 3027 21055 3030
rect 27613 3027 27679 3030
rect 5901 2954 5967 2957
rect 16389 2954 16455 2957
rect 5901 2952 16455 2954
rect 5901 2896 5906 2952
rect 5962 2896 16394 2952
rect 16450 2896 16455 2952
rect 5901 2894 16455 2896
rect 5901 2891 5967 2894
rect 16389 2891 16455 2894
rect 20437 2954 20503 2957
rect 26785 2954 26851 2957
rect 27245 2954 27311 2957
rect 20437 2952 25928 2954
rect 20437 2896 20442 2952
rect 20498 2896 25928 2952
rect 20437 2894 25928 2896
rect 20437 2891 20503 2894
rect 1393 2818 1459 2821
rect 4153 2818 4219 2821
rect 1393 2816 4219 2818
rect 1393 2760 1398 2816
rect 1454 2760 4158 2816
rect 4214 2760 4219 2816
rect 1393 2758 4219 2760
rect 1393 2755 1459 2758
rect 4153 2755 4219 2758
rect 8661 2818 8727 2821
rect 14733 2818 14799 2821
rect 8661 2816 14799 2818
rect 8661 2760 8666 2816
rect 8722 2760 14738 2816
rect 14794 2760 14799 2816
rect 8661 2758 14799 2760
rect 8661 2755 8727 2758
rect 14733 2755 14799 2758
rect 7984 2752 8300 2753
rect 7984 2688 7990 2752
rect 8054 2688 8070 2752
rect 8134 2688 8150 2752
rect 8214 2688 8230 2752
rect 8294 2688 8300 2752
rect 7984 2687 8300 2688
rect 15574 2752 15890 2753
rect 15574 2688 15580 2752
rect 15644 2688 15660 2752
rect 15724 2688 15740 2752
rect 15804 2688 15820 2752
rect 15884 2688 15890 2752
rect 15574 2687 15890 2688
rect 23164 2752 23480 2753
rect 23164 2688 23170 2752
rect 23234 2688 23250 2752
rect 23314 2688 23330 2752
rect 23394 2688 23410 2752
rect 23474 2688 23480 2752
rect 23164 2687 23480 2688
rect 1853 2682 1919 2685
rect 3785 2682 3851 2685
rect 5073 2682 5139 2685
rect 1853 2680 5139 2682
rect 1853 2624 1858 2680
rect 1914 2624 3790 2680
rect 3846 2624 5078 2680
rect 5134 2624 5139 2680
rect 1853 2622 5139 2624
rect 1853 2619 1919 2622
rect 3785 2619 3851 2622
rect 5073 2619 5139 2622
rect 20529 2682 20595 2685
rect 21817 2682 21883 2685
rect 24945 2682 25011 2685
rect 20529 2680 21883 2682
rect 20529 2624 20534 2680
rect 20590 2624 21822 2680
rect 21878 2624 21883 2680
rect 20529 2622 21883 2624
rect 20529 2619 20595 2622
rect 21817 2619 21883 2622
rect 23568 2680 25011 2682
rect 23568 2624 24950 2680
rect 25006 2624 25011 2680
rect 23568 2622 25011 2624
rect 25868 2682 25928 2894
rect 26785 2952 27311 2954
rect 26785 2896 26790 2952
rect 26846 2896 27250 2952
rect 27306 2896 27311 2952
rect 26785 2894 27311 2896
rect 26785 2891 26851 2894
rect 27245 2891 27311 2894
rect 26049 2818 26115 2821
rect 26969 2818 27035 2821
rect 26049 2816 27035 2818
rect 26049 2760 26054 2816
rect 26110 2760 26974 2816
rect 27030 2760 27035 2816
rect 26049 2758 27035 2760
rect 26049 2755 26115 2758
rect 26969 2755 27035 2758
rect 30754 2752 31070 2753
rect 30754 2688 30760 2752
rect 30824 2688 30840 2752
rect 30904 2688 30920 2752
rect 30984 2688 31000 2752
rect 31064 2688 31070 2752
rect 30754 2687 31070 2688
rect 26785 2682 26851 2685
rect 25868 2680 26851 2682
rect 25868 2624 26790 2680
rect 26846 2624 26851 2680
rect 25868 2622 26851 2624
rect 9489 2546 9555 2549
rect 23568 2546 23628 2622
rect 24945 2619 25011 2622
rect 26785 2619 26851 2622
rect 24669 2546 24735 2549
rect 9489 2544 23628 2546
rect 9489 2488 9494 2544
rect 9550 2488 23628 2544
rect 9489 2486 23628 2488
rect 23798 2544 24735 2546
rect 23798 2488 24674 2544
rect 24730 2488 24735 2544
rect 23798 2486 24735 2488
rect 9489 2483 9555 2486
rect 3233 2410 3299 2413
rect 3969 2410 4035 2413
rect 6545 2410 6611 2413
rect 23798 2410 23858 2486
rect 24669 2483 24735 2486
rect 3233 2408 4722 2410
rect 3233 2352 3238 2408
rect 3294 2352 3974 2408
rect 4030 2352 4722 2408
rect 3233 2350 4722 2352
rect 3233 2347 3299 2350
rect 3969 2347 4035 2350
rect 4662 2274 4722 2350
rect 6545 2408 23858 2410
rect 6545 2352 6550 2408
rect 6606 2352 23858 2408
rect 6545 2350 23858 2352
rect 24393 2410 24459 2413
rect 24853 2410 24919 2413
rect 24393 2408 24919 2410
rect 24393 2352 24398 2408
rect 24454 2352 24858 2408
rect 24914 2352 24919 2408
rect 24393 2350 24919 2352
rect 6545 2347 6611 2350
rect 24393 2347 24459 2350
rect 24853 2347 24919 2350
rect 9489 2274 9555 2277
rect 4662 2272 9555 2274
rect 4662 2216 9494 2272
rect 9550 2216 9555 2272
rect 4662 2214 9555 2216
rect 9489 2211 9555 2214
rect 16757 2274 16823 2277
rect 19241 2274 19307 2277
rect 16757 2272 19307 2274
rect 16757 2216 16762 2272
rect 16818 2216 19246 2272
rect 19302 2216 19307 2272
rect 16757 2214 19307 2216
rect 16757 2211 16823 2214
rect 19241 2211 19307 2214
rect 21081 2274 21147 2277
rect 26233 2274 26299 2277
rect 21081 2272 26299 2274
rect 21081 2216 21086 2272
rect 21142 2216 26238 2272
rect 26294 2216 26299 2272
rect 21081 2214 26299 2216
rect 21081 2211 21147 2214
rect 26233 2211 26299 2214
rect 4189 2208 4505 2209
rect 4189 2144 4195 2208
rect 4259 2144 4275 2208
rect 4339 2144 4355 2208
rect 4419 2144 4435 2208
rect 4499 2144 4505 2208
rect 4189 2143 4505 2144
rect 11779 2208 12095 2209
rect 11779 2144 11785 2208
rect 11849 2144 11865 2208
rect 11929 2144 11945 2208
rect 12009 2144 12025 2208
rect 12089 2144 12095 2208
rect 11779 2143 12095 2144
rect 19369 2208 19685 2209
rect 19369 2144 19375 2208
rect 19439 2144 19455 2208
rect 19519 2144 19535 2208
rect 19599 2144 19615 2208
rect 19679 2144 19685 2208
rect 19369 2143 19685 2144
rect 26959 2208 27275 2209
rect 26959 2144 26965 2208
rect 27029 2144 27045 2208
rect 27109 2144 27125 2208
rect 27189 2144 27205 2208
rect 27269 2144 27275 2208
rect 26959 2143 27275 2144
rect 9489 2140 9555 2141
rect 9438 2138 9444 2140
rect 9398 2078 9444 2138
rect 9508 2136 9555 2140
rect 9550 2080 9555 2136
rect 9438 2076 9444 2078
rect 9508 2076 9555 2080
rect 9489 2075 9555 2076
rect 21633 2138 21699 2141
rect 26417 2138 26483 2141
rect 26785 2138 26851 2141
rect 21633 2136 26851 2138
rect 21633 2080 21638 2136
rect 21694 2080 26422 2136
rect 26478 2080 26790 2136
rect 26846 2080 26851 2136
rect 21633 2078 26851 2080
rect 21633 2075 21699 2078
rect 26417 2075 26483 2078
rect 26785 2075 26851 2078
rect 2037 2002 2103 2005
rect 4521 2002 4587 2005
rect 2037 2000 4587 2002
rect 2037 1944 2042 2000
rect 2098 1944 4526 2000
rect 4582 1944 4587 2000
rect 2037 1942 4587 1944
rect 2037 1939 2103 1942
rect 4521 1939 4587 1942
rect 11237 2002 11303 2005
rect 11973 2002 12039 2005
rect 11237 2000 12039 2002
rect 11237 1944 11242 2000
rect 11298 1944 11978 2000
rect 12034 1944 12039 2000
rect 11237 1942 12039 1944
rect 11237 1939 11303 1942
rect 11973 1939 12039 1942
rect 15009 2002 15075 2005
rect 26693 2002 26759 2005
rect 15009 2000 26759 2002
rect 15009 1944 15014 2000
rect 15070 1944 26698 2000
rect 26754 1944 26759 2000
rect 15009 1942 26759 1944
rect 15009 1939 15075 1942
rect 26693 1939 26759 1942
rect 6269 1866 6335 1869
rect 10685 1866 10751 1869
rect 6269 1864 10751 1866
rect 6269 1808 6274 1864
rect 6330 1808 10690 1864
rect 10746 1808 10751 1864
rect 6269 1806 10751 1808
rect 6269 1803 6335 1806
rect 10685 1803 10751 1806
rect 12341 1866 12407 1869
rect 23565 1866 23631 1869
rect 12341 1864 23631 1866
rect 12341 1808 12346 1864
rect 12402 1808 23570 1864
rect 23626 1808 23631 1864
rect 12341 1806 23631 1808
rect 12341 1803 12407 1806
rect 23565 1803 23631 1806
rect 23749 1866 23815 1869
rect 28993 1866 29059 1869
rect 23749 1864 29059 1866
rect 23749 1808 23754 1864
rect 23810 1808 28998 1864
rect 29054 1808 29059 1864
rect 23749 1806 29059 1808
rect 23749 1803 23815 1806
rect 28993 1803 29059 1806
rect 20529 1730 20595 1733
rect 22921 1730 22987 1733
rect 20529 1728 22987 1730
rect 20529 1672 20534 1728
rect 20590 1672 22926 1728
rect 22982 1672 22987 1728
rect 20529 1670 22987 1672
rect 20529 1667 20595 1670
rect 22921 1667 22987 1670
rect 23749 1730 23815 1733
rect 26417 1730 26483 1733
rect 23749 1728 26483 1730
rect 23749 1672 23754 1728
rect 23810 1672 26422 1728
rect 26478 1672 26483 1728
rect 23749 1670 26483 1672
rect 23749 1667 23815 1670
rect 26417 1667 26483 1670
rect 7984 1664 8300 1665
rect 7984 1600 7990 1664
rect 8054 1600 8070 1664
rect 8134 1600 8150 1664
rect 8214 1600 8230 1664
rect 8294 1600 8300 1664
rect 7984 1599 8300 1600
rect 15574 1664 15890 1665
rect 15574 1600 15580 1664
rect 15644 1600 15660 1664
rect 15724 1600 15740 1664
rect 15804 1600 15820 1664
rect 15884 1600 15890 1664
rect 15574 1599 15890 1600
rect 23164 1664 23480 1665
rect 23164 1600 23170 1664
rect 23234 1600 23250 1664
rect 23314 1600 23330 1664
rect 23394 1600 23410 1664
rect 23474 1600 23480 1664
rect 23164 1599 23480 1600
rect 30754 1664 31070 1665
rect 30754 1600 30760 1664
rect 30824 1600 30840 1664
rect 30904 1600 30920 1664
rect 30984 1600 31000 1664
rect 31064 1600 31070 1664
rect 30754 1599 31070 1600
rect 3049 1594 3115 1597
rect 6637 1594 6703 1597
rect 3049 1592 6703 1594
rect 3049 1536 3054 1592
rect 3110 1536 6642 1592
rect 6698 1536 6703 1592
rect 3049 1534 6703 1536
rect 3049 1531 3115 1534
rect 6637 1531 6703 1534
rect 10593 1594 10659 1597
rect 11973 1594 12039 1597
rect 10593 1592 12039 1594
rect 10593 1536 10598 1592
rect 10654 1536 11978 1592
rect 12034 1536 12039 1592
rect 10593 1534 12039 1536
rect 10593 1531 10659 1534
rect 11973 1531 12039 1534
rect 16297 1594 16363 1597
rect 17401 1594 17467 1597
rect 20989 1594 21055 1597
rect 22645 1594 22711 1597
rect 24669 1594 24735 1597
rect 16297 1592 22711 1594
rect 16297 1536 16302 1592
rect 16358 1536 17406 1592
rect 17462 1536 20994 1592
rect 21050 1536 22650 1592
rect 22706 1536 22711 1592
rect 16297 1534 22711 1536
rect 16297 1531 16363 1534
rect 17401 1531 17467 1534
rect 20989 1531 21055 1534
rect 22645 1531 22711 1534
rect 23568 1592 24735 1594
rect 23568 1536 24674 1592
rect 24730 1536 24735 1592
rect 23568 1534 24735 1536
rect 4521 1458 4587 1461
rect 11329 1458 11395 1461
rect 4521 1456 11395 1458
rect 4521 1400 4526 1456
rect 4582 1400 11334 1456
rect 11390 1400 11395 1456
rect 4521 1398 11395 1400
rect 4521 1395 4587 1398
rect 11329 1395 11395 1398
rect 16205 1458 16271 1461
rect 23568 1458 23628 1534
rect 24669 1531 24735 1534
rect 16205 1456 23628 1458
rect 16205 1400 16210 1456
rect 16266 1400 23628 1456
rect 16205 1398 23628 1400
rect 26693 1458 26759 1461
rect 28625 1458 28691 1461
rect 30465 1458 30531 1461
rect 26693 1456 30531 1458
rect 26693 1400 26698 1456
rect 26754 1400 28630 1456
rect 28686 1400 30470 1456
rect 30526 1400 30531 1456
rect 26693 1398 30531 1400
rect 16205 1395 16271 1398
rect 26693 1395 26759 1398
rect 28625 1395 28691 1398
rect 30465 1395 30531 1398
rect 4245 1322 4311 1325
rect 28717 1322 28783 1325
rect 4245 1320 28783 1322
rect 4245 1264 4250 1320
rect 4306 1264 28722 1320
rect 28778 1264 28783 1320
rect 4245 1262 28783 1264
rect 4245 1259 4311 1262
rect 28717 1259 28783 1262
rect 5625 1186 5691 1189
rect 9397 1186 9463 1189
rect 5625 1184 9463 1186
rect 5625 1128 5630 1184
rect 5686 1128 9402 1184
rect 9458 1128 9463 1184
rect 5625 1126 9463 1128
rect 5625 1123 5691 1126
rect 9397 1123 9463 1126
rect 23473 1186 23539 1189
rect 26049 1186 26115 1189
rect 23473 1184 26115 1186
rect 23473 1128 23478 1184
rect 23534 1128 26054 1184
rect 26110 1128 26115 1184
rect 23473 1126 26115 1128
rect 23473 1123 23539 1126
rect 26049 1123 26115 1126
rect 4189 1120 4505 1121
rect 4189 1056 4195 1120
rect 4259 1056 4275 1120
rect 4339 1056 4355 1120
rect 4419 1056 4435 1120
rect 4499 1056 4505 1120
rect 4189 1055 4505 1056
rect 11779 1120 12095 1121
rect 11779 1056 11785 1120
rect 11849 1056 11865 1120
rect 11929 1056 11945 1120
rect 12009 1056 12025 1120
rect 12089 1056 12095 1120
rect 11779 1055 12095 1056
rect 19369 1120 19685 1121
rect 19369 1056 19375 1120
rect 19439 1056 19455 1120
rect 19519 1056 19535 1120
rect 19599 1056 19615 1120
rect 19679 1056 19685 1120
rect 19369 1055 19685 1056
rect 26959 1120 27275 1121
rect 26959 1056 26965 1120
rect 27029 1056 27045 1120
rect 27109 1056 27125 1120
rect 27189 1056 27205 1120
rect 27269 1056 27275 1120
rect 26959 1055 27275 1056
rect 21541 1050 21607 1053
rect 24945 1050 25011 1053
rect 21541 1048 25011 1050
rect 21541 992 21546 1048
rect 21602 992 24950 1048
rect 25006 992 25011 1048
rect 21541 990 25011 992
rect 21541 987 21607 990
rect 24945 987 25011 990
rect 12065 914 12131 917
rect 23657 914 23723 917
rect 12065 912 23723 914
rect 12065 856 12070 912
rect 12126 856 23662 912
rect 23718 856 23723 912
rect 12065 854 23723 856
rect 12065 851 12131 854
rect 23657 851 23723 854
rect 4981 778 5047 781
rect 29269 778 29335 781
rect 4981 776 29335 778
rect 4981 720 4986 776
rect 5042 720 29274 776
rect 29330 720 29335 776
rect 4981 718 29335 720
rect 4981 715 5047 718
rect 29269 715 29335 718
rect 12157 642 12223 645
rect 14457 642 14523 645
rect 12157 640 14523 642
rect 12157 584 12162 640
rect 12218 584 14462 640
rect 14518 584 14523 640
rect 12157 582 14523 584
rect 12157 579 12223 582
rect 14457 579 14523 582
rect 16481 642 16547 645
rect 18873 642 18939 645
rect 16481 640 18939 642
rect 16481 584 16486 640
rect 16542 584 18878 640
rect 18934 584 18939 640
rect 16481 582 18939 584
rect 16481 579 16547 582
rect 18873 579 18939 582
rect 7984 576 8300 577
rect 7984 512 7990 576
rect 8054 512 8070 576
rect 8134 512 8150 576
rect 8214 512 8230 576
rect 8294 512 8300 576
rect 7984 511 8300 512
rect 15574 576 15890 577
rect 15574 512 15580 576
rect 15644 512 15660 576
rect 15724 512 15740 576
rect 15804 512 15820 576
rect 15884 512 15890 576
rect 15574 511 15890 512
rect 23164 576 23480 577
rect 23164 512 23170 576
rect 23234 512 23250 576
rect 23314 512 23330 576
rect 23394 512 23410 576
rect 23474 512 23480 576
rect 23164 511 23480 512
rect 30754 576 31070 577
rect 30754 512 30760 576
rect 30824 512 30840 576
rect 30904 512 30920 576
rect 30984 512 31000 576
rect 31064 512 31070 576
rect 30754 511 31070 512
rect 20805 506 20871 509
rect 16622 504 20871 506
rect 16622 448 20810 504
rect 20866 448 20871 504
rect 16622 446 20871 448
rect 6913 370 6979 373
rect 16622 370 16682 446
rect 20805 443 20871 446
rect 6913 368 16682 370
rect 6913 312 6918 368
rect 6974 312 16682 368
rect 6913 310 16682 312
rect 20713 370 20779 373
rect 29361 370 29427 373
rect 20713 368 29427 370
rect 20713 312 20718 368
rect 20774 312 29366 368
rect 29422 312 29427 368
rect 20713 310 29427 312
rect 6913 307 6979 310
rect 20713 307 20779 310
rect 29361 307 29427 310
rect 6269 234 6335 237
rect 25681 234 25747 237
rect 6269 232 25747 234
rect 6269 176 6274 232
rect 6330 176 25686 232
rect 25742 176 25747 232
rect 6269 174 25747 176
rect 6269 171 6335 174
rect 25681 171 25747 174
rect 3785 98 3851 101
rect 18229 98 18295 101
rect 3785 96 18295 98
rect 3785 40 3790 96
rect 3846 40 18234 96
rect 18290 40 18295 96
rect 3785 38 18295 40
rect 3785 35 3851 38
rect 18229 35 18295 38
rect 18873 98 18939 101
rect 28073 98 28139 101
rect 18873 96 28139 98
rect 18873 40 18878 96
rect 18934 40 28078 96
rect 28134 40 28139 96
rect 18873 38 28139 40
rect 18873 35 18939 38
rect 28073 35 28139 38
<< via3 >>
rect 8892 22264 8956 22268
rect 8892 22208 8906 22264
rect 8906 22208 8956 22264
rect 8892 22204 8956 22208
rect 9628 22264 9692 22268
rect 9628 22208 9678 22264
rect 9678 22208 9692 22264
rect 9628 22204 9692 22208
rect 6868 22068 6932 22132
rect 25452 22068 25516 22132
rect 12388 21992 12452 21996
rect 12388 21936 12438 21992
rect 12438 21936 12452 21992
rect 12388 21932 12452 21936
rect 21956 21932 22020 21996
rect 23612 21992 23676 21996
rect 23612 21936 23626 21992
rect 23626 21936 23676 21992
rect 23612 21932 23676 21936
rect 4195 21788 4259 21792
rect 4195 21732 4199 21788
rect 4199 21732 4255 21788
rect 4255 21732 4259 21788
rect 4195 21728 4259 21732
rect 4275 21788 4339 21792
rect 4275 21732 4279 21788
rect 4279 21732 4335 21788
rect 4335 21732 4339 21788
rect 4275 21728 4339 21732
rect 4355 21788 4419 21792
rect 4355 21732 4359 21788
rect 4359 21732 4415 21788
rect 4415 21732 4419 21788
rect 4355 21728 4419 21732
rect 4435 21788 4499 21792
rect 4435 21732 4439 21788
rect 4439 21732 4495 21788
rect 4495 21732 4499 21788
rect 4435 21728 4499 21732
rect 11785 21788 11849 21792
rect 11785 21732 11789 21788
rect 11789 21732 11845 21788
rect 11845 21732 11849 21788
rect 11785 21728 11849 21732
rect 11865 21788 11929 21792
rect 11865 21732 11869 21788
rect 11869 21732 11925 21788
rect 11925 21732 11929 21788
rect 11865 21728 11929 21732
rect 11945 21788 12009 21792
rect 11945 21732 11949 21788
rect 11949 21732 12005 21788
rect 12005 21732 12009 21788
rect 11945 21728 12009 21732
rect 12025 21788 12089 21792
rect 12025 21732 12029 21788
rect 12029 21732 12085 21788
rect 12085 21732 12089 21788
rect 12025 21728 12089 21732
rect 19375 21788 19439 21792
rect 19375 21732 19379 21788
rect 19379 21732 19435 21788
rect 19435 21732 19439 21788
rect 19375 21728 19439 21732
rect 19455 21788 19519 21792
rect 19455 21732 19459 21788
rect 19459 21732 19515 21788
rect 19515 21732 19519 21788
rect 19455 21728 19519 21732
rect 19535 21788 19599 21792
rect 19535 21732 19539 21788
rect 19539 21732 19595 21788
rect 19595 21732 19599 21788
rect 19535 21728 19599 21732
rect 19615 21788 19679 21792
rect 19615 21732 19619 21788
rect 19619 21732 19675 21788
rect 19675 21732 19679 21788
rect 19615 21728 19679 21732
rect 26965 21788 27029 21792
rect 26965 21732 26969 21788
rect 26969 21732 27025 21788
rect 27025 21732 27029 21788
rect 26965 21728 27029 21732
rect 27045 21788 27109 21792
rect 27045 21732 27049 21788
rect 27049 21732 27105 21788
rect 27105 21732 27109 21788
rect 27045 21728 27109 21732
rect 27125 21788 27189 21792
rect 27125 21732 27129 21788
rect 27129 21732 27185 21788
rect 27185 21732 27189 21788
rect 27125 21728 27189 21732
rect 27205 21788 27269 21792
rect 27205 21732 27209 21788
rect 27209 21732 27265 21788
rect 27265 21732 27269 21788
rect 27205 21728 27269 21732
rect 11100 21524 11164 21588
rect 13124 21524 13188 21588
rect 16988 21524 17052 21588
rect 24900 21388 24964 21452
rect 7990 21244 8054 21248
rect 7990 21188 7994 21244
rect 7994 21188 8050 21244
rect 8050 21188 8054 21244
rect 7990 21184 8054 21188
rect 8070 21244 8134 21248
rect 8070 21188 8074 21244
rect 8074 21188 8130 21244
rect 8130 21188 8134 21244
rect 8070 21184 8134 21188
rect 8150 21244 8214 21248
rect 8150 21188 8154 21244
rect 8154 21188 8210 21244
rect 8210 21188 8214 21244
rect 8150 21184 8214 21188
rect 8230 21244 8294 21248
rect 8230 21188 8234 21244
rect 8234 21188 8290 21244
rect 8290 21188 8294 21244
rect 8230 21184 8294 21188
rect 15580 21244 15644 21248
rect 15580 21188 15584 21244
rect 15584 21188 15640 21244
rect 15640 21188 15644 21244
rect 15580 21184 15644 21188
rect 15660 21244 15724 21248
rect 15660 21188 15664 21244
rect 15664 21188 15720 21244
rect 15720 21188 15724 21244
rect 15660 21184 15724 21188
rect 15740 21244 15804 21248
rect 15740 21188 15744 21244
rect 15744 21188 15800 21244
rect 15800 21188 15804 21244
rect 15740 21184 15804 21188
rect 15820 21244 15884 21248
rect 15820 21188 15824 21244
rect 15824 21188 15880 21244
rect 15880 21188 15884 21244
rect 15820 21184 15884 21188
rect 23170 21244 23234 21248
rect 23170 21188 23174 21244
rect 23174 21188 23230 21244
rect 23230 21188 23234 21244
rect 23170 21184 23234 21188
rect 23250 21244 23314 21248
rect 23250 21188 23254 21244
rect 23254 21188 23310 21244
rect 23310 21188 23314 21244
rect 23250 21184 23314 21188
rect 23330 21244 23394 21248
rect 23330 21188 23334 21244
rect 23334 21188 23390 21244
rect 23390 21188 23394 21244
rect 23330 21184 23394 21188
rect 23410 21244 23474 21248
rect 23410 21188 23414 21244
rect 23414 21188 23470 21244
rect 23470 21188 23474 21244
rect 23410 21184 23474 21188
rect 30760 21244 30824 21248
rect 30760 21188 30764 21244
rect 30764 21188 30820 21244
rect 30820 21188 30824 21244
rect 30760 21184 30824 21188
rect 30840 21244 30904 21248
rect 30840 21188 30844 21244
rect 30844 21188 30900 21244
rect 30900 21188 30904 21244
rect 30840 21184 30904 21188
rect 30920 21244 30984 21248
rect 30920 21188 30924 21244
rect 30924 21188 30980 21244
rect 30980 21188 30984 21244
rect 30920 21184 30984 21188
rect 31000 21244 31064 21248
rect 31000 21188 31004 21244
rect 31004 21188 31060 21244
rect 31060 21188 31064 21244
rect 31000 21184 31064 21188
rect 26372 21116 26436 21180
rect 22876 20904 22940 20908
rect 22876 20848 22926 20904
rect 22926 20848 22940 20904
rect 22876 20844 22940 20848
rect 22508 20708 22572 20772
rect 24164 20708 24228 20772
rect 4195 20700 4259 20704
rect 4195 20644 4199 20700
rect 4199 20644 4255 20700
rect 4255 20644 4259 20700
rect 4195 20640 4259 20644
rect 4275 20700 4339 20704
rect 4275 20644 4279 20700
rect 4279 20644 4335 20700
rect 4335 20644 4339 20700
rect 4275 20640 4339 20644
rect 4355 20700 4419 20704
rect 4355 20644 4359 20700
rect 4359 20644 4415 20700
rect 4415 20644 4419 20700
rect 4355 20640 4419 20644
rect 4435 20700 4499 20704
rect 4435 20644 4439 20700
rect 4439 20644 4495 20700
rect 4495 20644 4499 20700
rect 4435 20640 4499 20644
rect 11785 20700 11849 20704
rect 11785 20644 11789 20700
rect 11789 20644 11845 20700
rect 11845 20644 11849 20700
rect 11785 20640 11849 20644
rect 11865 20700 11929 20704
rect 11865 20644 11869 20700
rect 11869 20644 11925 20700
rect 11925 20644 11929 20700
rect 11865 20640 11929 20644
rect 11945 20700 12009 20704
rect 11945 20644 11949 20700
rect 11949 20644 12005 20700
rect 12005 20644 12009 20700
rect 11945 20640 12009 20644
rect 12025 20700 12089 20704
rect 12025 20644 12029 20700
rect 12029 20644 12085 20700
rect 12085 20644 12089 20700
rect 12025 20640 12089 20644
rect 19375 20700 19439 20704
rect 19375 20644 19379 20700
rect 19379 20644 19435 20700
rect 19435 20644 19439 20700
rect 19375 20640 19439 20644
rect 19455 20700 19519 20704
rect 19455 20644 19459 20700
rect 19459 20644 19515 20700
rect 19515 20644 19519 20700
rect 19455 20640 19519 20644
rect 19535 20700 19599 20704
rect 19535 20644 19539 20700
rect 19539 20644 19595 20700
rect 19595 20644 19599 20700
rect 19535 20640 19599 20644
rect 19615 20700 19679 20704
rect 19615 20644 19619 20700
rect 19619 20644 19675 20700
rect 19675 20644 19679 20700
rect 19615 20640 19679 20644
rect 26965 20700 27029 20704
rect 26965 20644 26969 20700
rect 26969 20644 27025 20700
rect 27025 20644 27029 20700
rect 26965 20640 27029 20644
rect 27045 20700 27109 20704
rect 27045 20644 27049 20700
rect 27049 20644 27105 20700
rect 27105 20644 27109 20700
rect 27045 20640 27109 20644
rect 27125 20700 27189 20704
rect 27125 20644 27129 20700
rect 27129 20644 27185 20700
rect 27185 20644 27189 20700
rect 27125 20640 27189 20644
rect 27205 20700 27269 20704
rect 27205 20644 27209 20700
rect 27209 20644 27265 20700
rect 27265 20644 27269 20700
rect 27205 20640 27269 20644
rect 10364 20632 10428 20636
rect 10364 20576 10378 20632
rect 10378 20576 10428 20632
rect 10364 20572 10428 20576
rect 8892 20436 8956 20500
rect 10916 20436 10980 20500
rect 13676 20436 13740 20500
rect 16068 20496 16132 20500
rect 16068 20440 16118 20496
rect 16118 20440 16132 20496
rect 16068 20436 16132 20440
rect 14596 20360 14660 20364
rect 14596 20304 14610 20360
rect 14610 20304 14660 20360
rect 14596 20300 14660 20304
rect 7990 20156 8054 20160
rect 7990 20100 7994 20156
rect 7994 20100 8050 20156
rect 8050 20100 8054 20156
rect 7990 20096 8054 20100
rect 8070 20156 8134 20160
rect 8070 20100 8074 20156
rect 8074 20100 8130 20156
rect 8130 20100 8134 20156
rect 8070 20096 8134 20100
rect 8150 20156 8214 20160
rect 8150 20100 8154 20156
rect 8154 20100 8210 20156
rect 8210 20100 8214 20156
rect 8150 20096 8214 20100
rect 8230 20156 8294 20160
rect 8230 20100 8234 20156
rect 8234 20100 8290 20156
rect 8290 20100 8294 20156
rect 8230 20096 8294 20100
rect 15580 20156 15644 20160
rect 15580 20100 15584 20156
rect 15584 20100 15640 20156
rect 15640 20100 15644 20156
rect 15580 20096 15644 20100
rect 15660 20156 15724 20160
rect 15660 20100 15664 20156
rect 15664 20100 15720 20156
rect 15720 20100 15724 20156
rect 15660 20096 15724 20100
rect 15740 20156 15804 20160
rect 15740 20100 15744 20156
rect 15744 20100 15800 20156
rect 15800 20100 15804 20156
rect 15740 20096 15804 20100
rect 15820 20156 15884 20160
rect 15820 20100 15824 20156
rect 15824 20100 15880 20156
rect 15880 20100 15884 20156
rect 15820 20096 15884 20100
rect 23170 20156 23234 20160
rect 23170 20100 23174 20156
rect 23174 20100 23230 20156
rect 23230 20100 23234 20156
rect 23170 20096 23234 20100
rect 23250 20156 23314 20160
rect 23250 20100 23254 20156
rect 23254 20100 23310 20156
rect 23310 20100 23314 20156
rect 23250 20096 23314 20100
rect 23330 20156 23394 20160
rect 23330 20100 23334 20156
rect 23334 20100 23390 20156
rect 23390 20100 23394 20156
rect 23330 20096 23394 20100
rect 23410 20156 23474 20160
rect 23410 20100 23414 20156
rect 23414 20100 23470 20156
rect 23470 20100 23474 20156
rect 23410 20096 23474 20100
rect 30760 20156 30824 20160
rect 30760 20100 30764 20156
rect 30764 20100 30820 20156
rect 30820 20100 30824 20156
rect 30760 20096 30824 20100
rect 30840 20156 30904 20160
rect 30840 20100 30844 20156
rect 30844 20100 30900 20156
rect 30900 20100 30904 20156
rect 30840 20096 30904 20100
rect 30920 20156 30984 20160
rect 30920 20100 30924 20156
rect 30924 20100 30980 20156
rect 30980 20100 30984 20156
rect 30920 20096 30984 20100
rect 31000 20156 31064 20160
rect 31000 20100 31004 20156
rect 31004 20100 31060 20156
rect 31060 20100 31064 20156
rect 31000 20096 31064 20100
rect 9444 19756 9508 19820
rect 4195 19612 4259 19616
rect 4195 19556 4199 19612
rect 4199 19556 4255 19612
rect 4255 19556 4259 19612
rect 4195 19552 4259 19556
rect 4275 19612 4339 19616
rect 4275 19556 4279 19612
rect 4279 19556 4335 19612
rect 4335 19556 4339 19612
rect 4275 19552 4339 19556
rect 4355 19612 4419 19616
rect 4355 19556 4359 19612
rect 4359 19556 4415 19612
rect 4415 19556 4419 19612
rect 4355 19552 4419 19556
rect 4435 19612 4499 19616
rect 4435 19556 4439 19612
rect 4439 19556 4495 19612
rect 4495 19556 4499 19612
rect 4435 19552 4499 19556
rect 2084 19348 2148 19412
rect 6868 19348 6932 19412
rect 11785 19612 11849 19616
rect 11785 19556 11789 19612
rect 11789 19556 11845 19612
rect 11845 19556 11849 19612
rect 11785 19552 11849 19556
rect 11865 19612 11929 19616
rect 11865 19556 11869 19612
rect 11869 19556 11925 19612
rect 11925 19556 11929 19612
rect 11865 19552 11929 19556
rect 11945 19612 12009 19616
rect 11945 19556 11949 19612
rect 11949 19556 12005 19612
rect 12005 19556 12009 19612
rect 11945 19552 12009 19556
rect 12025 19612 12089 19616
rect 12025 19556 12029 19612
rect 12029 19556 12085 19612
rect 12085 19556 12089 19612
rect 12025 19552 12089 19556
rect 19375 19612 19439 19616
rect 19375 19556 19379 19612
rect 19379 19556 19435 19612
rect 19435 19556 19439 19612
rect 19375 19552 19439 19556
rect 19455 19612 19519 19616
rect 19455 19556 19459 19612
rect 19459 19556 19515 19612
rect 19515 19556 19519 19612
rect 19455 19552 19519 19556
rect 19535 19612 19599 19616
rect 19535 19556 19539 19612
rect 19539 19556 19595 19612
rect 19595 19556 19599 19612
rect 19535 19552 19599 19556
rect 19615 19612 19679 19616
rect 19615 19556 19619 19612
rect 19619 19556 19675 19612
rect 19675 19556 19679 19612
rect 19615 19552 19679 19556
rect 26965 19612 27029 19616
rect 26965 19556 26969 19612
rect 26969 19556 27025 19612
rect 27025 19556 27029 19612
rect 26965 19552 27029 19556
rect 27045 19612 27109 19616
rect 27045 19556 27049 19612
rect 27049 19556 27105 19612
rect 27105 19556 27109 19612
rect 27045 19552 27109 19556
rect 27125 19612 27189 19616
rect 27125 19556 27129 19612
rect 27129 19556 27185 19612
rect 27185 19556 27189 19612
rect 27125 19552 27189 19556
rect 27205 19612 27269 19616
rect 27205 19556 27209 19612
rect 27209 19556 27265 19612
rect 27265 19556 27269 19612
rect 27205 19552 27269 19556
rect 7052 19212 7116 19276
rect 11468 19212 11532 19276
rect 14228 19212 14292 19276
rect 16436 19272 16500 19276
rect 16436 19216 16450 19272
rect 16450 19216 16500 19272
rect 16436 19212 16500 19216
rect 15332 19136 15396 19140
rect 15332 19080 15382 19136
rect 15382 19080 15396 19136
rect 15332 19076 15396 19080
rect 7990 19068 8054 19072
rect 7990 19012 7994 19068
rect 7994 19012 8050 19068
rect 8050 19012 8054 19068
rect 7990 19008 8054 19012
rect 8070 19068 8134 19072
rect 8070 19012 8074 19068
rect 8074 19012 8130 19068
rect 8130 19012 8134 19068
rect 8070 19008 8134 19012
rect 8150 19068 8214 19072
rect 8150 19012 8154 19068
rect 8154 19012 8210 19068
rect 8210 19012 8214 19068
rect 8150 19008 8214 19012
rect 8230 19068 8294 19072
rect 8230 19012 8234 19068
rect 8234 19012 8290 19068
rect 8290 19012 8294 19068
rect 8230 19008 8294 19012
rect 15580 19068 15644 19072
rect 15580 19012 15584 19068
rect 15584 19012 15640 19068
rect 15640 19012 15644 19068
rect 15580 19008 15644 19012
rect 15660 19068 15724 19072
rect 15660 19012 15664 19068
rect 15664 19012 15720 19068
rect 15720 19012 15724 19068
rect 15660 19008 15724 19012
rect 15740 19068 15804 19072
rect 15740 19012 15744 19068
rect 15744 19012 15800 19068
rect 15800 19012 15804 19068
rect 15740 19008 15804 19012
rect 15820 19068 15884 19072
rect 15820 19012 15824 19068
rect 15824 19012 15880 19068
rect 15880 19012 15884 19068
rect 15820 19008 15884 19012
rect 23170 19068 23234 19072
rect 23170 19012 23174 19068
rect 23174 19012 23230 19068
rect 23230 19012 23234 19068
rect 23170 19008 23234 19012
rect 23250 19068 23314 19072
rect 23250 19012 23254 19068
rect 23254 19012 23310 19068
rect 23310 19012 23314 19068
rect 23250 19008 23314 19012
rect 23330 19068 23394 19072
rect 23330 19012 23334 19068
rect 23334 19012 23390 19068
rect 23390 19012 23394 19068
rect 23330 19008 23394 19012
rect 23410 19068 23474 19072
rect 23410 19012 23414 19068
rect 23414 19012 23470 19068
rect 23470 19012 23474 19068
rect 23410 19008 23474 19012
rect 30760 19068 30824 19072
rect 30760 19012 30764 19068
rect 30764 19012 30820 19068
rect 30820 19012 30824 19068
rect 30760 19008 30824 19012
rect 30840 19068 30904 19072
rect 30840 19012 30844 19068
rect 30844 19012 30900 19068
rect 30900 19012 30904 19068
rect 30840 19008 30904 19012
rect 30920 19068 30984 19072
rect 30920 19012 30924 19068
rect 30924 19012 30980 19068
rect 30980 19012 30984 19068
rect 30920 19008 30984 19012
rect 31000 19068 31064 19072
rect 31000 19012 31004 19068
rect 31004 19012 31060 19068
rect 31060 19012 31064 19068
rect 31000 19008 31064 19012
rect 5028 18940 5092 19004
rect 7604 18804 7668 18868
rect 7788 18668 7852 18732
rect 4195 18524 4259 18528
rect 4195 18468 4199 18524
rect 4199 18468 4255 18524
rect 4255 18468 4259 18524
rect 4195 18464 4259 18468
rect 4275 18524 4339 18528
rect 4275 18468 4279 18524
rect 4279 18468 4335 18524
rect 4335 18468 4339 18524
rect 4275 18464 4339 18468
rect 4355 18524 4419 18528
rect 4355 18468 4359 18524
rect 4359 18468 4415 18524
rect 4415 18468 4419 18524
rect 4355 18464 4419 18468
rect 4435 18524 4499 18528
rect 4435 18468 4439 18524
rect 4439 18468 4495 18524
rect 4495 18468 4499 18524
rect 4435 18464 4499 18468
rect 11785 18524 11849 18528
rect 11785 18468 11789 18524
rect 11789 18468 11845 18524
rect 11845 18468 11849 18524
rect 11785 18464 11849 18468
rect 11865 18524 11929 18528
rect 11865 18468 11869 18524
rect 11869 18468 11925 18524
rect 11925 18468 11929 18524
rect 11865 18464 11929 18468
rect 11945 18524 12009 18528
rect 11945 18468 11949 18524
rect 11949 18468 12005 18524
rect 12005 18468 12009 18524
rect 11945 18464 12009 18468
rect 12025 18524 12089 18528
rect 12025 18468 12029 18524
rect 12029 18468 12085 18524
rect 12085 18468 12089 18524
rect 12025 18464 12089 18468
rect 5396 18396 5460 18460
rect 19375 18524 19439 18528
rect 19375 18468 19379 18524
rect 19379 18468 19435 18524
rect 19435 18468 19439 18524
rect 19375 18464 19439 18468
rect 19455 18524 19519 18528
rect 19455 18468 19459 18524
rect 19459 18468 19515 18524
rect 19515 18468 19519 18524
rect 19455 18464 19519 18468
rect 19535 18524 19599 18528
rect 19535 18468 19539 18524
rect 19539 18468 19595 18524
rect 19595 18468 19599 18524
rect 19535 18464 19599 18468
rect 19615 18524 19679 18528
rect 19615 18468 19619 18524
rect 19619 18468 19675 18524
rect 19675 18468 19679 18524
rect 19615 18464 19679 18468
rect 26965 18524 27029 18528
rect 26965 18468 26969 18524
rect 26969 18468 27025 18524
rect 27025 18468 27029 18524
rect 26965 18464 27029 18468
rect 27045 18524 27109 18528
rect 27045 18468 27049 18524
rect 27049 18468 27105 18524
rect 27105 18468 27109 18524
rect 27045 18464 27109 18468
rect 27125 18524 27189 18528
rect 27125 18468 27129 18524
rect 27129 18468 27185 18524
rect 27185 18468 27189 18524
rect 27125 18464 27189 18468
rect 27205 18524 27269 18528
rect 27205 18468 27209 18524
rect 27209 18468 27265 18524
rect 27265 18468 27269 18524
rect 27205 18464 27269 18468
rect 4660 18124 4724 18188
rect 4844 18048 4908 18052
rect 4844 17992 4894 18048
rect 4894 17992 4908 18048
rect 4844 17988 4908 17992
rect 5948 17988 6012 18052
rect 8708 18048 8772 18052
rect 8708 17992 8722 18048
rect 8722 17992 8772 18048
rect 8708 17988 8772 17992
rect 12572 18124 12636 18188
rect 24716 18124 24780 18188
rect 14044 18048 14108 18052
rect 14044 17992 14058 18048
rect 14058 17992 14108 18048
rect 14044 17988 14108 17992
rect 7990 17980 8054 17984
rect 7990 17924 7994 17980
rect 7994 17924 8050 17980
rect 8050 17924 8054 17980
rect 7990 17920 8054 17924
rect 8070 17980 8134 17984
rect 8070 17924 8074 17980
rect 8074 17924 8130 17980
rect 8130 17924 8134 17980
rect 8070 17920 8134 17924
rect 8150 17980 8214 17984
rect 8150 17924 8154 17980
rect 8154 17924 8210 17980
rect 8210 17924 8214 17980
rect 8150 17920 8214 17924
rect 8230 17980 8294 17984
rect 8230 17924 8234 17980
rect 8234 17924 8290 17980
rect 8290 17924 8294 17980
rect 8230 17920 8294 17924
rect 15580 17980 15644 17984
rect 15580 17924 15584 17980
rect 15584 17924 15640 17980
rect 15640 17924 15644 17980
rect 15580 17920 15644 17924
rect 15660 17980 15724 17984
rect 15660 17924 15664 17980
rect 15664 17924 15720 17980
rect 15720 17924 15724 17980
rect 15660 17920 15724 17924
rect 15740 17980 15804 17984
rect 15740 17924 15744 17980
rect 15744 17924 15800 17980
rect 15800 17924 15804 17980
rect 15740 17920 15804 17924
rect 15820 17980 15884 17984
rect 15820 17924 15824 17980
rect 15824 17924 15880 17980
rect 15880 17924 15884 17980
rect 15820 17920 15884 17924
rect 23170 17980 23234 17984
rect 23170 17924 23174 17980
rect 23174 17924 23230 17980
rect 23230 17924 23234 17980
rect 23170 17920 23234 17924
rect 23250 17980 23314 17984
rect 23250 17924 23254 17980
rect 23254 17924 23310 17980
rect 23310 17924 23314 17980
rect 23250 17920 23314 17924
rect 23330 17980 23394 17984
rect 23330 17924 23334 17980
rect 23334 17924 23390 17980
rect 23390 17924 23394 17980
rect 23330 17920 23394 17924
rect 23410 17980 23474 17984
rect 23410 17924 23414 17980
rect 23414 17924 23470 17980
rect 23470 17924 23474 17980
rect 23410 17920 23474 17924
rect 30760 17980 30824 17984
rect 30760 17924 30764 17980
rect 30764 17924 30820 17980
rect 30820 17924 30824 17980
rect 30760 17920 30824 17924
rect 30840 17980 30904 17984
rect 30840 17924 30844 17980
rect 30844 17924 30900 17980
rect 30900 17924 30904 17980
rect 30840 17920 30904 17924
rect 30920 17980 30984 17984
rect 30920 17924 30924 17980
rect 30924 17924 30980 17980
rect 30980 17924 30984 17980
rect 30920 17920 30984 17924
rect 31000 17980 31064 17984
rect 31000 17924 31004 17980
rect 31004 17924 31060 17980
rect 31060 17924 31064 17980
rect 31000 17920 31064 17924
rect 4195 17436 4259 17440
rect 4195 17380 4199 17436
rect 4199 17380 4255 17436
rect 4255 17380 4259 17436
rect 4195 17376 4259 17380
rect 4275 17436 4339 17440
rect 4275 17380 4279 17436
rect 4279 17380 4335 17436
rect 4335 17380 4339 17436
rect 4275 17376 4339 17380
rect 4355 17436 4419 17440
rect 4355 17380 4359 17436
rect 4359 17380 4415 17436
rect 4415 17380 4419 17436
rect 4355 17376 4419 17380
rect 4435 17436 4499 17440
rect 4435 17380 4439 17436
rect 4439 17380 4495 17436
rect 4495 17380 4499 17436
rect 4435 17376 4499 17380
rect 11785 17436 11849 17440
rect 11785 17380 11789 17436
rect 11789 17380 11845 17436
rect 11845 17380 11849 17436
rect 11785 17376 11849 17380
rect 11865 17436 11929 17440
rect 11865 17380 11869 17436
rect 11869 17380 11925 17436
rect 11925 17380 11929 17436
rect 11865 17376 11929 17380
rect 11945 17436 12009 17440
rect 11945 17380 11949 17436
rect 11949 17380 12005 17436
rect 12005 17380 12009 17436
rect 11945 17376 12009 17380
rect 12025 17436 12089 17440
rect 12025 17380 12029 17436
rect 12029 17380 12085 17436
rect 12085 17380 12089 17436
rect 12025 17376 12089 17380
rect 19375 17436 19439 17440
rect 19375 17380 19379 17436
rect 19379 17380 19435 17436
rect 19435 17380 19439 17436
rect 19375 17376 19439 17380
rect 19455 17436 19519 17440
rect 19455 17380 19459 17436
rect 19459 17380 19515 17436
rect 19515 17380 19519 17436
rect 19455 17376 19519 17380
rect 19535 17436 19599 17440
rect 19535 17380 19539 17436
rect 19539 17380 19595 17436
rect 19595 17380 19599 17436
rect 19535 17376 19599 17380
rect 19615 17436 19679 17440
rect 19615 17380 19619 17436
rect 19619 17380 19675 17436
rect 19675 17380 19679 17436
rect 19615 17376 19679 17380
rect 26965 17436 27029 17440
rect 26965 17380 26969 17436
rect 26969 17380 27025 17436
rect 27025 17380 27029 17436
rect 26965 17376 27029 17380
rect 27045 17436 27109 17440
rect 27045 17380 27049 17436
rect 27049 17380 27105 17436
rect 27105 17380 27109 17436
rect 27045 17376 27109 17380
rect 27125 17436 27189 17440
rect 27125 17380 27129 17436
rect 27129 17380 27185 17436
rect 27185 17380 27189 17436
rect 27125 17376 27189 17380
rect 27205 17436 27269 17440
rect 27205 17380 27209 17436
rect 27209 17380 27265 17436
rect 27265 17380 27269 17436
rect 27205 17376 27269 17380
rect 10364 17308 10428 17372
rect 7990 16892 8054 16896
rect 7990 16836 7994 16892
rect 7994 16836 8050 16892
rect 8050 16836 8054 16892
rect 7990 16832 8054 16836
rect 8070 16892 8134 16896
rect 8070 16836 8074 16892
rect 8074 16836 8130 16892
rect 8130 16836 8134 16892
rect 8070 16832 8134 16836
rect 8150 16892 8214 16896
rect 8150 16836 8154 16892
rect 8154 16836 8210 16892
rect 8210 16836 8214 16892
rect 8150 16832 8214 16836
rect 8230 16892 8294 16896
rect 8230 16836 8234 16892
rect 8234 16836 8290 16892
rect 8290 16836 8294 16892
rect 8230 16832 8294 16836
rect 15580 16892 15644 16896
rect 15580 16836 15584 16892
rect 15584 16836 15640 16892
rect 15640 16836 15644 16892
rect 15580 16832 15644 16836
rect 15660 16892 15724 16896
rect 15660 16836 15664 16892
rect 15664 16836 15720 16892
rect 15720 16836 15724 16892
rect 15660 16832 15724 16836
rect 15740 16892 15804 16896
rect 15740 16836 15744 16892
rect 15744 16836 15800 16892
rect 15800 16836 15804 16892
rect 15740 16832 15804 16836
rect 15820 16892 15884 16896
rect 15820 16836 15824 16892
rect 15824 16836 15880 16892
rect 15880 16836 15884 16892
rect 15820 16832 15884 16836
rect 23170 16892 23234 16896
rect 23170 16836 23174 16892
rect 23174 16836 23230 16892
rect 23230 16836 23234 16892
rect 23170 16832 23234 16836
rect 23250 16892 23314 16896
rect 23250 16836 23254 16892
rect 23254 16836 23310 16892
rect 23310 16836 23314 16892
rect 23250 16832 23314 16836
rect 23330 16892 23394 16896
rect 23330 16836 23334 16892
rect 23334 16836 23390 16892
rect 23390 16836 23394 16892
rect 23330 16832 23394 16836
rect 23410 16892 23474 16896
rect 23410 16836 23414 16892
rect 23414 16836 23470 16892
rect 23470 16836 23474 16892
rect 23410 16832 23474 16836
rect 15148 16628 15212 16692
rect 30760 16892 30824 16896
rect 30760 16836 30764 16892
rect 30764 16836 30820 16892
rect 30820 16836 30824 16892
rect 30760 16832 30824 16836
rect 30840 16892 30904 16896
rect 30840 16836 30844 16892
rect 30844 16836 30900 16892
rect 30900 16836 30904 16892
rect 30840 16832 30904 16836
rect 30920 16892 30984 16896
rect 30920 16836 30924 16892
rect 30924 16836 30980 16892
rect 30980 16836 30984 16892
rect 30920 16832 30984 16836
rect 31000 16892 31064 16896
rect 31000 16836 31004 16892
rect 31004 16836 31060 16892
rect 31060 16836 31064 16892
rect 31000 16832 31064 16836
rect 6868 16492 6932 16556
rect 23980 16492 24044 16556
rect 4195 16348 4259 16352
rect 4195 16292 4199 16348
rect 4199 16292 4255 16348
rect 4255 16292 4259 16348
rect 4195 16288 4259 16292
rect 4275 16348 4339 16352
rect 4275 16292 4279 16348
rect 4279 16292 4335 16348
rect 4335 16292 4339 16348
rect 4275 16288 4339 16292
rect 4355 16348 4419 16352
rect 4355 16292 4359 16348
rect 4359 16292 4415 16348
rect 4415 16292 4419 16348
rect 4355 16288 4419 16292
rect 4435 16348 4499 16352
rect 4435 16292 4439 16348
rect 4439 16292 4495 16348
rect 4495 16292 4499 16348
rect 4435 16288 4499 16292
rect 11785 16348 11849 16352
rect 11785 16292 11789 16348
rect 11789 16292 11845 16348
rect 11845 16292 11849 16348
rect 11785 16288 11849 16292
rect 11865 16348 11929 16352
rect 11865 16292 11869 16348
rect 11869 16292 11925 16348
rect 11925 16292 11929 16348
rect 11865 16288 11929 16292
rect 11945 16348 12009 16352
rect 11945 16292 11949 16348
rect 11949 16292 12005 16348
rect 12005 16292 12009 16348
rect 11945 16288 12009 16292
rect 12025 16348 12089 16352
rect 12025 16292 12029 16348
rect 12029 16292 12085 16348
rect 12085 16292 12089 16348
rect 12025 16288 12089 16292
rect 19375 16348 19439 16352
rect 19375 16292 19379 16348
rect 19379 16292 19435 16348
rect 19435 16292 19439 16348
rect 19375 16288 19439 16292
rect 19455 16348 19519 16352
rect 19455 16292 19459 16348
rect 19459 16292 19515 16348
rect 19515 16292 19519 16348
rect 19455 16288 19519 16292
rect 19535 16348 19599 16352
rect 19535 16292 19539 16348
rect 19539 16292 19595 16348
rect 19595 16292 19599 16348
rect 19535 16288 19599 16292
rect 19615 16348 19679 16352
rect 19615 16292 19619 16348
rect 19619 16292 19675 16348
rect 19675 16292 19679 16348
rect 19615 16288 19679 16292
rect 26965 16348 27029 16352
rect 26965 16292 26969 16348
rect 26969 16292 27025 16348
rect 27025 16292 27029 16348
rect 26965 16288 27029 16292
rect 27045 16348 27109 16352
rect 27045 16292 27049 16348
rect 27049 16292 27105 16348
rect 27105 16292 27109 16348
rect 27045 16288 27109 16292
rect 27125 16348 27189 16352
rect 27125 16292 27129 16348
rect 27129 16292 27185 16348
rect 27185 16292 27189 16348
rect 27125 16288 27189 16292
rect 27205 16348 27269 16352
rect 27205 16292 27209 16348
rect 27209 16292 27265 16348
rect 27265 16292 27269 16348
rect 27205 16288 27269 16292
rect 27660 16220 27724 16284
rect 7990 15804 8054 15808
rect 7990 15748 7994 15804
rect 7994 15748 8050 15804
rect 8050 15748 8054 15804
rect 7990 15744 8054 15748
rect 8070 15804 8134 15808
rect 8070 15748 8074 15804
rect 8074 15748 8130 15804
rect 8130 15748 8134 15804
rect 8070 15744 8134 15748
rect 8150 15804 8214 15808
rect 8150 15748 8154 15804
rect 8154 15748 8210 15804
rect 8210 15748 8214 15804
rect 8150 15744 8214 15748
rect 8230 15804 8294 15808
rect 8230 15748 8234 15804
rect 8234 15748 8290 15804
rect 8290 15748 8294 15804
rect 8230 15744 8294 15748
rect 15580 15804 15644 15808
rect 15580 15748 15584 15804
rect 15584 15748 15640 15804
rect 15640 15748 15644 15804
rect 15580 15744 15644 15748
rect 15660 15804 15724 15808
rect 15660 15748 15664 15804
rect 15664 15748 15720 15804
rect 15720 15748 15724 15804
rect 15660 15744 15724 15748
rect 15740 15804 15804 15808
rect 15740 15748 15744 15804
rect 15744 15748 15800 15804
rect 15800 15748 15804 15804
rect 15740 15744 15804 15748
rect 15820 15804 15884 15808
rect 15820 15748 15824 15804
rect 15824 15748 15880 15804
rect 15880 15748 15884 15804
rect 15820 15744 15884 15748
rect 23170 15804 23234 15808
rect 23170 15748 23174 15804
rect 23174 15748 23230 15804
rect 23230 15748 23234 15804
rect 23170 15744 23234 15748
rect 23250 15804 23314 15808
rect 23250 15748 23254 15804
rect 23254 15748 23310 15804
rect 23310 15748 23314 15804
rect 23250 15744 23314 15748
rect 23330 15804 23394 15808
rect 23330 15748 23334 15804
rect 23334 15748 23390 15804
rect 23390 15748 23394 15804
rect 23330 15744 23394 15748
rect 23410 15804 23474 15808
rect 23410 15748 23414 15804
rect 23414 15748 23470 15804
rect 23470 15748 23474 15804
rect 23410 15744 23474 15748
rect 30760 15804 30824 15808
rect 30760 15748 30764 15804
rect 30764 15748 30820 15804
rect 30820 15748 30824 15804
rect 30760 15744 30824 15748
rect 30840 15804 30904 15808
rect 30840 15748 30844 15804
rect 30844 15748 30900 15804
rect 30900 15748 30904 15804
rect 30840 15744 30904 15748
rect 30920 15804 30984 15808
rect 30920 15748 30924 15804
rect 30924 15748 30980 15804
rect 30980 15748 30984 15804
rect 30920 15744 30984 15748
rect 31000 15804 31064 15808
rect 31000 15748 31004 15804
rect 31004 15748 31060 15804
rect 31060 15748 31064 15804
rect 31000 15744 31064 15748
rect 8524 15404 8588 15468
rect 4195 15260 4259 15264
rect 4195 15204 4199 15260
rect 4199 15204 4255 15260
rect 4255 15204 4259 15260
rect 4195 15200 4259 15204
rect 4275 15260 4339 15264
rect 4275 15204 4279 15260
rect 4279 15204 4335 15260
rect 4335 15204 4339 15260
rect 4275 15200 4339 15204
rect 4355 15260 4419 15264
rect 4355 15204 4359 15260
rect 4359 15204 4415 15260
rect 4415 15204 4419 15260
rect 4355 15200 4419 15204
rect 4435 15260 4499 15264
rect 4435 15204 4439 15260
rect 4439 15204 4495 15260
rect 4495 15204 4499 15260
rect 4435 15200 4499 15204
rect 11785 15260 11849 15264
rect 11785 15204 11789 15260
rect 11789 15204 11845 15260
rect 11845 15204 11849 15260
rect 11785 15200 11849 15204
rect 11865 15260 11929 15264
rect 11865 15204 11869 15260
rect 11869 15204 11925 15260
rect 11925 15204 11929 15260
rect 11865 15200 11929 15204
rect 11945 15260 12009 15264
rect 11945 15204 11949 15260
rect 11949 15204 12005 15260
rect 12005 15204 12009 15260
rect 11945 15200 12009 15204
rect 12025 15260 12089 15264
rect 12025 15204 12029 15260
rect 12029 15204 12085 15260
rect 12085 15204 12089 15260
rect 12025 15200 12089 15204
rect 19375 15260 19439 15264
rect 19375 15204 19379 15260
rect 19379 15204 19435 15260
rect 19435 15204 19439 15260
rect 19375 15200 19439 15204
rect 19455 15260 19519 15264
rect 19455 15204 19459 15260
rect 19459 15204 19515 15260
rect 19515 15204 19519 15260
rect 19455 15200 19519 15204
rect 19535 15260 19599 15264
rect 19535 15204 19539 15260
rect 19539 15204 19595 15260
rect 19595 15204 19599 15260
rect 19535 15200 19599 15204
rect 19615 15260 19679 15264
rect 19615 15204 19619 15260
rect 19619 15204 19675 15260
rect 19675 15204 19679 15260
rect 19615 15200 19679 15204
rect 26965 15260 27029 15264
rect 26965 15204 26969 15260
rect 26969 15204 27025 15260
rect 27025 15204 27029 15260
rect 26965 15200 27029 15204
rect 27045 15260 27109 15264
rect 27045 15204 27049 15260
rect 27049 15204 27105 15260
rect 27105 15204 27109 15260
rect 27045 15200 27109 15204
rect 27125 15260 27189 15264
rect 27125 15204 27129 15260
rect 27129 15204 27185 15260
rect 27185 15204 27189 15260
rect 27125 15200 27189 15204
rect 27205 15260 27269 15264
rect 27205 15204 27209 15260
rect 27209 15204 27265 15260
rect 27265 15204 27269 15260
rect 27205 15200 27269 15204
rect 7990 14716 8054 14720
rect 7990 14660 7994 14716
rect 7994 14660 8050 14716
rect 8050 14660 8054 14716
rect 7990 14656 8054 14660
rect 8070 14716 8134 14720
rect 8070 14660 8074 14716
rect 8074 14660 8130 14716
rect 8130 14660 8134 14716
rect 8070 14656 8134 14660
rect 8150 14716 8214 14720
rect 8150 14660 8154 14716
rect 8154 14660 8210 14716
rect 8210 14660 8214 14716
rect 8150 14656 8214 14660
rect 8230 14716 8294 14720
rect 8230 14660 8234 14716
rect 8234 14660 8290 14716
rect 8290 14660 8294 14716
rect 8230 14656 8294 14660
rect 15580 14716 15644 14720
rect 15580 14660 15584 14716
rect 15584 14660 15640 14716
rect 15640 14660 15644 14716
rect 15580 14656 15644 14660
rect 15660 14716 15724 14720
rect 15660 14660 15664 14716
rect 15664 14660 15720 14716
rect 15720 14660 15724 14716
rect 15660 14656 15724 14660
rect 15740 14716 15804 14720
rect 15740 14660 15744 14716
rect 15744 14660 15800 14716
rect 15800 14660 15804 14716
rect 15740 14656 15804 14660
rect 15820 14716 15884 14720
rect 15820 14660 15824 14716
rect 15824 14660 15880 14716
rect 15880 14660 15884 14716
rect 15820 14656 15884 14660
rect 23170 14716 23234 14720
rect 23170 14660 23174 14716
rect 23174 14660 23230 14716
rect 23230 14660 23234 14716
rect 23170 14656 23234 14660
rect 23250 14716 23314 14720
rect 23250 14660 23254 14716
rect 23254 14660 23310 14716
rect 23310 14660 23314 14716
rect 23250 14656 23314 14660
rect 23330 14716 23394 14720
rect 23330 14660 23334 14716
rect 23334 14660 23390 14716
rect 23390 14660 23394 14716
rect 23330 14656 23394 14660
rect 23410 14716 23474 14720
rect 23410 14660 23414 14716
rect 23414 14660 23470 14716
rect 23470 14660 23474 14716
rect 23410 14656 23474 14660
rect 30760 14716 30824 14720
rect 30760 14660 30764 14716
rect 30764 14660 30820 14716
rect 30820 14660 30824 14716
rect 30760 14656 30824 14660
rect 30840 14716 30904 14720
rect 30840 14660 30844 14716
rect 30844 14660 30900 14716
rect 30900 14660 30904 14716
rect 30840 14656 30904 14660
rect 30920 14716 30984 14720
rect 30920 14660 30924 14716
rect 30924 14660 30980 14716
rect 30980 14660 30984 14716
rect 30920 14656 30984 14660
rect 31000 14716 31064 14720
rect 31000 14660 31004 14716
rect 31004 14660 31060 14716
rect 31060 14660 31064 14716
rect 31000 14656 31064 14660
rect 2084 14316 2148 14380
rect 9444 14180 9508 14244
rect 4195 14172 4259 14176
rect 4195 14116 4199 14172
rect 4199 14116 4255 14172
rect 4255 14116 4259 14172
rect 4195 14112 4259 14116
rect 4275 14172 4339 14176
rect 4275 14116 4279 14172
rect 4279 14116 4335 14172
rect 4335 14116 4339 14172
rect 4275 14112 4339 14116
rect 4355 14172 4419 14176
rect 4355 14116 4359 14172
rect 4359 14116 4415 14172
rect 4415 14116 4419 14172
rect 4355 14112 4419 14116
rect 4435 14172 4499 14176
rect 4435 14116 4439 14172
rect 4439 14116 4495 14172
rect 4495 14116 4499 14172
rect 4435 14112 4499 14116
rect 11785 14172 11849 14176
rect 11785 14116 11789 14172
rect 11789 14116 11845 14172
rect 11845 14116 11849 14172
rect 11785 14112 11849 14116
rect 11865 14172 11929 14176
rect 11865 14116 11869 14172
rect 11869 14116 11925 14172
rect 11925 14116 11929 14172
rect 11865 14112 11929 14116
rect 11945 14172 12009 14176
rect 11945 14116 11949 14172
rect 11949 14116 12005 14172
rect 12005 14116 12009 14172
rect 11945 14112 12009 14116
rect 12025 14172 12089 14176
rect 12025 14116 12029 14172
rect 12029 14116 12085 14172
rect 12085 14116 12089 14172
rect 12025 14112 12089 14116
rect 19375 14172 19439 14176
rect 19375 14116 19379 14172
rect 19379 14116 19435 14172
rect 19435 14116 19439 14172
rect 19375 14112 19439 14116
rect 19455 14172 19519 14176
rect 19455 14116 19459 14172
rect 19459 14116 19515 14172
rect 19515 14116 19519 14172
rect 19455 14112 19519 14116
rect 19535 14172 19599 14176
rect 19535 14116 19539 14172
rect 19539 14116 19595 14172
rect 19595 14116 19599 14172
rect 19535 14112 19599 14116
rect 19615 14172 19679 14176
rect 19615 14116 19619 14172
rect 19619 14116 19675 14172
rect 19675 14116 19679 14172
rect 19615 14112 19679 14116
rect 26965 14172 27029 14176
rect 26965 14116 26969 14172
rect 26969 14116 27025 14172
rect 27025 14116 27029 14172
rect 26965 14112 27029 14116
rect 27045 14172 27109 14176
rect 27045 14116 27049 14172
rect 27049 14116 27105 14172
rect 27105 14116 27109 14172
rect 27045 14112 27109 14116
rect 27125 14172 27189 14176
rect 27125 14116 27129 14172
rect 27129 14116 27185 14172
rect 27185 14116 27189 14172
rect 27125 14112 27189 14116
rect 27205 14172 27269 14176
rect 27205 14116 27209 14172
rect 27209 14116 27265 14172
rect 27265 14116 27269 14172
rect 27205 14112 27269 14116
rect 7990 13628 8054 13632
rect 7990 13572 7994 13628
rect 7994 13572 8050 13628
rect 8050 13572 8054 13628
rect 7990 13568 8054 13572
rect 8070 13628 8134 13632
rect 8070 13572 8074 13628
rect 8074 13572 8130 13628
rect 8130 13572 8134 13628
rect 8070 13568 8134 13572
rect 8150 13628 8214 13632
rect 8150 13572 8154 13628
rect 8154 13572 8210 13628
rect 8210 13572 8214 13628
rect 8150 13568 8214 13572
rect 8230 13628 8294 13632
rect 8230 13572 8234 13628
rect 8234 13572 8290 13628
rect 8290 13572 8294 13628
rect 8230 13568 8294 13572
rect 8892 13636 8956 13700
rect 11100 13636 11164 13700
rect 15580 13628 15644 13632
rect 15580 13572 15584 13628
rect 15584 13572 15640 13628
rect 15640 13572 15644 13628
rect 15580 13568 15644 13572
rect 15660 13628 15724 13632
rect 15660 13572 15664 13628
rect 15664 13572 15720 13628
rect 15720 13572 15724 13628
rect 15660 13568 15724 13572
rect 15740 13628 15804 13632
rect 15740 13572 15744 13628
rect 15744 13572 15800 13628
rect 15800 13572 15804 13628
rect 15740 13568 15804 13572
rect 15820 13628 15884 13632
rect 15820 13572 15824 13628
rect 15824 13572 15880 13628
rect 15880 13572 15884 13628
rect 15820 13568 15884 13572
rect 23170 13628 23234 13632
rect 23170 13572 23174 13628
rect 23174 13572 23230 13628
rect 23230 13572 23234 13628
rect 23170 13568 23234 13572
rect 23250 13628 23314 13632
rect 23250 13572 23254 13628
rect 23254 13572 23310 13628
rect 23310 13572 23314 13628
rect 23250 13568 23314 13572
rect 23330 13628 23394 13632
rect 23330 13572 23334 13628
rect 23334 13572 23390 13628
rect 23390 13572 23394 13628
rect 23330 13568 23394 13572
rect 23410 13628 23474 13632
rect 23410 13572 23414 13628
rect 23414 13572 23470 13628
rect 23470 13572 23474 13628
rect 23410 13568 23474 13572
rect 30760 13628 30824 13632
rect 30760 13572 30764 13628
rect 30764 13572 30820 13628
rect 30820 13572 30824 13628
rect 30760 13568 30824 13572
rect 30840 13628 30904 13632
rect 30840 13572 30844 13628
rect 30844 13572 30900 13628
rect 30900 13572 30904 13628
rect 30840 13568 30904 13572
rect 30920 13628 30984 13632
rect 30920 13572 30924 13628
rect 30924 13572 30980 13628
rect 30980 13572 30984 13628
rect 30920 13568 30984 13572
rect 31000 13628 31064 13632
rect 31000 13572 31004 13628
rect 31004 13572 31060 13628
rect 31060 13572 31064 13628
rect 31000 13568 31064 13572
rect 8524 13364 8588 13428
rect 4195 13084 4259 13088
rect 4195 13028 4199 13084
rect 4199 13028 4255 13084
rect 4255 13028 4259 13084
rect 4195 13024 4259 13028
rect 4275 13084 4339 13088
rect 4275 13028 4279 13084
rect 4279 13028 4335 13084
rect 4335 13028 4339 13084
rect 4275 13024 4339 13028
rect 4355 13084 4419 13088
rect 4355 13028 4359 13084
rect 4359 13028 4415 13084
rect 4415 13028 4419 13084
rect 4355 13024 4419 13028
rect 4435 13084 4499 13088
rect 4435 13028 4439 13084
rect 4439 13028 4495 13084
rect 4495 13028 4499 13084
rect 4435 13024 4499 13028
rect 5028 13228 5092 13292
rect 11785 13084 11849 13088
rect 11785 13028 11789 13084
rect 11789 13028 11845 13084
rect 11845 13028 11849 13084
rect 11785 13024 11849 13028
rect 11865 13084 11929 13088
rect 11865 13028 11869 13084
rect 11869 13028 11925 13084
rect 11925 13028 11929 13084
rect 11865 13024 11929 13028
rect 11945 13084 12009 13088
rect 11945 13028 11949 13084
rect 11949 13028 12005 13084
rect 12005 13028 12009 13084
rect 11945 13024 12009 13028
rect 12025 13084 12089 13088
rect 12025 13028 12029 13084
rect 12029 13028 12085 13084
rect 12085 13028 12089 13084
rect 12025 13024 12089 13028
rect 19375 13084 19439 13088
rect 19375 13028 19379 13084
rect 19379 13028 19435 13084
rect 19435 13028 19439 13084
rect 19375 13024 19439 13028
rect 19455 13084 19519 13088
rect 19455 13028 19459 13084
rect 19459 13028 19515 13084
rect 19515 13028 19519 13084
rect 19455 13024 19519 13028
rect 19535 13084 19599 13088
rect 19535 13028 19539 13084
rect 19539 13028 19595 13084
rect 19595 13028 19599 13084
rect 19535 13024 19599 13028
rect 19615 13084 19679 13088
rect 19615 13028 19619 13084
rect 19619 13028 19675 13084
rect 19675 13028 19679 13084
rect 19615 13024 19679 13028
rect 26965 13084 27029 13088
rect 26965 13028 26969 13084
rect 26969 13028 27025 13084
rect 27025 13028 27029 13084
rect 26965 13024 27029 13028
rect 27045 13084 27109 13088
rect 27045 13028 27049 13084
rect 27049 13028 27105 13084
rect 27105 13028 27109 13084
rect 27045 13024 27109 13028
rect 27125 13084 27189 13088
rect 27125 13028 27129 13084
rect 27129 13028 27185 13084
rect 27185 13028 27189 13084
rect 27125 13024 27189 13028
rect 27205 13084 27269 13088
rect 27205 13028 27209 13084
rect 27209 13028 27265 13084
rect 27265 13028 27269 13084
rect 27205 13024 27269 13028
rect 27660 12684 27724 12748
rect 7990 12540 8054 12544
rect 7990 12484 7994 12540
rect 7994 12484 8050 12540
rect 8050 12484 8054 12540
rect 7990 12480 8054 12484
rect 8070 12540 8134 12544
rect 8070 12484 8074 12540
rect 8074 12484 8130 12540
rect 8130 12484 8134 12540
rect 8070 12480 8134 12484
rect 8150 12540 8214 12544
rect 8150 12484 8154 12540
rect 8154 12484 8210 12540
rect 8210 12484 8214 12540
rect 8150 12480 8214 12484
rect 8230 12540 8294 12544
rect 8230 12484 8234 12540
rect 8234 12484 8290 12540
rect 8290 12484 8294 12540
rect 8230 12480 8294 12484
rect 15580 12540 15644 12544
rect 15580 12484 15584 12540
rect 15584 12484 15640 12540
rect 15640 12484 15644 12540
rect 15580 12480 15644 12484
rect 15660 12540 15724 12544
rect 15660 12484 15664 12540
rect 15664 12484 15720 12540
rect 15720 12484 15724 12540
rect 15660 12480 15724 12484
rect 15740 12540 15804 12544
rect 15740 12484 15744 12540
rect 15744 12484 15800 12540
rect 15800 12484 15804 12540
rect 15740 12480 15804 12484
rect 15820 12540 15884 12544
rect 15820 12484 15824 12540
rect 15824 12484 15880 12540
rect 15880 12484 15884 12540
rect 15820 12480 15884 12484
rect 23170 12540 23234 12544
rect 23170 12484 23174 12540
rect 23174 12484 23230 12540
rect 23230 12484 23234 12540
rect 23170 12480 23234 12484
rect 23250 12540 23314 12544
rect 23250 12484 23254 12540
rect 23254 12484 23310 12540
rect 23310 12484 23314 12540
rect 23250 12480 23314 12484
rect 23330 12540 23394 12544
rect 23330 12484 23334 12540
rect 23334 12484 23390 12540
rect 23390 12484 23394 12540
rect 23330 12480 23394 12484
rect 23410 12540 23474 12544
rect 23410 12484 23414 12540
rect 23414 12484 23470 12540
rect 23470 12484 23474 12540
rect 23410 12480 23474 12484
rect 30760 12540 30824 12544
rect 30760 12484 30764 12540
rect 30764 12484 30820 12540
rect 30820 12484 30824 12540
rect 30760 12480 30824 12484
rect 30840 12540 30904 12544
rect 30840 12484 30844 12540
rect 30844 12484 30900 12540
rect 30900 12484 30904 12540
rect 30840 12480 30904 12484
rect 30920 12540 30984 12544
rect 30920 12484 30924 12540
rect 30924 12484 30980 12540
rect 30980 12484 30984 12540
rect 30920 12480 30984 12484
rect 31000 12540 31064 12544
rect 31000 12484 31004 12540
rect 31004 12484 31060 12540
rect 31060 12484 31064 12540
rect 31000 12480 31064 12484
rect 4195 11996 4259 12000
rect 4195 11940 4199 11996
rect 4199 11940 4255 11996
rect 4255 11940 4259 11996
rect 4195 11936 4259 11940
rect 4275 11996 4339 12000
rect 4275 11940 4279 11996
rect 4279 11940 4335 11996
rect 4335 11940 4339 11996
rect 4275 11936 4339 11940
rect 4355 11996 4419 12000
rect 4355 11940 4359 11996
rect 4359 11940 4415 11996
rect 4415 11940 4419 11996
rect 4355 11936 4419 11940
rect 4435 11996 4499 12000
rect 4435 11940 4439 11996
rect 4439 11940 4495 11996
rect 4495 11940 4499 11996
rect 4435 11936 4499 11940
rect 11785 11996 11849 12000
rect 11785 11940 11789 11996
rect 11789 11940 11845 11996
rect 11845 11940 11849 11996
rect 11785 11936 11849 11940
rect 11865 11996 11929 12000
rect 11865 11940 11869 11996
rect 11869 11940 11925 11996
rect 11925 11940 11929 11996
rect 11865 11936 11929 11940
rect 11945 11996 12009 12000
rect 11945 11940 11949 11996
rect 11949 11940 12005 11996
rect 12005 11940 12009 11996
rect 11945 11936 12009 11940
rect 12025 11996 12089 12000
rect 12025 11940 12029 11996
rect 12029 11940 12085 11996
rect 12085 11940 12089 11996
rect 12025 11936 12089 11940
rect 19375 11996 19439 12000
rect 19375 11940 19379 11996
rect 19379 11940 19435 11996
rect 19435 11940 19439 11996
rect 19375 11936 19439 11940
rect 19455 11996 19519 12000
rect 19455 11940 19459 11996
rect 19459 11940 19515 11996
rect 19515 11940 19519 11996
rect 19455 11936 19519 11940
rect 19535 11996 19599 12000
rect 19535 11940 19539 11996
rect 19539 11940 19595 11996
rect 19595 11940 19599 11996
rect 19535 11936 19599 11940
rect 19615 11996 19679 12000
rect 19615 11940 19619 11996
rect 19619 11940 19675 11996
rect 19675 11940 19679 11996
rect 19615 11936 19679 11940
rect 26965 11996 27029 12000
rect 26965 11940 26969 11996
rect 26969 11940 27025 11996
rect 27025 11940 27029 11996
rect 26965 11936 27029 11940
rect 27045 11996 27109 12000
rect 27045 11940 27049 11996
rect 27049 11940 27105 11996
rect 27105 11940 27109 11996
rect 27045 11936 27109 11940
rect 27125 11996 27189 12000
rect 27125 11940 27129 11996
rect 27129 11940 27185 11996
rect 27185 11940 27189 11996
rect 27125 11936 27189 11940
rect 27205 11996 27269 12000
rect 27205 11940 27209 11996
rect 27209 11940 27265 11996
rect 27265 11940 27269 11996
rect 27205 11936 27269 11940
rect 23980 11732 24044 11796
rect 15148 11596 15212 11660
rect 7990 11452 8054 11456
rect 7990 11396 7994 11452
rect 7994 11396 8050 11452
rect 8050 11396 8054 11452
rect 7990 11392 8054 11396
rect 8070 11452 8134 11456
rect 8070 11396 8074 11452
rect 8074 11396 8130 11452
rect 8130 11396 8134 11452
rect 8070 11392 8134 11396
rect 8150 11452 8214 11456
rect 8150 11396 8154 11452
rect 8154 11396 8210 11452
rect 8210 11396 8214 11452
rect 8150 11392 8214 11396
rect 8230 11452 8294 11456
rect 8230 11396 8234 11452
rect 8234 11396 8290 11452
rect 8290 11396 8294 11452
rect 8230 11392 8294 11396
rect 15580 11452 15644 11456
rect 15580 11396 15584 11452
rect 15584 11396 15640 11452
rect 15640 11396 15644 11452
rect 15580 11392 15644 11396
rect 15660 11452 15724 11456
rect 15660 11396 15664 11452
rect 15664 11396 15720 11452
rect 15720 11396 15724 11452
rect 15660 11392 15724 11396
rect 15740 11452 15804 11456
rect 15740 11396 15744 11452
rect 15744 11396 15800 11452
rect 15800 11396 15804 11452
rect 15740 11392 15804 11396
rect 15820 11452 15884 11456
rect 15820 11396 15824 11452
rect 15824 11396 15880 11452
rect 15880 11396 15884 11452
rect 15820 11392 15884 11396
rect 23170 11452 23234 11456
rect 23170 11396 23174 11452
rect 23174 11396 23230 11452
rect 23230 11396 23234 11452
rect 23170 11392 23234 11396
rect 23250 11452 23314 11456
rect 23250 11396 23254 11452
rect 23254 11396 23310 11452
rect 23310 11396 23314 11452
rect 23250 11392 23314 11396
rect 23330 11452 23394 11456
rect 23330 11396 23334 11452
rect 23334 11396 23390 11452
rect 23390 11396 23394 11452
rect 23330 11392 23394 11396
rect 23410 11452 23474 11456
rect 23410 11396 23414 11452
rect 23414 11396 23470 11452
rect 23470 11396 23474 11452
rect 23410 11392 23474 11396
rect 30760 11452 30824 11456
rect 30760 11396 30764 11452
rect 30764 11396 30820 11452
rect 30820 11396 30824 11452
rect 30760 11392 30824 11396
rect 30840 11452 30904 11456
rect 30840 11396 30844 11452
rect 30844 11396 30900 11452
rect 30900 11396 30904 11452
rect 30840 11392 30904 11396
rect 30920 11452 30984 11456
rect 30920 11396 30924 11452
rect 30924 11396 30980 11452
rect 30980 11396 30984 11452
rect 30920 11392 30984 11396
rect 31000 11452 31064 11456
rect 31000 11396 31004 11452
rect 31004 11396 31060 11452
rect 31060 11396 31064 11452
rect 31000 11392 31064 11396
rect 8524 11324 8588 11388
rect 10364 11052 10428 11116
rect 4195 10908 4259 10912
rect 4195 10852 4199 10908
rect 4199 10852 4255 10908
rect 4255 10852 4259 10908
rect 4195 10848 4259 10852
rect 4275 10908 4339 10912
rect 4275 10852 4279 10908
rect 4279 10852 4335 10908
rect 4335 10852 4339 10908
rect 4275 10848 4339 10852
rect 4355 10908 4419 10912
rect 4355 10852 4359 10908
rect 4359 10852 4415 10908
rect 4415 10852 4419 10908
rect 4355 10848 4419 10852
rect 4435 10908 4499 10912
rect 4435 10852 4439 10908
rect 4439 10852 4495 10908
rect 4495 10852 4499 10908
rect 4435 10848 4499 10852
rect 11785 10908 11849 10912
rect 11785 10852 11789 10908
rect 11789 10852 11845 10908
rect 11845 10852 11849 10908
rect 11785 10848 11849 10852
rect 11865 10908 11929 10912
rect 11865 10852 11869 10908
rect 11869 10852 11925 10908
rect 11925 10852 11929 10908
rect 11865 10848 11929 10852
rect 11945 10908 12009 10912
rect 11945 10852 11949 10908
rect 11949 10852 12005 10908
rect 12005 10852 12009 10908
rect 11945 10848 12009 10852
rect 12025 10908 12089 10912
rect 12025 10852 12029 10908
rect 12029 10852 12085 10908
rect 12085 10852 12089 10908
rect 12025 10848 12089 10852
rect 19375 10908 19439 10912
rect 19375 10852 19379 10908
rect 19379 10852 19435 10908
rect 19435 10852 19439 10908
rect 19375 10848 19439 10852
rect 19455 10908 19519 10912
rect 19455 10852 19459 10908
rect 19459 10852 19515 10908
rect 19515 10852 19519 10908
rect 19455 10848 19519 10852
rect 19535 10908 19599 10912
rect 19535 10852 19539 10908
rect 19539 10852 19595 10908
rect 19595 10852 19599 10908
rect 19535 10848 19599 10852
rect 19615 10908 19679 10912
rect 19615 10852 19619 10908
rect 19619 10852 19675 10908
rect 19675 10852 19679 10908
rect 19615 10848 19679 10852
rect 26965 10908 27029 10912
rect 26965 10852 26969 10908
rect 26969 10852 27025 10908
rect 27025 10852 27029 10908
rect 26965 10848 27029 10852
rect 27045 10908 27109 10912
rect 27045 10852 27049 10908
rect 27049 10852 27105 10908
rect 27105 10852 27109 10908
rect 27045 10848 27109 10852
rect 27125 10908 27189 10912
rect 27125 10852 27129 10908
rect 27129 10852 27185 10908
rect 27185 10852 27189 10908
rect 27125 10848 27189 10852
rect 27205 10908 27269 10912
rect 27205 10852 27209 10908
rect 27209 10852 27265 10908
rect 27265 10852 27269 10908
rect 27205 10848 27269 10852
rect 7990 10364 8054 10368
rect 7990 10308 7994 10364
rect 7994 10308 8050 10364
rect 8050 10308 8054 10364
rect 7990 10304 8054 10308
rect 8070 10364 8134 10368
rect 8070 10308 8074 10364
rect 8074 10308 8130 10364
rect 8130 10308 8134 10364
rect 8070 10304 8134 10308
rect 8150 10364 8214 10368
rect 8150 10308 8154 10364
rect 8154 10308 8210 10364
rect 8210 10308 8214 10364
rect 8150 10304 8214 10308
rect 8230 10364 8294 10368
rect 8230 10308 8234 10364
rect 8234 10308 8290 10364
rect 8290 10308 8294 10364
rect 8230 10304 8294 10308
rect 15580 10364 15644 10368
rect 15580 10308 15584 10364
rect 15584 10308 15640 10364
rect 15640 10308 15644 10364
rect 15580 10304 15644 10308
rect 15660 10364 15724 10368
rect 15660 10308 15664 10364
rect 15664 10308 15720 10364
rect 15720 10308 15724 10364
rect 15660 10304 15724 10308
rect 15740 10364 15804 10368
rect 15740 10308 15744 10364
rect 15744 10308 15800 10364
rect 15800 10308 15804 10364
rect 15740 10304 15804 10308
rect 15820 10364 15884 10368
rect 15820 10308 15824 10364
rect 15824 10308 15880 10364
rect 15880 10308 15884 10364
rect 15820 10304 15884 10308
rect 23170 10364 23234 10368
rect 23170 10308 23174 10364
rect 23174 10308 23230 10364
rect 23230 10308 23234 10364
rect 23170 10304 23234 10308
rect 23250 10364 23314 10368
rect 23250 10308 23254 10364
rect 23254 10308 23310 10364
rect 23310 10308 23314 10364
rect 23250 10304 23314 10308
rect 23330 10364 23394 10368
rect 23330 10308 23334 10364
rect 23334 10308 23390 10364
rect 23390 10308 23394 10364
rect 23330 10304 23394 10308
rect 23410 10364 23474 10368
rect 23410 10308 23414 10364
rect 23414 10308 23470 10364
rect 23470 10308 23474 10364
rect 23410 10304 23474 10308
rect 30760 10364 30824 10368
rect 30760 10308 30764 10364
rect 30764 10308 30820 10364
rect 30820 10308 30824 10364
rect 30760 10304 30824 10308
rect 30840 10364 30904 10368
rect 30840 10308 30844 10364
rect 30844 10308 30900 10364
rect 30900 10308 30904 10364
rect 30840 10304 30904 10308
rect 30920 10364 30984 10368
rect 30920 10308 30924 10364
rect 30924 10308 30980 10364
rect 30980 10308 30984 10364
rect 30920 10304 30984 10308
rect 31000 10364 31064 10368
rect 31000 10308 31004 10364
rect 31004 10308 31060 10364
rect 31060 10308 31064 10364
rect 31000 10304 31064 10308
rect 4195 9820 4259 9824
rect 4195 9764 4199 9820
rect 4199 9764 4255 9820
rect 4255 9764 4259 9820
rect 4195 9760 4259 9764
rect 4275 9820 4339 9824
rect 4275 9764 4279 9820
rect 4279 9764 4335 9820
rect 4335 9764 4339 9820
rect 4275 9760 4339 9764
rect 4355 9820 4419 9824
rect 4355 9764 4359 9820
rect 4359 9764 4415 9820
rect 4415 9764 4419 9820
rect 4355 9760 4419 9764
rect 4435 9820 4499 9824
rect 4435 9764 4439 9820
rect 4439 9764 4495 9820
rect 4495 9764 4499 9820
rect 4435 9760 4499 9764
rect 11785 9820 11849 9824
rect 11785 9764 11789 9820
rect 11789 9764 11845 9820
rect 11845 9764 11849 9820
rect 11785 9760 11849 9764
rect 11865 9820 11929 9824
rect 11865 9764 11869 9820
rect 11869 9764 11925 9820
rect 11925 9764 11929 9820
rect 11865 9760 11929 9764
rect 11945 9820 12009 9824
rect 11945 9764 11949 9820
rect 11949 9764 12005 9820
rect 12005 9764 12009 9820
rect 11945 9760 12009 9764
rect 12025 9820 12089 9824
rect 12025 9764 12029 9820
rect 12029 9764 12085 9820
rect 12085 9764 12089 9820
rect 12025 9760 12089 9764
rect 19375 9820 19439 9824
rect 19375 9764 19379 9820
rect 19379 9764 19435 9820
rect 19435 9764 19439 9820
rect 19375 9760 19439 9764
rect 19455 9820 19519 9824
rect 19455 9764 19459 9820
rect 19459 9764 19515 9820
rect 19515 9764 19519 9820
rect 19455 9760 19519 9764
rect 19535 9820 19599 9824
rect 19535 9764 19539 9820
rect 19539 9764 19595 9820
rect 19595 9764 19599 9820
rect 19535 9760 19599 9764
rect 19615 9820 19679 9824
rect 19615 9764 19619 9820
rect 19619 9764 19675 9820
rect 19675 9764 19679 9820
rect 19615 9760 19679 9764
rect 26965 9820 27029 9824
rect 26965 9764 26969 9820
rect 26969 9764 27025 9820
rect 27025 9764 27029 9820
rect 26965 9760 27029 9764
rect 27045 9820 27109 9824
rect 27045 9764 27049 9820
rect 27049 9764 27105 9820
rect 27105 9764 27109 9820
rect 27045 9760 27109 9764
rect 27125 9820 27189 9824
rect 27125 9764 27129 9820
rect 27129 9764 27185 9820
rect 27185 9764 27189 9820
rect 27125 9760 27189 9764
rect 27205 9820 27269 9824
rect 27205 9764 27209 9820
rect 27209 9764 27265 9820
rect 27265 9764 27269 9820
rect 27205 9760 27269 9764
rect 7990 9276 8054 9280
rect 7990 9220 7994 9276
rect 7994 9220 8050 9276
rect 8050 9220 8054 9276
rect 7990 9216 8054 9220
rect 8070 9276 8134 9280
rect 8070 9220 8074 9276
rect 8074 9220 8130 9276
rect 8130 9220 8134 9276
rect 8070 9216 8134 9220
rect 8150 9276 8214 9280
rect 8150 9220 8154 9276
rect 8154 9220 8210 9276
rect 8210 9220 8214 9276
rect 8150 9216 8214 9220
rect 8230 9276 8294 9280
rect 8230 9220 8234 9276
rect 8234 9220 8290 9276
rect 8290 9220 8294 9276
rect 8230 9216 8294 9220
rect 15580 9276 15644 9280
rect 15580 9220 15584 9276
rect 15584 9220 15640 9276
rect 15640 9220 15644 9276
rect 15580 9216 15644 9220
rect 15660 9276 15724 9280
rect 15660 9220 15664 9276
rect 15664 9220 15720 9276
rect 15720 9220 15724 9276
rect 15660 9216 15724 9220
rect 15740 9276 15804 9280
rect 15740 9220 15744 9276
rect 15744 9220 15800 9276
rect 15800 9220 15804 9276
rect 15740 9216 15804 9220
rect 15820 9276 15884 9280
rect 15820 9220 15824 9276
rect 15824 9220 15880 9276
rect 15880 9220 15884 9276
rect 15820 9216 15884 9220
rect 23170 9276 23234 9280
rect 23170 9220 23174 9276
rect 23174 9220 23230 9276
rect 23230 9220 23234 9276
rect 23170 9216 23234 9220
rect 23250 9276 23314 9280
rect 23250 9220 23254 9276
rect 23254 9220 23310 9276
rect 23310 9220 23314 9276
rect 23250 9216 23314 9220
rect 23330 9276 23394 9280
rect 23330 9220 23334 9276
rect 23334 9220 23390 9276
rect 23390 9220 23394 9276
rect 23330 9216 23394 9220
rect 23410 9276 23474 9280
rect 23410 9220 23414 9276
rect 23414 9220 23470 9276
rect 23470 9220 23474 9276
rect 23410 9216 23474 9220
rect 30760 9276 30824 9280
rect 30760 9220 30764 9276
rect 30764 9220 30820 9276
rect 30820 9220 30824 9276
rect 30760 9216 30824 9220
rect 30840 9276 30904 9280
rect 30840 9220 30844 9276
rect 30844 9220 30900 9276
rect 30900 9220 30904 9276
rect 30840 9216 30904 9220
rect 30920 9276 30984 9280
rect 30920 9220 30924 9276
rect 30924 9220 30980 9276
rect 30980 9220 30984 9276
rect 30920 9216 30984 9220
rect 31000 9276 31064 9280
rect 31000 9220 31004 9276
rect 31004 9220 31060 9276
rect 31060 9220 31064 9276
rect 31000 9216 31064 9220
rect 14044 8876 14108 8940
rect 4195 8732 4259 8736
rect 4195 8676 4199 8732
rect 4199 8676 4255 8732
rect 4255 8676 4259 8732
rect 4195 8672 4259 8676
rect 4275 8732 4339 8736
rect 4275 8676 4279 8732
rect 4279 8676 4335 8732
rect 4335 8676 4339 8732
rect 4275 8672 4339 8676
rect 4355 8732 4419 8736
rect 4355 8676 4359 8732
rect 4359 8676 4415 8732
rect 4415 8676 4419 8732
rect 4355 8672 4419 8676
rect 4435 8732 4499 8736
rect 4435 8676 4439 8732
rect 4439 8676 4495 8732
rect 4495 8676 4499 8732
rect 4435 8672 4499 8676
rect 11785 8732 11849 8736
rect 11785 8676 11789 8732
rect 11789 8676 11845 8732
rect 11845 8676 11849 8732
rect 11785 8672 11849 8676
rect 11865 8732 11929 8736
rect 11865 8676 11869 8732
rect 11869 8676 11925 8732
rect 11925 8676 11929 8732
rect 11865 8672 11929 8676
rect 11945 8732 12009 8736
rect 11945 8676 11949 8732
rect 11949 8676 12005 8732
rect 12005 8676 12009 8732
rect 11945 8672 12009 8676
rect 12025 8732 12089 8736
rect 12025 8676 12029 8732
rect 12029 8676 12085 8732
rect 12085 8676 12089 8732
rect 12025 8672 12089 8676
rect 19375 8732 19439 8736
rect 19375 8676 19379 8732
rect 19379 8676 19435 8732
rect 19435 8676 19439 8732
rect 19375 8672 19439 8676
rect 19455 8732 19519 8736
rect 19455 8676 19459 8732
rect 19459 8676 19515 8732
rect 19515 8676 19519 8732
rect 19455 8672 19519 8676
rect 19535 8732 19599 8736
rect 19535 8676 19539 8732
rect 19539 8676 19595 8732
rect 19595 8676 19599 8732
rect 19535 8672 19599 8676
rect 19615 8732 19679 8736
rect 19615 8676 19619 8732
rect 19619 8676 19675 8732
rect 19675 8676 19679 8732
rect 19615 8672 19679 8676
rect 26965 8732 27029 8736
rect 26965 8676 26969 8732
rect 26969 8676 27025 8732
rect 27025 8676 27029 8732
rect 26965 8672 27029 8676
rect 27045 8732 27109 8736
rect 27045 8676 27049 8732
rect 27049 8676 27105 8732
rect 27105 8676 27109 8732
rect 27045 8672 27109 8676
rect 27125 8732 27189 8736
rect 27125 8676 27129 8732
rect 27129 8676 27185 8732
rect 27185 8676 27189 8732
rect 27125 8672 27189 8676
rect 27205 8732 27269 8736
rect 27205 8676 27209 8732
rect 27209 8676 27265 8732
rect 27265 8676 27269 8732
rect 27205 8672 27269 8676
rect 7990 8188 8054 8192
rect 7990 8132 7994 8188
rect 7994 8132 8050 8188
rect 8050 8132 8054 8188
rect 7990 8128 8054 8132
rect 8070 8188 8134 8192
rect 8070 8132 8074 8188
rect 8074 8132 8130 8188
rect 8130 8132 8134 8188
rect 8070 8128 8134 8132
rect 8150 8188 8214 8192
rect 8150 8132 8154 8188
rect 8154 8132 8210 8188
rect 8210 8132 8214 8188
rect 8150 8128 8214 8132
rect 8230 8188 8294 8192
rect 8230 8132 8234 8188
rect 8234 8132 8290 8188
rect 8290 8132 8294 8188
rect 8230 8128 8294 8132
rect 15580 8188 15644 8192
rect 15580 8132 15584 8188
rect 15584 8132 15640 8188
rect 15640 8132 15644 8188
rect 15580 8128 15644 8132
rect 15660 8188 15724 8192
rect 15660 8132 15664 8188
rect 15664 8132 15720 8188
rect 15720 8132 15724 8188
rect 15660 8128 15724 8132
rect 15740 8188 15804 8192
rect 15740 8132 15744 8188
rect 15744 8132 15800 8188
rect 15800 8132 15804 8188
rect 15740 8128 15804 8132
rect 15820 8188 15884 8192
rect 15820 8132 15824 8188
rect 15824 8132 15880 8188
rect 15880 8132 15884 8188
rect 15820 8128 15884 8132
rect 23170 8188 23234 8192
rect 23170 8132 23174 8188
rect 23174 8132 23230 8188
rect 23230 8132 23234 8188
rect 23170 8128 23234 8132
rect 23250 8188 23314 8192
rect 23250 8132 23254 8188
rect 23254 8132 23310 8188
rect 23310 8132 23314 8188
rect 23250 8128 23314 8132
rect 23330 8188 23394 8192
rect 23330 8132 23334 8188
rect 23334 8132 23390 8188
rect 23390 8132 23394 8188
rect 23330 8128 23394 8132
rect 23410 8188 23474 8192
rect 23410 8132 23414 8188
rect 23414 8132 23470 8188
rect 23470 8132 23474 8188
rect 23410 8128 23474 8132
rect 30760 8188 30824 8192
rect 30760 8132 30764 8188
rect 30764 8132 30820 8188
rect 30820 8132 30824 8188
rect 30760 8128 30824 8132
rect 30840 8188 30904 8192
rect 30840 8132 30844 8188
rect 30844 8132 30900 8188
rect 30900 8132 30904 8188
rect 30840 8128 30904 8132
rect 30920 8188 30984 8192
rect 30920 8132 30924 8188
rect 30924 8132 30980 8188
rect 30980 8132 30984 8188
rect 30920 8128 30984 8132
rect 31000 8188 31064 8192
rect 31000 8132 31004 8188
rect 31004 8132 31060 8188
rect 31060 8132 31064 8188
rect 31000 8128 31064 8132
rect 4195 7644 4259 7648
rect 4195 7588 4199 7644
rect 4199 7588 4255 7644
rect 4255 7588 4259 7644
rect 4195 7584 4259 7588
rect 4275 7644 4339 7648
rect 4275 7588 4279 7644
rect 4279 7588 4335 7644
rect 4335 7588 4339 7644
rect 4275 7584 4339 7588
rect 4355 7644 4419 7648
rect 4355 7588 4359 7644
rect 4359 7588 4415 7644
rect 4415 7588 4419 7644
rect 4355 7584 4419 7588
rect 4435 7644 4499 7648
rect 4435 7588 4439 7644
rect 4439 7588 4495 7644
rect 4495 7588 4499 7644
rect 4435 7584 4499 7588
rect 11785 7644 11849 7648
rect 11785 7588 11789 7644
rect 11789 7588 11845 7644
rect 11845 7588 11849 7644
rect 11785 7584 11849 7588
rect 11865 7644 11929 7648
rect 11865 7588 11869 7644
rect 11869 7588 11925 7644
rect 11925 7588 11929 7644
rect 11865 7584 11929 7588
rect 11945 7644 12009 7648
rect 11945 7588 11949 7644
rect 11949 7588 12005 7644
rect 12005 7588 12009 7644
rect 11945 7584 12009 7588
rect 12025 7644 12089 7648
rect 12025 7588 12029 7644
rect 12029 7588 12085 7644
rect 12085 7588 12089 7644
rect 12025 7584 12089 7588
rect 12388 7788 12452 7852
rect 19375 7644 19439 7648
rect 19375 7588 19379 7644
rect 19379 7588 19435 7644
rect 19435 7588 19439 7644
rect 19375 7584 19439 7588
rect 19455 7644 19519 7648
rect 19455 7588 19459 7644
rect 19459 7588 19515 7644
rect 19515 7588 19519 7644
rect 19455 7584 19519 7588
rect 19535 7644 19599 7648
rect 19535 7588 19539 7644
rect 19539 7588 19595 7644
rect 19595 7588 19599 7644
rect 19535 7584 19599 7588
rect 19615 7644 19679 7648
rect 19615 7588 19619 7644
rect 19619 7588 19675 7644
rect 19675 7588 19679 7644
rect 19615 7584 19679 7588
rect 26965 7644 27029 7648
rect 26965 7588 26969 7644
rect 26969 7588 27025 7644
rect 27025 7588 27029 7644
rect 26965 7584 27029 7588
rect 27045 7644 27109 7648
rect 27045 7588 27049 7644
rect 27049 7588 27105 7644
rect 27105 7588 27109 7644
rect 27045 7584 27109 7588
rect 27125 7644 27189 7648
rect 27125 7588 27129 7644
rect 27129 7588 27185 7644
rect 27185 7588 27189 7644
rect 27125 7584 27189 7588
rect 27205 7644 27269 7648
rect 27205 7588 27209 7644
rect 27209 7588 27265 7644
rect 27265 7588 27269 7644
rect 27205 7584 27269 7588
rect 9444 7168 9508 7172
rect 9444 7112 9458 7168
rect 9458 7112 9508 7168
rect 9444 7108 9508 7112
rect 7990 7100 8054 7104
rect 7990 7044 7994 7100
rect 7994 7044 8050 7100
rect 8050 7044 8054 7100
rect 7990 7040 8054 7044
rect 8070 7100 8134 7104
rect 8070 7044 8074 7100
rect 8074 7044 8130 7100
rect 8130 7044 8134 7100
rect 8070 7040 8134 7044
rect 8150 7100 8214 7104
rect 8150 7044 8154 7100
rect 8154 7044 8210 7100
rect 8210 7044 8214 7100
rect 8150 7040 8214 7044
rect 8230 7100 8294 7104
rect 8230 7044 8234 7100
rect 8234 7044 8290 7100
rect 8290 7044 8294 7100
rect 8230 7040 8294 7044
rect 15580 7100 15644 7104
rect 15580 7044 15584 7100
rect 15584 7044 15640 7100
rect 15640 7044 15644 7100
rect 15580 7040 15644 7044
rect 15660 7100 15724 7104
rect 15660 7044 15664 7100
rect 15664 7044 15720 7100
rect 15720 7044 15724 7100
rect 15660 7040 15724 7044
rect 15740 7100 15804 7104
rect 15740 7044 15744 7100
rect 15744 7044 15800 7100
rect 15800 7044 15804 7100
rect 15740 7040 15804 7044
rect 15820 7100 15884 7104
rect 15820 7044 15824 7100
rect 15824 7044 15880 7100
rect 15880 7044 15884 7100
rect 15820 7040 15884 7044
rect 23170 7100 23234 7104
rect 23170 7044 23174 7100
rect 23174 7044 23230 7100
rect 23230 7044 23234 7100
rect 23170 7040 23234 7044
rect 23250 7100 23314 7104
rect 23250 7044 23254 7100
rect 23254 7044 23310 7100
rect 23310 7044 23314 7100
rect 23250 7040 23314 7044
rect 23330 7100 23394 7104
rect 23330 7044 23334 7100
rect 23334 7044 23390 7100
rect 23390 7044 23394 7100
rect 23330 7040 23394 7044
rect 23410 7100 23474 7104
rect 23410 7044 23414 7100
rect 23414 7044 23470 7100
rect 23470 7044 23474 7100
rect 23410 7040 23474 7044
rect 30760 7100 30824 7104
rect 30760 7044 30764 7100
rect 30764 7044 30820 7100
rect 30820 7044 30824 7100
rect 30760 7040 30824 7044
rect 30840 7100 30904 7104
rect 30840 7044 30844 7100
rect 30844 7044 30900 7100
rect 30900 7044 30904 7100
rect 30840 7040 30904 7044
rect 30920 7100 30984 7104
rect 30920 7044 30924 7100
rect 30924 7044 30980 7100
rect 30980 7044 30984 7100
rect 30920 7040 30984 7044
rect 31000 7100 31064 7104
rect 31000 7044 31004 7100
rect 31004 7044 31060 7100
rect 31060 7044 31064 7100
rect 31000 7040 31064 7044
rect 4195 6556 4259 6560
rect 4195 6500 4199 6556
rect 4199 6500 4255 6556
rect 4255 6500 4259 6556
rect 4195 6496 4259 6500
rect 4275 6556 4339 6560
rect 4275 6500 4279 6556
rect 4279 6500 4335 6556
rect 4335 6500 4339 6556
rect 4275 6496 4339 6500
rect 4355 6556 4419 6560
rect 4355 6500 4359 6556
rect 4359 6500 4415 6556
rect 4415 6500 4419 6556
rect 4355 6496 4419 6500
rect 4435 6556 4499 6560
rect 4435 6500 4439 6556
rect 4439 6500 4495 6556
rect 4495 6500 4499 6556
rect 4435 6496 4499 6500
rect 11785 6556 11849 6560
rect 11785 6500 11789 6556
rect 11789 6500 11845 6556
rect 11845 6500 11849 6556
rect 11785 6496 11849 6500
rect 11865 6556 11929 6560
rect 11865 6500 11869 6556
rect 11869 6500 11925 6556
rect 11925 6500 11929 6556
rect 11865 6496 11929 6500
rect 11945 6556 12009 6560
rect 11945 6500 11949 6556
rect 11949 6500 12005 6556
rect 12005 6500 12009 6556
rect 11945 6496 12009 6500
rect 12025 6556 12089 6560
rect 12025 6500 12029 6556
rect 12029 6500 12085 6556
rect 12085 6500 12089 6556
rect 12025 6496 12089 6500
rect 19375 6556 19439 6560
rect 19375 6500 19379 6556
rect 19379 6500 19435 6556
rect 19435 6500 19439 6556
rect 19375 6496 19439 6500
rect 19455 6556 19519 6560
rect 19455 6500 19459 6556
rect 19459 6500 19515 6556
rect 19515 6500 19519 6556
rect 19455 6496 19519 6500
rect 19535 6556 19599 6560
rect 19535 6500 19539 6556
rect 19539 6500 19595 6556
rect 19595 6500 19599 6556
rect 19535 6496 19599 6500
rect 19615 6556 19679 6560
rect 19615 6500 19619 6556
rect 19619 6500 19675 6556
rect 19675 6500 19679 6556
rect 19615 6496 19679 6500
rect 26965 6556 27029 6560
rect 26965 6500 26969 6556
rect 26969 6500 27025 6556
rect 27025 6500 27029 6556
rect 26965 6496 27029 6500
rect 27045 6556 27109 6560
rect 27045 6500 27049 6556
rect 27049 6500 27105 6556
rect 27105 6500 27109 6556
rect 27045 6496 27109 6500
rect 27125 6556 27189 6560
rect 27125 6500 27129 6556
rect 27129 6500 27185 6556
rect 27185 6500 27189 6556
rect 27125 6496 27189 6500
rect 27205 6556 27269 6560
rect 27205 6500 27209 6556
rect 27209 6500 27265 6556
rect 27265 6500 27269 6556
rect 27205 6496 27269 6500
rect 12204 6156 12268 6220
rect 7990 6012 8054 6016
rect 7990 5956 7994 6012
rect 7994 5956 8050 6012
rect 8050 5956 8054 6012
rect 7990 5952 8054 5956
rect 8070 6012 8134 6016
rect 8070 5956 8074 6012
rect 8074 5956 8130 6012
rect 8130 5956 8134 6012
rect 8070 5952 8134 5956
rect 8150 6012 8214 6016
rect 8150 5956 8154 6012
rect 8154 5956 8210 6012
rect 8210 5956 8214 6012
rect 8150 5952 8214 5956
rect 8230 6012 8294 6016
rect 8230 5956 8234 6012
rect 8234 5956 8290 6012
rect 8290 5956 8294 6012
rect 8230 5952 8294 5956
rect 15580 6012 15644 6016
rect 15580 5956 15584 6012
rect 15584 5956 15640 6012
rect 15640 5956 15644 6012
rect 15580 5952 15644 5956
rect 15660 6012 15724 6016
rect 15660 5956 15664 6012
rect 15664 5956 15720 6012
rect 15720 5956 15724 6012
rect 15660 5952 15724 5956
rect 15740 6012 15804 6016
rect 15740 5956 15744 6012
rect 15744 5956 15800 6012
rect 15800 5956 15804 6012
rect 15740 5952 15804 5956
rect 15820 6012 15884 6016
rect 15820 5956 15824 6012
rect 15824 5956 15880 6012
rect 15880 5956 15884 6012
rect 15820 5952 15884 5956
rect 23170 6012 23234 6016
rect 23170 5956 23174 6012
rect 23174 5956 23230 6012
rect 23230 5956 23234 6012
rect 23170 5952 23234 5956
rect 23250 6012 23314 6016
rect 23250 5956 23254 6012
rect 23254 5956 23310 6012
rect 23310 5956 23314 6012
rect 23250 5952 23314 5956
rect 23330 6012 23394 6016
rect 23330 5956 23334 6012
rect 23334 5956 23390 6012
rect 23390 5956 23394 6012
rect 23330 5952 23394 5956
rect 23410 6012 23474 6016
rect 23410 5956 23414 6012
rect 23414 5956 23470 6012
rect 23470 5956 23474 6012
rect 23410 5952 23474 5956
rect 30760 6012 30824 6016
rect 30760 5956 30764 6012
rect 30764 5956 30820 6012
rect 30820 5956 30824 6012
rect 30760 5952 30824 5956
rect 30840 6012 30904 6016
rect 30840 5956 30844 6012
rect 30844 5956 30900 6012
rect 30900 5956 30904 6012
rect 30840 5952 30904 5956
rect 30920 6012 30984 6016
rect 30920 5956 30924 6012
rect 30924 5956 30980 6012
rect 30980 5956 30984 6012
rect 30920 5952 30984 5956
rect 31000 6012 31064 6016
rect 31000 5956 31004 6012
rect 31004 5956 31060 6012
rect 31060 5956 31064 6012
rect 31000 5952 31064 5956
rect 4195 5468 4259 5472
rect 4195 5412 4199 5468
rect 4199 5412 4255 5468
rect 4255 5412 4259 5468
rect 4195 5408 4259 5412
rect 4275 5468 4339 5472
rect 4275 5412 4279 5468
rect 4279 5412 4335 5468
rect 4335 5412 4339 5468
rect 4275 5408 4339 5412
rect 4355 5468 4419 5472
rect 4355 5412 4359 5468
rect 4359 5412 4415 5468
rect 4415 5412 4419 5468
rect 4355 5408 4419 5412
rect 4435 5468 4499 5472
rect 4435 5412 4439 5468
rect 4439 5412 4495 5468
rect 4495 5412 4499 5468
rect 4435 5408 4499 5412
rect 11785 5468 11849 5472
rect 11785 5412 11789 5468
rect 11789 5412 11845 5468
rect 11845 5412 11849 5468
rect 11785 5408 11849 5412
rect 11865 5468 11929 5472
rect 11865 5412 11869 5468
rect 11869 5412 11925 5468
rect 11925 5412 11929 5468
rect 11865 5408 11929 5412
rect 11945 5468 12009 5472
rect 11945 5412 11949 5468
rect 11949 5412 12005 5468
rect 12005 5412 12009 5468
rect 11945 5408 12009 5412
rect 12025 5468 12089 5472
rect 12025 5412 12029 5468
rect 12029 5412 12085 5468
rect 12085 5412 12089 5468
rect 12025 5408 12089 5412
rect 19375 5468 19439 5472
rect 19375 5412 19379 5468
rect 19379 5412 19435 5468
rect 19435 5412 19439 5468
rect 19375 5408 19439 5412
rect 19455 5468 19519 5472
rect 19455 5412 19459 5468
rect 19459 5412 19515 5468
rect 19515 5412 19519 5468
rect 19455 5408 19519 5412
rect 19535 5468 19599 5472
rect 19535 5412 19539 5468
rect 19539 5412 19595 5468
rect 19595 5412 19599 5468
rect 19535 5408 19599 5412
rect 19615 5468 19679 5472
rect 19615 5412 19619 5468
rect 19619 5412 19675 5468
rect 19675 5412 19679 5468
rect 19615 5408 19679 5412
rect 26965 5468 27029 5472
rect 26965 5412 26969 5468
rect 26969 5412 27025 5468
rect 27025 5412 27029 5468
rect 26965 5408 27029 5412
rect 27045 5468 27109 5472
rect 27045 5412 27049 5468
rect 27049 5412 27105 5468
rect 27105 5412 27109 5468
rect 27045 5408 27109 5412
rect 27125 5468 27189 5472
rect 27125 5412 27129 5468
rect 27129 5412 27185 5468
rect 27185 5412 27189 5468
rect 27125 5408 27189 5412
rect 27205 5468 27269 5472
rect 27205 5412 27209 5468
rect 27209 5412 27265 5468
rect 27265 5412 27269 5468
rect 27205 5408 27269 5412
rect 7990 4924 8054 4928
rect 7990 4868 7994 4924
rect 7994 4868 8050 4924
rect 8050 4868 8054 4924
rect 7990 4864 8054 4868
rect 8070 4924 8134 4928
rect 8070 4868 8074 4924
rect 8074 4868 8130 4924
rect 8130 4868 8134 4924
rect 8070 4864 8134 4868
rect 8150 4924 8214 4928
rect 8150 4868 8154 4924
rect 8154 4868 8210 4924
rect 8210 4868 8214 4924
rect 8150 4864 8214 4868
rect 8230 4924 8294 4928
rect 8230 4868 8234 4924
rect 8234 4868 8290 4924
rect 8290 4868 8294 4924
rect 8230 4864 8294 4868
rect 15580 4924 15644 4928
rect 15580 4868 15584 4924
rect 15584 4868 15640 4924
rect 15640 4868 15644 4924
rect 15580 4864 15644 4868
rect 15660 4924 15724 4928
rect 15660 4868 15664 4924
rect 15664 4868 15720 4924
rect 15720 4868 15724 4924
rect 15660 4864 15724 4868
rect 15740 4924 15804 4928
rect 15740 4868 15744 4924
rect 15744 4868 15800 4924
rect 15800 4868 15804 4924
rect 15740 4864 15804 4868
rect 15820 4924 15884 4928
rect 15820 4868 15824 4924
rect 15824 4868 15880 4924
rect 15880 4868 15884 4924
rect 15820 4864 15884 4868
rect 23170 4924 23234 4928
rect 23170 4868 23174 4924
rect 23174 4868 23230 4924
rect 23230 4868 23234 4924
rect 23170 4864 23234 4868
rect 23250 4924 23314 4928
rect 23250 4868 23254 4924
rect 23254 4868 23310 4924
rect 23310 4868 23314 4924
rect 23250 4864 23314 4868
rect 23330 4924 23394 4928
rect 23330 4868 23334 4924
rect 23334 4868 23390 4924
rect 23390 4868 23394 4924
rect 23330 4864 23394 4868
rect 23410 4924 23474 4928
rect 23410 4868 23414 4924
rect 23414 4868 23470 4924
rect 23470 4868 23474 4924
rect 23410 4864 23474 4868
rect 30760 4924 30824 4928
rect 30760 4868 30764 4924
rect 30764 4868 30820 4924
rect 30820 4868 30824 4924
rect 30760 4864 30824 4868
rect 30840 4924 30904 4928
rect 30840 4868 30844 4924
rect 30844 4868 30900 4924
rect 30900 4868 30904 4924
rect 30840 4864 30904 4868
rect 30920 4924 30984 4928
rect 30920 4868 30924 4924
rect 30924 4868 30980 4924
rect 30980 4868 30984 4924
rect 30920 4864 30984 4868
rect 31000 4924 31064 4928
rect 31000 4868 31004 4924
rect 31004 4868 31060 4924
rect 31060 4868 31064 4924
rect 31000 4864 31064 4868
rect 4195 4380 4259 4384
rect 4195 4324 4199 4380
rect 4199 4324 4255 4380
rect 4255 4324 4259 4380
rect 4195 4320 4259 4324
rect 4275 4380 4339 4384
rect 4275 4324 4279 4380
rect 4279 4324 4335 4380
rect 4335 4324 4339 4380
rect 4275 4320 4339 4324
rect 4355 4380 4419 4384
rect 4355 4324 4359 4380
rect 4359 4324 4415 4380
rect 4415 4324 4419 4380
rect 4355 4320 4419 4324
rect 4435 4380 4499 4384
rect 4435 4324 4439 4380
rect 4439 4324 4495 4380
rect 4495 4324 4499 4380
rect 4435 4320 4499 4324
rect 11785 4380 11849 4384
rect 11785 4324 11789 4380
rect 11789 4324 11845 4380
rect 11845 4324 11849 4380
rect 11785 4320 11849 4324
rect 11865 4380 11929 4384
rect 11865 4324 11869 4380
rect 11869 4324 11925 4380
rect 11925 4324 11929 4380
rect 11865 4320 11929 4324
rect 11945 4380 12009 4384
rect 11945 4324 11949 4380
rect 11949 4324 12005 4380
rect 12005 4324 12009 4380
rect 11945 4320 12009 4324
rect 12025 4380 12089 4384
rect 12025 4324 12029 4380
rect 12029 4324 12085 4380
rect 12085 4324 12089 4380
rect 12025 4320 12089 4324
rect 19375 4380 19439 4384
rect 19375 4324 19379 4380
rect 19379 4324 19435 4380
rect 19435 4324 19439 4380
rect 19375 4320 19439 4324
rect 19455 4380 19519 4384
rect 19455 4324 19459 4380
rect 19459 4324 19515 4380
rect 19515 4324 19519 4380
rect 19455 4320 19519 4324
rect 19535 4380 19599 4384
rect 19535 4324 19539 4380
rect 19539 4324 19595 4380
rect 19595 4324 19599 4380
rect 19535 4320 19599 4324
rect 19615 4380 19679 4384
rect 19615 4324 19619 4380
rect 19619 4324 19675 4380
rect 19675 4324 19679 4380
rect 19615 4320 19679 4324
rect 26965 4380 27029 4384
rect 26965 4324 26969 4380
rect 26969 4324 27025 4380
rect 27025 4324 27029 4380
rect 26965 4320 27029 4324
rect 27045 4380 27109 4384
rect 27045 4324 27049 4380
rect 27049 4324 27105 4380
rect 27105 4324 27109 4380
rect 27045 4320 27109 4324
rect 27125 4380 27189 4384
rect 27125 4324 27129 4380
rect 27129 4324 27185 4380
rect 27185 4324 27189 4380
rect 27125 4320 27189 4324
rect 27205 4380 27269 4384
rect 27205 4324 27209 4380
rect 27209 4324 27265 4380
rect 27265 4324 27269 4380
rect 27205 4320 27269 4324
rect 8524 3980 8588 4044
rect 7990 3836 8054 3840
rect 7990 3780 7994 3836
rect 7994 3780 8050 3836
rect 8050 3780 8054 3836
rect 7990 3776 8054 3780
rect 8070 3836 8134 3840
rect 8070 3780 8074 3836
rect 8074 3780 8130 3836
rect 8130 3780 8134 3836
rect 8070 3776 8134 3780
rect 8150 3836 8214 3840
rect 8150 3780 8154 3836
rect 8154 3780 8210 3836
rect 8210 3780 8214 3836
rect 8150 3776 8214 3780
rect 8230 3836 8294 3840
rect 8230 3780 8234 3836
rect 8234 3780 8290 3836
rect 8290 3780 8294 3836
rect 8230 3776 8294 3780
rect 15580 3836 15644 3840
rect 15580 3780 15584 3836
rect 15584 3780 15640 3836
rect 15640 3780 15644 3836
rect 15580 3776 15644 3780
rect 15660 3836 15724 3840
rect 15660 3780 15664 3836
rect 15664 3780 15720 3836
rect 15720 3780 15724 3836
rect 15660 3776 15724 3780
rect 15740 3836 15804 3840
rect 15740 3780 15744 3836
rect 15744 3780 15800 3836
rect 15800 3780 15804 3836
rect 15740 3776 15804 3780
rect 15820 3836 15884 3840
rect 15820 3780 15824 3836
rect 15824 3780 15880 3836
rect 15880 3780 15884 3836
rect 15820 3776 15884 3780
rect 23170 3836 23234 3840
rect 23170 3780 23174 3836
rect 23174 3780 23230 3836
rect 23230 3780 23234 3836
rect 23170 3776 23234 3780
rect 23250 3836 23314 3840
rect 23250 3780 23254 3836
rect 23254 3780 23310 3836
rect 23310 3780 23314 3836
rect 23250 3776 23314 3780
rect 23330 3836 23394 3840
rect 23330 3780 23334 3836
rect 23334 3780 23390 3836
rect 23390 3780 23394 3836
rect 23330 3776 23394 3780
rect 23410 3836 23474 3840
rect 23410 3780 23414 3836
rect 23414 3780 23470 3836
rect 23470 3780 23474 3836
rect 23410 3776 23474 3780
rect 30760 3836 30824 3840
rect 30760 3780 30764 3836
rect 30764 3780 30820 3836
rect 30820 3780 30824 3836
rect 30760 3776 30824 3780
rect 30840 3836 30904 3840
rect 30840 3780 30844 3836
rect 30844 3780 30900 3836
rect 30900 3780 30904 3836
rect 30840 3776 30904 3780
rect 30920 3836 30984 3840
rect 30920 3780 30924 3836
rect 30924 3780 30980 3836
rect 30980 3780 30984 3836
rect 30920 3776 30984 3780
rect 31000 3836 31064 3840
rect 31000 3780 31004 3836
rect 31004 3780 31060 3836
rect 31060 3780 31064 3836
rect 31000 3776 31064 3780
rect 4195 3292 4259 3296
rect 4195 3236 4199 3292
rect 4199 3236 4255 3292
rect 4255 3236 4259 3292
rect 4195 3232 4259 3236
rect 4275 3292 4339 3296
rect 4275 3236 4279 3292
rect 4279 3236 4335 3292
rect 4335 3236 4339 3292
rect 4275 3232 4339 3236
rect 4355 3292 4419 3296
rect 4355 3236 4359 3292
rect 4359 3236 4415 3292
rect 4415 3236 4419 3292
rect 4355 3232 4419 3236
rect 4435 3292 4499 3296
rect 4435 3236 4439 3292
rect 4439 3236 4495 3292
rect 4495 3236 4499 3292
rect 4435 3232 4499 3236
rect 11785 3292 11849 3296
rect 11785 3236 11789 3292
rect 11789 3236 11845 3292
rect 11845 3236 11849 3292
rect 11785 3232 11849 3236
rect 11865 3292 11929 3296
rect 11865 3236 11869 3292
rect 11869 3236 11925 3292
rect 11925 3236 11929 3292
rect 11865 3232 11929 3236
rect 11945 3292 12009 3296
rect 11945 3236 11949 3292
rect 11949 3236 12005 3292
rect 12005 3236 12009 3292
rect 11945 3232 12009 3236
rect 12025 3292 12089 3296
rect 12025 3236 12029 3292
rect 12029 3236 12085 3292
rect 12085 3236 12089 3292
rect 12025 3232 12089 3236
rect 19375 3292 19439 3296
rect 19375 3236 19379 3292
rect 19379 3236 19435 3292
rect 19435 3236 19439 3292
rect 19375 3232 19439 3236
rect 19455 3292 19519 3296
rect 19455 3236 19459 3292
rect 19459 3236 19515 3292
rect 19515 3236 19519 3292
rect 19455 3232 19519 3236
rect 19535 3292 19599 3296
rect 19535 3236 19539 3292
rect 19539 3236 19595 3292
rect 19595 3236 19599 3292
rect 19535 3232 19599 3236
rect 19615 3292 19679 3296
rect 19615 3236 19619 3292
rect 19619 3236 19675 3292
rect 19675 3236 19679 3292
rect 19615 3232 19679 3236
rect 26965 3292 27029 3296
rect 26965 3236 26969 3292
rect 26969 3236 27025 3292
rect 27025 3236 27029 3292
rect 26965 3232 27029 3236
rect 27045 3292 27109 3296
rect 27045 3236 27049 3292
rect 27049 3236 27105 3292
rect 27105 3236 27109 3292
rect 27045 3232 27109 3236
rect 27125 3292 27189 3296
rect 27125 3236 27129 3292
rect 27129 3236 27185 3292
rect 27185 3236 27189 3292
rect 27125 3232 27189 3236
rect 27205 3292 27269 3296
rect 27205 3236 27209 3292
rect 27209 3236 27265 3292
rect 27265 3236 27269 3292
rect 27205 3232 27269 3236
rect 7990 2748 8054 2752
rect 7990 2692 7994 2748
rect 7994 2692 8050 2748
rect 8050 2692 8054 2748
rect 7990 2688 8054 2692
rect 8070 2748 8134 2752
rect 8070 2692 8074 2748
rect 8074 2692 8130 2748
rect 8130 2692 8134 2748
rect 8070 2688 8134 2692
rect 8150 2748 8214 2752
rect 8150 2692 8154 2748
rect 8154 2692 8210 2748
rect 8210 2692 8214 2748
rect 8150 2688 8214 2692
rect 8230 2748 8294 2752
rect 8230 2692 8234 2748
rect 8234 2692 8290 2748
rect 8290 2692 8294 2748
rect 8230 2688 8294 2692
rect 15580 2748 15644 2752
rect 15580 2692 15584 2748
rect 15584 2692 15640 2748
rect 15640 2692 15644 2748
rect 15580 2688 15644 2692
rect 15660 2748 15724 2752
rect 15660 2692 15664 2748
rect 15664 2692 15720 2748
rect 15720 2692 15724 2748
rect 15660 2688 15724 2692
rect 15740 2748 15804 2752
rect 15740 2692 15744 2748
rect 15744 2692 15800 2748
rect 15800 2692 15804 2748
rect 15740 2688 15804 2692
rect 15820 2748 15884 2752
rect 15820 2692 15824 2748
rect 15824 2692 15880 2748
rect 15880 2692 15884 2748
rect 15820 2688 15884 2692
rect 23170 2748 23234 2752
rect 23170 2692 23174 2748
rect 23174 2692 23230 2748
rect 23230 2692 23234 2748
rect 23170 2688 23234 2692
rect 23250 2748 23314 2752
rect 23250 2692 23254 2748
rect 23254 2692 23310 2748
rect 23310 2692 23314 2748
rect 23250 2688 23314 2692
rect 23330 2748 23394 2752
rect 23330 2692 23334 2748
rect 23334 2692 23390 2748
rect 23390 2692 23394 2748
rect 23330 2688 23394 2692
rect 23410 2748 23474 2752
rect 23410 2692 23414 2748
rect 23414 2692 23470 2748
rect 23470 2692 23474 2748
rect 23410 2688 23474 2692
rect 30760 2748 30824 2752
rect 30760 2692 30764 2748
rect 30764 2692 30820 2748
rect 30820 2692 30824 2748
rect 30760 2688 30824 2692
rect 30840 2748 30904 2752
rect 30840 2692 30844 2748
rect 30844 2692 30900 2748
rect 30900 2692 30904 2748
rect 30840 2688 30904 2692
rect 30920 2748 30984 2752
rect 30920 2692 30924 2748
rect 30924 2692 30980 2748
rect 30980 2692 30984 2748
rect 30920 2688 30984 2692
rect 31000 2748 31064 2752
rect 31000 2692 31004 2748
rect 31004 2692 31060 2748
rect 31060 2692 31064 2748
rect 31000 2688 31064 2692
rect 4195 2204 4259 2208
rect 4195 2148 4199 2204
rect 4199 2148 4255 2204
rect 4255 2148 4259 2204
rect 4195 2144 4259 2148
rect 4275 2204 4339 2208
rect 4275 2148 4279 2204
rect 4279 2148 4335 2204
rect 4335 2148 4339 2204
rect 4275 2144 4339 2148
rect 4355 2204 4419 2208
rect 4355 2148 4359 2204
rect 4359 2148 4415 2204
rect 4415 2148 4419 2204
rect 4355 2144 4419 2148
rect 4435 2204 4499 2208
rect 4435 2148 4439 2204
rect 4439 2148 4495 2204
rect 4495 2148 4499 2204
rect 4435 2144 4499 2148
rect 11785 2204 11849 2208
rect 11785 2148 11789 2204
rect 11789 2148 11845 2204
rect 11845 2148 11849 2204
rect 11785 2144 11849 2148
rect 11865 2204 11929 2208
rect 11865 2148 11869 2204
rect 11869 2148 11925 2204
rect 11925 2148 11929 2204
rect 11865 2144 11929 2148
rect 11945 2204 12009 2208
rect 11945 2148 11949 2204
rect 11949 2148 12005 2204
rect 12005 2148 12009 2204
rect 11945 2144 12009 2148
rect 12025 2204 12089 2208
rect 12025 2148 12029 2204
rect 12029 2148 12085 2204
rect 12085 2148 12089 2204
rect 12025 2144 12089 2148
rect 19375 2204 19439 2208
rect 19375 2148 19379 2204
rect 19379 2148 19435 2204
rect 19435 2148 19439 2204
rect 19375 2144 19439 2148
rect 19455 2204 19519 2208
rect 19455 2148 19459 2204
rect 19459 2148 19515 2204
rect 19515 2148 19519 2204
rect 19455 2144 19519 2148
rect 19535 2204 19599 2208
rect 19535 2148 19539 2204
rect 19539 2148 19595 2204
rect 19595 2148 19599 2204
rect 19535 2144 19599 2148
rect 19615 2204 19679 2208
rect 19615 2148 19619 2204
rect 19619 2148 19675 2204
rect 19675 2148 19679 2204
rect 19615 2144 19679 2148
rect 26965 2204 27029 2208
rect 26965 2148 26969 2204
rect 26969 2148 27025 2204
rect 27025 2148 27029 2204
rect 26965 2144 27029 2148
rect 27045 2204 27109 2208
rect 27045 2148 27049 2204
rect 27049 2148 27105 2204
rect 27105 2148 27109 2204
rect 27045 2144 27109 2148
rect 27125 2204 27189 2208
rect 27125 2148 27129 2204
rect 27129 2148 27185 2204
rect 27185 2148 27189 2204
rect 27125 2144 27189 2148
rect 27205 2204 27269 2208
rect 27205 2148 27209 2204
rect 27209 2148 27265 2204
rect 27265 2148 27269 2204
rect 27205 2144 27269 2148
rect 9444 2136 9508 2140
rect 9444 2080 9494 2136
rect 9494 2080 9508 2136
rect 9444 2076 9508 2080
rect 7990 1660 8054 1664
rect 7990 1604 7994 1660
rect 7994 1604 8050 1660
rect 8050 1604 8054 1660
rect 7990 1600 8054 1604
rect 8070 1660 8134 1664
rect 8070 1604 8074 1660
rect 8074 1604 8130 1660
rect 8130 1604 8134 1660
rect 8070 1600 8134 1604
rect 8150 1660 8214 1664
rect 8150 1604 8154 1660
rect 8154 1604 8210 1660
rect 8210 1604 8214 1660
rect 8150 1600 8214 1604
rect 8230 1660 8294 1664
rect 8230 1604 8234 1660
rect 8234 1604 8290 1660
rect 8290 1604 8294 1660
rect 8230 1600 8294 1604
rect 15580 1660 15644 1664
rect 15580 1604 15584 1660
rect 15584 1604 15640 1660
rect 15640 1604 15644 1660
rect 15580 1600 15644 1604
rect 15660 1660 15724 1664
rect 15660 1604 15664 1660
rect 15664 1604 15720 1660
rect 15720 1604 15724 1660
rect 15660 1600 15724 1604
rect 15740 1660 15804 1664
rect 15740 1604 15744 1660
rect 15744 1604 15800 1660
rect 15800 1604 15804 1660
rect 15740 1600 15804 1604
rect 15820 1660 15884 1664
rect 15820 1604 15824 1660
rect 15824 1604 15880 1660
rect 15880 1604 15884 1660
rect 15820 1600 15884 1604
rect 23170 1660 23234 1664
rect 23170 1604 23174 1660
rect 23174 1604 23230 1660
rect 23230 1604 23234 1660
rect 23170 1600 23234 1604
rect 23250 1660 23314 1664
rect 23250 1604 23254 1660
rect 23254 1604 23310 1660
rect 23310 1604 23314 1660
rect 23250 1600 23314 1604
rect 23330 1660 23394 1664
rect 23330 1604 23334 1660
rect 23334 1604 23390 1660
rect 23390 1604 23394 1660
rect 23330 1600 23394 1604
rect 23410 1660 23474 1664
rect 23410 1604 23414 1660
rect 23414 1604 23470 1660
rect 23470 1604 23474 1660
rect 23410 1600 23474 1604
rect 30760 1660 30824 1664
rect 30760 1604 30764 1660
rect 30764 1604 30820 1660
rect 30820 1604 30824 1660
rect 30760 1600 30824 1604
rect 30840 1660 30904 1664
rect 30840 1604 30844 1660
rect 30844 1604 30900 1660
rect 30900 1604 30904 1660
rect 30840 1600 30904 1604
rect 30920 1660 30984 1664
rect 30920 1604 30924 1660
rect 30924 1604 30980 1660
rect 30980 1604 30984 1660
rect 30920 1600 30984 1604
rect 31000 1660 31064 1664
rect 31000 1604 31004 1660
rect 31004 1604 31060 1660
rect 31060 1604 31064 1660
rect 31000 1600 31064 1604
rect 4195 1116 4259 1120
rect 4195 1060 4199 1116
rect 4199 1060 4255 1116
rect 4255 1060 4259 1116
rect 4195 1056 4259 1060
rect 4275 1116 4339 1120
rect 4275 1060 4279 1116
rect 4279 1060 4335 1116
rect 4335 1060 4339 1116
rect 4275 1056 4339 1060
rect 4355 1116 4419 1120
rect 4355 1060 4359 1116
rect 4359 1060 4415 1116
rect 4415 1060 4419 1116
rect 4355 1056 4419 1060
rect 4435 1116 4499 1120
rect 4435 1060 4439 1116
rect 4439 1060 4495 1116
rect 4495 1060 4499 1116
rect 4435 1056 4499 1060
rect 11785 1116 11849 1120
rect 11785 1060 11789 1116
rect 11789 1060 11845 1116
rect 11845 1060 11849 1116
rect 11785 1056 11849 1060
rect 11865 1116 11929 1120
rect 11865 1060 11869 1116
rect 11869 1060 11925 1116
rect 11925 1060 11929 1116
rect 11865 1056 11929 1060
rect 11945 1116 12009 1120
rect 11945 1060 11949 1116
rect 11949 1060 12005 1116
rect 12005 1060 12009 1116
rect 11945 1056 12009 1060
rect 12025 1116 12089 1120
rect 12025 1060 12029 1116
rect 12029 1060 12085 1116
rect 12085 1060 12089 1116
rect 12025 1056 12089 1060
rect 19375 1116 19439 1120
rect 19375 1060 19379 1116
rect 19379 1060 19435 1116
rect 19435 1060 19439 1116
rect 19375 1056 19439 1060
rect 19455 1116 19519 1120
rect 19455 1060 19459 1116
rect 19459 1060 19515 1116
rect 19515 1060 19519 1116
rect 19455 1056 19519 1060
rect 19535 1116 19599 1120
rect 19535 1060 19539 1116
rect 19539 1060 19595 1116
rect 19595 1060 19599 1116
rect 19535 1056 19599 1060
rect 19615 1116 19679 1120
rect 19615 1060 19619 1116
rect 19619 1060 19675 1116
rect 19675 1060 19679 1116
rect 19615 1056 19679 1060
rect 26965 1116 27029 1120
rect 26965 1060 26969 1116
rect 26969 1060 27025 1116
rect 27025 1060 27029 1116
rect 26965 1056 27029 1060
rect 27045 1116 27109 1120
rect 27045 1060 27049 1116
rect 27049 1060 27105 1116
rect 27105 1060 27109 1116
rect 27045 1056 27109 1060
rect 27125 1116 27189 1120
rect 27125 1060 27129 1116
rect 27129 1060 27185 1116
rect 27185 1060 27189 1116
rect 27125 1056 27189 1060
rect 27205 1116 27269 1120
rect 27205 1060 27209 1116
rect 27209 1060 27265 1116
rect 27265 1060 27269 1116
rect 27205 1056 27269 1060
rect 7990 572 8054 576
rect 7990 516 7994 572
rect 7994 516 8050 572
rect 8050 516 8054 572
rect 7990 512 8054 516
rect 8070 572 8134 576
rect 8070 516 8074 572
rect 8074 516 8130 572
rect 8130 516 8134 572
rect 8070 512 8134 516
rect 8150 572 8214 576
rect 8150 516 8154 572
rect 8154 516 8210 572
rect 8210 516 8214 572
rect 8150 512 8214 516
rect 8230 572 8294 576
rect 8230 516 8234 572
rect 8234 516 8290 572
rect 8290 516 8294 572
rect 8230 512 8294 516
rect 15580 572 15644 576
rect 15580 516 15584 572
rect 15584 516 15640 572
rect 15640 516 15644 572
rect 15580 512 15644 516
rect 15660 572 15724 576
rect 15660 516 15664 572
rect 15664 516 15720 572
rect 15720 516 15724 572
rect 15660 512 15724 516
rect 15740 572 15804 576
rect 15740 516 15744 572
rect 15744 516 15800 572
rect 15800 516 15804 572
rect 15740 512 15804 516
rect 15820 572 15884 576
rect 15820 516 15824 572
rect 15824 516 15880 572
rect 15880 516 15884 572
rect 15820 512 15884 516
rect 23170 572 23234 576
rect 23170 516 23174 572
rect 23174 516 23230 572
rect 23230 516 23234 572
rect 23170 512 23234 516
rect 23250 572 23314 576
rect 23250 516 23254 572
rect 23254 516 23310 572
rect 23310 516 23314 572
rect 23250 512 23314 516
rect 23330 572 23394 576
rect 23330 516 23334 572
rect 23334 516 23390 572
rect 23390 516 23394 572
rect 23330 512 23394 516
rect 23410 572 23474 576
rect 23410 516 23414 572
rect 23414 516 23470 572
rect 23470 516 23474 572
rect 23410 512 23474 516
rect 30760 572 30824 576
rect 30760 516 30764 572
rect 30764 516 30820 572
rect 30820 516 30824 572
rect 30760 512 30824 516
rect 30840 572 30904 576
rect 30840 516 30844 572
rect 30844 516 30900 572
rect 30900 516 30904 572
rect 30840 512 30904 516
rect 30920 572 30984 576
rect 30920 516 30924 572
rect 30924 516 30980 572
rect 30980 516 30984 572
rect 30920 512 30984 516
rect 31000 572 31064 576
rect 31000 516 31004 572
rect 31004 516 31060 572
rect 31060 516 31064 572
rect 31000 512 31064 516
<< metal4 >>
rect 4294 22130 4354 22304
rect 4478 22174 4722 22234
rect 4478 22130 4538 22174
rect 4294 22070 4538 22130
rect 4187 21792 4507 21808
rect 4187 21728 4195 21792
rect 4259 21728 4275 21792
rect 4339 21728 4355 21792
rect 4419 21728 4435 21792
rect 4499 21728 4507 21792
rect 4187 20704 4507 21728
rect 4187 20640 4195 20704
rect 4259 20640 4275 20704
rect 4339 20640 4355 20704
rect 4419 20640 4435 20704
rect 4499 20640 4507 20704
rect 4187 19616 4507 20640
rect 4187 19552 4195 19616
rect 4259 19552 4275 19616
rect 4339 19552 4355 19616
rect 4419 19552 4435 19616
rect 4499 19552 4507 19616
rect 2083 19412 2149 19413
rect 2083 19348 2084 19412
rect 2148 19348 2149 19412
rect 2083 19347 2149 19348
rect 2086 14381 2146 19347
rect 4187 18528 4507 19552
rect 4187 18464 4195 18528
rect 4259 18464 4275 18528
rect 4339 18464 4355 18528
rect 4419 18464 4435 18528
rect 4499 18464 4507 18528
rect 4187 17440 4507 18464
rect 4662 18189 4722 22174
rect 4659 18188 4725 18189
rect 4659 18124 4660 18188
rect 4724 18124 4725 18188
rect 4659 18123 4725 18124
rect 4846 18053 4906 22304
rect 5027 19004 5093 19005
rect 5027 18940 5028 19004
rect 5092 18940 5093 19004
rect 5027 18939 5093 18940
rect 4843 18052 4909 18053
rect 4843 17988 4844 18052
rect 4908 17988 4909 18052
rect 4843 17987 4909 17988
rect 4187 17376 4195 17440
rect 4259 17376 4275 17440
rect 4339 17376 4355 17440
rect 4419 17376 4435 17440
rect 4499 17376 4507 17440
rect 4187 16352 4507 17376
rect 4187 16288 4195 16352
rect 4259 16288 4275 16352
rect 4339 16288 4355 16352
rect 4419 16288 4435 16352
rect 4499 16288 4507 16352
rect 4187 15264 4507 16288
rect 4187 15200 4195 15264
rect 4259 15200 4275 15264
rect 4339 15200 4355 15264
rect 4419 15200 4435 15264
rect 4499 15200 4507 15264
rect 2083 14380 2149 14381
rect 2083 14316 2084 14380
rect 2148 14316 2149 14380
rect 2083 14315 2149 14316
rect 4187 14176 4507 15200
rect 4187 14112 4195 14176
rect 4259 14112 4275 14176
rect 4339 14112 4355 14176
rect 4419 14112 4435 14176
rect 4499 14112 4507 14176
rect 4187 13088 4507 14112
rect 5030 13293 5090 18939
rect 5398 18461 5458 22304
rect 5395 18460 5461 18461
rect 5395 18396 5396 18460
rect 5460 18396 5461 18460
rect 5395 18395 5461 18396
rect 5950 18053 6010 22304
rect 6502 22130 6562 22304
rect 6867 22132 6933 22133
rect 6867 22130 6868 22132
rect 6502 22070 6868 22130
rect 6867 22068 6868 22070
rect 6932 22068 6933 22132
rect 6867 22067 6933 22068
rect 6867 19412 6933 19413
rect 6867 19348 6868 19412
rect 6932 19348 6933 19412
rect 6867 19347 6933 19348
rect 5947 18052 6013 18053
rect 5947 17988 5948 18052
rect 6012 17988 6013 18052
rect 5947 17987 6013 17988
rect 6870 16557 6930 19347
rect 7054 19277 7114 22304
rect 7051 19276 7117 19277
rect 7051 19212 7052 19276
rect 7116 19212 7117 19276
rect 7051 19211 7117 19212
rect 7606 18869 7666 22304
rect 7790 22174 8034 22234
rect 7603 18868 7669 18869
rect 7603 18804 7604 18868
rect 7668 18804 7669 18868
rect 7603 18803 7669 18804
rect 7790 18733 7850 22174
rect 7974 22130 8034 22174
rect 8158 22130 8218 22304
rect 7974 22070 8218 22130
rect 7982 21248 8302 21808
rect 7982 21184 7990 21248
rect 8054 21184 8070 21248
rect 8134 21184 8150 21248
rect 8214 21184 8230 21248
rect 8294 21184 8302 21248
rect 7982 20160 8302 21184
rect 7982 20096 7990 20160
rect 8054 20096 8070 20160
rect 8134 20096 8150 20160
rect 8214 20096 8230 20160
rect 8294 20096 8302 20160
rect 7982 19072 8302 20096
rect 7982 19008 7990 19072
rect 8054 19008 8070 19072
rect 8134 19008 8150 19072
rect 8214 19008 8230 19072
rect 8294 19008 8302 19072
rect 7787 18732 7853 18733
rect 7787 18668 7788 18732
rect 7852 18668 7853 18732
rect 7787 18667 7853 18668
rect 7982 17984 8302 19008
rect 8710 18053 8770 22304
rect 8891 22268 8957 22269
rect 8891 22204 8892 22268
rect 8956 22234 8957 22268
rect 8956 22204 9138 22234
rect 8891 22203 9138 22204
rect 8894 22174 9138 22203
rect 9078 22130 9138 22174
rect 9262 22130 9322 22304
rect 9627 22268 9693 22269
rect 9627 22204 9628 22268
rect 9692 22204 9693 22268
rect 9627 22203 9693 22204
rect 9078 22070 9322 22130
rect 9630 22130 9690 22203
rect 9814 22130 9874 22304
rect 9630 22070 9874 22130
rect 10366 20637 10426 22304
rect 10363 20636 10429 20637
rect 10363 20572 10364 20636
rect 10428 20572 10429 20636
rect 10363 20571 10429 20572
rect 10918 20501 10978 22304
rect 11099 21588 11165 21589
rect 11099 21524 11100 21588
rect 11164 21524 11165 21588
rect 11099 21523 11165 21524
rect 8891 20500 8957 20501
rect 8891 20436 8892 20500
rect 8956 20436 8957 20500
rect 8891 20435 8957 20436
rect 10915 20500 10981 20501
rect 10915 20436 10916 20500
rect 10980 20436 10981 20500
rect 10915 20435 10981 20436
rect 8707 18052 8773 18053
rect 8707 17988 8708 18052
rect 8772 17988 8773 18052
rect 8707 17987 8773 17988
rect 7982 17920 7990 17984
rect 8054 17920 8070 17984
rect 8134 17920 8150 17984
rect 8214 17920 8230 17984
rect 8294 17920 8302 17984
rect 7982 16896 8302 17920
rect 7982 16832 7990 16896
rect 8054 16832 8070 16896
rect 8134 16832 8150 16896
rect 8214 16832 8230 16896
rect 8294 16832 8302 16896
rect 6867 16556 6933 16557
rect 6867 16492 6868 16556
rect 6932 16492 6933 16556
rect 6867 16491 6933 16492
rect 7982 15808 8302 16832
rect 7982 15744 7990 15808
rect 8054 15744 8070 15808
rect 8134 15744 8150 15808
rect 8214 15744 8230 15808
rect 8294 15744 8302 15808
rect 7982 14720 8302 15744
rect 8523 15468 8589 15469
rect 8523 15404 8524 15468
rect 8588 15404 8589 15468
rect 8523 15403 8589 15404
rect 7982 14656 7990 14720
rect 8054 14656 8070 14720
rect 8134 14656 8150 14720
rect 8214 14656 8230 14720
rect 8294 14656 8302 14720
rect 7982 13632 8302 14656
rect 7982 13568 7990 13632
rect 8054 13568 8070 13632
rect 8134 13568 8150 13632
rect 8214 13568 8230 13632
rect 8294 13568 8302 13632
rect 5027 13292 5093 13293
rect 5027 13228 5028 13292
rect 5092 13228 5093 13292
rect 5027 13227 5093 13228
rect 4187 13024 4195 13088
rect 4259 13024 4275 13088
rect 4339 13024 4355 13088
rect 4419 13024 4435 13088
rect 4499 13024 4507 13088
rect 4187 12000 4507 13024
rect 4187 11936 4195 12000
rect 4259 11936 4275 12000
rect 4339 11936 4355 12000
rect 4419 11936 4435 12000
rect 4499 11936 4507 12000
rect 4187 10912 4507 11936
rect 4187 10848 4195 10912
rect 4259 10848 4275 10912
rect 4339 10848 4355 10912
rect 4419 10848 4435 10912
rect 4499 10848 4507 10912
rect 4187 9824 4507 10848
rect 4187 9760 4195 9824
rect 4259 9760 4275 9824
rect 4339 9760 4355 9824
rect 4419 9760 4435 9824
rect 4499 9760 4507 9824
rect 4187 8736 4507 9760
rect 4187 8672 4195 8736
rect 4259 8672 4275 8736
rect 4339 8672 4355 8736
rect 4419 8672 4435 8736
rect 4499 8672 4507 8736
rect 4187 7648 4507 8672
rect 4187 7584 4195 7648
rect 4259 7584 4275 7648
rect 4339 7584 4355 7648
rect 4419 7584 4435 7648
rect 4499 7584 4507 7648
rect 4187 6560 4507 7584
rect 4187 6496 4195 6560
rect 4259 6496 4275 6560
rect 4339 6496 4355 6560
rect 4419 6496 4435 6560
rect 4499 6496 4507 6560
rect 4187 5472 4507 6496
rect 4187 5408 4195 5472
rect 4259 5408 4275 5472
rect 4339 5408 4355 5472
rect 4419 5408 4435 5472
rect 4499 5408 4507 5472
rect 4187 4384 4507 5408
rect 4187 4320 4195 4384
rect 4259 4320 4275 4384
rect 4339 4320 4355 4384
rect 4419 4320 4435 4384
rect 4499 4320 4507 4384
rect 4187 3296 4507 4320
rect 4187 3232 4195 3296
rect 4259 3232 4275 3296
rect 4339 3232 4355 3296
rect 4419 3232 4435 3296
rect 4499 3232 4507 3296
rect 4187 2208 4507 3232
rect 4187 2144 4195 2208
rect 4259 2144 4275 2208
rect 4339 2144 4355 2208
rect 4419 2144 4435 2208
rect 4499 2144 4507 2208
rect 4187 1120 4507 2144
rect 4187 1056 4195 1120
rect 4259 1056 4275 1120
rect 4339 1056 4355 1120
rect 4419 1056 4435 1120
rect 4499 1056 4507 1120
rect 4187 496 4507 1056
rect 7982 12544 8302 13568
rect 8526 13429 8586 15403
rect 8894 13701 8954 20435
rect 9443 19820 9509 19821
rect 9443 19756 9444 19820
rect 9508 19756 9509 19820
rect 9443 19755 9509 19756
rect 9446 14245 9506 19755
rect 10363 17372 10429 17373
rect 10363 17308 10364 17372
rect 10428 17308 10429 17372
rect 10363 17307 10429 17308
rect 9443 14244 9509 14245
rect 9443 14180 9444 14244
rect 9508 14180 9509 14244
rect 9443 14179 9509 14180
rect 8891 13700 8957 13701
rect 8891 13636 8892 13700
rect 8956 13636 8957 13700
rect 8891 13635 8957 13636
rect 8523 13428 8589 13429
rect 8523 13364 8524 13428
rect 8588 13364 8589 13428
rect 8523 13363 8589 13364
rect 7982 12480 7990 12544
rect 8054 12480 8070 12544
rect 8134 12480 8150 12544
rect 8214 12480 8230 12544
rect 8294 12480 8302 12544
rect 7982 11456 8302 12480
rect 7982 11392 7990 11456
rect 8054 11392 8070 11456
rect 8134 11392 8150 11456
rect 8214 11392 8230 11456
rect 8294 11392 8302 11456
rect 7982 10368 8302 11392
rect 8523 11388 8589 11389
rect 8523 11324 8524 11388
rect 8588 11324 8589 11388
rect 8523 11323 8589 11324
rect 7982 10304 7990 10368
rect 8054 10304 8070 10368
rect 8134 10304 8150 10368
rect 8214 10304 8230 10368
rect 8294 10304 8302 10368
rect 7982 9280 8302 10304
rect 7982 9216 7990 9280
rect 8054 9216 8070 9280
rect 8134 9216 8150 9280
rect 8214 9216 8230 9280
rect 8294 9216 8302 9280
rect 7982 8192 8302 9216
rect 7982 8128 7990 8192
rect 8054 8128 8070 8192
rect 8134 8128 8150 8192
rect 8214 8128 8230 8192
rect 8294 8128 8302 8192
rect 7982 7104 8302 8128
rect 7982 7040 7990 7104
rect 8054 7040 8070 7104
rect 8134 7040 8150 7104
rect 8214 7040 8230 7104
rect 8294 7040 8302 7104
rect 7982 6016 8302 7040
rect 7982 5952 7990 6016
rect 8054 5952 8070 6016
rect 8134 5952 8150 6016
rect 8214 5952 8230 6016
rect 8294 5952 8302 6016
rect 7982 4928 8302 5952
rect 7982 4864 7990 4928
rect 8054 4864 8070 4928
rect 8134 4864 8150 4928
rect 8214 4864 8230 4928
rect 8294 4864 8302 4928
rect 7982 3840 8302 4864
rect 8526 4045 8586 11323
rect 10366 11117 10426 17307
rect 11102 13701 11162 21523
rect 11470 19277 11530 22304
rect 12022 22130 12082 22304
rect 12022 22070 12450 22130
rect 12390 21997 12450 22070
rect 12387 21996 12453 21997
rect 12387 21932 12388 21996
rect 12452 21932 12453 21996
rect 12387 21931 12453 21932
rect 11777 21792 12097 21808
rect 11777 21728 11785 21792
rect 11849 21728 11865 21792
rect 11929 21728 11945 21792
rect 12009 21728 12025 21792
rect 12089 21728 12097 21792
rect 11777 20704 12097 21728
rect 11777 20640 11785 20704
rect 11849 20640 11865 20704
rect 11929 20640 11945 20704
rect 12009 20640 12025 20704
rect 12089 20640 12097 20704
rect 11777 19616 12097 20640
rect 11777 19552 11785 19616
rect 11849 19552 11865 19616
rect 11929 19552 11945 19616
rect 12009 19552 12025 19616
rect 12089 19552 12097 19616
rect 11467 19276 11533 19277
rect 11467 19212 11468 19276
rect 11532 19212 11533 19276
rect 11467 19211 11533 19212
rect 11777 18528 12097 19552
rect 11777 18464 11785 18528
rect 11849 18464 11865 18528
rect 11929 18464 11945 18528
rect 12009 18464 12025 18528
rect 12089 18464 12097 18528
rect 11777 17440 12097 18464
rect 12574 18189 12634 22304
rect 13126 21589 13186 22304
rect 13123 21588 13189 21589
rect 13123 21524 13124 21588
rect 13188 21524 13189 21588
rect 13123 21523 13189 21524
rect 13678 20501 13738 22304
rect 13675 20500 13741 20501
rect 13675 20436 13676 20500
rect 13740 20436 13741 20500
rect 13675 20435 13741 20436
rect 14230 19277 14290 22304
rect 14782 20770 14842 22304
rect 14598 20710 14842 20770
rect 14598 20365 14658 20710
rect 14595 20364 14661 20365
rect 14595 20300 14596 20364
rect 14660 20300 14661 20364
rect 14595 20299 14661 20300
rect 14227 19276 14293 19277
rect 14227 19212 14228 19276
rect 14292 19212 14293 19276
rect 14227 19211 14293 19212
rect 15334 19141 15394 22304
rect 15886 22130 15946 22304
rect 15886 22070 16130 22130
rect 15572 21248 15892 21808
rect 15572 21184 15580 21248
rect 15644 21184 15660 21248
rect 15724 21184 15740 21248
rect 15804 21184 15820 21248
rect 15884 21184 15892 21248
rect 15572 20160 15892 21184
rect 16070 20501 16130 22070
rect 16067 20500 16133 20501
rect 16067 20436 16068 20500
rect 16132 20436 16133 20500
rect 16067 20435 16133 20436
rect 15572 20096 15580 20160
rect 15644 20096 15660 20160
rect 15724 20096 15740 20160
rect 15804 20096 15820 20160
rect 15884 20096 15892 20160
rect 15331 19140 15397 19141
rect 15331 19076 15332 19140
rect 15396 19076 15397 19140
rect 15331 19075 15397 19076
rect 15572 19072 15892 20096
rect 16438 19277 16498 22304
rect 16990 21589 17050 22304
rect 17542 22104 17602 22304
rect 18094 22104 18154 22304
rect 18646 22104 18706 22304
rect 19198 22104 19258 22304
rect 19750 22104 19810 22304
rect 20302 22104 20362 22304
rect 20854 22104 20914 22304
rect 21406 22104 21466 22304
rect 21958 21997 22018 22304
rect 21955 21996 22021 21997
rect 21955 21932 21956 21996
rect 22020 21932 22021 21996
rect 21955 21931 22021 21932
rect 19367 21792 19687 21808
rect 19367 21728 19375 21792
rect 19439 21728 19455 21792
rect 19519 21728 19535 21792
rect 19599 21728 19615 21792
rect 19679 21728 19687 21792
rect 16987 21588 17053 21589
rect 16987 21524 16988 21588
rect 17052 21524 17053 21588
rect 16987 21523 17053 21524
rect 19367 20704 19687 21728
rect 22510 20773 22570 22304
rect 23062 21994 23122 22304
rect 23614 21997 23674 22304
rect 22878 21934 23122 21994
rect 23611 21996 23677 21997
rect 22878 20909 22938 21934
rect 23611 21932 23612 21996
rect 23676 21932 23677 21996
rect 23611 21931 23677 21932
rect 23162 21248 23482 21808
rect 23162 21184 23170 21248
rect 23234 21184 23250 21248
rect 23314 21184 23330 21248
rect 23394 21184 23410 21248
rect 23474 21184 23482 21248
rect 22875 20908 22941 20909
rect 22875 20844 22876 20908
rect 22940 20844 22941 20908
rect 22875 20843 22941 20844
rect 22507 20772 22573 20773
rect 22507 20708 22508 20772
rect 22572 20708 22573 20772
rect 22507 20707 22573 20708
rect 19367 20640 19375 20704
rect 19439 20640 19455 20704
rect 19519 20640 19535 20704
rect 19599 20640 19615 20704
rect 19679 20640 19687 20704
rect 19367 19616 19687 20640
rect 19367 19552 19375 19616
rect 19439 19552 19455 19616
rect 19519 19552 19535 19616
rect 19599 19552 19615 19616
rect 19679 19552 19687 19616
rect 16435 19276 16501 19277
rect 16435 19212 16436 19276
rect 16500 19212 16501 19276
rect 16435 19211 16501 19212
rect 15572 19008 15580 19072
rect 15644 19008 15660 19072
rect 15724 19008 15740 19072
rect 15804 19008 15820 19072
rect 15884 19008 15892 19072
rect 12571 18188 12637 18189
rect 12571 18124 12572 18188
rect 12636 18124 12637 18188
rect 12571 18123 12637 18124
rect 14043 18052 14109 18053
rect 14043 17988 14044 18052
rect 14108 17988 14109 18052
rect 14043 17987 14109 17988
rect 11777 17376 11785 17440
rect 11849 17376 11865 17440
rect 11929 17376 11945 17440
rect 12009 17376 12025 17440
rect 12089 17376 12097 17440
rect 11777 16352 12097 17376
rect 11777 16288 11785 16352
rect 11849 16288 11865 16352
rect 11929 16288 11945 16352
rect 12009 16288 12025 16352
rect 12089 16288 12097 16352
rect 11777 15264 12097 16288
rect 11777 15200 11785 15264
rect 11849 15200 11865 15264
rect 11929 15200 11945 15264
rect 12009 15200 12025 15264
rect 12089 15200 12097 15264
rect 11777 14176 12097 15200
rect 11777 14112 11785 14176
rect 11849 14112 11865 14176
rect 11929 14112 11945 14176
rect 12009 14112 12025 14176
rect 12089 14112 12097 14176
rect 11099 13700 11165 13701
rect 11099 13636 11100 13700
rect 11164 13636 11165 13700
rect 11099 13635 11165 13636
rect 11777 13088 12097 14112
rect 11777 13024 11785 13088
rect 11849 13024 11865 13088
rect 11929 13024 11945 13088
rect 12009 13024 12025 13088
rect 12089 13024 12097 13088
rect 11777 12000 12097 13024
rect 11777 11936 11785 12000
rect 11849 11936 11865 12000
rect 11929 11936 11945 12000
rect 12009 11936 12025 12000
rect 12089 11936 12097 12000
rect 10363 11116 10429 11117
rect 10363 11052 10364 11116
rect 10428 11052 10429 11116
rect 10363 11051 10429 11052
rect 11777 10912 12097 11936
rect 11777 10848 11785 10912
rect 11849 10848 11865 10912
rect 11929 10848 11945 10912
rect 12009 10848 12025 10912
rect 12089 10848 12097 10912
rect 11777 9824 12097 10848
rect 11777 9760 11785 9824
rect 11849 9760 11865 9824
rect 11929 9760 11945 9824
rect 12009 9760 12025 9824
rect 12089 9760 12097 9824
rect 11777 8736 12097 9760
rect 14046 8941 14106 17987
rect 15572 17984 15892 19008
rect 15572 17920 15580 17984
rect 15644 17920 15660 17984
rect 15724 17920 15740 17984
rect 15804 17920 15820 17984
rect 15884 17920 15892 17984
rect 15572 16896 15892 17920
rect 15572 16832 15580 16896
rect 15644 16832 15660 16896
rect 15724 16832 15740 16896
rect 15804 16832 15820 16896
rect 15884 16832 15892 16896
rect 15147 16692 15213 16693
rect 15147 16628 15148 16692
rect 15212 16628 15213 16692
rect 15147 16627 15213 16628
rect 15150 11661 15210 16627
rect 15572 15808 15892 16832
rect 15572 15744 15580 15808
rect 15644 15744 15660 15808
rect 15724 15744 15740 15808
rect 15804 15744 15820 15808
rect 15884 15744 15892 15808
rect 15572 14720 15892 15744
rect 15572 14656 15580 14720
rect 15644 14656 15660 14720
rect 15724 14656 15740 14720
rect 15804 14656 15820 14720
rect 15884 14656 15892 14720
rect 15572 13632 15892 14656
rect 15572 13568 15580 13632
rect 15644 13568 15660 13632
rect 15724 13568 15740 13632
rect 15804 13568 15820 13632
rect 15884 13568 15892 13632
rect 15572 12544 15892 13568
rect 15572 12480 15580 12544
rect 15644 12480 15660 12544
rect 15724 12480 15740 12544
rect 15804 12480 15820 12544
rect 15884 12480 15892 12544
rect 15147 11660 15213 11661
rect 15147 11596 15148 11660
rect 15212 11596 15213 11660
rect 15147 11595 15213 11596
rect 15572 11456 15892 12480
rect 15572 11392 15580 11456
rect 15644 11392 15660 11456
rect 15724 11392 15740 11456
rect 15804 11392 15820 11456
rect 15884 11392 15892 11456
rect 15572 10368 15892 11392
rect 15572 10304 15580 10368
rect 15644 10304 15660 10368
rect 15724 10304 15740 10368
rect 15804 10304 15820 10368
rect 15884 10304 15892 10368
rect 15572 9280 15892 10304
rect 15572 9216 15580 9280
rect 15644 9216 15660 9280
rect 15724 9216 15740 9280
rect 15804 9216 15820 9280
rect 15884 9216 15892 9280
rect 14043 8940 14109 8941
rect 14043 8876 14044 8940
rect 14108 8876 14109 8940
rect 14043 8875 14109 8876
rect 11777 8672 11785 8736
rect 11849 8672 11865 8736
rect 11929 8672 11945 8736
rect 12009 8672 12025 8736
rect 12089 8672 12097 8736
rect 11777 7648 12097 8672
rect 15572 8192 15892 9216
rect 15572 8128 15580 8192
rect 15644 8128 15660 8192
rect 15724 8128 15740 8192
rect 15804 8128 15820 8192
rect 15884 8128 15892 8192
rect 12387 7852 12453 7853
rect 12387 7850 12388 7852
rect 11777 7584 11785 7648
rect 11849 7584 11865 7648
rect 11929 7584 11945 7648
rect 12009 7584 12025 7648
rect 12089 7584 12097 7648
rect 9443 7172 9509 7173
rect 9443 7108 9444 7172
rect 9508 7108 9509 7172
rect 9443 7107 9509 7108
rect 8523 4044 8589 4045
rect 8523 3980 8524 4044
rect 8588 3980 8589 4044
rect 8523 3979 8589 3980
rect 7982 3776 7990 3840
rect 8054 3776 8070 3840
rect 8134 3776 8150 3840
rect 8214 3776 8230 3840
rect 8294 3776 8302 3840
rect 7982 2752 8302 3776
rect 7982 2688 7990 2752
rect 8054 2688 8070 2752
rect 8134 2688 8150 2752
rect 8214 2688 8230 2752
rect 8294 2688 8302 2752
rect 7982 1664 8302 2688
rect 9446 2141 9506 7107
rect 11777 6560 12097 7584
rect 11777 6496 11785 6560
rect 11849 6496 11865 6560
rect 11929 6496 11945 6560
rect 12009 6496 12025 6560
rect 12089 6496 12097 6560
rect 11777 5472 12097 6496
rect 12206 7790 12388 7850
rect 12206 6221 12266 7790
rect 12387 7788 12388 7790
rect 12452 7788 12453 7852
rect 12387 7787 12453 7788
rect 15572 7104 15892 8128
rect 15572 7040 15580 7104
rect 15644 7040 15660 7104
rect 15724 7040 15740 7104
rect 15804 7040 15820 7104
rect 15884 7040 15892 7104
rect 12203 6220 12269 6221
rect 12203 6156 12204 6220
rect 12268 6156 12269 6220
rect 12203 6155 12269 6156
rect 11777 5408 11785 5472
rect 11849 5408 11865 5472
rect 11929 5408 11945 5472
rect 12009 5408 12025 5472
rect 12089 5408 12097 5472
rect 11777 4384 12097 5408
rect 11777 4320 11785 4384
rect 11849 4320 11865 4384
rect 11929 4320 11945 4384
rect 12009 4320 12025 4384
rect 12089 4320 12097 4384
rect 11777 3296 12097 4320
rect 11777 3232 11785 3296
rect 11849 3232 11865 3296
rect 11929 3232 11945 3296
rect 12009 3232 12025 3296
rect 12089 3232 12097 3296
rect 11777 2208 12097 3232
rect 11777 2144 11785 2208
rect 11849 2144 11865 2208
rect 11929 2144 11945 2208
rect 12009 2144 12025 2208
rect 12089 2144 12097 2208
rect 9443 2140 9509 2141
rect 9443 2076 9444 2140
rect 9508 2076 9509 2140
rect 9443 2075 9509 2076
rect 7982 1600 7990 1664
rect 8054 1600 8070 1664
rect 8134 1600 8150 1664
rect 8214 1600 8230 1664
rect 8294 1600 8302 1664
rect 7982 576 8302 1600
rect 7982 512 7990 576
rect 8054 512 8070 576
rect 8134 512 8150 576
rect 8214 512 8230 576
rect 8294 512 8302 576
rect 7982 496 8302 512
rect 11777 1120 12097 2144
rect 11777 1056 11785 1120
rect 11849 1056 11865 1120
rect 11929 1056 11945 1120
rect 12009 1056 12025 1120
rect 12089 1056 12097 1120
rect 11777 496 12097 1056
rect 15572 6016 15892 7040
rect 15572 5952 15580 6016
rect 15644 5952 15660 6016
rect 15724 5952 15740 6016
rect 15804 5952 15820 6016
rect 15884 5952 15892 6016
rect 15572 4928 15892 5952
rect 15572 4864 15580 4928
rect 15644 4864 15660 4928
rect 15724 4864 15740 4928
rect 15804 4864 15820 4928
rect 15884 4864 15892 4928
rect 15572 3840 15892 4864
rect 15572 3776 15580 3840
rect 15644 3776 15660 3840
rect 15724 3776 15740 3840
rect 15804 3776 15820 3840
rect 15884 3776 15892 3840
rect 15572 2752 15892 3776
rect 15572 2688 15580 2752
rect 15644 2688 15660 2752
rect 15724 2688 15740 2752
rect 15804 2688 15820 2752
rect 15884 2688 15892 2752
rect 15572 1664 15892 2688
rect 15572 1600 15580 1664
rect 15644 1600 15660 1664
rect 15724 1600 15740 1664
rect 15804 1600 15820 1664
rect 15884 1600 15892 1664
rect 15572 576 15892 1600
rect 15572 512 15580 576
rect 15644 512 15660 576
rect 15724 512 15740 576
rect 15804 512 15820 576
rect 15884 512 15892 576
rect 15572 496 15892 512
rect 19367 18528 19687 19552
rect 19367 18464 19375 18528
rect 19439 18464 19455 18528
rect 19519 18464 19535 18528
rect 19599 18464 19615 18528
rect 19679 18464 19687 18528
rect 19367 17440 19687 18464
rect 19367 17376 19375 17440
rect 19439 17376 19455 17440
rect 19519 17376 19535 17440
rect 19599 17376 19615 17440
rect 19679 17376 19687 17440
rect 19367 16352 19687 17376
rect 19367 16288 19375 16352
rect 19439 16288 19455 16352
rect 19519 16288 19535 16352
rect 19599 16288 19615 16352
rect 19679 16288 19687 16352
rect 19367 15264 19687 16288
rect 19367 15200 19375 15264
rect 19439 15200 19455 15264
rect 19519 15200 19535 15264
rect 19599 15200 19615 15264
rect 19679 15200 19687 15264
rect 19367 14176 19687 15200
rect 19367 14112 19375 14176
rect 19439 14112 19455 14176
rect 19519 14112 19535 14176
rect 19599 14112 19615 14176
rect 19679 14112 19687 14176
rect 19367 13088 19687 14112
rect 19367 13024 19375 13088
rect 19439 13024 19455 13088
rect 19519 13024 19535 13088
rect 19599 13024 19615 13088
rect 19679 13024 19687 13088
rect 19367 12000 19687 13024
rect 19367 11936 19375 12000
rect 19439 11936 19455 12000
rect 19519 11936 19535 12000
rect 19599 11936 19615 12000
rect 19679 11936 19687 12000
rect 19367 10912 19687 11936
rect 19367 10848 19375 10912
rect 19439 10848 19455 10912
rect 19519 10848 19535 10912
rect 19599 10848 19615 10912
rect 19679 10848 19687 10912
rect 19367 9824 19687 10848
rect 19367 9760 19375 9824
rect 19439 9760 19455 9824
rect 19519 9760 19535 9824
rect 19599 9760 19615 9824
rect 19679 9760 19687 9824
rect 19367 8736 19687 9760
rect 19367 8672 19375 8736
rect 19439 8672 19455 8736
rect 19519 8672 19535 8736
rect 19599 8672 19615 8736
rect 19679 8672 19687 8736
rect 19367 7648 19687 8672
rect 19367 7584 19375 7648
rect 19439 7584 19455 7648
rect 19519 7584 19535 7648
rect 19599 7584 19615 7648
rect 19679 7584 19687 7648
rect 19367 6560 19687 7584
rect 19367 6496 19375 6560
rect 19439 6496 19455 6560
rect 19519 6496 19535 6560
rect 19599 6496 19615 6560
rect 19679 6496 19687 6560
rect 19367 5472 19687 6496
rect 19367 5408 19375 5472
rect 19439 5408 19455 5472
rect 19519 5408 19535 5472
rect 19599 5408 19615 5472
rect 19679 5408 19687 5472
rect 19367 4384 19687 5408
rect 19367 4320 19375 4384
rect 19439 4320 19455 4384
rect 19519 4320 19535 4384
rect 19599 4320 19615 4384
rect 19679 4320 19687 4384
rect 19367 3296 19687 4320
rect 19367 3232 19375 3296
rect 19439 3232 19455 3296
rect 19519 3232 19535 3296
rect 19599 3232 19615 3296
rect 19679 3232 19687 3296
rect 19367 2208 19687 3232
rect 19367 2144 19375 2208
rect 19439 2144 19455 2208
rect 19519 2144 19535 2208
rect 19599 2144 19615 2208
rect 19679 2144 19687 2208
rect 19367 1120 19687 2144
rect 19367 1056 19375 1120
rect 19439 1056 19455 1120
rect 19519 1056 19535 1120
rect 19599 1056 19615 1120
rect 19679 1056 19687 1120
rect 19367 496 19687 1056
rect 23162 20160 23482 21184
rect 24166 20773 24226 22304
rect 24163 20772 24229 20773
rect 24163 20708 24164 20772
rect 24228 20708 24229 20772
rect 24163 20707 24229 20708
rect 23162 20096 23170 20160
rect 23234 20096 23250 20160
rect 23314 20096 23330 20160
rect 23394 20096 23410 20160
rect 23474 20096 23482 20160
rect 23162 19072 23482 20096
rect 23162 19008 23170 19072
rect 23234 19008 23250 19072
rect 23314 19008 23330 19072
rect 23394 19008 23410 19072
rect 23474 19008 23482 19072
rect 23162 17984 23482 19008
rect 24718 18189 24778 22304
rect 24902 22174 25146 22234
rect 24902 21453 24962 22174
rect 25086 22130 25146 22174
rect 25270 22130 25330 22304
rect 25086 22070 25330 22130
rect 25451 22132 25517 22133
rect 25451 22068 25452 22132
rect 25516 22130 25517 22132
rect 25822 22130 25882 22304
rect 25516 22070 25882 22130
rect 25516 22068 25517 22070
rect 25451 22067 25517 22068
rect 24899 21452 24965 21453
rect 24899 21388 24900 21452
rect 24964 21388 24965 21452
rect 24899 21387 24965 21388
rect 26374 21181 26434 22304
rect 26926 22104 26986 22304
rect 27478 22104 27538 22304
rect 26957 21792 27277 21808
rect 26957 21728 26965 21792
rect 27029 21728 27045 21792
rect 27109 21728 27125 21792
rect 27189 21728 27205 21792
rect 27269 21728 27277 21792
rect 26371 21180 26437 21181
rect 26371 21116 26372 21180
rect 26436 21116 26437 21180
rect 26371 21115 26437 21116
rect 26957 20704 27277 21728
rect 26957 20640 26965 20704
rect 27029 20640 27045 20704
rect 27109 20640 27125 20704
rect 27189 20640 27205 20704
rect 27269 20640 27277 20704
rect 26957 19616 27277 20640
rect 26957 19552 26965 19616
rect 27029 19552 27045 19616
rect 27109 19552 27125 19616
rect 27189 19552 27205 19616
rect 27269 19552 27277 19616
rect 26957 18528 27277 19552
rect 26957 18464 26965 18528
rect 27029 18464 27045 18528
rect 27109 18464 27125 18528
rect 27189 18464 27205 18528
rect 27269 18464 27277 18528
rect 24715 18188 24781 18189
rect 24715 18124 24716 18188
rect 24780 18124 24781 18188
rect 24715 18123 24781 18124
rect 23162 17920 23170 17984
rect 23234 17920 23250 17984
rect 23314 17920 23330 17984
rect 23394 17920 23410 17984
rect 23474 17920 23482 17984
rect 23162 16896 23482 17920
rect 23162 16832 23170 16896
rect 23234 16832 23250 16896
rect 23314 16832 23330 16896
rect 23394 16832 23410 16896
rect 23474 16832 23482 16896
rect 23162 15808 23482 16832
rect 26957 17440 27277 18464
rect 26957 17376 26965 17440
rect 27029 17376 27045 17440
rect 27109 17376 27125 17440
rect 27189 17376 27205 17440
rect 27269 17376 27277 17440
rect 23979 16556 24045 16557
rect 23979 16492 23980 16556
rect 24044 16492 24045 16556
rect 23979 16491 24045 16492
rect 23162 15744 23170 15808
rect 23234 15744 23250 15808
rect 23314 15744 23330 15808
rect 23394 15744 23410 15808
rect 23474 15744 23482 15808
rect 23162 14720 23482 15744
rect 23162 14656 23170 14720
rect 23234 14656 23250 14720
rect 23314 14656 23330 14720
rect 23394 14656 23410 14720
rect 23474 14656 23482 14720
rect 23162 13632 23482 14656
rect 23162 13568 23170 13632
rect 23234 13568 23250 13632
rect 23314 13568 23330 13632
rect 23394 13568 23410 13632
rect 23474 13568 23482 13632
rect 23162 12544 23482 13568
rect 23162 12480 23170 12544
rect 23234 12480 23250 12544
rect 23314 12480 23330 12544
rect 23394 12480 23410 12544
rect 23474 12480 23482 12544
rect 23162 11456 23482 12480
rect 23982 11797 24042 16491
rect 26957 16352 27277 17376
rect 26957 16288 26965 16352
rect 27029 16288 27045 16352
rect 27109 16288 27125 16352
rect 27189 16288 27205 16352
rect 27269 16288 27277 16352
rect 26957 15264 27277 16288
rect 30752 21248 31072 21808
rect 30752 21184 30760 21248
rect 30824 21184 30840 21248
rect 30904 21184 30920 21248
rect 30984 21184 31000 21248
rect 31064 21184 31072 21248
rect 30752 20160 31072 21184
rect 30752 20096 30760 20160
rect 30824 20096 30840 20160
rect 30904 20096 30920 20160
rect 30984 20096 31000 20160
rect 31064 20096 31072 20160
rect 30752 19072 31072 20096
rect 30752 19008 30760 19072
rect 30824 19008 30840 19072
rect 30904 19008 30920 19072
rect 30984 19008 31000 19072
rect 31064 19008 31072 19072
rect 30752 17984 31072 19008
rect 30752 17920 30760 17984
rect 30824 17920 30840 17984
rect 30904 17920 30920 17984
rect 30984 17920 31000 17984
rect 31064 17920 31072 17984
rect 30752 16896 31072 17920
rect 30752 16832 30760 16896
rect 30824 16832 30840 16896
rect 30904 16832 30920 16896
rect 30984 16832 31000 16896
rect 31064 16832 31072 16896
rect 27659 16284 27725 16285
rect 27659 16220 27660 16284
rect 27724 16220 27725 16284
rect 27659 16219 27725 16220
rect 26957 15200 26965 15264
rect 27029 15200 27045 15264
rect 27109 15200 27125 15264
rect 27189 15200 27205 15264
rect 27269 15200 27277 15264
rect 26957 14176 27277 15200
rect 26957 14112 26965 14176
rect 27029 14112 27045 14176
rect 27109 14112 27125 14176
rect 27189 14112 27205 14176
rect 27269 14112 27277 14176
rect 26957 13088 27277 14112
rect 26957 13024 26965 13088
rect 27029 13024 27045 13088
rect 27109 13024 27125 13088
rect 27189 13024 27205 13088
rect 27269 13024 27277 13088
rect 26957 12000 27277 13024
rect 27662 12749 27722 16219
rect 30752 15808 31072 16832
rect 30752 15744 30760 15808
rect 30824 15744 30840 15808
rect 30904 15744 30920 15808
rect 30984 15744 31000 15808
rect 31064 15744 31072 15808
rect 30752 14720 31072 15744
rect 30752 14656 30760 14720
rect 30824 14656 30840 14720
rect 30904 14656 30920 14720
rect 30984 14656 31000 14720
rect 31064 14656 31072 14720
rect 30752 13632 31072 14656
rect 30752 13568 30760 13632
rect 30824 13568 30840 13632
rect 30904 13568 30920 13632
rect 30984 13568 31000 13632
rect 31064 13568 31072 13632
rect 27659 12748 27725 12749
rect 27659 12684 27660 12748
rect 27724 12684 27725 12748
rect 27659 12683 27725 12684
rect 26957 11936 26965 12000
rect 27029 11936 27045 12000
rect 27109 11936 27125 12000
rect 27189 11936 27205 12000
rect 27269 11936 27277 12000
rect 23979 11796 24045 11797
rect 23979 11732 23980 11796
rect 24044 11732 24045 11796
rect 23979 11731 24045 11732
rect 23162 11392 23170 11456
rect 23234 11392 23250 11456
rect 23314 11392 23330 11456
rect 23394 11392 23410 11456
rect 23474 11392 23482 11456
rect 23162 10368 23482 11392
rect 23162 10304 23170 10368
rect 23234 10304 23250 10368
rect 23314 10304 23330 10368
rect 23394 10304 23410 10368
rect 23474 10304 23482 10368
rect 23162 9280 23482 10304
rect 23162 9216 23170 9280
rect 23234 9216 23250 9280
rect 23314 9216 23330 9280
rect 23394 9216 23410 9280
rect 23474 9216 23482 9280
rect 23162 8192 23482 9216
rect 23162 8128 23170 8192
rect 23234 8128 23250 8192
rect 23314 8128 23330 8192
rect 23394 8128 23410 8192
rect 23474 8128 23482 8192
rect 23162 7104 23482 8128
rect 23162 7040 23170 7104
rect 23234 7040 23250 7104
rect 23314 7040 23330 7104
rect 23394 7040 23410 7104
rect 23474 7040 23482 7104
rect 23162 6016 23482 7040
rect 23162 5952 23170 6016
rect 23234 5952 23250 6016
rect 23314 5952 23330 6016
rect 23394 5952 23410 6016
rect 23474 5952 23482 6016
rect 23162 4928 23482 5952
rect 23162 4864 23170 4928
rect 23234 4864 23250 4928
rect 23314 4864 23330 4928
rect 23394 4864 23410 4928
rect 23474 4864 23482 4928
rect 23162 3840 23482 4864
rect 23162 3776 23170 3840
rect 23234 3776 23250 3840
rect 23314 3776 23330 3840
rect 23394 3776 23410 3840
rect 23474 3776 23482 3840
rect 23162 2752 23482 3776
rect 23162 2688 23170 2752
rect 23234 2688 23250 2752
rect 23314 2688 23330 2752
rect 23394 2688 23410 2752
rect 23474 2688 23482 2752
rect 23162 1664 23482 2688
rect 23162 1600 23170 1664
rect 23234 1600 23250 1664
rect 23314 1600 23330 1664
rect 23394 1600 23410 1664
rect 23474 1600 23482 1664
rect 23162 576 23482 1600
rect 23162 512 23170 576
rect 23234 512 23250 576
rect 23314 512 23330 576
rect 23394 512 23410 576
rect 23474 512 23482 576
rect 23162 496 23482 512
rect 26957 10912 27277 11936
rect 26957 10848 26965 10912
rect 27029 10848 27045 10912
rect 27109 10848 27125 10912
rect 27189 10848 27205 10912
rect 27269 10848 27277 10912
rect 26957 9824 27277 10848
rect 26957 9760 26965 9824
rect 27029 9760 27045 9824
rect 27109 9760 27125 9824
rect 27189 9760 27205 9824
rect 27269 9760 27277 9824
rect 26957 8736 27277 9760
rect 26957 8672 26965 8736
rect 27029 8672 27045 8736
rect 27109 8672 27125 8736
rect 27189 8672 27205 8736
rect 27269 8672 27277 8736
rect 26957 7648 27277 8672
rect 26957 7584 26965 7648
rect 27029 7584 27045 7648
rect 27109 7584 27125 7648
rect 27189 7584 27205 7648
rect 27269 7584 27277 7648
rect 26957 6560 27277 7584
rect 26957 6496 26965 6560
rect 27029 6496 27045 6560
rect 27109 6496 27125 6560
rect 27189 6496 27205 6560
rect 27269 6496 27277 6560
rect 26957 5472 27277 6496
rect 26957 5408 26965 5472
rect 27029 5408 27045 5472
rect 27109 5408 27125 5472
rect 27189 5408 27205 5472
rect 27269 5408 27277 5472
rect 26957 4384 27277 5408
rect 26957 4320 26965 4384
rect 27029 4320 27045 4384
rect 27109 4320 27125 4384
rect 27189 4320 27205 4384
rect 27269 4320 27277 4384
rect 26957 3296 27277 4320
rect 26957 3232 26965 3296
rect 27029 3232 27045 3296
rect 27109 3232 27125 3296
rect 27189 3232 27205 3296
rect 27269 3232 27277 3296
rect 26957 2208 27277 3232
rect 26957 2144 26965 2208
rect 27029 2144 27045 2208
rect 27109 2144 27125 2208
rect 27189 2144 27205 2208
rect 27269 2144 27277 2208
rect 26957 1120 27277 2144
rect 26957 1056 26965 1120
rect 27029 1056 27045 1120
rect 27109 1056 27125 1120
rect 27189 1056 27205 1120
rect 27269 1056 27277 1120
rect 26957 496 27277 1056
rect 30752 12544 31072 13568
rect 30752 12480 30760 12544
rect 30824 12480 30840 12544
rect 30904 12480 30920 12544
rect 30984 12480 31000 12544
rect 31064 12480 31072 12544
rect 30752 11456 31072 12480
rect 30752 11392 30760 11456
rect 30824 11392 30840 11456
rect 30904 11392 30920 11456
rect 30984 11392 31000 11456
rect 31064 11392 31072 11456
rect 30752 10368 31072 11392
rect 30752 10304 30760 10368
rect 30824 10304 30840 10368
rect 30904 10304 30920 10368
rect 30984 10304 31000 10368
rect 31064 10304 31072 10368
rect 30752 9280 31072 10304
rect 30752 9216 30760 9280
rect 30824 9216 30840 9280
rect 30904 9216 30920 9280
rect 30984 9216 31000 9280
rect 31064 9216 31072 9280
rect 30752 8192 31072 9216
rect 30752 8128 30760 8192
rect 30824 8128 30840 8192
rect 30904 8128 30920 8192
rect 30984 8128 31000 8192
rect 31064 8128 31072 8192
rect 30752 7104 31072 8128
rect 30752 7040 30760 7104
rect 30824 7040 30840 7104
rect 30904 7040 30920 7104
rect 30984 7040 31000 7104
rect 31064 7040 31072 7104
rect 30752 6016 31072 7040
rect 30752 5952 30760 6016
rect 30824 5952 30840 6016
rect 30904 5952 30920 6016
rect 30984 5952 31000 6016
rect 31064 5952 31072 6016
rect 30752 4928 31072 5952
rect 30752 4864 30760 4928
rect 30824 4864 30840 4928
rect 30904 4864 30920 4928
rect 30984 4864 31000 4928
rect 31064 4864 31072 4928
rect 30752 3840 31072 4864
rect 30752 3776 30760 3840
rect 30824 3776 30840 3840
rect 30904 3776 30920 3840
rect 30984 3776 31000 3840
rect 31064 3776 31072 3840
rect 30752 2752 31072 3776
rect 30752 2688 30760 2752
rect 30824 2688 30840 2752
rect 30904 2688 30920 2752
rect 30984 2688 31000 2752
rect 31064 2688 31072 2752
rect 30752 1664 31072 2688
rect 30752 1600 30760 1664
rect 30824 1600 30840 1664
rect 30904 1600 30920 1664
rect 30984 1600 31000 1664
rect 31064 1600 31072 1664
rect 30752 576 31072 1600
rect 30752 512 30760 576
rect 30824 512 30840 576
rect 30904 512 30920 576
rect 30984 512 31000 576
rect 31064 512 31072 576
rect 30752 496 31072 512
use sky130_fd_sc_hd__inv_2  _05_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28612 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _06_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 21252 0 1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _07_
timestamp 1693170804
transform 1 0 23828 0 1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _08_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 23828 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _09_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 23184 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _10_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 18676 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _11_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 19136 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 11224 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _21_
timestamp 1693170804
transform 1 0 13432 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _22_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8096 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _23_
timestamp 1693170804
transform 1 0 12880 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _24_
timestamp 1693170804
transform 1 0 3312 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _25_
timestamp 1693170804
transform 1 0 2024 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _26_
timestamp 1693170804
transform 1 0 1472 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _27_
timestamp 1693170804
transform 1 0 8004 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 15364 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1693170804
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1693170804
transform 1 0 25024 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1693170804
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1693170804
transform 1 0 25484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1693170804
transform 1 0 29900 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1693170804
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1693170804
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1693170804
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1693170804
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1693170804
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1693170804
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1693170804
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1693170804
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1693170804
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1693170804
transform 1 0 25116 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1693170804
transform 1 0 1104 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1693170804
transform 1 0 19780 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1693170804
transform 1 0 5888 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1693170804
transform 1 0 5244 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1693170804
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1693170804
transform 1 0 4876 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1693170804
transform 1 0 1840 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1693170804
transform 1 0 3772 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1693170804
transform 1 0 2208 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1693170804
transform 1 0 3404 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__mux2i_2  ct.cw.cc_test_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28980 0 1 20128
box -38 -48 1050 592
use sky130_ht_sc_tt05__mux2i_2  ct.cw.cc_test_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699069426
transform 1 0 28980 0 1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__maj3_2  ct.cw.cc_test_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 29532 0 -1 16864
box -38 -48 866 592
use sky130_ht_sc_tt05__maj3_2  ct.cw.cc_test_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699069426
transform 1 0 28060 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dlrtp_1  ct.cw.cc_test_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28980 0 1 19040
box -38 -48 1234 592
use sky130_ht_sc_tt05__dlrtp_1  ct.cw.cc_test_5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699069426
transform 1 0 28980 0 1 17952
box -38 -48 1418 592
use sky130_fd_sc_hd__dfrtp_1  ct.cw.cc_test_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28612 0 -1 17952
box -38 -48 1878 592
use sky130_ht_sc_tt05__dfrtp_1  ct.cw.cc_test_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1699069426
transform 1 0 28612 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[0\].bits\[0\].cc_flop $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28612 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[0\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 16836 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[0\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[0\].cc_clkbuf
timestamp 1693170804
transform 1 0 28980 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[1\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[1\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 6164 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[1\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 14260 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[1\].cc_clkbuf
timestamp 1693170804
transform 1 0 29532 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[2\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[2\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[2\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 26772 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[2\].cc_clkbuf
timestamp 1693170804
transform 1 0 29992 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[3\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 16836 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[3\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[3\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 26864 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[3\].cc_clkbuf
timestamp 1693170804
transform 1 0 25760 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[4\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 26404 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[4\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 21988 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[4\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[4\].cc_clkbuf
timestamp 1693170804
transform 1 0 26036 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[5\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 26864 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[5\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 26864 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[5\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 26404 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[5\].cc_clkbuf
timestamp 1693170804
transform 1 0 23828 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[6\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 21804 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[6\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 23828 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[6\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 24380 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[6\].cc_clkbuf
timestamp 1693170804
transform 1 0 22540 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[7\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[7\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[7\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[7\].cc_clkbuf
timestamp 1693170804
transform 1 0 21252 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[8\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 18676 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[8\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 18676 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[8\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 19136 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[8\].cc_clkbuf
timestamp 1693170804
transform 1 0 20424 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[9\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 16928 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[9\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 16928 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[9\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 18676 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[9\].cc_clkbuf
timestamp 1693170804
transform 1 0 17848 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[10\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 16100 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[10\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 15824 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[10\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 15916 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[10\].cc_clkbuf
timestamp 1693170804
transform 1 0 16192 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[11\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 14260 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[11\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 16100 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[11\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 14260 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[11\].cc_clkbuf
timestamp 1693170804
transform 1 0 13708 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[0\].cc_scanflop $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 13524 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 12144 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 15732 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 8464 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8280 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 3128 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11868 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[0\].cc_clkbuf
timestamp 1693170804
transform 1 0 13524 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[0\].rs_mbuf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 7728 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 10856 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 10764 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 8464 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 10672 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 5888 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 13892 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 5428 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 12052 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 14168 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[1\].cc_clkbuf
timestamp 1693170804
transform 1 0 10948 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[1\].rs_mbuf
timestamp 1693170804
transform 1 0 5152 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 6164 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 28152 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 5888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 5980 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3036 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[2\].bits\[5\].rs_cbuf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9568 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[2\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10120 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 2576 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[2\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 9844 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[2\].cc_clkbuf
timestamp 1693170804
transform 1 0 4600 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[2\].rs_mbuf
timestamp 1693170804
transform 1 0 920 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16376 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 5888 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 7912 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 16376 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 2392 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 6532 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 828 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10396 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 10948 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[3\].cc_clkbuf
timestamp 1693170804
transform 1 0 3220 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[3\].rs_mbuf
timestamp 1693170804
transform 1 0 1104 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 4600 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 11500 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 8740 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 828 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[4\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 9752 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[4\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 9016 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[4\].cc_clkbuf
timestamp 1693170804
transform 1 0 1656 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[4\].rs_mbuf
timestamp 1693170804
transform 1 0 3220 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 3128 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3772 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 4324 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 14996 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 16744 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10488 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[5\].cc_clkbuf
timestamp 1693170804
transform 1 0 3220 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[5\].rs_mbuf
timestamp 1693170804
transform 1 0 3220 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5152 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 6256 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 9384 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 8464 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[6\].cc_clkbuf
timestamp 1693170804
transform 1 0 5796 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[6\].rs_mbuf
timestamp 1693170804
transform 1 0 9016 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 11500 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 10304 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 12696 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 11776 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 12972 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11776 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[7\].cc_clkbuf
timestamp 1693170804
transform 1 0 10948 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[7\].rs_mbuf
timestamp 1693170804
transform 1 0 11868 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 14168 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 13616 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 14536 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 15732 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 13892 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 14536 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 15732 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 14168 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 13984 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 13984 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 14168 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[8\].cc_clkbuf
timestamp 1693170804
transform 1 0 13524 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[8\].rs_mbuf
timestamp 1693170804
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 17020 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 18952 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 19228 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 17020 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 18676 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 16928 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 19136 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 19136 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 16928 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 16928 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 16376 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[9\].cc_clkbuf
timestamp 1693170804
transform 1 0 16100 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[9\].rs_mbuf
timestamp 1693170804
transform 1 0 18676 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 19596 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 19320 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 19596 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 19596 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 20148 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 20424 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 18952 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 20332 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 19228 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 20332 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 19504 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[10\].cc_clkbuf
timestamp 1693170804
transform 1 0 18676 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[10\].rs_mbuf
timestamp 1693170804
transform 1 0 19780 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 23000 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 23736 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 22724 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 24656 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 23552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 24656 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 25576 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 24380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[11\].cc_clkbuf
timestamp 1693170804
transform 1 0 22540 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[11\].rs_mbuf
timestamp 1693170804
transform 1 0 23184 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 26036 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 26036 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 25668 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 25852 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 27692 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 28612 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 21896 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 30176 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[12\].cc_clkbuf
timestamp 1693170804
transform 1 0 26404 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[12\].rs_mbuf
timestamp 1693170804
transform 1 0 27140 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 24472 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 23920 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 24196 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 23184 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 27324 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 28336 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 28428 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 29532 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[13\].cc_clkbuf
timestamp 1693170804
transform 1 0 28980 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[13\].rs_mbuf
timestamp 1693170804
transform 1 0 25760 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 22816 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 22172 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 21896 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 28612 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 29532 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 27968 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 29808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[14\].cc_clkbuf
timestamp 1693170804
transform 1 0 28980 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[14\].rs_mbuf
timestamp 1693170804
transform 1 0 25668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 20332 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 20792 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 19780 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 19872 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 20056 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 24656 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 27784 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 30268 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 27784 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[15\].cc_clkbuf
timestamp 1693170804
transform 1 0 26036 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[15\].rs_mbuf
timestamp 1693170804
transform 1 0 29532 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 19596 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 18952 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18032 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 18676 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 26312 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 28520 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 28244 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[16\].cc_clkbuf
timestamp 1693170804
transform 1 0 24104 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[16\].rs_mbuf
timestamp 1693170804
transform 1 0 17480 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 17204 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16928 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16836 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 17020 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 19964 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 21896 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 23092 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 24564 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 26036 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 26036 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 25944 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[17\].cc_clkbuf
timestamp 1693170804
transform 1 0 17848 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[17\].rs_mbuf
timestamp 1693170804
transform 1 0 19044 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16560 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 16836 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 19044 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 25668 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 22632 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 22908 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 23368 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[18\].cc_clkbuf
timestamp 1693170804
transform 1 0 20608 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[18\].rs_mbuf
timestamp 1693170804
transform 1 0 20240 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 17204 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18032 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 17756 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 17480 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 18032 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 20424 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 21712 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 21988 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[19\].cc_clkbuf
timestamp 1693170804
transform 1 0 17480 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[19\].rs_mbuf
timestamp 1693170804
transform 1 0 18032 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 24012 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 28428 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 27508 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26220 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 27968 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 30084 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 27968 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 27876 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[20\].cc_clkbuf
timestamp 1693170804
transform 1 0 23092 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[20\].rs_mbuf
timestamp 1693170804
transform 1 0 26404 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3772 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 1012 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__dlymetal6s2s_1  ct.oc.frame\[21\].bits\[1\].rs_cbuf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28980 0 1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 28152 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 18952 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[21\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 18952 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[21\].cc_clkbuf
timestamp 1693170804
transform 1 0 27232 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[21\].rs_mbuf
timestamp 1693170804
transform 1 0 27324 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 29440 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 26496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26312 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 25944 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 26312 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26036 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 28520 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 16744 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 27048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[22\].cc_clkbuf
timestamp 1693170804
transform 1 0 27232 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[22\].rs_mbuf
timestamp 1693170804
transform 1 0 26680 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[23\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 28888 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[23\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 29164 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 25208 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 24564 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 24012 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 25668 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 24012 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 25944 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 18952 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 28612 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 25484 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[23\].cc_clkbuf
timestamp 1693170804
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[23\].rs_mbuf
timestamp 1693170804
transform 1 0 24656 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 24104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 22172 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 23368 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 23092 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 22172 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 23092 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 24380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[24\].cc_clkbuf
timestamp 1693170804
transform 1 0 23460 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[24\].rs_mbuf
timestamp 1693170804
transform 1 0 23092 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 23368 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 26036 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 21528 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 20792 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 21804 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[25\].cc_clkbuf
timestamp 1693170804
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[25\].rs_mbuf
timestamp 1693170804
transform 1 0 20608 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18400 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 20240 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 18400 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 20608 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 18400 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 23092 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 21804 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[26\].cc_clkbuf
timestamp 1693170804
transform 1 0 21252 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[26\].rs_mbuf
timestamp 1693170804
transform 1 0 18400 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16192 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 18676 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 16192 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 13708 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 16192 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 17204 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 16192 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 16192 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 16928 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 16192 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 20608 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 16284 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[27\].cc_clkbuf
timestamp 1693170804
transform 1 0 15456 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[27\].rs_mbuf
timestamp 1693170804
transform 1 0 16192 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13892 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 11316 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13984 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 13708 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 14076 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 13984 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 13800 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 14076 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 13616 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[28\].cc_clkbuf
timestamp 1693170804
transform 1 0 14904 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[28\].rs_mbuf
timestamp 1693170804
transform 1 0 13524 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 12052 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 11500 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 11040 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 11316 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 9844 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[29\].cc_clkbuf
timestamp 1693170804
transform 1 0 12880 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[29\].rs_mbuf
timestamp 1693170804
transform 1 0 12328 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 9568 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 10120 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 9292 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[30\].cc_clkbuf
timestamp 1693170804
transform 1 0 10948 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[30\].rs_mbuf
timestamp 1693170804
transform 1 0 10948 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 25760 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 24380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 8648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 5520 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 8004 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 2668 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10856 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10212 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[31\].cc_clkbuf
timestamp 1693170804
transform 1 0 8464 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[31\].rs_mbuf
timestamp 1693170804
transform 1 0 8372 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[32\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16376 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[32\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 24656 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 5980 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 8924 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 5980 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[32\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 16928 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[32\].cc_clkbuf
timestamp 1693170804
transform 1 0 5888 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[32\].rs_mbuf
timestamp 1693170804
transform 1 0 8372 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 11500 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 8648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 1104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[33\].cc_clkbuf
timestamp 1693170804
transform 1 0 5796 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[33\].rs_mbuf
timestamp 1693170804
transform 1 0 3312 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 15732 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 12696 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 17480 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 6348 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 12604 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 12052 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[34\].cc_clkbuf
timestamp 1693170804
transform 1 0 2944 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[34\].rs_mbuf
timestamp 1693170804
transform 1 0 8004 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 1012 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 9108 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 1012 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 3588 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 1012 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 3588 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 2392 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 828 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[35\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 17756 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[35\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 16836 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[35\].cc_clkbuf
timestamp 1693170804
transform 1 0 3220 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[35\].rs_mbuf
timestamp 1693170804
transform 1 0 3220 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6164 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 7912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 6164 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 6440 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 5704 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8464 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[36\].cc_clkbuf
timestamp 1693170804
transform 1 0 7728 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[36\].rs_mbuf
timestamp 1693170804
transform 1 0 6716 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 14352 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 14076 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 14352 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 16560 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 17204 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11040 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 11316 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10672 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[37\].cc_clkbuf
timestamp 1693170804
transform 1 0 10948 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[37\].rs_mbuf
timestamp 1693170804
transform 1 0 13524 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 15732 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 14628 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 10948 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10028 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 10764 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 10948 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10304 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[38\].cc_clkbuf
timestamp 1693170804
transform 1 0 11684 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[38\].rs_mbuf
timestamp 1693170804
transform 1 0 12880 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 12420 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 12420 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 12236 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 12512 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 12880 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 12604 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 9752 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 9476 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[39\].cc_clkbuf
timestamp 1693170804
transform 1 0 11868 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[39\].rs_mbuf
timestamp 1693170804
transform 1 0 13524 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 9660 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 9660 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 10212 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 11500 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 9660 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 7544 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 7268 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 7728 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[40\].cc_clkbuf
timestamp 1693170804
transform 1 0 9476 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[40\].rs_mbuf
timestamp 1693170804
transform 1 0 8924 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 9016 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 6256 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6808 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6808 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 9016 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 6716 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 7728 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[41\].cc_clkbuf
timestamp 1693170804
transform 1 0 7728 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[41\].rs_mbuf
timestamp 1693170804
transform 1 0 5888 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 6072 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 1196 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 3312 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[42\].cc_clkbuf
timestamp 1693170804
transform 1 0 4600 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[42\].rs_mbuf
timestamp 1693170804
transform 1 0 3680 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 1472 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 1472 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 12144 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 19228 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 1012 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 4324 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[43\].cc_clkbuf
timestamp 1693170804
transform 1 0 5796 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[43\].rs_mbuf
timestamp 1693170804
transform 1 0 5152 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dlclkp_4  ct.ro.cc_clock_gate $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 18768 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_4  ct.ro.cc_clock_inv $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 20424 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  ct.ro.cc_ring_osc_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 21252 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  ct.ro.cc_ring_osc_1
timestamp 1693170804
transform 1 0 16376 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  ct.ro.cc_ring_osc_2
timestamp 1693170804
transform 1 0 18676 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[1\].cc_div_flop $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 18952 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[2\].cc_div_flop
timestamp 1693170804
transform 1 0 19320 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[3\].cc_div_flop
timestamp 1693170804
transform 1 0 21252 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[4\].cc_div_flop
timestamp 1693170804
transform 1 0 23460 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[5\].cc_div_flop
timestamp 1693170804
transform 1 0 22172 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[6\].cc_div_flop
timestamp 1693170804
transform 1 0 21528 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[7\].cc_div_flop
timestamp 1693170804
transform 1 0 23828 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2i_2  cw.cc_test_0
timestamp 1693170804
transform 1 0 17848 0 -1 21216
box -38 -48 1050 592
use sky130_ht_sc_tt05__mux2i_2  cw.cc_test_1
timestamp 1699069426
transform 1 0 17572 0 1 17952
box -38 -48 1050 592
use sky130_fd_sc_hd__maj3_2  cw.cc_test_2
timestamp 1693170804
transform 1 0 16100 0 -1 20128
box -38 -48 866 592
use sky130_ht_sc_tt05__maj3_2  cw.cc_test_3
timestamp 1699069426
transform 1 0 16100 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dlrtp_1  cw.cc_test_4
timestamp 1693170804
transform 1 0 10948 0 -1 20128
box -38 -48 1234 592
use sky130_ht_sc_tt05__dlrtp_1  cw.cc_test_5
timestamp 1699069426
transform 1 0 14352 0 -1 20128
box -38 -48 1418 592
use sky130_fd_sc_hd__dfrtp_1  cw.cc_test_6
timestamp 1693170804
transform 1 0 14260 0 1 20128
box -38 -48 1878 592
use sky130_ht_sc_tt05__dfrtp_1  cw.cc_test_7
timestamp 1699069426
transform 1 0 14076 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_4  fanout5
timestamp 1693170804
transform 1 0 8372 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 12236 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout7
timestamp 1693170804
transform 1 0 10672 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout8
timestamp 1693170804
transform 1 0 28980 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout9
timestamp 1693170804
transform 1 0 29164 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout10
timestamp 1693170804
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout11
timestamp 1693170804
transform 1 0 12972 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout12
timestamp 1693170804
transform 1 0 10948 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 1693170804
transform 1 0 29532 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1693170804
transform 1 0 29532 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout15
timestamp 1693170804
transform 1 0 8924 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 1693170804
transform 1 0 13156 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout17
timestamp 1693170804
transform 1 0 11224 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 1693170804
transform 1 0 30084 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 1693170804
transform 1 0 29716 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout20
timestamp 1693170804
transform 1 0 8372 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout21
timestamp 1693170804
transform 1 0 14076 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1693170804
transform 1 0 13616 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1693170804
transform 1 0 30084 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1693170804
transform 1 0 29992 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout25
timestamp 1693170804
transform 1 0 16284 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp 1693170804
transform 1 0 16100 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 1693170804
transform 1 0 13524 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1693170804
transform 1 0 28612 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout29
timestamp 1693170804
transform 1 0 28244 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout30
timestamp 1693170804
transform 1 0 30176 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 1693170804
transform 1 0 15732 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout32
timestamp 1693170804
transform 1 0 5152 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 1693170804
transform 1 0 4784 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout34
timestamp 1693170804
transform 1 0 28980 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout35
timestamp 1693170804
transform 1 0 26588 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout36
timestamp 1693170804
transform 1 0 16836 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 1693170804
transform 1 0 15364 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout38
timestamp 1693170804
transform 1 0 17664 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout39
timestamp 1693170804
transform 1 0 29532 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 1693170804
transform 1 0 25944 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 1693170804
transform 1 0 26956 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1693170804
transform 1 0 17388 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp 1693170804
transform 1 0 16468 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout44
timestamp 1693170804
transform 1 0 20424 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 1693170804
transform 1 0 25116 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout46
timestamp 1693170804
transform 1 0 26312 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 1693170804
transform 1 0 30268 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout48
timestamp 1693170804
transform 1 0 14352 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout49
timestamp 1693170804
transform 1 0 13156 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout50
timestamp 1693170804
transform 1 0 8096 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 1693170804
transform 1 0 28980 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout52
timestamp 1693170804
transform 1 0 25668 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout53
timestamp 1693170804
transform 1 0 30084 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 828 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3220 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_33
timestamp 1693170804
transform 1 0 3588 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3956 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_45
timestamp 1693170804
transform 1 0 4692 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_49
timestamp 1693170804
transform 1 0 5060 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_312 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 29256 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_324
timestamp 1693170804
transform 1 0 30360 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 1380 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_13
timestamp 1693170804
transform 1 0 1748 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_16
timestamp 1693170804
transform 1 0 2024 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_63
timestamp 1693170804
transform 1 0 6348 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_116
timestamp 1693170804
transform 1 0 11224 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_169
timestamp 1693170804
transform 1 0 16100 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1693170804
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_317
timestamp 1693170804
transform 1 0 29716 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_321 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 30084 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 1693170804
transform 1 0 828 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_56
timestamp 1693170804
transform 1 0 5704 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_91
timestamp 1693170804
transform 1 0 8924 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 1693170804
transform 1 0 13524 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1693170804
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1693170804
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_315
timestamp 1693170804
transform 1 0 29532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_3
timestamp 1693170804
transform 1 0 828 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_87
timestamp 1693170804
transform 1 0 8556 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_119
timestamp 1693170804
transform 1 0 11500 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_169
timestamp 1693170804
transform 1 0 16100 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_255
timestamp 1693170804
transform 1 0 24012 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_296
timestamp 1693170804
transform 1 0 27784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_322
timestamp 1693170804
transform 1 0 30176 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_326
timestamp 1693170804
transform 1 0 30544 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_3
timestamp 1693170804
transform 1 0 828 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_29
timestamp 1693170804
transform 1 0 3220 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1693170804
transform 1 0 8372 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1693170804
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1693170804
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1693170804
transform 1 0 28244 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1693170804
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_319
timestamp 1693170804
transform 1 0 29900 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_3
timestamp 1693170804
transform 1 0 828 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1693170804
transform 1 0 5796 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_149
timestamp 1693170804
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_169
timestamp 1693170804
transform 1 0 16100 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_234
timestamp 1693170804
transform 1 0 22080 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_277
timestamp 1693170804
transform 1 0 26036 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_281
timestamp 1693170804
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_285
timestamp 1693170804
transform 1 0 26772 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_321
timestamp 1693170804
transform 1 0 30084 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 1693170804
transform 1 0 828 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1693170804
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_94
timestamp 1693170804
transform 1 0 9200 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_141
timestamp 1693170804
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1693170804
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1693170804
transform 1 0 23644 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_265
timestamp 1693170804
transform 1 0 24932 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_269
timestamp 1693170804
transform 1 0 25300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_273
timestamp 1693170804
transform 1 0 25668 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_303
timestamp 1693170804
transform 1 0 28428 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1693170804
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_312
timestamp 1693170804
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_324
timestamp 1693170804
transform 1 0 30360 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_27
timestamp 1693170804
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 1693170804
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_83
timestamp 1693170804
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_119
timestamp 1693170804
transform 1 0 11500 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_169
timestamp 1693170804
transform 1 0 16100 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_234
timestamp 1693170804
transform 1 0 22080 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_259
timestamp 1693170804
transform 1 0 24380 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_264
timestamp 1693170804
transform 1 0 24840 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_268
timestamp 1693170804
transform 1 0 25208 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_281
timestamp 1693170804
transform 1 0 26404 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_285
timestamp 1693170804
transform 1 0 26772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_289
timestamp 1693170804
transform 1 0 27140 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_297
timestamp 1693170804
transform 1 0 27876 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_322
timestamp 1693170804
transform 1 0 30176 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_326
timestamp 1693170804
transform 1 0 30544 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1693170804
transform 1 0 828 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_35
timestamp 1693170804
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_91
timestamp 1693170804
transform 1 0 8924 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_141
timestamp 1693170804
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_194
timestamp 1693170804
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1693170804
transform 1 0 23644 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_277
timestamp 1693170804
transform 1 0 26036 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_283
timestamp 1693170804
transform 1 0 26588 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1693170804
transform 1 0 28980 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_321
timestamp 1693170804
transform 1 0 30084 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_3
timestamp 1693170804
transform 1 0 828 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_108
timestamp 1693170804
transform 1 0 10488 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 1693170804
transform 1 0 10948 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_169
timestamp 1693170804
transform 1 0 16100 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1693170804
transform 1 0 26220 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_315
timestamp 1693170804
transform 1 0 29532 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 1693170804
transform 1 0 828 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_53
timestamp 1693170804
transform 1 0 5428 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_115
timestamp 1693170804
transform 1 0 11132 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_174
timestamp 1693170804
transform 1 0 16560 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_248
timestamp 1693170804
transform 1 0 23368 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_253
timestamp 1693170804
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_279
timestamp 1693170804
transform 1 0 26220 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_312
timestamp 1693170804
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_324
timestamp 1693170804
transform 1 0 30360 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1693170804
transform 1 0 828 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_84
timestamp 1693170804
transform 1 0 8280 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_113
timestamp 1693170804
transform 1 0 10948 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1693170804
transform 1 0 21068 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_228
timestamp 1693170804
transform 1 0 21528 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_254
timestamp 1693170804
transform 1 0 23920 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1693170804
transform 1 0 26220 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_284
timestamp 1693170804
transform 1 0 26680 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_320
timestamp 1693170804
transform 1 0 29992 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_326
timestamp 1693170804
transform 1 0 30544 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 1693170804
transform 1 0 828 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1693170804
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1693170804
transform 1 0 8372 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_180
timestamp 1693170804
transform 1 0 17112 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_221
timestamp 1693170804
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_225
timestamp 1693170804
transform 1 0 21252 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_253
timestamp 1693170804
transform 1 0 23828 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_306
timestamp 1693170804
transform 1 0 28704 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_315
timestamp 1693170804
transform 1 0 29532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_3
timestamp 1693170804
transform 1 0 828 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_60
timestamp 1693170804
transform 1 0 6072 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_119
timestamp 1693170804
transform 1 0 11500 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_169
timestamp 1693170804
transform 1 0 16100 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_189
timestamp 1693170804
transform 1 0 17940 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_214
timestamp 1693170804
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_219
timestamp 1693170804
transform 1 0 20700 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_252
timestamp 1693170804
transform 1 0 23736 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_287
timestamp 1693170804
transform 1 0 26956 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_320
timestamp 1693170804
transform 1 0 29992 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 1693170804
transform 1 0 828 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_29
timestamp 1693170804
transform 1 0 3220 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_91
timestamp 1693170804
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_96
timestamp 1693170804
transform 1 0 9384 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_171
timestamp 1693170804
transform 1 0 16284 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1693170804
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_283
timestamp 1693170804
transform 1 0 26588 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 1693170804
transform 1 0 828 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_60
timestamp 1693170804
transform 1 0 6072 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_172
timestamp 1693170804
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_204
timestamp 1693170804
transform 1 0 19320 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_212
timestamp 1693170804
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_220
timestamp 1693170804
transform 1 0 20792 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_228
timestamp 1693170804
transform 1 0 21528 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_232
timestamp 1693170804
transform 1 0 21896 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_236
timestamp 1693170804
transform 1 0 22264 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1693170804
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_324
timestamp 1693170804
transform 1 0 30360 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 1693170804
transform 1 0 828 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_29
timestamp 1693170804
transform 1 0 3220 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 1693170804
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1693170804
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_165
timestamp 1693170804
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_245
timestamp 1693170804
transform 1 0 23092 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1693170804
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1693170804
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1693170804
transform 1 0 28980 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_321
timestamp 1693170804
transform 1 0 30084 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_326
timestamp 1693170804
transform 1 0 30544 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 1693170804
transform 1 0 828 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1693170804
transform 1 0 5796 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_172
timestamp 1693170804
transform 1 0 16376 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_205
timestamp 1693170804
transform 1 0 19412 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_214
timestamp 1693170804
transform 1 0 20240 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_249
timestamp 1693170804
transform 1 0 23460 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_3
timestamp 1693170804
transform 1 0 828 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_53
timestamp 1693170804
transform 1 0 5428 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_89
timestamp 1693170804
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_97
timestamp 1693170804
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_135
timestamp 1693170804
transform 1 0 12972 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_165
timestamp 1693170804
transform 1 0 15732 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_169
timestamp 1693170804
transform 1 0 16100 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_248
timestamp 1693170804
transform 1 0 23368 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_256
timestamp 1693170804
transform 1 0 24104 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_260
timestamp 1693170804
transform 1 0 24472 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_304
timestamp 1693170804
transform 1 0 28520 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_325
timestamp 1693170804
transform 1 0 30452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_3
timestamp 1693170804
transform 1 0 828 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_8
timestamp 1693170804
transform 1 0 1288 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_40
timestamp 1693170804
transform 1 0 4232 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_66
timestamp 1693170804
transform 1 0 6624 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_95
timestamp 1693170804
transform 1 0 9292 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_103
timestamp 1693170804
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1693170804
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_128
timestamp 1693170804
transform 1 0 12328 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_159
timestamp 1693170804
transform 1 0 15180 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_163
timestamp 1693170804
transform 1 0 15548 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1693170804
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_169
timestamp 1693170804
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_173
timestamp 1693170804
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_210
timestamp 1693170804
transform 1 0 19872 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_222
timestamp 1693170804
transform 1 0 20976 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_228
timestamp 1693170804
transform 1 0 21528 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_3
timestamp 1693170804
transform 1 0 828 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_29
timestamp 1693170804
transform 1 0 3220 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_91
timestamp 1693170804
transform 1 0 8924 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_165
timestamp 1693170804
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_221
timestamp 1693170804
transform 1 0 20884 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_227
timestamp 1693170804
transform 1 0 21436 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_321
timestamp 1693170804
transform 1 0 30084 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1693170804
transform 1 0 828 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_63
timestamp 1693170804
transform 1 0 6348 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_125
timestamp 1693170804
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_163
timestamp 1693170804
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_175
timestamp 1693170804
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_182
timestamp 1693170804
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_214
timestamp 1693170804
transform 1 0 20240 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1693170804
transform 1 0 21068 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1693170804
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_3
timestamp 1693170804
transform 1 0 828 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_29
timestamp 1693170804
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_91
timestamp 1693170804
transform 1 0 8924 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_98
timestamp 1693170804
transform 1 0 9568 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_129
timestamp 1693170804
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_151
timestamp 1693170804
transform 1 0 14444 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_179
timestamp 1693170804
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_183
timestamp 1693170804
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_187
timestamp 1693170804
transform 1 0 17756 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1693170804
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_203
timestamp 1693170804
transform 1 0 19228 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_239
timestamp 1693170804
transform 1 0 22540 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_245
timestamp 1693170804
transform 1 0 23092 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_283
timestamp 1693170804
transform 1 0 26588 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_321
timestamp 1693170804
transform 1 0 30084 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp 1693170804
transform 1 0 828 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1693170804
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1693170804
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_128
timestamp 1693170804
transform 1 0 12328 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_153
timestamp 1693170804
transform 1 0 14628 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_177
timestamp 1693170804
transform 1 0 16836 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_203
timestamp 1693170804
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_207
timestamp 1693170804
transform 1 0 19596 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_211
timestamp 1693170804
transform 1 0 19964 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_219
timestamp 1693170804
transform 1 0 20700 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1693170804
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_225
timestamp 1693170804
transform 1 0 21252 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_324
timestamp 1693170804
transform 1 0 30360 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_3
timestamp 1693170804
transform 1 0 828 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_29
timestamp 1693170804
transform 1 0 3220 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_85
timestamp 1693170804
transform 1 0 8372 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_95
timestamp 1693170804
transform 1 0 9292 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1693170804
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1693170804
transform 1 0 13524 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_206
timestamp 1693170804
transform 1 0 19504 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_234
timestamp 1693170804
transform 1 0 22080 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_238
timestamp 1693170804
transform 1 0 22448 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_247
timestamp 1693170804
transform 1 0 23276 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_253
timestamp 1693170804
transform 1 0 23828 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_318
timestamp 1693170804
transform 1 0 29808 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_326
timestamp 1693170804
transform 1 0 30544 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_3
timestamp 1693170804
transform 1 0 828 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_37
timestamp 1693170804
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_60
timestamp 1693170804
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_98
timestamp 1693170804
transform 1 0 9568 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_119
timestamp 1693170804
transform 1 0 11500 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_273
timestamp 1693170804
transform 1 0 25668 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_3
timestamp 1693170804
transform 1 0 828 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_35
timestamp 1693170804
transform 1 0 3772 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_112
timestamp 1693170804
transform 1 0 10856 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_151
timestamp 1693170804
transform 1 0 14444 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_176
timestamp 1693170804
transform 1 0 16744 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_203
timestamp 1693170804
transform 1 0 19228 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_231
timestamp 1693170804
transform 1 0 21804 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_321
timestamp 1693170804
transform 1 0 30084 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_325
timestamp 1693170804
transform 1 0 30452 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_3
timestamp 1693170804
transform 1 0 828 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_7
timestamp 1693170804
transform 1 0 1196 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_63
timestamp 1693170804
transform 1 0 6348 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_143
timestamp 1693170804
transform 1 0 13708 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_178
timestamp 1693170804
transform 1 0 16928 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_203
timestamp 1693170804
transform 1 0 19228 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_281
timestamp 1693170804
transform 1 0 26404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_326
timestamp 1693170804
transform 1 0 30544 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_3
timestamp 1693170804
transform 1 0 828 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_59
timestamp 1693170804
transform 1 0 5980 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_112
timestamp 1693170804
transform 1 0 10856 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_147
timestamp 1693170804
transform 1 0 14076 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_206
timestamp 1693170804
transform 1 0 19504 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1693170804
transform 1 0 23552 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1693170804
transform 1 0 28796 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_309
timestamp 1693170804
transform 1 0 28980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_3
timestamp 1693170804
transform 1 0 828 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_31
timestamp 1693170804
transform 1 0 3404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1693170804
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_119
timestamp 1693170804
transform 1 0 11500 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_255
timestamp 1693170804
transform 1 0 24012 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_3
timestamp 1693170804
transform 1 0 828 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_35
timestamp 1693170804
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_115
timestamp 1693170804
transform 1 0 11132 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_141
timestamp 1693170804
transform 1 0 13524 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_245
timestamp 1693170804
transform 1 0 23092 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_326
timestamp 1693170804
transform 1 0 30544 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_3
timestamp 1693170804
transform 1 0 828 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_31
timestamp 1693170804
transform 1 0 3404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_57
timestamp 1693170804
transform 1 0 5796 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_169
timestamp 1693170804
transform 1 0 16100 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_176
timestamp 1693170804
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_249
timestamp 1693170804
transform 1 0 23460 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_325
timestamp 1693170804
transform 1 0 30452 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_3
timestamp 1693170804
transform 1 0 828 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_35
timestamp 1693170804
transform 1 0 3772 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 1693170804
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_135
timestamp 1693170804
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_165
timestamp 1693170804
transform 1 0 15732 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_197
timestamp 1693170804
transform 1 0 18676 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_248
timestamp 1693170804
transform 1 0 23368 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_18
timestamp 1693170804
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_57
timestamp 1693170804
transform 1 0 5796 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1693170804
transform 1 0 20976 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_231
timestamp 1693170804
transform 1 0 21804 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_326
timestamp 1693170804
transform 1 0 30544 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_3
timestamp 1693170804
transform 1 0 828 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_77
timestamp 1693170804
transform 1 0 7636 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_109
timestamp 1693170804
transform 1 0 10580 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_165
timestamp 1693170804
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_226
timestamp 1693170804
transform 1 0 21344 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_322
timestamp 1693170804
transform 1 0 30176 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_51
timestamp 1693170804
transform 1 0 5244 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_57
timestamp 1693170804
transform 1 0 5796 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_110
timestamp 1693170804
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_234
timestamp 1693170804
transform 1 0 22080 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_278
timestamp 1693170804
transform 1 0 26128 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_300
timestamp 1693170804
transform 1 0 28152 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_326
timestamp 1693170804
transform 1 0 30544 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1693170804
transform 1 0 3036 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_29
timestamp 1693170804
transform 1 0 3220 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_85
timestamp 1693170804
transform 1 0 8372 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_141
timestamp 1693170804
transform 1 0 13524 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_194
timestamp 1693170804
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_202
timestamp 1693170804
transform 1 0 19136 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_283
timestamp 1693170804
transform 1 0 26588 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_326
timestamp 1693170804
transform 1 0 30544 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_3
timestamp 1693170804
transform 1 0 828 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_60
timestamp 1693170804
transform 1 0 6072 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_83
timestamp 1693170804
transform 1 0 8188 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1693170804
transform 1 0 10764 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_146
timestamp 1693170804
transform 1 0 13984 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_199
timestamp 1693170804
transform 1 0 18860 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1693170804
transform 1 0 26220 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_3
timestamp 1693170804
transform 1 0 828 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_147
timestamp 1693170804
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_325
timestamp 1693170804
transform 1 0 30452 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1693170804
transform 1 0 23460 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1693170804
transform 1 0 23092 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1693170804
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1693170804
transform 1 0 26404 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_39
timestamp 1693170804
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1693170804
transform -1 0 30912 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_40
timestamp 1693170804
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1693170804
transform -1 0 30912 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_41
timestamp 1693170804
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1693170804
transform -1 0 30912 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_42
timestamp 1693170804
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1693170804
transform -1 0 30912 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_43
timestamp 1693170804
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1693170804
transform -1 0 30912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_44
timestamp 1693170804
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1693170804
transform -1 0 30912 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_45
timestamp 1693170804
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1693170804
transform -1 0 30912 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_46
timestamp 1693170804
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1693170804
transform -1 0 30912 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_47
timestamp 1693170804
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1693170804
transform -1 0 30912 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_48
timestamp 1693170804
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1693170804
transform -1 0 30912 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_49
timestamp 1693170804
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1693170804
transform -1 0 30912 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_50
timestamp 1693170804
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1693170804
transform -1 0 30912 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_51
timestamp 1693170804
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1693170804
transform -1 0 30912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_52
timestamp 1693170804
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1693170804
transform -1 0 30912 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_53
timestamp 1693170804
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1693170804
transform -1 0 30912 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_54
timestamp 1693170804
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1693170804
transform -1 0 30912 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_55
timestamp 1693170804
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1693170804
transform -1 0 30912 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_56
timestamp 1693170804
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1693170804
transform -1 0 30912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_57
timestamp 1693170804
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1693170804
transform -1 0 30912 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_58
timestamp 1693170804
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1693170804
transform -1 0 30912 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_59
timestamp 1693170804
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1693170804
transform -1 0 30912 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_60
timestamp 1693170804
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1693170804
transform -1 0 30912 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_61
timestamp 1693170804
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1693170804
transform -1 0 30912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_62
timestamp 1693170804
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1693170804
transform -1 0 30912 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_63
timestamp 1693170804
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1693170804
transform -1 0 30912 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_64
timestamp 1693170804
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1693170804
transform -1 0 30912 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_65
timestamp 1693170804
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1693170804
transform -1 0 30912 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_66
timestamp 1693170804
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1693170804
transform -1 0 30912 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_67
timestamp 1693170804
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1693170804
transform -1 0 30912 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_68
timestamp 1693170804
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1693170804
transform -1 0 30912 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_69
timestamp 1693170804
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1693170804
transform -1 0 30912 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_70
timestamp 1693170804
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1693170804
transform -1 0 30912 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_71
timestamp 1693170804
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1693170804
transform -1 0 30912 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_72
timestamp 1693170804
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1693170804
transform -1 0 30912 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_73
timestamp 1693170804
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1693170804
transform -1 0 30912 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_74
timestamp 1693170804
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1693170804
transform -1 0 30912 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_75
timestamp 1693170804
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1693170804
transform -1 0 30912 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_76
timestamp 1693170804
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1693170804
transform -1 0 30912 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_77
timestamp 1693170804
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1693170804
transform -1 0 30912 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp 1693170804
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp 1693170804
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_81
timestamp 1693170804
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82
timestamp 1693170804
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_83
timestamp 1693170804
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 1693170804
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1693170804
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1693170804
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1693170804
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1693170804
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_89
timestamp 1693170804
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_90
timestamp 1693170804
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_91
timestamp 1693170804
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1693170804
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1693170804
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_94
timestamp 1693170804
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_95
timestamp 1693170804
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1693170804
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1693170804
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1693170804
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1693170804
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1693170804
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1693170804
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1693170804
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1693170804
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_104
timestamp 1693170804
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1693170804
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1693170804
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1693170804
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_108
timestamp 1693170804
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_109
timestamp 1693170804
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_110
timestamp 1693170804
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1693170804
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_112
timestamp 1693170804
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_113
timestamp 1693170804
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_114
timestamp 1693170804
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_115
timestamp 1693170804
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_116
timestamp 1693170804
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_117
timestamp 1693170804
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_118
timestamp 1693170804
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_119
timestamp 1693170804
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_120
timestamp 1693170804
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_121
timestamp 1693170804
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_122
timestamp 1693170804
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_123
timestamp 1693170804
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_124
timestamp 1693170804
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_125
timestamp 1693170804
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_126
timestamp 1693170804
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_127
timestamp 1693170804
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_128
timestamp 1693170804
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_129
timestamp 1693170804
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_130
timestamp 1693170804
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_131
timestamp 1693170804
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_132
timestamp 1693170804
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_133
timestamp 1693170804
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_134
timestamp 1693170804
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_135
timestamp 1693170804
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_136
timestamp 1693170804
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_137
timestamp 1693170804
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_138
timestamp 1693170804
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_139
timestamp 1693170804
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_140
timestamp 1693170804
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 1693170804
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_142
timestamp 1693170804
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 1693170804
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp 1693170804
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp 1693170804
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp 1693170804
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp 1693170804
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp 1693170804
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_149
timestamp 1693170804
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_150
timestamp 1693170804
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_151
timestamp 1693170804
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_152
timestamp 1693170804
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_153
timestamp 1693170804
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_154
timestamp 1693170804
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_155
timestamp 1693170804
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_156
timestamp 1693170804
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_157
timestamp 1693170804
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_158
timestamp 1693170804
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_159
timestamp 1693170804
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_160
timestamp 1693170804
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_161
timestamp 1693170804
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_162
timestamp 1693170804
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp 1693170804
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_164
timestamp 1693170804
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_165
timestamp 1693170804
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_166
timestamp 1693170804
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_167
timestamp 1693170804
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_168
timestamp 1693170804
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_169
timestamp 1693170804
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_170
timestamp 1693170804
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_171
timestamp 1693170804
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_172
timestamp 1693170804
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_173
timestamp 1693170804
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_174
timestamp 1693170804
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_175
timestamp 1693170804
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_176
timestamp 1693170804
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_177
timestamp 1693170804
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_178
timestamp 1693170804
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_179
timestamp 1693170804
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_180
timestamp 1693170804
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_181
timestamp 1693170804
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_182
timestamp 1693170804
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_183
timestamp 1693170804
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_184
timestamp 1693170804
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 1693170804
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_186
timestamp 1693170804
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_187
timestamp 1693170804
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_188
timestamp 1693170804
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_189
timestamp 1693170804
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_190
timestamp 1693170804
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_191
timestamp 1693170804
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_192
timestamp 1693170804
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_193
timestamp 1693170804
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_194
timestamp 1693170804
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_195
timestamp 1693170804
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_196
timestamp 1693170804
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_197
timestamp 1693170804
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_198
timestamp 1693170804
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_199
timestamp 1693170804
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_200
timestamp 1693170804
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_201
timestamp 1693170804
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_202
timestamp 1693170804
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_203
timestamp 1693170804
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_204
timestamp 1693170804
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_205
timestamp 1693170804
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_206
timestamp 1693170804
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_207
timestamp 1693170804
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_208
timestamp 1693170804
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp 1693170804
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_210
timestamp 1693170804
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_211
timestamp 1693170804
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_212
timestamp 1693170804
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_213
timestamp 1693170804
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp 1693170804
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_215
timestamp 1693170804
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_216
timestamp 1693170804
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_217
timestamp 1693170804
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_218
timestamp 1693170804
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp 1693170804
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp 1693170804
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_221
timestamp 1693170804
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_222
timestamp 1693170804
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_223
timestamp 1693170804
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp 1693170804
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp 1693170804
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_226
timestamp 1693170804
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_227
timestamp 1693170804
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_228
timestamp 1693170804
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp 1693170804
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp 1693170804
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp 1693170804
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_232
timestamp 1693170804
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_233
timestamp 1693170804
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp 1693170804
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp 1693170804
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp 1693170804
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_237
timestamp 1693170804
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_238
timestamp 1693170804
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp 1693170804
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp 1693170804
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp 1693170804
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp 1693170804
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_243
timestamp 1693170804
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp 1693170804
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp 1693170804
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp 1693170804
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp 1693170804
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_248
timestamp 1693170804
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp 1693170804
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp 1693170804
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp 1693170804
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp 1693170804
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 1693170804
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp 1693170804
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp 1693170804
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp 1693170804
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp 1693170804
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 1693170804
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp 1693170804
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp 1693170804
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp 1693170804
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp 1693170804
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 1693170804
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 1693170804
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1693170804
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp 1693170804
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp 1693170804
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 1693170804
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 1693170804
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp 1693170804
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp 1693170804
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp 1693170804
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 1693170804
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 1693170804
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1693170804
transform 1 0 28888 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp 1693170804
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp 1693170804
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 1693170804
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 1693170804
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1693170804
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp 1693170804
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp 1693170804
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 1693170804
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 1693170804
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1693170804
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 1693170804
transform 1 0 28888 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp 1693170804
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 1693170804
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 1693170804
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1693170804
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 1693170804
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp 1693170804
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 1693170804
transform 1 0 5704 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 1693170804
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1693170804
transform 1 0 10856 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 1693170804
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 1693170804
transform 1 0 16008 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_298
timestamp 1693170804
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp 1693170804
transform 1 0 21160 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_300
timestamp 1693170804
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp 1693170804
transform 1 0 26312 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_302
timestamp 1693170804
transform 1 0 28888 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 20792 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_55
timestamp 1693170804
transform 1 0 21068 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_56
timestamp 1693170804
transform 1 0 18676 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_57
timestamp 1693170804
transform 1 0 16100 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_58
timestamp 1693170804
transform 1 0 6532 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_59
timestamp 1693170804
transform 1 0 10028 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_60
timestamp 1693170804
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_61
timestamp 1693170804
transform 1 0 9292 0 1 12512
box -38 -48 314 592
<< labels >>
flabel metal4 s 7982 496 8302 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15572 496 15892 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 23162 496 23482 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 30752 496 31072 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4187 496 4507 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11777 496 12097 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19367 496 19687 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26957 496 27277 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26926 22104 26986 22304 0 FreeSans 480 90 0 0 clk
port 2 nsew signal input
flabel metal4 s 27478 22104 27538 22304 0 FreeSans 480 90 0 0 ena
port 3 nsew signal input
flabel metal4 s 26374 22104 26434 22304 0 FreeSans 480 90 0 0 rst_n
port 4 nsew signal input
flabel metal4 s 25822 22104 25882 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 5 nsew signal input
flabel metal4 s 25270 22104 25330 22304 0 FreeSans 480 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal4 s 24718 22104 24778 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal4 s 24166 22104 24226 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal4 s 23614 22104 23674 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal4 s 23062 22104 23122 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal4 s 22510 22104 22570 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal4 s 21958 22104 22018 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal4 s 21406 22104 21466 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal4 s 20854 22104 20914 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal4 s 20302 22104 20362 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal4 s 19750 22104 19810 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal4 s 19198 22104 19258 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal4 s 18646 22104 18706 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal4 s 18094 22104 18154 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal4 s 17542 22104 17602 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal4 s 8158 22104 8218 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 21 nsew signal tristate
flabel metal4 s 7606 22104 7666 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 22 nsew signal tristate
flabel metal4 s 7054 22104 7114 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 23 nsew signal tristate
flabel metal4 s 6502 22104 6562 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 24 nsew signal tristate
flabel metal4 s 5950 22104 6010 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 25 nsew signal tristate
flabel metal4 s 5398 22104 5458 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 26 nsew signal tristate
flabel metal4 s 4846 22104 4906 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 27 nsew signal tristate
flabel metal4 s 4294 22104 4354 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 28 nsew signal tristate
flabel metal4 s 12574 22104 12634 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 29 nsew signal tristate
flabel metal4 s 12022 22104 12082 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 30 nsew signal tristate
flabel metal4 s 11470 22104 11530 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 31 nsew signal tristate
flabel metal4 s 10918 22104 10978 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 32 nsew signal tristate
flabel metal4 s 10366 22104 10426 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 33 nsew signal tristate
flabel metal4 s 9814 22104 9874 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 34 nsew signal tristate
flabel metal4 s 9262 22104 9322 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 35 nsew signal tristate
flabel metal4 s 8710 22104 8770 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 36 nsew signal tristate
flabel metal4 s 16990 22104 17050 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 37 nsew signal tristate
flabel metal4 s 16438 22104 16498 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 38 nsew signal tristate
flabel metal4 s 15886 22104 15946 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 39 nsew signal tristate
flabel metal4 s 15334 22104 15394 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 40 nsew signal tristate
flabel metal4 s 14782 22104 14842 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 41 nsew signal tristate
flabel metal4 s 14230 22104 14290 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 42 nsew signal tristate
flabel metal4 s 13678 22104 13738 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 43 nsew signal tristate
flabel metal4 s 13126 22104 13186 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 44 nsew signal tristate
rlabel via1 15812 21216 15812 21216 0 VGND
rlabel metal1 15732 21760 15732 21760 0 VPWR
rlabel metal2 28750 20740 28750 20740 0 _00_
rlabel metal1 24104 19278 24104 19278 0 _01_
rlabel metal2 24334 20026 24334 20026 0 _02_
rlabel metal1 23874 19210 23874 19210 0 _03_
rlabel metal1 19182 20570 19182 20570 0 _04_
rlabel metal1 29854 16660 29854 16660 0 ct.cw.source\[0\]
rlabel metal1 19274 14994 19274 14994 0 ct.cw.source\[1\]
rlabel metal1 21298 14586 21298 14586 0 ct.cw.source\[2\]
rlabel metal2 2070 15249 2070 15249 0 ct.cw.target\[0\]
rlabel via2 15502 11203 15502 11203 0 ct.cw.target\[1\]
rlabel metal2 17020 13260 17020 13260 0 ct.cw.target\[2\]
rlabel metal1 2116 12818 2116 12818 0 ct.cw.target\[3\]
rlabel metal2 1886 11594 1886 11594 0 ct.cw.target\[4\]
rlabel metal1 14536 17714 14536 17714 0 ct.cw.target\[5\]
rlabel via2 2162 10659 2162 10659 0 ct.cw.target\[6\]
rlabel metal1 13386 18224 13386 18224 0 ct.cw.target\[7\]
rlabel metal1 29440 13158 29440 13158 0 ct.ic.data_chain\[10\]
rlabel metal1 27692 10642 27692 10642 0 ct.ic.data_chain\[11\]
rlabel metal2 18630 21794 18630 21794 0 ct.ic.data_chain\[12\]
rlabel metal1 28382 13362 28382 13362 0 ct.ic.data_chain\[13\]
rlabel metal2 28658 13838 28658 13838 0 ct.ic.data_chain\[14\]
rlabel metal1 27508 20910 27508 20910 0 ct.ic.data_chain\[15\]
rlabel metal1 22632 14994 22632 14994 0 ct.ic.data_chain\[16\]
rlabel metal1 28474 14450 28474 14450 0 ct.ic.data_chain\[17\]
rlabel metal1 25024 16218 25024 16218 0 ct.ic.data_chain\[18\]
rlabel metal1 25714 17170 25714 17170 0 ct.ic.data_chain\[19\]
rlabel metal1 26404 19890 26404 19890 0 ct.ic.data_chain\[20\]
rlabel metal2 21022 16252 21022 16252 0 ct.ic.data_chain\[21\]
rlabel metal2 22034 17935 22034 17935 0 ct.ic.data_chain\[22\]
rlabel metal1 21298 15538 21298 15538 0 ct.ic.data_chain\[23\]
rlabel metal1 19780 16626 19780 16626 0 ct.ic.data_chain\[24\]
rlabel metal1 19780 21454 19780 21454 0 ct.ic.data_chain\[25\]
rlabel metal1 20240 15470 20240 15470 0 ct.ic.data_chain\[26\]
rlabel metal1 18814 18802 18814 18802 0 ct.ic.data_chain\[27\]
rlabel metal1 18814 19890 18814 19890 0 ct.ic.data_chain\[28\]
rlabel metal1 19688 17714 19688 17714 0 ct.ic.data_chain\[29\]
rlabel metal1 17388 18802 17388 18802 0 ct.ic.data_chain\[30\]
rlabel metal2 17250 19108 17250 19108 0 ct.ic.data_chain\[31\]
rlabel metal1 18906 19278 18906 19278 0 ct.ic.data_chain\[32\]
rlabel metal1 16192 20434 16192 20434 0 ct.ic.data_chain\[33\]
rlabel metal1 16330 18258 16330 18258 0 ct.ic.data_chain\[34\]
rlabel metal1 16054 18938 16054 18938 0 ct.ic.data_chain\[35\]
rlabel metal1 29486 9010 29486 9010 0 ct.ic.data_chain\[3\]
rlabel metal2 16238 15555 16238 15555 0 ct.ic.data_chain\[4\]
rlabel metal1 19642 14450 19642 14450 0 ct.ic.data_chain\[5\]
rlabel metal1 28888 10030 28888 10030 0 ct.ic.data_chain\[6\]
rlabel metal1 19320 13362 19320 13362 0 ct.ic.data_chain\[7\]
rlabel metal3 15065 16660 15065 16660 0 ct.ic.data_chain\[8\]
rlabel metal1 18492 21658 18492 21658 0 ct.ic.data_chain\[9\]
rlabel metal1 28612 21454 28612 21454 0 ct.ic.trig_chain\[0\]
rlabel metal1 16928 18734 16928 18734 0 ct.ic.trig_chain\[10\]
rlabel metal1 16146 20298 16146 20298 0 ct.ic.trig_chain\[11\]
rlabel metal1 14490 21522 14490 21522 0 ct.ic.trig_chain\[12\]
rlabel metal2 19458 14399 19458 14399 0 ct.ic.trig_chain\[1\]
rlabel metal1 14214 17646 14214 17646 0 ct.ic.trig_chain\[2\]
rlabel metal1 30084 20434 30084 20434 0 ct.ic.trig_chain\[3\]
rlabel metal2 21666 21913 21666 21913 0 ct.ic.trig_chain\[4\]
rlabel metal2 23598 14841 23598 14841 0 ct.ic.trig_chain\[5\]
rlabel metal1 26680 19822 26680 19822 0 ct.ic.trig_chain\[6\]
rlabel metal1 23230 18394 23230 18394 0 ct.ic.trig_chain\[7\]
rlabel metal1 20286 18870 20286 18870 0 ct.ic.trig_chain\[8\]
rlabel metal1 18354 19822 18354 19822 0 ct.ic.trig_chain\[9\]
rlabel metal3 13340 18156 13340 18156 0 ct.oc.capture_buffer\[0\]
rlabel metal1 26358 18802 26358 18802 0 ct.oc.capture_buffer\[100\]
rlabel metal1 29670 18394 29670 18394 0 ct.oc.capture_buffer\[101\]
rlabel metal1 28244 18326 28244 18326 0 ct.oc.capture_buffer\[102\]
rlabel metal1 29854 15130 29854 15130 0 ct.oc.capture_buffer\[103\]
rlabel metal1 24932 13838 24932 13838 0 ct.oc.capture_buffer\[104\]
rlabel metal1 26864 13362 26864 13362 0 ct.oc.capture_buffer\[105\]
rlabel metal1 27140 13838 27140 13838 0 ct.oc.capture_buffer\[106\]
rlabel metal1 23506 12886 23506 12886 0 ct.oc.capture_buffer\[107\]
rlabel metal1 28566 14042 28566 14042 0 ct.oc.capture_buffer\[108\]
rlabel metal1 29210 14042 29210 14042 0 ct.oc.capture_buffer\[109\]
rlabel metal1 12466 20536 12466 20536 0 ct.oc.capture_buffer\[10\]
rlabel metal1 29670 14042 29670 14042 0 ct.oc.capture_buffer\[110\]
rlabel metal1 29854 14586 29854 14586 0 ct.oc.capture_buffer\[111\]
rlabel metal1 24564 12818 24564 12818 0 ct.oc.capture_buffer\[112\]
rlabel metal1 24242 13362 24242 13362 0 ct.oc.capture_buffer\[113\]
rlabel metal1 21942 13396 21942 13396 0 ct.oc.capture_buffer\[114\]
rlabel metal1 23828 12614 23828 12614 0 ct.oc.capture_buffer\[115\]
rlabel metal2 28658 12240 28658 12240 0 ct.oc.capture_buffer\[116\]
rlabel metal1 28520 12750 28520 12750 0 ct.oc.capture_buffer\[117\]
rlabel metal1 28244 14926 28244 14926 0 ct.oc.capture_buffer\[118\]
rlabel metal2 29854 14212 29854 14212 0 ct.oc.capture_buffer\[119\]
rlabel metal1 11224 20366 11224 20366 0 ct.oc.capture_buffer\[11\]
rlabel metal1 20976 12410 20976 12410 0 ct.oc.capture_buffer\[120\]
rlabel metal1 20516 12614 20516 12614 0 ct.oc.capture_buffer\[121\]
rlabel metal1 20378 12954 20378 12954 0 ct.oc.capture_buffer\[122\]
rlabel metal2 22310 11492 22310 11492 0 ct.oc.capture_buffer\[123\]
rlabel metal1 25116 11662 25116 11662 0 ct.oc.capture_buffer\[124\]
rlabel metal1 28934 11322 28934 11322 0 ct.oc.capture_buffer\[125\]
rlabel metal1 29440 6834 29440 6834 0 ct.oc.capture_buffer\[126\]
rlabel metal1 29348 7922 29348 7922 0 ct.oc.capture_buffer\[127\]
rlabel metal1 19596 10574 19596 10574 0 ct.oc.capture_buffer\[128\]
rlabel metal1 19366 12614 19366 12614 0 ct.oc.capture_buffer\[129\]
rlabel metal2 13938 15793 13938 15793 0 ct.oc.capture_buffer\[12\]
rlabel metal1 18768 12274 18768 12274 0 ct.oc.capture_buffer\[130\]
rlabel metal1 21620 10574 21620 10574 0 ct.oc.capture_buffer\[131\]
rlabel metal1 24380 10778 24380 10778 0 ct.oc.capture_buffer\[132\]
rlabel metal2 26358 9894 26358 9894 0 ct.oc.capture_buffer\[133\]
rlabel metal1 27876 8942 27876 8942 0 ct.oc.capture_buffer\[134\]
rlabel metal2 28290 9860 28290 9860 0 ct.oc.capture_buffer\[135\]
rlabel metal2 17986 9962 17986 9962 0 ct.oc.capture_buffer\[136\]
rlabel metal1 16882 11186 16882 11186 0 ct.oc.capture_buffer\[137\]
rlabel metal1 17112 11730 17112 11730 0 ct.oc.capture_buffer\[138\]
rlabel metal1 21620 10098 21620 10098 0 ct.oc.capture_buffer\[139\]
rlabel metal1 11868 13226 11868 13226 0 ct.oc.capture_buffer\[13\]
rlabel metal1 22908 10778 22908 10778 0 ct.oc.capture_buffer\[140\]
rlabel metal1 25714 8602 25714 8602 0 ct.oc.capture_buffer\[141\]
rlabel metal1 26404 9146 26404 9146 0 ct.oc.capture_buffer\[142\]
rlabel metal1 24794 10030 24794 10030 0 ct.oc.capture_buffer\[143\]
rlabel metal2 17158 9724 17158 9724 0 ct.oc.capture_buffer\[144\]
rlabel metal2 19458 9350 19458 9350 0 ct.oc.capture_buffer\[145\]
rlabel metal1 17710 8942 17710 8942 0 ct.oc.capture_buffer\[146\]
rlabel metal1 19136 8398 19136 8398 0 ct.oc.capture_buffer\[147\]
rlabel metal1 21482 9146 21482 9146 0 ct.oc.capture_buffer\[148\]
rlabel metal2 25714 9316 25714 9316 0 ct.oc.capture_buffer\[149\]
rlabel metal1 14168 15062 14168 15062 0 ct.oc.capture_buffer\[14\]
rlabel metal1 24564 8466 24564 8466 0 ct.oc.capture_buffer\[150\]
rlabel metal2 23690 9180 23690 9180 0 ct.oc.capture_buffer\[151\]
rlabel metal2 17250 7514 17250 7514 0 ct.oc.capture_buffer\[152\]
rlabel metal1 17802 6324 17802 6324 0 ct.oc.capture_buffer\[153\]
rlabel metal2 17526 7174 17526 7174 0 ct.oc.capture_buffer\[154\]
rlabel metal1 18400 6426 18400 6426 0 ct.oc.capture_buffer\[155\]
rlabel metal2 20470 8194 20470 8194 0 ct.oc.capture_buffer\[156\]
rlabel metal2 21574 7276 21574 7276 0 ct.oc.capture_buffer\[157\]
rlabel metal1 22264 7378 22264 7378 0 ct.oc.capture_buffer\[158\]
rlabel metal1 21988 7922 21988 7922 0 ct.oc.capture_buffer\[159\]
rlabel metal1 11868 13158 11868 13158 0 ct.oc.capture_buffer\[15\]
rlabel metal1 24150 6426 24150 6426 0 ct.oc.capture_buffer\[160\]
rlabel metal2 28474 7616 28474 7616 0 ct.oc.capture_buffer\[161\]
rlabel metal1 27508 6290 27508 6290 0 ct.oc.capture_buffer\[162\]
rlabel metal1 26726 6970 26726 6970 0 ct.oc.capture_buffer\[163\]
rlabel metal1 29440 4658 29440 4658 0 ct.oc.capture_buffer\[164\]
rlabel metal1 29026 7446 29026 7446 0 ct.oc.capture_buffer\[165\]
rlabel metal1 28244 5202 28244 5202 0 ct.oc.capture_buffer\[166\]
rlabel metal2 28658 5644 28658 5644 0 ct.oc.capture_buffer\[167\]
rlabel via2 4554 4131 4554 4131 0 ct.oc.capture_buffer\[168\]
rlabel metal1 2277 2414 2277 2414 0 ct.oc.capture_buffer\[169\]
rlabel metal1 7958 21318 7958 21318 0 ct.oc.capture_buffer\[16\]
rlabel metal2 12374 1496 12374 1496 0 ct.oc.capture_buffer\[170\]
rlabel metal2 20654 4420 20654 4420 0 ct.oc.capture_buffer\[171\]
rlabel metal1 27416 850 27416 850 0 ct.oc.capture_buffer\[172\]
rlabel metal2 20194 4692 20194 4692 0 ct.oc.capture_buffer\[173\]
rlabel metal2 18630 10132 18630 10132 0 ct.oc.capture_buffer\[174\]
rlabel metal2 15042 1377 15042 1377 0 ct.oc.capture_buffer\[175\]
rlabel via2 4002 2397 4002 2397 0 ct.oc.capture_buffer\[176\]
rlabel metal1 4876 1938 4876 1938 0 ct.oc.capture_buffer\[177\]
rlabel metal1 24472 374 24472 374 0 ct.oc.capture_buffer\[178\]
rlabel metal1 27048 1870 27048 1870 0 ct.oc.capture_buffer\[179\]
rlabel metal1 7314 17850 7314 17850 0 ct.oc.capture_buffer\[17\]
rlabel metal1 26680 4114 26680 4114 0 ct.oc.capture_buffer\[180\]
rlabel metal1 26772 3026 26772 3026 0 ct.oc.capture_buffer\[181\]
rlabel via2 4278 1309 4278 1309 0 ct.oc.capture_buffer\[182\]
rlabel metal1 19090 3638 19090 3638 0 ct.oc.capture_buffer\[183\]
rlabel metal2 28382 850 28382 850 0 ct.oc.capture_buffer\[184\]
rlabel metal2 20746 391 20746 391 0 ct.oc.capture_buffer\[185\]
rlabel metal1 25070 2482 25070 2482 0 ct.oc.capture_buffer\[186\]
rlabel metal1 25438 4794 25438 4794 0 ct.oc.capture_buffer\[187\]
rlabel metal1 25714 5644 25714 5644 0 ct.oc.capture_buffer\[188\]
rlabel metal2 25990 6324 25990 6324 0 ct.oc.capture_buffer\[189\]
rlabel via1 12466 22083 12466 22083 0 ct.oc.capture_buffer\[18\]
rlabel metal1 20516 782 20516 782 0 ct.oc.capture_buffer\[190\]
rlabel metal1 27094 1326 27094 1326 0 ct.oc.capture_buffer\[191\]
rlabel metal1 24564 1938 24564 1938 0 ct.oc.capture_buffer\[192\]
rlabel metal2 24610 1564 24610 1564 0 ct.oc.capture_buffer\[193\]
rlabel metal2 22954 3740 22954 3740 0 ct.oc.capture_buffer\[194\]
rlabel metal1 24334 5134 24334 5134 0 ct.oc.capture_buffer\[195\]
rlabel metal1 23276 4998 23276 4998 0 ct.oc.capture_buffer\[196\]
rlabel metal2 22954 5372 22954 5372 0 ct.oc.capture_buffer\[197\]
rlabel metal1 25944 986 25944 986 0 ct.oc.capture_buffer\[198\]
rlabel metal1 24564 3026 24564 3026 0 ct.oc.capture_buffer\[199\]
rlabel metal1 9338 17646 9338 17646 0 ct.oc.capture_buffer\[19\]
rlabel metal1 10902 18598 10902 18598 0 ct.oc.capture_buffer\[1\]
rlabel metal2 23138 1836 23138 1836 0 ct.oc.capture_buffer\[200\]
rlabel metal1 23414 1258 23414 1258 0 ct.oc.capture_buffer\[201\]
rlabel metal1 21620 4114 21620 4114 0 ct.oc.capture_buffer\[202\]
rlabel metal1 21620 6290 21620 6290 0 ct.oc.capture_buffer\[203\]
rlabel metal1 21620 5746 21620 5746 0 ct.oc.capture_buffer\[204\]
rlabel metal1 21436 5134 21436 5134 0 ct.oc.capture_buffer\[205\]
rlabel metal2 26082 476 26082 476 0 ct.oc.capture_buffer\[206\]
rlabel metal1 21758 3026 21758 3026 0 ct.oc.capture_buffer\[207\]
rlabel metal1 20194 1530 20194 1530 0 ct.oc.capture_buffer\[208\]
rlabel metal1 21114 918 21114 918 0 ct.oc.capture_buffer\[209\]
rlabel metal1 6026 13260 6026 13260 0 ct.oc.capture_buffer\[20\]
rlabel metal1 20081 4114 20081 4114 0 ct.oc.capture_buffer\[210\]
rlabel metal1 19872 6290 19872 6290 0 ct.oc.capture_buffer\[211\]
rlabel metal1 19918 5678 19918 5678 0 ct.oc.capture_buffer\[212\]
rlabel metal1 20010 5202 20010 5202 0 ct.oc.capture_buffer\[213\]
rlabel metal2 19182 2244 19182 2244 0 ct.oc.capture_buffer\[214\]
rlabel metal1 20056 3026 20056 3026 0 ct.oc.capture_buffer\[215\]
rlabel metal1 16514 986 16514 986 0 ct.oc.capture_buffer\[216\]
rlabel metal1 17848 986 17848 986 0 ct.oc.capture_buffer\[217\]
rlabel metal1 16652 4046 16652 4046 0 ct.oc.capture_buffer\[218\]
rlabel metal1 17112 4658 17112 4658 0 ct.oc.capture_buffer\[219\]
rlabel metal2 5382 17816 5382 17816 0 ct.oc.capture_buffer\[21\]
rlabel metal1 16928 5746 16928 5746 0 ct.oc.capture_buffer\[220\]
rlabel metal2 16974 5644 16974 5644 0 ct.oc.capture_buffer\[221\]
rlabel metal2 20654 1734 20654 1734 0 ct.oc.capture_buffer\[222\]
rlabel metal1 17710 2074 17710 2074 0 ct.oc.capture_buffer\[223\]
rlabel metal2 13570 1394 13570 1394 0 ct.oc.capture_buffer\[224\]
rlabel metal1 14490 1326 14490 1326 0 ct.oc.capture_buffer\[225\]
rlabel metal2 14766 3604 14766 3604 0 ct.oc.capture_buffer\[226\]
rlabel metal1 14168 4658 14168 4658 0 ct.oc.capture_buffer\[227\]
rlabel metal1 14536 5746 14536 5746 0 ct.oc.capture_buffer\[228\]
rlabel metal1 14674 5202 14674 5202 0 ct.oc.capture_buffer\[229\]
rlabel metal2 1702 21505 1702 21505 0 ct.oc.capture_buffer\[22\]
rlabel metal2 14582 1802 14582 1802 0 ct.oc.capture_buffer\[230\]
rlabel metal1 14260 2074 14260 2074 0 ct.oc.capture_buffer\[231\]
rlabel metal2 10626 1275 10626 1275 0 ct.oc.capture_buffer\[232\]
rlabel metal2 5474 476 5474 476 0 ct.oc.capture_buffer\[233\]
rlabel metal1 12190 3638 12190 3638 0 ct.oc.capture_buffer\[234\]
rlabel metal1 12052 5746 12052 5746 0 ct.oc.capture_buffer\[235\]
rlabel metal1 11822 5134 11822 5134 0 ct.oc.capture_buffer\[236\]
rlabel metal2 13570 5372 13570 5372 0 ct.oc.capture_buffer\[237\]
rlabel metal1 12282 2414 12282 2414 0 ct.oc.capture_buffer\[238\]
rlabel metal1 11684 2958 11684 2958 0 ct.oc.capture_buffer\[239\]
rlabel metal1 9798 13158 9798 13158 0 ct.oc.capture_buffer\[23\]
rlabel metal1 9752 1938 9752 1938 0 ct.oc.capture_buffer\[240\]
rlabel metal1 10212 1326 10212 1326 0 ct.oc.capture_buffer\[241\]
rlabel metal2 9430 3740 9430 3740 0 ct.oc.capture_buffer\[242\]
rlabel metal1 10350 4590 10350 4590 0 ct.oc.capture_buffer\[243\]
rlabel metal1 10856 4114 10856 4114 0 ct.oc.capture_buffer\[244\]
rlabel metal1 10396 4794 10396 4794 0 ct.oc.capture_buffer\[245\]
rlabel metal1 8648 9690 8648 9690 0 ct.oc.capture_buffer\[246\]
rlabel metal1 9798 2992 9798 2992 0 ct.oc.capture_buffer\[247\]
rlabel metal1 20746 5066 20746 5066 0 ct.oc.capture_buffer\[248\]
rlabel metal1 13202 952 13202 952 0 ct.oc.capture_buffer\[249\]
rlabel metal1 16100 15334 16100 15334 0 ct.oc.capture_buffer\[24\]
rlabel metal1 7406 3570 7406 3570 0 ct.oc.capture_buffer\[250\]
rlabel metal1 6532 5134 6532 5134 0 ct.oc.capture_buffer\[251\]
rlabel metal2 2714 1530 2714 1530 0 ct.oc.capture_buffer\[252\]
rlabel metal1 8464 4522 8464 4522 0 ct.oc.capture_buffer\[253\]
rlabel metal1 7912 1326 7912 1326 0 ct.oc.capture_buffer\[254\]
rlabel metal1 7498 3026 7498 3026 0 ct.oc.capture_buffer\[255\]
rlabel metal2 16606 6681 16606 6681 0 ct.oc.capture_buffer\[256\]
rlabel metal1 2162 1870 2162 1870 0 ct.oc.capture_buffer\[257\]
rlabel via2 6578 2397 6578 2397 0 ct.oc.capture_buffer\[258\]
rlabel metal1 6256 5746 6256 5746 0 ct.oc.capture_buffer\[259\]
rlabel metal2 16698 15776 16698 15776 0 ct.oc.capture_buffer\[25\]
rlabel metal1 8648 4250 8648 4250 0 ct.oc.capture_buffer\[260\]
rlabel metal2 6762 3876 6762 3876 0 ct.oc.capture_buffer\[261\]
rlabel metal2 20194 6987 20194 6987 0 ct.oc.capture_buffer\[262\]
rlabel metal1 4968 3026 4968 3026 0 ct.oc.capture_buffer\[263\]
rlabel metal1 12466 10642 12466 10642 0 ct.oc.capture_buffer\[264\]
rlabel metal2 1702 17085 1702 17085 0 ct.oc.capture_buffer\[265\]
rlabel metal1 4830 3502 4830 3502 0 ct.oc.capture_buffer\[266\]
rlabel metal1 1058 1258 1058 1258 0 ct.oc.capture_buffer\[267\]
rlabel metal1 4646 4658 4646 4658 0 ct.oc.capture_buffer\[268\]
rlabel metal1 4830 5746 4830 5746 0 ct.oc.capture_buffer\[269\]
rlabel metal1 7222 18802 7222 18802 0 ct.oc.capture_buffer\[26\]
rlabel metal1 4416 7922 4416 7922 0 ct.oc.capture_buffer\[270\]
rlabel metal2 2070 3553 2070 3553 0 ct.oc.capture_buffer\[271\]
rlabel metal1 14490 18190 14490 18190 0 ct.oc.capture_buffer\[272\]
rlabel metal2 1702 13396 1702 13396 0 ct.oc.capture_buffer\[273\]
rlabel metal2 1702 3009 1702 3009 0 ct.oc.capture_buffer\[274\]
rlabel metal1 3956 6222 3956 6222 0 ct.oc.capture_buffer\[275\]
rlabel metal2 2070 5729 2070 5729 0 ct.oc.capture_buffer\[276\]
rlabel metal2 1978 6273 1978 6273 0 ct.oc.capture_buffer\[277\]
rlabel via2 12098 11339 12098 11339 0 ct.oc.capture_buffer\[278\]
rlabel metal2 5474 10659 5474 10659 0 ct.oc.capture_buffer\[279\]
rlabel metal2 14858 13804 14858 13804 0 ct.oc.capture_buffer\[27\]
rlabel metal2 1794 8381 1794 8381 0 ct.oc.capture_buffer\[280\]
rlabel metal1 2346 8398 2346 8398 0 ct.oc.capture_buffer\[281\]
rlabel metal1 2208 7854 2208 7854 0 ct.oc.capture_buffer\[282\]
rlabel metal1 3588 2074 3588 2074 0 ct.oc.capture_buffer\[283\]
rlabel metal1 2162 6630 2162 6630 0 ct.oc.capture_buffer\[284\]
rlabel metal1 2346 1190 2346 1190 0 ct.oc.capture_buffer\[285\]
rlabel metal2 9476 4658 9476 4658 0 ct.oc.capture_buffer\[286\]
rlabel metal2 1702 6749 1702 6749 0 ct.oc.capture_buffer\[287\]
rlabel metal1 7452 7514 7452 7514 0 ct.oc.capture_buffer\[288\]
rlabel metal2 3266 4352 3266 4352 0 ct.oc.capture_buffer\[289\]
rlabel metal1 6256 14246 6256 14246 0 ct.oc.capture_buffer\[28\]
rlabel metal1 6256 6290 6256 6290 0 ct.oc.capture_buffer\[290\]
rlabel metal1 4600 7378 4600 7378 0 ct.oc.capture_buffer\[291\]
rlabel metal1 1909 5542 1909 5542 0 ct.oc.capture_buffer\[292\]
rlabel metal1 8648 6630 8648 6630 0 ct.oc.capture_buffer\[293\]
rlabel metal2 9154 7514 9154 7514 0 ct.oc.capture_buffer\[294\]
rlabel metal1 8878 5338 8878 5338 0 ct.oc.capture_buffer\[295\]
rlabel metal2 16146 7378 16146 7378 0 ct.oc.capture_buffer\[296\]
rlabel metal1 14904 7310 14904 7310 0 ct.oc.capture_buffer\[297\]
rlabel metal2 14582 7990 14582 7990 0 ct.oc.capture_buffer\[298\]
rlabel metal1 15732 6290 15732 6290 0 ct.oc.capture_buffer\[299\]
rlabel via2 1610 20349 1610 20349 0 ct.oc.capture_buffer\[29\]
rlabel metal1 11776 20978 11776 20978 0 ct.oc.capture_buffer\[2\]
rlabel metal1 15870 6766 15870 6766 0 ct.oc.capture_buffer\[300\]
rlabel metal1 11776 7310 11776 7310 0 ct.oc.capture_buffer\[301\]
rlabel metal1 11730 6222 11730 6222 0 ct.oc.capture_buffer\[302\]
rlabel metal2 12098 6868 12098 6868 0 ct.oc.capture_buffer\[303\]
rlabel metal1 14904 8466 14904 8466 0 ct.oc.capture_buffer\[304\]
rlabel metal1 14628 9010 14628 9010 0 ct.oc.capture_buffer\[305\]
rlabel metal1 15042 10030 15042 10030 0 ct.oc.capture_buffer\[306\]
rlabel metal1 14076 9486 14076 9486 0 ct.oc.capture_buffer\[307\]
rlabel metal1 14490 10642 14490 10642 0 ct.oc.capture_buffer\[308\]
rlabel metal1 10488 8806 10488 8806 0 ct.oc.capture_buffer\[309\]
rlabel metal1 10948 13158 10948 13158 0 ct.oc.capture_buffer\[30\]
rlabel metal1 11086 9146 11086 9146 0 ct.oc.capture_buffer\[310\]
rlabel metal1 11684 9010 11684 9010 0 ct.oc.capture_buffer\[311\]
rlabel metal1 13984 11186 13984 11186 0 ct.oc.capture_buffer\[312\]
rlabel metal1 12558 12410 12558 12410 0 ct.oc.capture_buffer\[313\]
rlabel metal1 13248 12274 13248 12274 0 ct.oc.capture_buffer\[314\]
rlabel metal1 13662 12886 13662 12886 0 ct.oc.capture_buffer\[315\]
rlabel metal1 12190 11730 12190 11730 0 ct.oc.capture_buffer\[316\]
rlabel metal1 9798 9112 9798 9112 0 ct.oc.capture_buffer\[317\]
rlabel metal1 9982 10098 9982 10098 0 ct.oc.capture_buffer\[318\]
rlabel metal1 10488 8466 10488 8466 0 ct.oc.capture_buffer\[319\]
rlabel metal1 11546 13498 11546 13498 0 ct.oc.capture_buffer\[31\]
rlabel metal1 10994 12172 10994 12172 0 ct.oc.capture_buffer\[320\]
rlabel metal1 9890 12206 9890 12206 0 ct.oc.capture_buffer\[321\]
rlabel metal2 10258 13260 10258 13260 0 ct.oc.capture_buffer\[322\]
rlabel metal1 10212 11730 10212 11730 0 ct.oc.capture_buffer\[323\]
rlabel metal1 10672 10642 10672 10642 0 ct.oc.capture_buffer\[324\]
rlabel metal1 7958 9010 7958 9010 0 ct.oc.capture_buffer\[325\]
rlabel metal1 7682 8602 7682 8602 0 ct.oc.capture_buffer\[326\]
rlabel viali 6854 9484 6854 9484 0 ct.oc.capture_buffer\[327\]
rlabel metal1 7866 12818 7866 12818 0 ct.oc.capture_buffer\[328\]
rlabel metal2 6210 12852 6210 12852 0 ct.oc.capture_buffer\[329\]
rlabel metal1 5060 17102 5060 17102 0 ct.oc.capture_buffer\[32\]
rlabel metal1 7820 11866 7820 11866 0 ct.oc.capture_buffer\[330\]
rlabel metal1 8326 13294 8326 13294 0 ct.oc.capture_buffer\[331\]
rlabel metal1 7636 11186 7636 11186 0 ct.oc.capture_buffer\[332\]
rlabel metal1 5796 8058 5796 8058 0 ct.oc.capture_buffer\[333\]
rlabel metal2 5474 8194 5474 8194 0 ct.oc.capture_buffer\[334\]
rlabel metal2 3266 7072 3266 7072 0 ct.oc.capture_buffer\[335\]
rlabel metal1 4830 11730 4830 11730 0 ct.oc.capture_buffer\[336\]
rlabel metal1 5244 13906 5244 13906 0 ct.oc.capture_buffer\[337\]
rlabel metal1 4692 13294 4692 13294 0 ct.oc.capture_buffer\[338\]
rlabel metal2 4646 13634 4646 13634 0 ct.oc.capture_buffer\[339\]
rlabel metal1 5198 14246 5198 14246 0 ct.oc.capture_buffer\[33\]
rlabel metal1 1518 14280 1518 14280 0 ct.oc.capture_buffer\[340\]
rlabel metal1 3496 13974 3496 13974 0 ct.oc.capture_buffer\[341\]
rlabel metal1 4094 10030 4094 10030 0 ct.oc.capture_buffer\[342\]
rlabel metal1 4922 8942 4922 8942 0 ct.oc.capture_buffer\[343\]
rlabel metal2 2254 13481 2254 13481 0 ct.oc.capture_buffer\[344\]
rlabel metal1 2208 11186 2208 11186 0 ct.oc.capture_buffer\[345\]
rlabel metal1 11132 12954 11132 12954 0 ct.oc.capture_buffer\[346\]
rlabel metal2 2162 13209 2162 13209 0 ct.oc.capture_buffer\[347\]
rlabel metal1 2024 12206 2024 12206 0 ct.oc.capture_buffer\[348\]
rlabel metal1 1012 1530 1012 1530 0 ct.oc.capture_buffer\[349\]
rlabel metal3 13156 18428 13156 18428 0 ct.oc.capture_buffer\[34\]
rlabel metal1 2231 10574 2231 10574 0 ct.oc.capture_buffer\[350\]
rlabel metal1 1656 9486 1656 9486 0 ct.oc.capture_buffer\[351\]
rlabel via2 11546 13243 11546 13243 0 ct.oc.capture_buffer\[35\]
rlabel metal2 2438 17340 2438 17340 0 ct.oc.capture_buffer\[36\]
rlabel metal1 8142 13974 8142 13974 0 ct.oc.capture_buffer\[37\]
rlabel metal3 1863 19380 1863 19380 0 ct.oc.capture_buffer\[38\]
rlabel metal2 1978 17153 1978 17153 0 ct.oc.capture_buffer\[39\]
rlabel metal2 13110 19482 13110 19482 0 ct.oc.capture_buffer\[3\]
rlabel metal2 4278 15878 4278 15878 0 ct.oc.capture_buffer\[40\]
rlabel metal2 4094 14756 4094 14756 0 ct.oc.capture_buffer\[41\]
rlabel metal1 3956 16626 3956 16626 0 ct.oc.capture_buffer\[42\]
rlabel metal1 4462 14586 4462 14586 0 ct.oc.capture_buffer\[43\]
rlabel metal1 2254 15470 2254 15470 0 ct.oc.capture_buffer\[44\]
rlabel metal1 2208 14926 2208 14926 0 ct.oc.capture_buffer\[45\]
rlabel metal2 2162 16269 2162 16269 0 ct.oc.capture_buffer\[46\]
rlabel metal2 2530 18938 2530 18938 0 ct.oc.capture_buffer\[47\]
rlabel metal1 6532 13838 6532 13838 0 ct.oc.capture_buffer\[48\]
rlabel metal1 5474 14552 5474 14552 0 ct.oc.capture_buffer\[49\]
rlabel via2 16146 15419 16146 15419 0 ct.oc.capture_buffer\[4\]
rlabel metal1 6578 14586 6578 14586 0 ct.oc.capture_buffer\[50\]
rlabel metal1 5014 14586 5014 14586 0 ct.oc.capture_buffer\[51\]
rlabel metal2 9430 15861 9430 15861 0 ct.oc.capture_buffer\[52\]
rlabel metal1 9384 14042 9384 14042 0 ct.oc.capture_buffer\[53\]
rlabel metal1 8924 15538 8924 15538 0 ct.oc.capture_buffer\[54\]
rlabel metal1 8740 14042 8740 14042 0 ct.oc.capture_buffer\[55\]
rlabel metal1 10718 14314 10718 14314 0 ct.oc.capture_buffer\[56\]
rlabel metal2 12742 14994 12742 14994 0 ct.oc.capture_buffer\[57\]
rlabel metal2 12466 14484 12466 14484 0 ct.oc.capture_buffer\[58\]
rlabel metal1 11960 14450 11960 14450 0 ct.oc.capture_buffer\[59\]
rlabel metal1 3358 17850 3358 17850 0 ct.oc.capture_buffer\[5\]
rlabel metal1 12788 14042 12788 14042 0 ct.oc.capture_buffer\[60\]
rlabel metal2 10994 16456 10994 16456 0 ct.oc.capture_buffer\[61\]
rlabel metal1 11730 17748 11730 17748 0 ct.oc.capture_buffer\[62\]
rlabel metal1 10948 15130 10948 15130 0 ct.oc.capture_buffer\[63\]
rlabel metal1 14628 13838 14628 13838 0 ct.oc.capture_buffer\[64\]
rlabel metal1 15548 12818 15548 12818 0 ct.oc.capture_buffer\[65\]
rlabel metal2 13938 14246 13938 14246 0 ct.oc.capture_buffer\[66\]
rlabel metal1 15594 12410 15594 12410 0 ct.oc.capture_buffer\[67\]
rlabel metal1 14766 16014 14766 16014 0 ct.oc.capture_buffer\[68\]
rlabel metal1 14536 16626 14536 16626 0 ct.oc.capture_buffer\[69\]
rlabel metal3 8165 19788 8165 19788 0 ct.oc.capture_buffer\[6\]
rlabel metal1 16698 15470 16698 15470 0 ct.oc.capture_buffer\[70\]
rlabel metal2 14582 15759 14582 15759 0 ct.oc.capture_buffer\[71\]
rlabel metal2 18998 14756 18998 14756 0 ct.oc.capture_buffer\[72\]
rlabel metal1 18216 13906 18216 13906 0 ct.oc.capture_buffer\[73\]
rlabel metal1 18262 13362 18262 13362 0 ct.oc.capture_buffer\[74\]
rlabel metal1 18446 14382 18446 14382 0 ct.oc.capture_buffer\[75\]
rlabel metal1 18676 16762 18676 16762 0 ct.oc.capture_buffer\[76\]
rlabel metal1 16928 16014 16928 16014 0 ct.oc.capture_buffer\[77\]
rlabel metal1 17388 16626 17388 16626 0 ct.oc.capture_buffer\[78\]
rlabel metal2 16422 17238 16422 17238 0 ct.oc.capture_buffer\[79\]
rlabel metal2 9154 21862 9154 21862 0 ct.oc.capture_buffer\[7\]
rlabel metal1 19826 15130 19826 15130 0 ct.oc.capture_buffer\[80\]
rlabel metal1 20010 14042 20010 14042 0 ct.oc.capture_buffer\[81\]
rlabel metal1 21068 13226 21068 13226 0 ct.oc.capture_buffer\[82\]
rlabel metal1 21160 13158 21160 13158 0 ct.oc.capture_buffer\[83\]
rlabel metal2 18998 17408 18998 17408 0 ct.oc.capture_buffer\[84\]
rlabel metal1 21068 17102 21068 17102 0 ct.oc.capture_buffer\[85\]
rlabel viali 22034 16559 22034 16559 0 ct.oc.capture_buffer\[86\]
rlabel metal2 19550 16949 19550 16949 0 ct.oc.capture_buffer\[87\]
rlabel metal2 23046 14824 23046 14824 0 ct.oc.capture_buffer\[88\]
rlabel metal1 24196 14450 24196 14450 0 ct.oc.capture_buffer\[89\]
rlabel metal2 10902 18020 10902 18020 0 ct.oc.capture_buffer\[8\]
rlabel metal1 23920 15538 23920 15538 0 ct.oc.capture_buffer\[90\]
rlabel metal1 22862 14042 22862 14042 0 ct.oc.capture_buffer\[91\]
rlabel metal1 23598 17816 23598 17816 0 ct.oc.capture_buffer\[92\]
rlabel metal1 24564 17714 24564 17714 0 ct.oc.capture_buffer\[93\]
rlabel metal1 25530 17306 25530 17306 0 ct.oc.capture_buffer\[94\]
rlabel metal1 24932 16626 24932 16626 0 ct.oc.capture_buffer\[95\]
rlabel metal1 26312 15130 26312 15130 0 ct.oc.capture_buffer\[96\]
rlabel metal1 26266 15674 26266 15674 0 ct.oc.capture_buffer\[97\]
rlabel metal1 27554 15674 27554 15674 0 ct.oc.capture_buffer\[98\]
rlabel metal2 30406 17680 30406 17680 0 ct.oc.capture_buffer\[99\]
rlabel metal1 11454 18258 11454 18258 0 ct.oc.capture_buffer\[9\]
rlabel metal2 13478 18224 13478 18224 0 ct.oc.data_chain\[0\]
rlabel metal1 25461 19346 25461 19346 0 ct.oc.data_chain\[100\]
rlabel metal1 25208 20842 25208 20842 0 ct.oc.data_chain\[101\]
rlabel metal2 23598 18921 23598 18921 0 ct.oc.data_chain\[102\]
rlabel via1 24611 16560 24611 16560 0 ct.oc.data_chain\[103\]
rlabel metal1 26726 14042 26726 14042 0 ct.oc.data_chain\[104\]
rlabel metal1 27439 16082 27439 16082 0 ct.oc.data_chain\[105\]
rlabel metal1 26979 17170 26979 17170 0 ct.oc.data_chain\[106\]
rlabel metal1 27025 18734 27025 18734 0 ct.oc.data_chain\[107\]
rlabel metal2 29210 17391 29210 17391 0 ct.oc.data_chain\[108\]
rlabel metal1 27393 21522 27393 21522 0 ct.oc.data_chain\[109\]
rlabel metal2 10534 20740 10534 20740 0 ct.oc.data_chain\[10\]
rlabel metal2 22034 20332 22034 20332 0 ct.oc.data_chain\[110\]
rlabel viali 22403 18736 22403 18736 0 ct.oc.data_chain\[111\]
rlabel metal1 25369 13906 25369 13906 0 ct.oc.data_chain\[112\]
rlabel metal1 26685 13294 26685 13294 0 ct.oc.data_chain\[113\]
rlabel metal1 27049 13906 27049 13906 0 ct.oc.data_chain\[114\]
rlabel metal1 25668 12410 25668 12410 0 ct.oc.data_chain\[115\]
rlabel via1 27922 16559 27922 16559 0 ct.oc.data_chain\[116\]
rlabel metal1 28842 12954 28842 12954 0 ct.oc.data_chain\[117\]
rlabel metal1 28888 15130 28888 15130 0 ct.oc.data_chain\[118\]
rlabel metal1 27899 20434 27899 20434 0 ct.oc.data_chain\[119\]
rlabel metal2 12190 19788 12190 19788 0 ct.oc.data_chain\[11\]
rlabel metal1 24289 12800 24289 12800 0 ct.oc.data_chain\[120\]
rlabel metal1 23368 12410 23368 12410 0 ct.oc.data_chain\[121\]
rlabel viali 22403 13294 22403 13294 0 ct.oc.data_chain\[122\]
rlabel metal1 23782 11866 23782 11866 0 ct.oc.data_chain\[123\]
rlabel metal1 26772 11866 26772 11866 0 ct.oc.data_chain\[124\]
rlabel metal1 27508 12818 27508 12818 0 ct.oc.data_chain\[125\]
rlabel metal1 27462 6698 27462 6698 0 ct.oc.data_chain\[126\]
rlabel metal2 28704 15470 28704 15470 0 ct.oc.data_chain\[127\]
rlabel via1 20839 12818 20839 12818 0 ct.oc.data_chain\[128\]
rlabel metal1 21252 11866 21252 11866 0 ct.oc.data_chain\[129\]
rlabel viali 8982 19840 8982 19840 0 ct.oc.data_chain\[12\]
rlabel metal1 20287 13906 20287 13906 0 ct.oc.data_chain\[130\]
rlabel metal1 22425 11730 22425 11730 0 ct.oc.data_chain\[131\]
rlabel metal1 25461 11730 25461 11730 0 ct.oc.data_chain\[132\]
rlabel metal1 28198 11050 28198 11050 0 ct.oc.data_chain\[133\]
rlabel via1 28291 6766 28291 6766 0 ct.oc.data_chain\[134\]
rlabel metal1 28405 7854 28405 7854 0 ct.oc.data_chain\[135\]
rlabel viali 19194 10624 19194 10624 0 ct.oc.data_chain\[136\]
rlabel metal1 19091 11730 19091 11730 0 ct.oc.data_chain\[137\]
rlabel metal1 18492 11866 18492 11866 0 ct.oc.data_chain\[138\]
rlabel metal1 21758 10608 21758 10608 0 ct.oc.data_chain\[139\]
rlabel metal1 7636 19278 7636 19278 0 ct.oc.data_chain\[13\]
rlabel metal1 24565 11120 24565 11120 0 ct.oc.data_chain\[140\]
rlabel metal1 26818 10506 26818 10506 0 ct.oc.data_chain\[141\]
rlabel metal1 27025 8942 27025 8942 0 ct.oc.data_chain\[142\]
rlabel viali 26911 10030 26911 10030 0 ct.oc.data_chain\[143\]
rlabel metal1 17825 10030 17825 10030 0 ct.oc.data_chain\[144\]
rlabel metal1 18193 11118 18193 11118 0 ct.oc.data_chain\[145\]
rlabel metal2 17848 8806 17848 8806 0 ct.oc.data_chain\[146\]
rlabel metal1 21160 8602 21160 8602 0 ct.oc.data_chain\[147\]
rlabel metal1 22517 11118 22517 11118 0 ct.oc.data_chain\[148\]
rlabel metal1 25415 10642 25415 10642 0 ct.oc.data_chain\[149\]
rlabel viali 6624 20433 6624 20433 0 ct.oc.data_chain\[14\]
rlabel metal1 26545 9517 26545 9517 0 ct.oc.data_chain\[150\]
rlabel metal1 24795 10098 24795 10098 0 ct.oc.data_chain\[151\]
rlabel metal2 18262 8823 18262 8823 0 ct.oc.data_chain\[152\]
rlabel metal2 19642 9044 19642 9044 0 ct.oc.data_chain\[153\]
rlabel metal2 19826 8228 19826 8228 0 ct.oc.data_chain\[154\]
rlabel metal1 19481 8466 19481 8466 0 ct.oc.data_chain\[155\]
rlabel metal2 21758 9078 21758 9078 0 ct.oc.data_chain\[156\]
rlabel metal1 24243 9554 24243 9554 0 ct.oc.data_chain\[157\]
rlabel metal1 24059 8466 24059 8466 0 ct.oc.data_chain\[158\]
rlabel metal1 23529 8942 23529 8942 0 ct.oc.data_chain\[159\]
rlabel viali 8881 21521 8881 21521 0 ct.oc.data_chain\[15\]
rlabel metal1 17894 8364 17894 8364 0 ct.oc.data_chain\[160\]
rlabel metal1 21574 8024 21574 8024 0 ct.oc.data_chain\[161\]
rlabel metal2 21758 7004 21758 7004 0 ct.oc.data_chain\[162\]
rlabel metal2 18722 7276 18722 7276 0 ct.oc.data_chain\[163\]
rlabel metal1 23690 8500 23690 8500 0 ct.oc.data_chain\[164\]
rlabel metal1 29624 2618 29624 2618 0 ct.oc.data_chain\[165\]
rlabel viali 22080 7377 22080 7377 0 ct.oc.data_chain\[166\]
rlabel via2 22034 7837 22034 7837 0 ct.oc.data_chain\[167\]
rlabel metal2 16422 5032 16422 5032 0 ct.oc.data_chain\[168\]
rlabel metal2 15962 5712 15962 5712 0 ct.oc.data_chain\[169\]
rlabel metal1 9269 18734 9269 18734 0 ct.oc.data_chain\[16\]
rlabel metal1 13340 986 13340 986 0 ct.oc.data_chain\[170\]
rlabel metal1 21390 3570 21390 3570 0 ct.oc.data_chain\[171\]
rlabel via1 28543 4590 28543 4590 0 ct.oc.data_chain\[172\]
rlabel metal2 21022 3757 21022 3757 0 ct.oc.data_chain\[173\]
rlabel metal2 20562 9860 20562 9860 0 ct.oc.data_chain\[174\]
rlabel metal2 18906 340 18906 340 0 ct.oc.data_chain\[175\]
rlabel metal1 4876 2618 4876 2618 0 ct.oc.data_chain\[176\]
rlabel metal2 1702 2244 1702 2244 0 ct.oc.data_chain\[177\]
rlabel via2 12098 867 12098 867 0 ct.oc.data_chain\[178\]
rlabel metal1 20838 3502 20838 3502 0 ct.oc.data_chain\[179\]
rlabel metal1 10995 18258 10995 18258 0 ct.oc.data_chain\[17\]
rlabel metal2 27554 2346 27554 2346 0 ct.oc.data_chain\[180\]
rlabel metal2 26818 2737 26818 2737 0 ct.oc.data_chain\[181\]
rlabel metal1 16745 10642 16745 10642 0 ct.oc.data_chain\[182\]
rlabel viali 14352 849 14352 849 0 ct.oc.data_chain\[183\]
rlabel metal2 18262 357 18262 357 0 ct.oc.data_chain\[184\]
rlabel viali 4003 1936 4003 1936 0 ct.oc.data_chain\[185\]
rlabel metal1 22793 850 22793 850 0 ct.oc.data_chain\[186\]
rlabel metal1 27301 1938 27301 1938 0 ct.oc.data_chain\[187\]
rlabel metal1 26313 4114 26313 4114 0 ct.oc.data_chain\[188\]
rlabel metal1 26545 2992 26545 2992 0 ct.oc.data_chain\[189\]
rlabel metal1 9637 20434 9637 20434 0 ct.oc.data_chain\[18\]
rlabel metal3 16652 408 16652 408 0 ct.oc.data_chain\[190\]
rlabel via2 17250 3485 17250 3485 0 ct.oc.data_chain\[191\]
rlabel metal1 20746 1224 20746 1224 0 ct.oc.data_chain\[192\]
rlabel metal2 25714 425 25714 425 0 ct.oc.data_chain\[193\]
rlabel metal1 24646 2449 24646 2449 0 ct.oc.data_chain\[194\]
rlabel metal1 26404 5338 26404 5338 0 ct.oc.data_chain\[195\]
rlabel metal1 24725 6290 24725 6290 0 ct.oc.data_chain\[196\]
rlabel metal1 24380 4794 24380 4794 0 ct.oc.data_chain\[197\]
rlabel metal1 20079 850 20079 850 0 ct.oc.data_chain\[198\]
rlabel metal1 26913 1363 26913 1363 0 ct.oc.data_chain\[199\]
rlabel metal1 11133 20434 11133 20434 0 ct.oc.data_chain\[19\]
rlabel metal2 13570 20502 13570 20502 0 ct.oc.data_chain\[1\]
rlabel viali 24335 1920 24335 1920 0 ct.oc.data_chain\[200\]
rlabel metal1 23967 850 23967 850 0 ct.oc.data_chain\[201\]
rlabel viali 22681 3503 22681 3503 0 ct.oc.data_chain\[202\]
rlabel metal1 24243 5202 24243 5202 0 ct.oc.data_chain\[203\]
rlabel viali 23967 5678 23967 5678 0 ct.oc.data_chain\[204\]
rlabel viali 22679 4592 22679 4592 0 ct.oc.data_chain\[205\]
rlabel via1 23967 1326 23967 1326 0 ct.oc.data_chain\[206\]
rlabel metal1 23691 3026 23691 3026 0 ct.oc.data_chain\[207\]
rlabel metal1 21115 1938 21115 1938 0 ct.oc.data_chain\[208\]
rlabel viali 21759 1344 21759 1344 0 ct.oc.data_chain\[209\]
rlabel metal1 5566 19822 5566 19822 0 ct.oc.data_chain\[20\]
rlabel metal1 21115 4114 21115 4114 0 ct.oc.data_chain\[210\]
rlabel metal1 21115 6290 21115 6290 0 ct.oc.data_chain\[211\]
rlabel via1 21759 5678 21759 5678 0 ct.oc.data_chain\[212\]
rlabel metal1 21115 5202 21115 5202 0 ct.oc.data_chain\[213\]
rlabel viali 21761 2415 21761 2415 0 ct.oc.data_chain\[214\]
rlabel metal1 21115 3026 21115 3026 0 ct.oc.data_chain\[215\]
rlabel metal1 18723 1938 18723 1938 0 ct.oc.data_chain\[216\]
rlabel viali 18907 1326 18907 1326 0 ct.oc.data_chain\[217\]
rlabel metal1 18769 4114 18769 4114 0 ct.oc.data_chain\[218\]
rlabel metal1 19091 6290 19091 6290 0 ct.oc.data_chain\[219\]
rlabel metal1 5521 19346 5521 19346 0 ct.oc.data_chain\[21\]
rlabel metal1 18909 5713 18909 5713 0 ct.oc.data_chain\[220\]
rlabel metal1 18769 5202 18769 5202 0 ct.oc.data_chain\[221\]
rlabel viali 18907 2432 18907 2432 0 ct.oc.data_chain\[222\]
rlabel metal1 18815 3026 18815 3026 0 ct.oc.data_chain\[223\]
rlabel viali 16607 1920 16607 1920 0 ct.oc.data_chain\[224\]
rlabel metal1 16331 1326 16331 1326 0 ct.oc.data_chain\[225\]
rlabel metal1 16423 4114 16423 4114 0 ct.oc.data_chain\[226\]
rlabel metal1 16701 4625 16701 4625 0 ct.oc.data_chain\[227\]
rlabel metal1 16701 5713 16701 5713 0 ct.oc.data_chain\[228\]
rlabel metal1 16423 5202 16423 5202 0 ct.oc.data_chain\[229\]
rlabel metal1 5107 21522 5107 21522 0 ct.oc.data_chain\[22\]
rlabel metal1 16331 2414 16331 2414 0 ct.oc.data_chain\[230\]
rlabel metal1 16515 3026 16515 3026 0 ct.oc.data_chain\[231\]
rlabel metal1 13893 1938 13893 1938 0 ct.oc.data_chain\[232\]
rlabel viali 14307 1326 14307 1326 0 ct.oc.data_chain\[233\]
rlabel via1 14491 4114 14491 4114 0 ct.oc.data_chain\[234\]
rlabel via1 14307 4590 14307 4590 0 ct.oc.data_chain\[235\]
rlabel metal1 13846 5338 13846 5338 0 ct.oc.data_chain\[236\]
rlabel metal1 14493 5167 14493 5167 0 ct.oc.data_chain\[237\]
rlabel viali 14307 2414 14307 2414 0 ct.oc.data_chain\[238\]
rlabel metal1 13985 3026 13985 3026 0 ct.oc.data_chain\[239\]
rlabel metal1 4485 20434 4485 20434 0 ct.oc.data_chain\[23\]
rlabel metal1 11455 1938 11455 1938 0 ct.oc.data_chain\[240\]
rlabel metal1 11918 1326 11918 1326 0 ct.oc.data_chain\[241\]
rlabel metal2 12558 3434 12558 3434 0 ct.oc.data_chain\[242\]
rlabel metal1 11454 4454 11454 4454 0 ct.oc.data_chain\[243\]
rlabel via1 11731 5202 11731 5202 0 ct.oc.data_chain\[244\]
rlabel metal1 12053 4608 12053 4608 0 ct.oc.data_chain\[245\]
rlabel metal1 12101 2451 12101 2451 0 ct.oc.data_chain\[246\]
rlabel metal1 11455 3026 11455 3026 0 ct.oc.data_chain\[247\]
rlabel metal1 8879 1938 8879 1938 0 ct.oc.data_chain\[248\]
rlabel metal1 9269 1326 9269 1326 0 ct.oc.data_chain\[249\]
rlabel viali 9157 17169 9157 17169 0 ct.oc.data_chain\[24\]
rlabel metal1 9157 3537 9157 3537 0 ct.oc.data_chain\[250\]
rlabel viali 9157 4591 9157 4591 0 ct.oc.data_chain\[251\]
rlabel metal1 10489 4114 10489 4114 0 ct.oc.data_chain\[252\]
rlabel metal2 9706 5100 9706 5100 0 ct.oc.data_chain\[253\]
rlabel metal1 8832 1530 8832 1530 0 ct.oc.data_chain\[254\]
rlabel metal1 8879 3026 8879 3026 0 ct.oc.data_chain\[255\]
rlabel metal1 6303 1870 6303 1870 0 ct.oc.data_chain\[256\]
rlabel metal1 8695 850 8695 850 0 ct.oc.data_chain\[257\]
rlabel metal1 7360 2618 7360 2618 0 ct.oc.data_chain\[258\]
rlabel metal1 7153 5202 7153 5202 0 ct.oc.data_chain\[259\]
rlabel metal1 8925 18258 8925 18258 0 ct.oc.data_chain\[25\]
rlabel metal2 7866 5270 7866 5270 0 ct.oc.data_chain\[260\]
rlabel metal1 8741 6290 8741 6290 0 ct.oc.data_chain\[261\]
rlabel metal1 4968 986 4968 986 0 ct.oc.data_chain\[262\]
rlabel metal1 6303 3026 6303 3026 0 ct.oc.data_chain\[263\]
rlabel metal1 4554 10234 4554 10234 0 ct.oc.data_chain\[264\]
rlabel metal1 1909 1938 1909 1938 0 ct.oc.data_chain\[265\]
rlabel via1 6303 2414 6303 2414 0 ct.oc.data_chain\[266\]
rlabel metal1 6118 5338 6118 5338 0 ct.oc.data_chain\[267\]
rlabel viali 6487 4592 6487 4592 0 ct.oc.data_chain\[268\]
rlabel metal1 6027 4114 6027 4114 0 ct.oc.data_chain\[269\]
rlabel metal1 8741 19346 8741 19346 0 ct.oc.data_chain\[26\]
rlabel viali 1462 841 1462 841 0 ct.oc.data_chain\[270\]
rlabel metal1 4003 3026 4003 3026 0 ct.oc.data_chain\[271\]
rlabel via2 4002 8483 4002 8483 0 ct.oc.data_chain\[272\]
rlabel viali 1462 16567 1462 16567 0 ct.oc.data_chain\[273\]
rlabel metal1 3036 3162 3036 3162 0 ct.oc.data_chain\[274\]
rlabel metal1 4761 5202 4761 5202 0 ct.oc.data_chain\[275\]
rlabel metal1 3819 4590 3819 4590 0 ct.oc.data_chain\[276\]
rlabel metal1 3542 5338 3542 5338 0 ct.oc.data_chain\[277\]
rlabel metal1 3266 11594 3266 11594 0 ct.oc.data_chain\[278\]
rlabel metal1 1978 3536 1978 3536 0 ct.oc.data_chain\[279\]
rlabel metal1 9157 17681 9157 17681 0 ct.oc.data_chain\[27\]
rlabel via3 14053 18020 14053 18020 0 ct.oc.data_chain\[280\]
rlabel metal1 1748 13906 1748 13906 0 ct.oc.data_chain\[281\]
rlabel viali 1472 3017 1472 3017 0 ct.oc.data_chain\[282\]
rlabel metal1 4439 6290 4439 6290 0 ct.oc.data_chain\[283\]
rlabel metal1 1978 5712 1978 5712 0 ct.oc.data_chain\[284\]
rlabel metal2 2162 6188 2162 6188 0 ct.oc.data_chain\[285\]
rlabel metal1 2116 4794 2116 4794 0 ct.oc.data_chain\[286\]
rlabel metal1 2162 4080 2162 4080 0 ct.oc.data_chain\[287\]
rlabel metal1 1702 8976 1702 8976 0 ct.oc.data_chain\[288\]
rlabel metal1 2323 8466 2323 8466 0 ct.oc.data_chain\[289\]
rlabel metal1 4025 19346 4025 19346 0 ct.oc.data_chain\[28\]
rlabel metal1 1633 7854 1633 7854 0 ct.oc.data_chain\[290\]
rlabel metal1 3841 6766 3841 6766 0 ct.oc.data_chain\[291\]
rlabel metal1 2162 6800 2162 6800 0 ct.oc.data_chain\[292\]
rlabel metal1 2116 7378 2116 7378 0 ct.oc.data_chain\[293\]
rlabel metal2 1518 4522 1518 4522 0 ct.oc.data_chain\[294\]
rlabel metal2 10258 7242 10258 7242 0 ct.oc.data_chain\[295\]
rlabel metal2 13478 8007 13478 8007 0 ct.oc.data_chain\[296\]
rlabel metal2 15226 6409 15226 6409 0 ct.oc.data_chain\[297\]
rlabel metal2 15318 7021 15318 7021 0 ct.oc.data_chain\[298\]
rlabel metal2 16238 6579 16238 6579 0 ct.oc.data_chain\[299\]
rlabel viali 3590 19824 3590 19824 0 ct.oc.data_chain\[29\]
rlabel metal2 11178 20400 11178 20400 0 ct.oc.data_chain\[2\]
rlabel via2 13754 6851 13754 6851 0 ct.oc.data_chain\[300\]
rlabel metal1 10718 7446 10718 7446 0 ct.oc.data_chain\[301\]
rlabel metal2 11178 6596 11178 6596 0 ct.oc.data_chain\[302\]
rlabel metal2 13202 7344 13202 7344 0 ct.oc.data_chain\[303\]
rlabel metal1 12213 7854 12213 7854 0 ct.oc.data_chain\[304\]
rlabel metal1 15065 7378 15065 7378 0 ct.oc.data_chain\[305\]
rlabel metal1 14835 7854 14835 7854 0 ct.oc.data_chain\[306\]
rlabel metal1 14973 6290 14973 6290 0 ct.oc.data_chain\[307\]
rlabel metal1 14421 6766 14421 6766 0 ct.oc.data_chain\[308\]
rlabel metal2 12374 8636 12374 8636 0 ct.oc.data_chain\[309\]
rlabel metal1 3266 21590 3266 21590 0 ct.oc.data_chain\[30\]
rlabel metal2 12466 7820 12466 7820 0 ct.oc.data_chain\[310\]
rlabel metal2 12834 7786 12834 7786 0 ct.oc.data_chain\[311\]
rlabel metal1 14145 8466 14145 8466 0 ct.oc.data_chain\[312\]
rlabel metal2 14214 12818 14214 12818 0 ct.oc.data_chain\[313\]
rlabel metal1 14145 10030 14145 10030 0 ct.oc.data_chain\[314\]
rlabel metal1 14559 9554 14559 9554 0 ct.oc.data_chain\[315\]
rlabel metal1 13709 10642 13709 10642 0 ct.oc.data_chain\[316\]
rlabel metal1 10672 9622 10672 9622 0 ct.oc.data_chain\[317\]
rlabel metal1 10948 9894 10948 9894 0 ct.oc.data_chain\[318\]
rlabel viali 11455 8944 11455 8944 0 ct.oc.data_chain\[319\]
rlabel metal2 3082 21522 3082 21522 0 ct.oc.data_chain\[31\]
rlabel metal1 12929 11152 12929 11152 0 ct.oc.data_chain\[320\]
rlabel metal1 10764 12410 10764 12410 0 ct.oc.data_chain\[321\]
rlabel metal1 12835 12206 12835 12206 0 ct.oc.data_chain\[322\]
rlabel viali 14076 11729 14076 11729 0 ct.oc.data_chain\[323\]
rlabel viali 11733 11721 11733 11721 0 ct.oc.data_chain\[324\]
rlabel metal1 9269 9554 9269 9554 0 ct.oc.data_chain\[325\]
rlabel metal1 9157 10065 9157 10065 0 ct.oc.data_chain\[326\]
rlabel metal1 9615 8466 9615 8466 0 ct.oc.data_chain\[327\]
rlabel metal1 8234 12716 8234 12716 0 ct.oc.data_chain\[328\]
rlabel metal1 9157 12241 9157 12241 0 ct.oc.data_chain\[329\]
rlabel metal1 6303 17170 6303 17170 0 ct.oc.data_chain\[32\]
rlabel metal2 9706 14195 9706 14195 0 ct.oc.data_chain\[330\]
rlabel metal1 9201 11730 9201 11730 0 ct.oc.data_chain\[331\]
rlabel metal1 10029 10642 10029 10642 0 ct.oc.data_chain\[332\]
rlabel via1 8051 8942 8051 8942 0 ct.oc.data_chain\[333\]
rlabel metal1 7061 10030 7061 10030 0 ct.oc.data_chain\[334\]
rlabel via1 6579 9554 6579 9554 0 ct.oc.data_chain\[335\]
rlabel metal1 5981 12818 5981 12818 0 ct.oc.data_chain\[336\]
rlabel metal1 6440 14042 6440 14042 0 ct.oc.data_chain\[337\]
rlabel metal2 5658 13821 5658 13821 0 ct.oc.data_chain\[338\]
rlabel metal1 6624 12954 6624 12954 0 ct.oc.data_chain\[339\]
rlabel viali 6949 17647 6949 17647 0 ct.oc.data_chain\[33\]
rlabel metal1 7225 11153 7225 11153 0 ct.oc.data_chain\[340\]
rlabel metal1 5935 10642 5935 10642 0 ct.oc.data_chain\[341\]
rlabel metal1 5566 10030 5566 10030 0 ct.oc.data_chain\[342\]
rlabel metal1 5981 11730 5981 11730 0 ct.oc.data_chain\[343\]
rlabel metal1 3726 12954 3726 12954 0 ct.oc.data_chain\[344\]
rlabel metal1 4462 13906 4462 13906 0 ct.oc.data_chain\[345\]
rlabel metal1 3819 13294 3819 13294 0 ct.oc.data_chain\[346\]
rlabel metal1 4325 12818 4325 12818 0 ct.oc.data_chain\[347\]
rlabel viali 4014 12208 4014 12208 0 ct.oc.data_chain\[348\]
rlabel metal1 3451 9554 3451 9554 0 ct.oc.data_chain\[349\]
rlabel metal1 6164 18394 6164 18394 0 ct.oc.data_chain\[34\]
rlabel via1 3727 10030 3727 10030 0 ct.oc.data_chain\[350\]
rlabel viali 3729 8951 3729 8951 0 ct.oc.data_chain\[351\]
rlabel metal1 6119 18258 6119 18258 0 ct.oc.data_chain\[35\]
rlabel viali 2899 18736 2899 18736 0 ct.oc.data_chain\[36\]
rlabel metal2 2806 19142 2806 19142 0 ct.oc.data_chain\[37\]
rlabel metal1 3589 21522 3589 21522 0 ct.oc.data_chain\[38\]
rlabel metal1 4094 19142 4094 19142 0 ct.oc.data_chain\[39\]
rlabel metal2 13018 19890 13018 19890 0 ct.oc.data_chain\[3\]
rlabel metal1 4853 17170 4853 17170 0 ct.oc.data_chain\[40\]
rlabel metal1 6118 14858 6118 14858 0 ct.oc.data_chain\[41\]
rlabel via1 4371 18258 4371 18258 0 ct.oc.data_chain\[42\]
rlabel viali 4005 17655 4005 17655 0 ct.oc.data_chain\[43\]
rlabel metal2 3174 16966 3174 16966 0 ct.oc.data_chain\[44\]
rlabel metal1 1610 17680 1610 17680 0 ct.oc.data_chain\[45\]
rlabel metal1 1518 19856 1518 19856 0 ct.oc.data_chain\[46\]
rlabel metal2 2070 17782 2070 17782 0 ct.oc.data_chain\[47\]
rlabel metal1 5037 15470 5037 15470 0 ct.oc.data_chain\[48\]
rlabel metal1 5267 14994 5267 14994 0 ct.oc.data_chain\[49\]
rlabel metal1 3729 20298 3729 20298 0 ct.oc.data_chain\[4\]
rlabel viali 4005 16559 4005 16559 0 ct.oc.data_chain\[50\]
rlabel metal1 5221 16082 5221 16082 0 ct.oc.data_chain\[51\]
rlabel metal1 1978 15504 1978 15504 0 ct.oc.data_chain\[52\]
rlabel metal2 3542 15283 3542 15283 0 ct.oc.data_chain\[53\]
rlabel metal1 2116 17170 2116 17170 0 ct.oc.data_chain\[54\]
rlabel metal1 1426 16073 1426 16073 0 ct.oc.data_chain\[55\]
rlabel metal1 10074 13872 10074 13872 0 ct.oc.data_chain\[56\]
rlabel metal2 13110 15776 13110 15776 0 ct.oc.data_chain\[57\]
rlabel metal1 9338 14960 9338 14960 0 ct.oc.data_chain\[58\]
rlabel metal2 12374 14144 12374 14144 0 ct.oc.data_chain\[59\]
rlabel metal2 8786 21488 8786 21488 0 ct.oc.data_chain\[5\]
rlabel metal2 13018 16813 13018 16813 0 ct.oc.data_chain\[60\]
rlabel metal2 12834 16711 12834 16711 0 ct.oc.data_chain\[61\]
rlabel metal2 13662 17289 13662 17289 0 ct.oc.data_chain\[62\]
rlabel metal2 13110 16592 13110 16592 0 ct.oc.data_chain\[63\]
rlabel metal1 13662 15402 13662 15402 0 ct.oc.data_chain\[64\]
rlabel via1 11731 16080 11731 16080 0 ct.oc.data_chain\[65\]
rlabel metal2 15410 14824 15410 14824 0 ct.oc.data_chain\[66\]
rlabel metal1 13754 14484 13754 14484 0 ct.oc.data_chain\[67\]
rlabel metal1 15686 15878 15686 15878 0 ct.oc.data_chain\[68\]
rlabel metal1 12213 16558 12213 16558 0 ct.oc.data_chain\[69\]
rlabel metal1 1610 21080 1610 21080 0 ct.oc.data_chain\[6\]
rlabel metal1 13938 17578 13938 17578 0 ct.oc.data_chain\[70\]
rlabel metal2 13478 16422 13478 16422 0 ct.oc.data_chain\[71\]
rlabel metal1 15571 13906 15571 13906 0 ct.oc.data_chain\[72\]
rlabel metal1 15157 12818 15157 12818 0 ct.oc.data_chain\[73\]
rlabel viali 14352 14383 14352 14383 0 ct.oc.data_chain\[74\]
rlabel metal1 15939 14994 15939 14994 0 ct.oc.data_chain\[75\]
rlabel metal1 15387 16082 15387 16082 0 ct.oc.data_chain\[76\]
rlabel viali 14307 16560 14307 16560 0 ct.oc.data_chain\[77\]
rlabel metal1 15571 17170 15571 17170 0 ct.oc.data_chain\[78\]
rlabel metal1 15387 15470 15387 15470 0 ct.oc.data_chain\[79\]
rlabel metal1 8418 16694 8418 16694 0 ct.oc.data_chain\[7\]
rlabel metal1 17641 15470 17641 15470 0 ct.oc.data_chain\[80\]
rlabel metal1 21206 14314 21206 14314 0 ct.oc.data_chain\[81\]
rlabel metal2 21298 13770 21298 13770 0 ct.oc.data_chain\[82\]
rlabel metal1 20838 15504 20838 15504 0 ct.oc.data_chain\[83\]
rlabel via2 17894 17187 17894 17187 0 ct.oc.data_chain\[84\]
rlabel metal2 17894 16303 17894 16303 0 ct.oc.data_chain\[85\]
rlabel metal1 21229 16762 21229 16762 0 ct.oc.data_chain\[86\]
rlabel metal2 17526 18020 17526 18020 0 ct.oc.data_chain\[87\]
rlabel metal1 21574 15946 21574 15946 0 ct.oc.data_chain\[88\]
rlabel metal1 21114 14926 21114 14926 0 ct.oc.data_chain\[89\]
rlabel metal1 13617 19346 13617 19346 0 ct.oc.data_chain\[8\]
rlabel metal2 21942 14858 21942 14858 0 ct.oc.data_chain\[90\]
rlabel metal1 21942 15504 21942 15504 0 ct.oc.data_chain\[91\]
rlabel via1 21759 17646 21759 17646 0 ct.oc.data_chain\[92\]
rlabel metal1 21482 17170 21482 17170 0 ct.oc.data_chain\[93\]
rlabel metal1 21804 16593 21804 16593 0 ct.oc.data_chain\[94\]
rlabel metal2 22862 17374 22862 17374 0 ct.oc.data_chain\[95\]
rlabel viali 24335 16080 24335 16080 0 ct.oc.data_chain\[96\]
rlabel metal1 24265 14382 24265 14382 0 ct.oc.data_chain\[97\]
rlabel metal1 24357 15470 24357 15470 0 ct.oc.data_chain\[98\]
rlabel metal1 24587 14994 24587 14994 0 ct.oc.data_chain\[99\]
rlabel via1 12651 19822 12651 19822 0 ct.oc.data_chain\[9\]
rlabel metal2 12466 19193 12466 19193 0 ct.oc.mode_buffer\[0\]
rlabel via1 21645 15470 21645 15470 0 ct.oc.mode_buffer\[10\]
rlabel via1 25165 18054 25165 18054 0 ct.oc.mode_buffer\[11\]
rlabel metal1 26935 21454 26935 21454 0 ct.oc.mode_buffer\[12\]
rlabel via1 28845 20026 28845 20026 0 ct.oc.mode_buffer\[13\]
rlabel metal1 27327 14790 27327 14790 0 ct.oc.mode_buffer\[14\]
rlabel metal1 29762 11798 29762 11798 0 ct.oc.mode_buffer\[15\]
rlabel metal1 20292 10438 20292 10438 0 ct.oc.mode_buffer\[16\]
rlabel metal1 17253 11322 17253 11322 0 ct.oc.mode_buffer\[17\]
rlabel metal1 23163 9010 23163 9010 0 ct.oc.mode_buffer\[18\]
rlabel metal1 18357 8058 18357 8058 0 ct.oc.mode_buffer\[19\]
rlabel metal1 11319 20230 11319 20230 0 ct.oc.mode_buffer\[1\]
rlabel metal1 28361 3570 28361 3570 0 ct.oc.mode_buffer\[20\]
rlabel metal2 2070 2295 2070 2295 0 ct.oc.mode_buffer\[21\]
rlabel metal2 13570 2176 13570 2176 0 ct.oc.mode_buffer\[22\]
rlabel metal1 7590 408 7590 408 0 ct.oc.mode_buffer\[23\]
rlabel metal1 23991 1394 23991 1394 0 ct.oc.mode_buffer\[24\]
rlabel metal1 21669 5882 21669 5882 0 ct.oc.mode_buffer\[25\]
rlabel via1 18793 2482 18793 2482 0 ct.oc.mode_buffer\[26\]
rlabel metal1 16655 2618 16655 2618 0 ct.oc.mode_buffer\[27\]
rlabel via1 14193 2414 14193 2414 0 ct.oc.mode_buffer\[28\]
rlabel metal1 11825 4998 11825 4998 0 ct.oc.mode_buffer\[29\]
rlabel via1 1429 21318 1429 21318 0 ct.oc.mode_buffer\[2\]
rlabel metal1 9111 2618 9111 2618 0 ct.oc.mode_buffer\[30\]
rlabel metal1 7593 1530 7593 1530 0 ct.oc.mode_buffer\[31\]
rlabel metal1 4695 10438 4695 10438 0 ct.oc.mode_buffer\[32\]
rlabel metal1 2165 16762 2165 16762 0 ct.oc.mode_buffer\[33\]
rlabel via1 1429 13702 1429 13702 0 ct.oc.mode_buffer\[34\]
rlabel metal1 1221 4590 1221 4590 0 ct.oc.mode_buffer\[35\]
rlabel metal1 5112 7174 5112 7174 0 ct.oc.mode_buffer\[36\]
rlabel metal1 13846 7208 13846 7208 0 ct.oc.mode_buffer\[37\]
rlabel via1 13917 10030 13917 10030 0 ct.oc.mode_buffer\[38\]
rlabel metal1 13846 12818 13846 12818 0 ct.oc.mode_buffer\[39\]
rlabel metal1 1380 18870 1380 18870 0 ct.oc.mode_buffer\[3\]
rlabel metal2 9614 13158 9614 13158 0 ct.oc.mode_buffer\[40\]
rlabel via1 7201 13294 7201 13294 0 ct.oc.mode_buffer\[41\]
rlabel metal1 3913 9350 3913 9350 0 ct.oc.mode_buffer\[42\]
rlabel via1 1429 9350 1429 9350 0 ct.oc.mode_buffer\[43\]
rlabel metal1 1889 17850 1889 17850 0 ct.oc.mode_buffer\[4\]
rlabel via1 1429 15878 1429 15878 0 ct.oc.mode_buffer\[5\]
rlabel metal1 6535 14790 6535 14790 0 ct.oc.mode_buffer\[6\]
rlabel via1 12169 18734 12169 18734 0 ct.oc.mode_buffer\[7\]
rlabel metal1 14996 13294 14996 13294 0 ct.oc.mode_buffer\[8\]
rlabel metal1 17391 16762 17391 16762 0 ct.oc.mode_buffer\[9\]
rlabel metal1 17158 15470 17158 15470 0 ct.oc.trig_chain\[10\]
rlabel metal1 19182 16048 19182 16048 0 ct.oc.trig_chain\[11\]
rlabel metal1 24702 18292 24702 18292 0 ct.oc.trig_chain\[12\]
rlabel metal1 29118 14824 29118 14824 0 ct.oc.trig_chain\[13\]
rlabel metal1 28428 19890 28428 19890 0 ct.oc.trig_chain\[14\]
rlabel metal1 26772 14926 26772 14926 0 ct.oc.trig_chain\[15\]
rlabel metal1 26634 8466 26634 8466 0 ct.oc.trig_chain\[16\]
rlabel metal2 26450 9520 26450 9520 0 ct.oc.trig_chain\[17\]
rlabel metal1 16790 11118 16790 11118 0 ct.oc.trig_chain\[18\]
rlabel metal1 17756 7310 17756 7310 0 ct.oc.trig_chain\[19\]
rlabel metal1 8464 19890 8464 19890 0 ct.oc.trig_chain\[1\]
rlabel metal1 17940 7922 17940 7922 0 ct.oc.trig_chain\[20\]
rlabel metal1 23920 7854 23920 7854 0 ct.oc.trig_chain\[21\]
rlabel metal2 1886 2567 1886 2567 0 ct.oc.trig_chain\[22\]
rlabel metal1 3266 2346 3266 2346 0 ct.oc.trig_chain\[23\]
rlabel metal2 5842 408 5842 408 0 ct.oc.trig_chain\[24\]
rlabel metal2 23874 2244 23874 2244 0 ct.oc.trig_chain\[25\]
rlabel metal1 21114 2482 21114 2482 0 ct.oc.trig_chain\[26\]
rlabel metal1 18538 1326 18538 1326 0 ct.oc.trig_chain\[27\]
rlabel metal1 16192 2482 16192 2482 0 ct.oc.trig_chain\[28\]
rlabel metal1 13938 2414 13938 2414 0 ct.oc.trig_chain\[29\]
rlabel metal2 10810 16388 10810 16388 0 ct.oc.trig_chain\[2\]
rlabel metal2 12098 3740 12098 3740 0 ct.oc.trig_chain\[30\]
rlabel metal1 10120 4114 10120 4114 0 ct.oc.trig_chain\[31\]
rlabel metal1 8188 5678 8188 5678 0 ct.oc.trig_chain\[32\]
rlabel metal1 3404 10438 3404 10438 0 ct.oc.trig_chain\[33\]
rlabel metal2 920 16626 920 16626 0 ct.oc.trig_chain\[34\]
rlabel metal1 1104 13838 1104 13838 0 ct.oc.trig_chain\[35\]
rlabel metal1 920 6222 920 6222 0 ct.oc.trig_chain\[36\]
rlabel metal1 11086 8024 11086 8024 0 ct.oc.trig_chain\[37\]
rlabel metal2 13846 7072 13846 7072 0 ct.oc.trig_chain\[38\]
rlabel metal2 13570 10336 13570 10336 0 ct.oc.trig_chain\[39\]
rlabel metal1 966 21590 966 21590 0 ct.oc.trig_chain\[3\]
rlabel metal2 12512 12274 12512 12274 0 ct.oc.trig_chain\[40\]
rlabel metal1 8050 10506 8050 10506 0 ct.oc.trig_chain\[41\]
rlabel metal2 6854 13872 6854 13872 0 ct.oc.trig_chain\[42\]
rlabel metal1 3312 9486 3312 9486 0 ct.oc.trig_chain\[43\]
rlabel metal1 1426 13294 1426 13294 0 ct.oc.trig_chain\[44\]
rlabel metal1 1518 18802 1518 18802 0 ct.oc.trig_chain\[4\]
rlabel metal1 920 19346 920 19346 0 ct.oc.trig_chain\[5\]
rlabel metal1 1334 15402 1334 15402 0 ct.oc.trig_chain\[6\]
rlabel metal1 8694 15402 8694 15402 0 ct.oc.trig_chain\[7\]
rlabel metal1 11776 18734 11776 18734 0 ct.oc.trig_chain\[8\]
rlabel metal1 14214 13770 14214 13770 0 ct.oc.trig_chain\[9\]
rlabel metal1 20424 18258 20424 18258 0 ct.ro.counter\[0\]
rlabel metal2 21298 21284 21298 21284 0 ct.ro.counter\[1\]
rlabel metal2 21574 20876 21574 20876 0 ct.ro.counter\[2\]
rlabel metal2 22218 21284 22218 21284 0 ct.ro.counter\[3\]
rlabel metal2 24058 21420 24058 21420 0 ct.ro.counter\[4\]
rlabel metal1 23920 21522 23920 21522 0 ct.ro.counter\[5\]
rlabel metal1 24150 20230 24150 20230 0 ct.ro.counter\[6\]
rlabel metal1 25576 20230 25576 20230 0 ct.ro.counter\[7\]
rlabel metal2 20562 20400 20562 20400 0 ct.ro.counter_n\[0\]
rlabel metal1 20148 20910 20148 20910 0 ct.ro.counter_n\[1\]
rlabel metal1 21160 20366 21160 20366 0 ct.ro.counter_n\[2\]
rlabel metal1 23322 20944 23322 20944 0 ct.ro.counter_n\[3\]
rlabel metal1 23690 20910 23690 20910 0 ct.ro.counter_n\[4\]
rlabel metal1 21574 20332 21574 20332 0 ct.ro.counter_n\[5\]
rlabel metal1 23598 20400 23598 20400 0 ct.ro.counter_n\[6\]
rlabel metal1 25898 20400 25898 20400 0 ct.ro.counter_n\[7\]
rlabel metal1 19136 18122 19136 18122 0 ct.ro.gate
rlabel metal1 19826 18265 19826 18265 0 ct.ro.ring\[0\]
rlabel metal1 16698 21522 16698 21522 0 ct.ro.ring\[1\]
rlabel metal1 17756 21522 17756 21522 0 ct.ro.ring\[2\]
rlabel metal1 23920 18054 23920 18054 0 net1
rlabel metal1 16882 6834 16882 6834 0 net10
rlabel metal1 5750 10098 5750 10098 0 net11
rlabel metal1 12328 9486 12328 9486 0 net12
rlabel metal1 29302 1904 29302 1904 0 net13
rlabel metal1 18998 17102 18998 17102 0 net14
rlabel metal2 12650 8109 12650 8109 0 net15
rlabel metal1 13570 6222 13570 6222 0 net16
rlabel metal1 13018 9078 13018 9078 0 net17
rlabel metal2 18630 6392 18630 6392 0 net18
rlabel metal1 18630 17680 18630 17680 0 net19
rlabel metal1 23046 18326 23046 18326 0 net2
rlabel metal1 1196 13362 1196 13362 0 net20
rlabel metal1 14214 6222 14214 6222 0 net21
rlabel metal1 14122 17238 14122 17238 0 net22
rlabel metal1 21666 9010 21666 9010 0 net23
rlabel metal1 30498 17306 30498 17306 0 net24
rlabel metal2 2070 1564 2070 1564 0 net25
rlabel metal1 4508 14450 4508 14450 0 net26
rlabel metal1 13478 20876 13478 20876 0 net27
rlabel metal1 19734 9010 19734 9010 0 net28
rlabel metal2 30406 16422 30406 16422 0 net29
rlabel metal2 21114 20842 21114 20842 0 net3
rlabel metal1 13570 14858 13570 14858 0 net30
rlabel metal3 19780 3128 19780 3128 0 net31
rlabel metal1 8142 21046 8142 21046 0 net32
rlabel metal1 13386 21488 13386 21488 0 net33
rlabel metal1 27738 7990 27738 7990 0 net34
rlabel metal1 16698 12920 16698 12920 0 net35
rlabel metal1 16652 6834 16652 6834 0 net36
rlabel metal1 6486 13396 6486 13396 0 net37
rlabel metal2 11132 19652 11132 19652 0 net38
rlabel metal1 21482 748 21482 748 0 net39
rlabel metal1 24518 19414 24518 19414 0 net4
rlabel metal1 19182 12852 19182 12852 0 net40
rlabel metal2 17802 18003 17802 18003 0 net41
rlabel metal2 12650 10404 12650 10404 0 net42
rlabel metal1 5244 21454 5244 21454 0 net43
rlabel metal1 21068 19210 21068 19210 0 net44
rlabel metal2 21114 1479 21114 1479 0 net45
rlabel metal2 17066 10540 17066 10540 0 net46
rlabel metal1 30498 14960 30498 14960 0 net47
rlabel metal1 13616 2958 13616 2958 0 net48
rlabel metal1 13156 9894 13156 9894 0 net49
rlabel metal1 16882 7344 16882 7344 0 net5
rlabel metal1 1058 20978 1058 20978 0 net50
rlabel metal1 20654 2414 20654 2414 0 net51
rlabel metal2 19642 19788 19642 19788 0 net52
rlabel metal2 18998 20876 18998 20876 0 net53
rlabel metal2 20838 18989 20838 18989 0 net54
rlabel metal2 21114 18921 21114 18921 0 net55
rlabel metal2 18722 17391 18722 17391 0 net56
rlabel metal1 16146 21590 16146 21590 0 net57
rlabel metal2 6578 15759 6578 15759 0 net58
rlabel metal2 8602 14705 8602 14705 0 net59
rlabel metal1 10810 4046 10810 4046 0 net6
rlabel metal2 9338 13294 9338 13294 0 net60
rlabel metal2 7682 13243 7682 13243 0 net61
rlabel metal1 11178 19482 11178 19482 0 net7
rlabel metal1 18538 1802 18538 1802 0 net8
rlabel metal1 16606 16694 16606 16694 0 net9
rlabel metal1 25031 20978 25031 20978 0 rst_n
rlabel metal2 18446 21454 18446 21454 0 ui_in[0]
rlabel metal1 18722 21012 18722 21012 0 ui_in[1]
rlabel metal1 17710 18088 17710 18088 0 ui_in[2]
rlabel metal4 24196 21457 24196 21457 0 ui_in[3]
rlabel metal1 18768 20434 18768 20434 0 ui_in[4]
rlabel metal4 23092 22069 23092 22069 0 ui_in[5]
rlabel metal4 22540 21457 22540 21457 0 ui_in[6]
rlabel metal4 21988 22069 21988 22069 0 ui_in[7]
rlabel metal4 12604 20165 12604 20165 0 uio_out[0]
rlabel metal2 12466 21539 12466 21539 0 uio_out[1]
rlabel metal2 8326 19584 8326 19584 0 uio_out[2]
rlabel metal2 12558 20519 12558 20519 0 uio_out[3]
rlabel via2 10350 20587 10350 20587 0 uio_out[4]
rlabel metal4 9844 22137 9844 22137 0 uio_out[5]
rlabel metal2 1978 21658 1978 21658 0 uio_out[6]
rlabel metal1 8510 16762 8510 16762 0 uio_out[7]
rlabel metal1 18400 21114 18400 21114 0 uo_out[0]
rlabel metal1 18032 18258 18032 18258 0 uo_out[1]
rlabel metal1 16468 20026 16468 20026 0 uo_out[2]
rlabel metal1 16100 18666 16100 18666 0 uo_out[3]
rlabel metal4 14812 21457 14812 21457 0 uo_out[4]
rlabel metal1 15502 19686 15502 19686 0 uo_out[5]
rlabel metal1 14950 20570 14950 20570 0 uo_out[6]
rlabel metal1 15594 21114 15594 21114 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 31464 22304
<< end >>
