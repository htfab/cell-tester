magic
tech sky130A
magscale 1 2
timestamp 1698890999
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1931 203
rect 29 -17 63 21
<< scnmos >>
rect 81 47 111 177
rect 165 47 195 177
rect 353 47 383 177
rect 437 47 467 177
rect 533 47 563 177
rect 617 47 647 177
rect 781 47 811 177
rect 865 47 895 177
rect 1617 47 1647 177
rect 1701 47 1731 177
rect 1785 47 1815 177
rect 1053 47 1083 177
rect 1149 47 1179 177
rect 1233 47 1263 177
rect 1329 47 1359 177
rect 1413 47 1443 177
<< scpmoshvt >>
rect 81 297 111 497
rect 165 297 195 497
rect 353 297 383 497
rect 437 297 467 497
rect 533 297 563 497
rect 617 297 647 497
rect 781 297 811 497
rect 865 297 895 497
rect 1617 297 1647 497
rect 1701 297 1731 497
rect 1785 297 1815 497
rect 1053 297 1083 497
rect 1149 297 1179 497
rect 1233 297 1263 497
rect 1329 297 1359 497
rect 1413 297 1443 497
<< ndiff >>
rect 811 47 865 177
rect 1565 47 1617 59
rect 1565 59 1573 93
rect 1607 59 1617 93
rect 1565 93 1617 177
rect 301 47 353 59
rect 301 59 309 93
rect 343 59 353 93
rect 301 93 353 127
rect 301 127 309 161
rect 343 127 353 161
rect 301 161 353 177
rect 29 47 81 67
rect 29 67 37 101
rect 71 67 81 101
rect 29 101 81 177
rect 111 47 165 59
rect 111 59 121 93
rect 155 59 165 93
rect 111 93 165 177
rect 195 47 247 67
rect 195 67 205 101
rect 239 67 247 101
rect 195 101 247 177
rect 383 47 437 177
rect 467 47 533 127
rect 467 127 489 161
rect 523 127 533 161
rect 467 161 533 177
rect 563 47 617 59
rect 563 59 573 93
rect 607 59 617 93
rect 563 93 617 177
rect 647 47 781 59
rect 647 59 657 93
rect 691 59 781 93
rect 647 93 781 177
rect 1001 47 1053 59
rect 1001 59 1009 93
rect 1043 59 1053 93
rect 1001 93 1053 177
rect 895 47 947 59
rect 895 59 905 93
rect 939 59 947 93
rect 895 93 947 177
rect 1647 47 1701 177
rect 1731 47 1785 59
rect 1731 59 1741 93
rect 1775 59 1785 93
rect 1731 93 1785 177
rect 1815 47 1867 59
rect 1815 59 1825 93
rect 1859 59 1867 93
rect 1815 93 1867 177
rect 1083 47 1149 67
rect 1083 67 1093 101
rect 1127 67 1149 101
rect 1083 101 1149 177
rect 1179 47 1233 127
rect 1179 127 1189 161
rect 1223 127 1233 161
rect 1179 161 1233 177
rect 1263 47 1329 59
rect 1263 59 1285 93
rect 1319 59 1329 93
rect 1263 93 1329 177
rect 1359 47 1413 59
rect 1359 59 1369 93
rect 1403 59 1413 93
rect 1359 93 1413 177
rect 1443 47 1511 59
rect 1443 59 1469 93
rect 1503 59 1511 93
rect 1443 93 1511 177
<< pdiff >>
rect 1359 297 1413 497
rect 1443 297 1511 451
rect 1443 451 1469 485
rect 1503 451 1511 485
rect 1443 485 1511 497
rect 1001 297 1053 443
rect 1001 443 1009 477
rect 1043 443 1053 477
rect 1001 477 1053 497
rect 1565 297 1617 383
rect 1565 383 1573 417
rect 1607 383 1617 417
rect 1565 417 1617 451
rect 1565 451 1573 485
rect 1607 451 1617 485
rect 1565 485 1617 497
rect 301 297 353 383
rect 301 383 309 417
rect 343 383 353 417
rect 301 417 353 451
rect 301 451 309 485
rect 343 451 353 485
rect 301 485 353 497
rect 29 297 81 375
rect 29 375 37 409
rect 71 375 81 409
rect 29 409 81 443
rect 29 443 37 477
rect 71 443 81 477
rect 29 477 81 497
rect 111 297 165 451
rect 111 451 121 485
rect 155 451 165 485
rect 111 485 165 497
rect 195 297 247 443
rect 195 443 205 477
rect 239 443 247 477
rect 195 477 247 497
rect 383 297 437 443
rect 383 443 393 477
rect 427 443 437 477
rect 383 477 437 497
rect 467 297 533 443
rect 467 443 489 477
rect 523 443 533 477
rect 467 477 533 497
rect 563 297 617 451
rect 563 451 573 485
rect 607 451 617 485
rect 563 485 617 497
rect 811 297 865 451
rect 811 451 821 485
rect 855 451 865 485
rect 811 485 865 497
rect 895 297 947 443
rect 895 443 905 477
rect 939 443 947 477
rect 895 477 947 497
rect 1647 297 1701 443
rect 1647 443 1657 477
rect 1691 443 1701 477
rect 1647 477 1701 497
rect 1731 297 1785 451
rect 1731 451 1741 485
rect 1775 451 1785 485
rect 1731 485 1785 497
rect 1815 297 1867 451
rect 1815 451 1825 485
rect 1859 451 1867 485
rect 1815 485 1867 497
rect 1083 297 1149 443
rect 1083 443 1105 477
rect 1139 443 1149 477
rect 1083 477 1149 497
rect 1179 297 1233 443
rect 1179 443 1189 477
rect 1223 443 1233 477
rect 1179 477 1233 497
rect 1263 297 1329 451
rect 1263 451 1285 485
rect 1319 451 1329 485
rect 1263 485 1329 497
rect 647 297 781 443
rect 647 443 737 477
rect 771 443 781 477
rect 647 477 781 497
<< ndiffc >>
rect 309 127 343 161
rect 489 127 523 161
rect 1189 127 1223 161
rect 1093 67 1127 101
rect 37 67 71 101
rect 205 67 239 101
rect 905 59 939 93
rect 1469 59 1503 93
rect 1573 59 1607 93
rect 657 59 691 93
rect 309 59 343 93
rect 573 59 607 93
rect 121 59 155 93
rect 1741 59 1775 93
rect 1285 59 1319 93
rect 1009 59 1043 93
rect 1825 59 1859 93
rect 1369 59 1403 93
<< pdiffc >>
rect 1285 451 1319 485
rect 121 451 155 485
rect 309 451 343 485
rect 573 451 607 485
rect 821 451 855 485
rect 1469 451 1503 485
rect 1573 451 1607 485
rect 1741 451 1775 485
rect 1825 451 1859 485
rect 905 443 939 477
rect 1105 443 1139 477
rect 1009 443 1043 477
rect 205 443 239 477
rect 393 443 427 477
rect 489 443 523 477
rect 737 443 771 477
rect 37 443 71 477
rect 1657 443 1691 477
rect 1189 443 1223 477
rect 1573 383 1607 417
rect 309 383 343 417
rect 37 375 71 409
<< poly >>
rect 617 497 647 523
rect 353 497 383 523
rect 1233 497 1263 523
rect 1701 497 1731 523
rect 81 497 111 523
rect 533 497 563 523
rect 1149 497 1179 523
rect 165 497 195 523
rect 1413 497 1443 523
rect 1053 497 1083 523
rect 1329 497 1359 523
rect 865 497 895 523
rect 1617 497 1647 523
rect 1785 497 1815 523
rect 781 497 811 523
rect 437 497 467 523
rect 81 177 111 199
rect 57 199 111 215
rect 57 215 67 249
rect 101 215 111 249
rect 57 249 111 265
rect 81 265 111 297
rect 865 177 895 199
rect 853 199 907 215
rect 853 215 863 249
rect 897 215 907 249
rect 853 249 907 265
rect 865 265 895 297
rect 1617 177 1647 199
rect 1509 199 1647 215
rect 1509 215 1519 249
rect 1553 215 1647 249
rect 1509 249 1647 265
rect 1617 265 1647 297
rect 781 177 811 199
rect 757 199 811 215
rect 757 215 767 249
rect 801 215 811 249
rect 757 249 811 265
rect 781 265 811 297
rect 617 177 647 199
rect 617 199 671 215
rect 617 215 627 249
rect 661 215 671 249
rect 617 249 671 265
rect 617 265 647 297
rect 533 177 563 199
rect 521 199 575 215
rect 521 215 531 249
rect 565 215 575 249
rect 521 249 575 265
rect 533 265 563 297
rect 437 177 467 199
rect 425 199 479 215
rect 425 215 435 249
rect 469 215 479 249
rect 425 249 479 265
rect 437 265 467 297
rect 353 177 383 199
rect 313 199 383 215
rect 313 215 323 249
rect 357 215 383 249
rect 313 249 383 265
rect 353 265 383 297
rect 1413 177 1443 199
rect 1413 199 1467 215
rect 1413 215 1423 249
rect 1457 215 1467 249
rect 1413 249 1467 265
rect 1413 265 1443 297
rect 1233 177 1263 199
rect 1221 199 1275 215
rect 1221 215 1231 249
rect 1265 215 1275 249
rect 1221 249 1275 265
rect 1233 265 1263 297
rect 1149 177 1179 199
rect 1125 199 1179 215
rect 1125 215 1135 249
rect 1169 215 1179 249
rect 1125 249 1179 265
rect 1149 265 1179 297
rect 1053 177 1083 199
rect 949 199 1083 215
rect 949 215 959 249
rect 993 215 1083 249
rect 949 249 1083 265
rect 1053 265 1083 297
rect 1785 177 1815 199
rect 1785 199 1839 215
rect 1785 215 1795 249
rect 1829 215 1839 249
rect 1785 249 1839 265
rect 1785 265 1815 297
rect 1701 177 1731 199
rect 1689 199 1743 215
rect 1689 215 1699 249
rect 1733 215 1743 249
rect 1689 249 1743 265
rect 1701 265 1731 297
rect 165 177 195 199
rect 153 199 207 215
rect 153 215 163 249
rect 197 215 207 249
rect 153 249 207 265
rect 165 265 195 297
rect 1329 177 1359 199
rect 1317 199 1371 215
rect 1317 215 1327 249
rect 1361 215 1371 249
rect 1317 249 1371 265
rect 1329 265 1359 297
rect 81 21 111 47
rect 865 21 895 47
rect 781 21 811 47
rect 617 21 647 47
rect 533 21 563 47
rect 437 21 467 47
rect 353 21 383 47
rect 1413 21 1443 47
rect 1329 21 1359 47
rect 1233 21 1263 47
rect 1149 21 1179 47
rect 1053 21 1083 47
rect 1785 21 1815 47
rect 1701 21 1731 47
rect 1617 21 1647 47
rect 165 21 195 47
<< polycont >>
rect 627 215 661 249
rect 1231 215 1265 249
rect 67 215 101 249
rect 1423 215 1457 249
rect 163 215 197 249
rect 1519 215 1553 249
rect 1795 215 1829 249
rect 863 215 897 249
rect 1135 215 1169 249
rect 959 215 993 249
rect 767 215 801 249
rect 531 215 565 249
rect 1327 215 1361 249
rect 435 215 469 249
rect 1699 215 1733 249
rect 323 215 357 249
<< locali >>
rect 121 485 155 527
rect 63 527 121 561
rect 155 527 213 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 37 477 71 493
rect 1093 101 1127 127
rect 1029 127 1127 161
rect 1029 161 1063 215
rect 801 215 803 249
rect 1029 215 1063 249
rect 767 249 803 265
rect 1029 249 1063 265
rect 769 265 803 299
rect 1029 265 1063 299
rect 769 299 1063 333
rect 1029 333 1063 357
rect 1029 357 1111 391
rect 1077 391 1111 427
rect 1077 427 1223 443
rect 1077 443 1105 477
rect 1139 443 1189 477
rect 1105 477 1223 493
rect 393 427 523 443
rect 427 443 489 477
rect 393 477 523 493
rect 905 477 939 493
rect 1657 477 1691 493
rect 737 477 771 493
rect 523 127 991 161
rect 697 161 731 199
rect 957 161 991 199
rect 697 199 731 215
rect 957 199 993 215
rect 697 215 731 249
rect 957 215 959 249
rect 697 249 731 265
rect 959 249 993 265
rect 697 265 731 299
rect 669 299 731 333
rect 669 333 703 451
rect 607 451 703 485
rect 1223 127 1535 161
rect 1501 161 1535 199
rect 1501 199 1553 215
rect 1501 215 1519 249
rect 1501 249 1553 265
rect 1501 265 1535 357
rect 1393 357 1535 391
rect 1393 391 1427 451
rect 1319 451 1427 485
rect 1859 59 1903 93
rect 1869 93 1903 451
rect 1859 451 1903 485
rect 1809 451 1825 485
rect 1269 451 1285 485
rect 557 451 573 485
rect 189 443 205 477
rect 239 67 267 101
rect 233 101 267 215
rect 233 215 267 249
rect 419 215 435 249
rect 233 249 267 299
rect 421 249 455 299
rect 233 299 455 333
rect 233 333 267 357
rect 421 333 455 357
rect 233 357 267 391
rect 421 357 581 391
rect 233 391 267 443
rect 239 443 267 477
rect 1741 435 1775 451
rect 121 435 155 451
rect 309 417 343 451
rect 1009 427 1043 443
rect 737 375 939 409
rect 737 409 771 443
rect 905 409 939 443
rect 37 409 71 443
rect 1327 199 1361 215
rect 1169 215 1179 249
rect 1317 215 1327 249
rect 1135 249 1179 265
rect 1317 249 1361 265
rect 1145 265 1179 357
rect 1317 265 1351 357
rect 1145 357 1317 391
rect 1573 367 1607 383
rect 309 367 343 383
rect 37 101 71 143
rect 37 143 195 177
rect 161 177 195 199
rect 161 199 197 215
rect 161 215 163 249
rect 161 249 197 265
rect 161 265 195 289
rect 155 289 195 323
rect 161 323 195 359
rect 37 359 71 367
rect 161 359 195 367
rect 37 367 195 375
rect 71 375 195 401
rect 531 199 565 215
rect 529 215 531 249
rect 529 249 565 265
rect 529 265 563 289
rect 523 289 563 323
rect 1423 199 1457 215
rect 1409 215 1423 249
rect 1409 249 1457 265
rect 1409 265 1443 289
rect 1231 199 1265 215
rect 1225 215 1231 249
rect 1225 249 1265 265
rect 1225 265 1259 289
rect 1607 59 1707 93
rect 1673 93 1707 143
rect 1673 143 1819 177
rect 1785 177 1819 199
rect 1785 199 1829 215
rect 1785 215 1795 249
rect 1785 249 1829 265
rect 1785 265 1819 289
rect 1811 289 1819 323
rect 1785 323 1819 357
rect 1657 357 1819 391
rect 1657 391 1691 443
rect 29 215 67 249
rect 29 249 63 323
rect 891 249 897 255
rect 863 255 897 265
rect 305 215 323 249
rect 305 249 339 255
rect 1593 153 1627 215
rect 1593 215 1699 221
rect 1593 221 1685 249
rect 469 215 485 249
rect 101 215 117 249
rect 1733 215 1749 249
rect 357 215 373 249
rect 1135 199 1169 215
rect 767 199 801 215
rect 863 199 897 215
rect 309 161 343 177
rect 1173 127 1189 161
rect 473 127 489 161
rect 309 93 343 127
rect 1741 93 1775 109
rect 121 93 155 109
rect 189 67 205 101
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 1403 59 1419 93
rect 691 59 707 93
rect 557 59 573 93
rect 1809 59 1825 93
rect 1557 59 1573 93
rect 1319 59 1369 93
rect 1269 59 1285 93
rect 607 59 657 93
rect 37 51 71 67
rect 1093 51 1127 67
rect 0 527 29 561
rect 309 485 343 527
rect 339 527 397 561
rect 247 527 305 561
rect 805 451 821 485
rect 855 451 871 485
rect 805 485 871 527
rect 799 527 857 561
rect 707 527 765 561
rect 615 527 673 561
rect 523 527 581 561
rect 431 527 489 561
rect 1009 477 1043 527
rect 983 527 1041 561
rect 891 527 949 561
rect 1573 417 1607 435
rect 1469 435 1607 451
rect 1503 451 1573 485
rect 1469 485 1607 527
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1351 527 1409 561
rect 1259 527 1317 561
rect 1167 527 1225 561
rect 1075 527 1133 561
rect 1741 485 1775 527
rect 1719 527 1777 561
rect 1627 527 1685 561
rect 627 199 661 215
rect 601 215 627 249
rect 601 249 661 265
rect 601 265 635 357
rect 615 357 635 391
rect 1719 -17 1777 17
rect 1741 17 1775 59
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1453 17 1519 59
rect 1453 59 1469 93
rect 1503 59 1519 93
rect 1351 -17 1409 17
rect 1259 -17 1317 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 889 17 1059 59
rect 889 59 905 93
rect 939 59 1009 93
rect 1043 59 1059 93
rect 799 -17 857 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 339 -17 397 17
rect 309 17 343 59
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 121 17 155 59
rect 0 -17 29 17
<< viali >>
rect 1869 527 1903 561
rect 581 527 615 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 857 527 891 561
rect 1225 527 1259 561
rect 673 527 707 561
rect 1777 527 1811 561
rect 121 527 155 561
rect 305 527 339 561
rect 949 527 983 561
rect 397 527 431 561
rect 29 527 63 561
rect 765 527 799 561
rect 213 527 247 561
rect 1317 527 1351 561
rect 489 527 523 561
rect 1133 527 1167 561
rect 1685 527 1719 561
rect 1593 527 1627 561
rect 1041 527 1075 561
rect 1317 357 1351 391
rect 581 357 615 391
rect 1225 289 1259 323
rect 1777 289 1811 323
rect 121 289 155 323
rect 1409 289 1443 323
rect 489 289 523 323
rect 857 221 891 255
rect 1685 221 1719 255
rect 1317 -17 1351 17
rect 1685 -17 1719 17
rect 857 -17 891 17
rect 489 -17 523 17
rect 305 -17 339 17
rect 1133 -17 1167 17
rect 949 -17 983 17
rect 29 -17 63 17
rect 765 -17 799 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 397 -17 431 17
rect 1225 -17 1259 17
rect 1041 -17 1075 17
rect 673 -17 707 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 581 -17 615 17
rect 1593 -17 1627 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 496 1932 527
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 561 1932 592
rect 569 351 627 357
rect 1305 351 1363 357
rect 569 357 581 360
rect 615 357 627 360
rect 1305 357 1317 360
rect 1351 357 1363 360
rect 569 360 581 388
rect 615 360 1317 388
rect 1351 360 1363 388
rect 569 388 581 391
rect 615 388 627 391
rect 1305 388 1317 391
rect 1351 388 1363 391
rect 569 391 627 397
rect 1305 391 1363 397
rect 109 283 167 289
rect 477 283 535 289
rect 1213 283 1271 289
rect 109 289 121 292
rect 155 289 167 292
rect 477 289 489 292
rect 523 289 535 292
rect 1213 289 1225 292
rect 1259 289 1271 292
rect 109 292 121 320
rect 155 292 489 320
rect 523 292 1225 320
rect 1259 292 1271 320
rect 109 320 121 323
rect 155 320 167 323
rect 477 320 489 323
rect 523 320 535 323
rect 1213 320 1225 323
rect 1259 320 1271 323
rect 109 323 167 329
rect 477 323 535 329
rect 1213 323 1271 329
rect 1397 283 1455 289
rect 1765 283 1823 289
rect 1397 289 1409 292
rect 1443 289 1455 292
rect 1765 289 1777 292
rect 1811 289 1823 292
rect 1397 292 1409 320
rect 1443 292 1777 320
rect 1811 292 1823 320
rect 1397 320 1409 323
rect 1443 320 1455 323
rect 1765 320 1777 323
rect 1811 320 1823 323
rect 1397 323 1455 329
rect 1765 323 1823 329
rect 845 215 903 221
rect 1673 215 1731 221
rect 845 221 857 224
rect 891 221 903 224
rect 1673 221 1685 224
rect 1719 221 1731 224
rect 845 224 857 252
rect 891 224 1685 252
rect 1719 224 1731 252
rect 845 252 857 255
rect 891 252 903 255
rect 1673 252 1685 255
rect 1719 252 1731 255
rect 845 255 903 261
rect 1673 255 1731 261
rect 0 -48 1932 -17
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 17 1932 48
<< labels >>
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 CLK
port 5 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 CLK
port 5 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 D
port 6 nsew signal input
flabel locali s 1593 153 1627 187 0 FreeSans 200 0 0 0 RESET_B
port 7 nsew signal input
flabel locali s 1869 85 1903 119 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1869 153 1903 187 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1869 221 1903 255 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1869 289 1903 323 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1869 357 1903 391 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1869 425 1903 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 1 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 2 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 -48 1932 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 1 VPWR
port 4 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 dfrtp_1
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ht_sc_tt05.gds
string GDS_START 24132
string GDS_END 38260
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
