VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ht_sc_tt05__mux2i_2
  CLASS CORE ;
  FOREIGN sky130_ht_sc_tt05__mux2i_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.060 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 5.060 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 5.055 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 5.250 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 5.060 2.960 ;
    END
  END VPWR
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.014 ;
    PORT
      LAYER li1 ;
        RECT 2.445 1.075 3.535 1.275 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.170 ;
    ANTENNAGATEAREA 0.852 ;
    PORT
      LAYER li1 ;
        RECT 4.255 0.995 4.425 1.105 ;
        RECT 4.255 1.105 4.475 1.325 ;
        RECT 4.285 1.325 4.475 1.615 ;
    END
  END A1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.308 ;
    PORT
      LAYER li1 ;
        RECT 0.595 0.765 0.785 0.995 ;
        RECT 0.445 0.995 0.785 1.275 ;
        RECT 0.445 1.275 0.615 1.325 ;
    END
  END S
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.170 ;
    PORT
      LAYER li1 ;
        RECT 2.715 0.295 4.965 0.465 ;
        RECT 4.795 0.465 4.965 1.785 ;
        RECT 4.735 1.785 4.965 2.255 ;
        RECT 2.715 2.255 4.965 2.425 ;
    END
  END Y
  OBS
      LAYER li1 ;
        RECT 2.275 2.175 2.445 2.255 ;
        RECT 0.515 2.255 0.845 2.635 ;
        RECT 1.355 2.255 1.685 2.635 ;
        RECT 2.275 2.255 2.445 2.635 ;
        RECT 0.000 2.635 5.060 2.805 ;
        RECT 1.855 1.835 2.965 1.915 ;
        RECT 1.855 1.915 4.355 2.005 ;
        RECT 1.855 2.005 2.025 2.085 ;
        RECT 2.795 2.005 4.355 2.085 ;
        RECT 1.855 2.085 2.025 2.465 ;
        RECT 0.095 0.255 0.345 0.585 ;
        RECT 0.095 0.585 0.265 1.075 ;
        RECT 0.095 1.075 0.265 1.155 ;
        RECT 1.435 1.075 1.955 1.155 ;
        RECT 0.095 1.155 0.265 1.245 ;
        RECT 1.015 1.155 1.955 1.245 ;
        RECT 0.095 1.245 0.265 1.325 ;
        RECT 1.015 1.245 1.605 1.325 ;
        RECT 0.095 1.325 0.265 1.495 ;
        RECT 1.015 1.325 1.185 1.495 ;
        RECT 0.095 1.495 1.185 1.665 ;
        RECT 0.095 1.665 0.265 2.135 ;
        RECT 0.095 2.135 0.345 2.465 ;
        RECT 1.435 1.495 3.465 1.665 ;
        RECT 1.435 1.665 1.605 1.745 ;
        RECT 3.135 1.665 3.465 1.745 ;
        RECT 1.435 1.745 1.605 1.835 ;
        RECT 0.935 1.835 1.605 2.005 ;
        RECT 1.015 0.555 1.245 0.965 ;
        RECT 3.815 0.635 4.355 0.805 ;
        RECT 3.815 0.805 4.005 0.935 ;
        RECT 1.855 0.255 2.025 0.635 ;
        RECT 1.855 0.635 2.025 0.715 ;
        RECT 3.135 0.635 3.465 0.715 ;
        RECT 1.855 0.715 3.465 0.885 ;
        RECT 0.000 -0.085 5.060 0.085 ;
        RECT 0.595 0.085 0.765 0.545 ;
        RECT 1.435 0.085 1.605 0.545 ;
        RECT 2.275 0.085 2.445 0.545 ;
        RECT 1.435 0.545 1.605 0.885 ;
      LAYER mcon ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 3.825 0.765 3.995 0.935 ;
        RECT 1.065 0.765 1.235 0.935 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
      LAYER met1 ;
        RECT 1.005 0.735 1.295 0.780 ;
        RECT 3.765 0.735 4.055 0.780 ;
        RECT 1.005 0.780 4.055 0.920 ;
        RECT 1.005 0.920 1.295 0.965 ;
        RECT 3.765 0.920 4.055 0.965 ;
  END
END sky130_ht_sc_tt05__mux2i_2
MACRO sky130_ht_sc_tt05__maj3_2
  CLASS CORE ;
  FOREIGN sky130_ht_sc_tt05__maj3_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.140 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.140 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 4.135 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 4.330 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.140 2.960 ;
    END
  END VPWR
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.842 ;
    PORT
      LAYER li1 ;
        RECT 1.055 0.995 1.225 1.105 ;
        RECT 1.055 1.105 1.695 1.275 ;
        RECT 1.055 1.275 1.225 1.325 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.842 ;
    PORT
      LAYER li1 ;
        RECT 1.895 0.995 2.065 1.105 ;
        RECT 1.895 1.105 2.155 1.275 ;
        RECT 1.895 1.275 2.065 1.325 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.850 ;
    ANTENNAGATEAREA 0.416 ;
    PORT
      LAYER li1 ;
        RECT 0.435 0.995 0.745 1.105 ;
        RECT 2.535 0.995 2.705 1.105 ;
        RECT 0.435 1.105 0.775 1.325 ;
        RECT 2.445 1.105 2.705 1.325 ;
        RECT 0.605 1.325 0.775 1.575 ;
        RECT 2.445 1.325 2.615 1.575 ;
        RECT 0.605 1.575 2.615 1.745 ;
    END
  END C
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.502 ;
    PORT
      LAYER li1 ;
        RECT 3.285 0.295 3.615 0.805 ;
        RECT 3.445 0.805 3.615 1.575 ;
        RECT 3.285 1.575 3.615 2.425 ;
    END
  END X
  OBS
      LAYER li1 ;
        RECT 3.785 1.495 3.955 1.915 ;
        RECT 2.705 1.915 3.035 2.255 ;
        RECT 3.785 1.915 3.955 2.255 ;
        RECT 0.985 2.255 1.315 2.635 ;
        RECT 2.705 2.255 3.035 2.635 ;
        RECT 3.785 2.255 3.955 2.635 ;
        RECT 0.000 2.635 4.140 2.805 ;
        RECT 0.085 0.295 0.435 0.635 ;
        RECT 1.825 0.295 2.155 0.635 ;
        RECT 0.085 0.635 3.115 0.805 ;
        RECT 0.085 0.805 0.255 0.995 ;
        RECT 2.945 0.805 3.115 0.995 ;
        RECT 0.085 0.995 0.255 1.245 ;
        RECT 2.945 0.995 3.225 1.245 ;
        RECT 0.085 1.245 0.255 1.325 ;
        RECT 3.055 1.245 3.225 1.325 ;
        RECT 0.085 1.325 0.255 1.915 ;
        RECT 0.085 1.915 2.155 2.085 ;
        RECT 0.085 2.085 0.435 2.425 ;
        RECT 1.825 2.085 2.155 2.425 ;
        RECT 0.000 -0.085 4.140 0.085 ;
        RECT 0.985 0.085 1.315 0.465 ;
        RECT 2.705 0.085 3.035 0.465 ;
        RECT 3.785 0.085 3.955 0.465 ;
        RECT 3.785 0.465 3.955 0.885 ;
      LAYER mcon ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
      LAYER met1 ;
  END
END sky130_ht_sc_tt05__maj3_2
MACRO sky130_ht_sc_tt05__dlrtp_1
  CLASS CORE ;
  FOREIGN sky130_ht_sc_tt05__dlrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.900 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.900 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 6.895 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 7.090 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.900 2.960 ;
    END
  END VPWR
  PIN GATE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.090 ;
    ANTENNAGATEAREA 0.476 ;
    PORT
      LAYER li1 ;
        RECT 0.155 0.995 0.325 1.105 ;
        RECT 0.145 1.105 0.325 1.325 ;
        RECT 0.145 1.325 0.315 1.615 ;
    END
  END GATE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.449 ;
    PORT
      LAYER li1 ;
        RECT 1.515 1.075 1.845 1.275 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.059 ;
    ANTENNAGATEAREA 0.416 ;
    PORT
      LAYER li1 ;
        RECT 5.665 0.425 5.835 1.075 ;
        RECT 5.665 1.075 6.005 1.245 ;
        RECT 5.665 1.245 5.835 1.275 ;
    END
  END RESET_B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365 0.295 6.815 0.595 ;
        RECT 6.645 0.595 6.815 1.785 ;
        RECT 6.365 1.785 6.815 2.425 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 2.025 1.835 2.195 2.175 ;
        RECT 2.025 2.175 2.195 2.255 ;
        RECT 4.545 2.175 5.235 2.255 ;
        RECT 6.025 2.175 6.195 2.255 ;
        RECT 0.525 2.255 0.855 2.635 ;
        RECT 2.025 2.255 2.195 2.635 ;
        RECT 4.545 2.255 5.235 2.635 ;
        RECT 6.025 2.255 6.195 2.635 ;
        RECT 0.000 2.635 6.900 2.805 ;
        RECT 1.545 0.255 1.715 0.715 ;
        RECT 1.545 0.715 2.195 0.885 ;
        RECT 2.025 0.885 2.195 0.995 ;
        RECT 2.025 0.995 2.405 1.325 ;
        RECT 2.025 1.325 2.195 1.445 ;
        RECT 1.545 1.445 2.195 1.615 ;
        RECT 1.545 1.615 1.715 2.465 ;
        RECT 1.025 1.755 1.255 2.465 ;
        RECT 0.105 0.635 0.775 0.805 ;
        RECT 0.605 0.805 0.775 0.995 ;
        RECT 0.605 0.995 0.985 1.325 ;
        RECT 0.605 1.325 0.795 1.615 ;
        RECT 0.605 1.615 0.775 1.875 ;
        RECT 0.105 1.875 0.775 2.045 ;
        RECT 0.185 2.045 0.355 2.465 ;
        RECT 3.025 0.295 3.355 0.715 ;
        RECT 3.025 0.715 4.455 0.885 ;
        RECT 4.285 0.885 4.455 1.445 ;
        RECT 4.285 1.445 4.475 1.615 ;
        RECT 4.285 1.615 4.455 1.785 ;
        RECT 4.205 1.785 4.455 1.955 ;
        RECT 4.205 1.955 4.375 2.255 ;
        RECT 3.565 2.255 4.375 2.425 ;
        RECT 5.465 2.255 5.795 2.425 ;
        RECT 4.885 0.295 5.315 0.465 ;
        RECT 4.885 0.465 5.055 0.715 ;
        RECT 4.705 0.715 5.055 0.885 ;
        RECT 4.705 0.885 4.875 0.995 ;
        RECT 4.695 0.995 4.875 1.075 ;
        RECT 6.295 0.995 6.465 1.075 ;
        RECT 4.695 1.075 4.875 1.325 ;
        RECT 6.285 1.075 6.465 1.325 ;
        RECT 4.705 1.325 4.875 1.445 ;
        RECT 6.285 1.325 6.455 1.445 ;
        RECT 4.705 1.445 4.875 1.615 ;
        RECT 5.665 1.445 6.455 1.615 ;
        RECT 4.705 1.615 4.875 1.785 ;
        RECT 5.665 1.615 5.835 1.785 ;
        RECT 4.705 1.785 5.835 1.955 ;
        RECT 2.445 0.425 2.755 0.595 ;
        RECT 2.585 0.595 2.755 1.075 ;
        RECT 2.585 1.075 3.025 1.245 ;
        RECT 3.775 1.075 4.105 1.245 ;
        RECT 2.585 1.245 2.755 1.785 ;
        RECT 3.865 1.245 4.035 1.785 ;
        RECT 2.445 1.785 4.035 1.955 ;
        RECT 5.135 1.075 5.465 1.245 ;
        RECT 5.205 1.245 5.375 1.445 ;
        RECT 5.205 1.445 5.395 1.615 ;
        RECT 3.235 1.075 3.565 1.275 ;
        RECT 3.365 1.275 3.555 1.615 ;
        RECT 1.025 0.255 1.255 0.625 ;
        RECT 0.000 -0.085 6.900 0.085 ;
        RECT 0.525 0.085 0.855 0.465 ;
        RECT 1.945 0.085 2.275 0.465 ;
        RECT 4.545 0.085 4.715 0.465 ;
        RECT 6.025 0.085 6.195 0.465 ;
        RECT 4.545 0.465 4.715 0.545 ;
        RECT 6.025 0.465 6.195 0.545 ;
      LAYER mcon ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 1.065 1.785 1.235 1.955 ;
        RECT 2.445 1.785 2.615 1.955 ;
        RECT 3.365 1.445 3.535 1.615 ;
        RECT 4.285 1.445 4.455 1.615 ;
        RECT 5.205 1.445 5.375 1.615 ;
        RECT 0.605 1.445 0.775 1.615 ;
        RECT 2.445 0.425 2.615 0.595 ;
        RECT 1.065 0.425 1.235 0.595 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 6.585 -0.085 6.755 0.085 ;
      LAYER met1 ;
        RECT 1.005 1.755 1.295 1.800 ;
        RECT 2.385 1.755 2.675 1.800 ;
        RECT 1.005 1.800 2.675 1.940 ;
        RECT 1.005 1.940 1.295 1.985 ;
        RECT 2.385 1.940 2.675 1.985 ;
        RECT 0.545 1.415 0.835 1.460 ;
        RECT 3.305 1.415 3.595 1.460 ;
        RECT 0.545 1.460 3.595 1.600 ;
        RECT 0.545 1.600 0.835 1.645 ;
        RECT 3.305 1.600 3.595 1.645 ;
        RECT 4.225 1.415 4.515 1.460 ;
        RECT 5.145 1.415 5.435 1.460 ;
        RECT 4.225 1.460 5.435 1.600 ;
        RECT 4.225 1.600 4.515 1.645 ;
        RECT 5.145 1.600 5.435 1.645 ;
        RECT 1.005 0.395 1.295 0.440 ;
        RECT 2.385 0.395 2.675 0.440 ;
        RECT 1.005 0.440 2.675 0.580 ;
        RECT 1.005 0.580 1.295 0.625 ;
        RECT 2.385 0.580 2.675 0.625 ;
  END
END sky130_ht_sc_tt05__dlrtp_1
MACRO sky130_ht_sc_tt05__dfrtp_1
  CLASS CORE ;
  FOREIGN sky130_ht_sc_tt05__dfrtp_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.660 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.660 0.240 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.005 0.105 9.655 1.015 ;
        RECT 0.145 -0.085 0.315 0.105 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 1.305 9.850 2.910 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.660 2.960 ;
    END
  END VPWR
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.090 ;
    PORT
      LAYER li1 ;
        RECT 0.145 1.075 0.585 1.245 ;
        RECT 0.145 1.245 0.315 1.615 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.469 ;
    PORT
      LAYER li1 ;
        RECT 1.535 0.995 1.705 1.075 ;
        RECT 1.525 1.075 1.705 1.275 ;
        RECT 1.535 1.275 1.705 1.325 ;
    END
  END D
  PIN RESET_B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.510 ;
    PORT
      LAYER li1 ;
        RECT 8.025 1.075 8.805 1.245 ;
        RECT 8.025 1.245 8.195 1.275 ;
        RECT 8.425 1.245 8.595 1.275 ;
        RECT 8.025 1.275 8.195 1.495 ;
        RECT 7.965 1.495 8.195 1.665 ;
        RECT 7.965 1.665 8.135 1.955 ;
    END
  END RESET_B
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.105 0.295 9.515 0.465 ;
        RECT 9.345 0.465 9.515 0.635 ;
        RECT 9.345 0.635 9.575 0.805 ;
        RECT 9.405 0.805 9.575 1.575 ;
        RECT 9.345 1.575 9.575 1.745 ;
        RECT 9.345 1.745 9.515 2.255 ;
        RECT 9.105 2.255 9.515 2.425 ;
    END
  END Q
  OBS
      LAYER li1 ;
        RECT 1.545 1.835 1.715 2.135 ;
        RECT 1.545 2.135 1.715 2.175 ;
        RECT 5.105 2.135 5.275 2.175 ;
        RECT 0.605 2.175 0.775 2.255 ;
        RECT 1.545 2.175 1.715 2.255 ;
        RECT 5.105 2.175 5.275 2.255 ;
        RECT 7.405 2.175 8.095 2.255 ;
        RECT 8.765 2.175 8.935 2.255 ;
        RECT 0.605 2.255 0.775 2.635 ;
        RECT 1.545 2.255 1.715 2.635 ;
        RECT 4.085 2.255 4.415 2.635 ;
        RECT 5.105 2.255 5.275 2.635 ;
        RECT 7.405 2.255 8.095 2.635 ;
        RECT 8.765 2.255 8.935 2.635 ;
        RECT 0.000 2.635 9.660 2.805 ;
        RECT 7.845 0.295 8.595 0.465 ;
        RECT 8.425 0.465 8.595 0.715 ;
        RECT 8.425 0.715 9.155 0.885 ;
        RECT 8.985 0.885 9.155 0.995 ;
        RECT 8.985 0.995 9.205 1.325 ;
        RECT 8.985 1.325 9.155 1.445 ;
        RECT 8.885 1.445 9.155 1.615 ;
        RECT 8.985 1.615 9.155 1.785 ;
        RECT 8.345 1.785 9.155 1.955 ;
        RECT 8.345 1.955 8.515 2.465 ;
        RECT 0.145 0.255 0.355 0.625 ;
        RECT 0.185 0.625 0.355 0.715 ;
        RECT 0.185 0.715 0.975 0.885 ;
        RECT 0.805 0.885 0.975 0.995 ;
        RECT 0.805 0.995 0.985 1.325 ;
        RECT 0.805 1.325 0.975 1.445 ;
        RECT 0.605 1.445 0.975 1.615 ;
        RECT 0.605 1.615 0.775 1.795 ;
        RECT 0.185 1.795 0.355 1.835 ;
        RECT 0.605 1.795 0.775 1.835 ;
        RECT 0.185 1.835 0.775 2.005 ;
        RECT 0.185 2.005 0.355 2.465 ;
        RECT 2.845 0.295 3.715 0.465 ;
        RECT 3.545 0.465 3.715 0.635 ;
        RECT 3.545 0.635 5.015 0.805 ;
        RECT 3.545 0.805 3.715 0.995 ;
        RECT 4.845 0.805 5.015 0.995 ;
        RECT 3.545 0.995 3.715 1.245 ;
        RECT 4.845 0.995 5.025 1.245 ;
        RECT 3.545 1.245 3.715 1.325 ;
        RECT 4.855 1.245 5.025 1.325 ;
        RECT 3.545 1.325 3.715 1.495 ;
        RECT 3.405 1.495 3.715 1.665 ;
        RECT 3.405 1.665 3.575 2.135 ;
        RECT 2.505 2.135 2.675 2.215 ;
        RECT 3.405 2.135 3.575 2.215 ;
        RECT 2.505 2.215 3.575 2.385 ;
        RECT 2.505 2.385 2.675 2.465 ;
        RECT 3.745 1.875 4.755 2.045 ;
        RECT 3.745 2.045 3.915 2.465 ;
        RECT 4.585 2.045 4.755 2.465 ;
        RECT 5.525 0.255 5.695 0.635 ;
        RECT 5.205 0.635 5.695 0.805 ;
        RECT 5.205 0.805 5.375 0.995 ;
        RECT 3.895 0.995 4.065 1.075 ;
        RECT 5.205 0.995 5.375 1.075 ;
        RECT 3.895 1.075 4.075 1.325 ;
        RECT 5.205 1.075 5.375 1.325 ;
        RECT 3.905 1.325 4.075 1.495 ;
        RECT 5.205 1.325 5.375 1.495 ;
        RECT 3.905 1.495 5.375 1.665 ;
        RECT 5.205 1.665 5.375 1.785 ;
        RECT 5.205 1.785 5.615 1.955 ;
        RECT 5.445 1.955 5.615 2.135 ;
        RECT 5.445 2.135 6.175 2.385 ;
        RECT 5.585 2.385 6.175 2.465 ;
        RECT 0.945 0.335 1.335 0.505 ;
        RECT 1.165 0.505 1.335 1.785 ;
        RECT 1.025 1.785 1.335 1.955 ;
        RECT 1.025 1.955 1.195 2.465 ;
        RECT 1.945 0.295 2.275 0.635 ;
        RECT 1.885 0.635 2.275 0.805 ;
        RECT 1.885 0.805 2.055 1.915 ;
        RECT 1.885 1.915 2.275 2.085 ;
        RECT 1.945 2.085 2.275 2.425 ;
        RECT 5.925 0.295 6.255 0.635 ;
        RECT 5.925 0.635 7.735 0.805 ;
        RECT 7.565 0.805 7.735 0.995 ;
        RECT 7.565 0.995 7.825 1.325 ;
        RECT 7.565 1.325 7.735 1.785 ;
        RECT 7.025 1.785 7.735 1.955 ;
        RECT 7.025 1.955 7.195 2.255 ;
        RECT 6.405 2.255 7.195 2.425 ;
        RECT 5.735 0.995 5.905 1.075 ;
        RECT 6.695 0.995 6.865 1.075 ;
        RECT 5.735 1.075 5.955 1.325 ;
        RECT 6.645 1.075 6.865 1.325 ;
        RECT 5.785 1.325 5.955 1.785 ;
        RECT 6.645 1.325 6.815 1.785 ;
        RECT 5.785 1.785 6.815 1.955 ;
        RECT 2.235 0.995 2.405 1.075 ;
        RECT 3.195 0.995 3.365 1.075 ;
        RECT 2.235 1.075 2.415 1.325 ;
        RECT 3.065 1.075 3.365 1.325 ;
        RECT 2.245 1.325 2.415 1.495 ;
        RECT 3.065 1.325 3.235 1.495 ;
        RECT 2.245 1.495 3.235 1.665 ;
        RECT 2.905 1.665 3.075 1.955 ;
        RECT 6.215 0.995 6.385 1.075 ;
        RECT 6.125 1.075 6.385 1.325 ;
        RECT 6.125 1.325 6.295 1.615 ;
        RECT 7.175 0.995 7.345 1.075 ;
        RECT 7.045 1.075 7.345 1.325 ;
        RECT 7.045 1.325 7.215 1.615 ;
        RECT 2.445 0.425 2.615 0.635 ;
        RECT 2.445 0.635 2.875 0.805 ;
        RECT 2.705 0.805 2.875 0.995 ;
        RECT 2.705 0.995 2.885 1.245 ;
        RECT 2.715 1.245 2.885 1.325 ;
        RECT 4.375 0.995 4.545 1.105 ;
        RECT 4.285 1.105 4.545 1.275 ;
        RECT 4.375 1.275 4.545 1.325 ;
        RECT 0.000 -0.085 9.660 0.085 ;
        RECT 0.605 0.085 0.775 0.465 ;
        RECT 1.545 0.085 1.715 0.465 ;
        RECT 4.505 0.085 5.355 0.465 ;
        RECT 7.325 0.085 7.655 0.465 ;
        RECT 8.765 0.085 8.935 0.465 ;
        RECT 0.605 0.465 0.775 0.545 ;
        RECT 1.545 0.465 1.715 0.545 ;
        RECT 8.765 0.465 8.935 0.545 ;
      LAYER mcon ;
        RECT 9.345 2.635 9.515 2.805 ;
        RECT 3.365 2.635 3.535 2.805 ;
        RECT 0.145 2.635 0.315 2.805 ;
        RECT 5.205 2.635 5.375 2.805 ;
        RECT 7.505 2.635 7.675 2.805 ;
        RECT 1.065 2.635 1.235 2.805 ;
        RECT 6.125 2.635 6.295 2.805 ;
        RECT 8.885 2.635 9.055 2.805 ;
        RECT 7.045 2.635 7.215 2.805 ;
        RECT 4.745 2.635 4.915 2.805 ;
        RECT 2.905 2.635 3.075 2.805 ;
        RECT 1.525 2.635 1.695 2.805 ;
        RECT 4.285 2.635 4.455 2.805 ;
        RECT 1.985 2.635 2.155 2.805 ;
        RECT 7.965 2.635 8.135 2.805 ;
        RECT 5.665 2.635 5.835 2.805 ;
        RECT 6.585 2.635 6.755 2.805 ;
        RECT 2.445 2.635 2.615 2.805 ;
        RECT 8.425 2.635 8.595 2.805 ;
        RECT 0.605 2.635 0.775 2.805 ;
        RECT 3.825 2.635 3.995 2.805 ;
        RECT 2.905 1.785 3.075 1.955 ;
        RECT 6.585 1.785 6.755 1.955 ;
        RECT 1.065 1.785 1.235 1.955 ;
        RECT 8.885 1.445 9.055 1.615 ;
        RECT 7.045 1.445 7.215 1.615 ;
        RECT 6.125 1.445 6.295 1.615 ;
        RECT 0.605 1.445 0.775 1.615 ;
        RECT 4.285 1.105 4.455 1.275 ;
        RECT 8.425 1.105 8.595 1.275 ;
        RECT 2.445 0.425 2.615 0.595 ;
        RECT 0.145 0.425 0.315 0.595 ;
        RECT 6.585 -0.085 6.755 0.085 ;
        RECT 8.425 -0.085 8.595 0.085 ;
        RECT 4.285 -0.085 4.455 0.085 ;
        RECT 2.445 -0.085 2.615 0.085 ;
        RECT 1.985 -0.085 2.155 0.085 ;
        RECT 1.525 -0.085 1.695 0.085 ;
        RECT 0.605 -0.085 0.775 0.085 ;
        RECT 4.745 -0.085 4.915 0.085 ;
        RECT 7.965 -0.085 8.135 0.085 ;
        RECT 0.145 -0.085 0.315 0.085 ;
        RECT 1.065 -0.085 1.235 0.085 ;
        RECT 3.365 -0.085 3.535 0.085 ;
        RECT 6.125 -0.085 6.295 0.085 ;
        RECT 5.205 -0.085 5.375 0.085 ;
        RECT 2.905 -0.085 3.075 0.085 ;
        RECT 7.045 -0.085 7.215 0.085 ;
        RECT 7.505 -0.085 7.675 0.085 ;
        RECT 5.665 -0.085 5.835 0.085 ;
        RECT 3.825 -0.085 3.995 0.085 ;
        RECT 8.885 -0.085 9.055 0.085 ;
        RECT 9.345 -0.085 9.515 0.085 ;
      LAYER met1 ;
        RECT 1.005 1.755 1.295 1.800 ;
        RECT 2.845 1.755 3.135 1.800 ;
        RECT 6.525 1.755 6.815 1.800 ;
        RECT 1.005 1.800 6.815 1.940 ;
        RECT 1.005 1.940 1.295 1.985 ;
        RECT 2.845 1.940 3.135 1.985 ;
        RECT 6.525 1.940 6.815 1.985 ;
        RECT 0.545 1.415 0.835 1.460 ;
        RECT 6.065 1.415 6.355 1.460 ;
        RECT 0.545 1.460 6.355 1.600 ;
        RECT 0.545 1.600 0.835 1.645 ;
        RECT 6.065 1.600 6.355 1.645 ;
        RECT 6.985 1.415 7.275 1.460 ;
        RECT 8.825 1.415 9.115 1.460 ;
        RECT 6.985 1.460 9.115 1.600 ;
        RECT 6.985 1.600 7.275 1.645 ;
        RECT 8.825 1.600 9.115 1.645 ;
        RECT 4.225 1.075 4.515 1.120 ;
        RECT 8.365 1.075 8.655 1.120 ;
        RECT 4.225 1.120 8.655 1.260 ;
        RECT 4.225 1.260 4.515 1.305 ;
        RECT 8.365 1.260 8.655 1.305 ;
        RECT 0.085 0.395 0.375 0.440 ;
        RECT 2.385 0.395 2.675 0.440 ;
        RECT 0.085 0.440 2.675 0.580 ;
        RECT 0.085 0.580 0.375 0.625 ;
        RECT 2.385 0.580 2.675 0.625 ;
  END
END sky130_ht_sc_tt05__dfrtp_1
