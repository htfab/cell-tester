magic
tech sky130A
magscale 1 2
timestamp 1699069691
<< nwell >>
rect 514 21477 30950 21798
rect 514 20389 30950 20955
rect 514 19301 30950 19867
rect 514 18213 30950 18779
rect 514 17125 30950 17691
rect 514 16037 30950 16603
rect 514 14949 30950 15515
rect 514 13861 30950 14427
rect 514 12773 30950 13339
rect 514 11685 30950 12251
rect 514 10597 30950 11163
rect 514 9509 30950 10075
rect 514 8421 30950 8987
rect 514 7333 30950 7899
rect 514 6245 30950 6811
rect 514 5157 30950 5723
rect 514 4069 30950 4635
rect 514 2981 30950 3547
rect 514 1893 30950 2459
rect 514 805 30950 1371
<< obsli1 >>
rect 552 527 30912 21777
<< obsm1 >>
rect 552 8 31450 22296
<< obsm2 >>
rect 848 2 31446 22302
<< obsm3 >>
rect 1025 35 31451 22269
<< metal4 >>
rect 4294 22104 4354 22304
rect 4846 22104 4906 22304
rect 5398 22104 5458 22304
rect 5950 22104 6010 22304
rect 6502 22104 6562 22304
rect 7054 22104 7114 22304
rect 7606 22104 7666 22304
rect 8158 22104 8218 22304
rect 8710 22104 8770 22304
rect 9262 22104 9322 22304
rect 9814 22104 9874 22304
rect 10366 22104 10426 22304
rect 10918 22104 10978 22304
rect 11470 22104 11530 22304
rect 12022 22104 12082 22304
rect 12574 22104 12634 22304
rect 13126 22104 13186 22304
rect 13678 22104 13738 22304
rect 14230 22104 14290 22304
rect 14782 22104 14842 22304
rect 15334 22104 15394 22304
rect 15886 22104 15946 22304
rect 16438 22104 16498 22304
rect 16990 22104 17050 22304
rect 17542 22104 17602 22304
rect 18094 22104 18154 22304
rect 18646 22104 18706 22304
rect 19198 22104 19258 22304
rect 19750 22104 19810 22304
rect 20302 22104 20362 22304
rect 20854 22104 20914 22304
rect 21406 22104 21466 22304
rect 21958 22104 22018 22304
rect 22510 22104 22570 22304
rect 23062 22104 23122 22304
rect 23614 22104 23674 22304
rect 24166 22104 24226 22304
rect 24718 22104 24778 22304
rect 25270 22104 25330 22304
rect 25822 22104 25882 22304
rect 26374 22104 26434 22304
rect 26926 22104 26986 22304
rect 27478 22104 27538 22304
rect 4187 496 4507 21808
rect 7982 496 8302 21808
rect 11777 496 12097 21808
rect 15572 496 15892 21808
rect 19367 496 19687 21808
rect 23162 496 23482 21808
rect 26957 496 27277 21808
rect 30752 496 31072 21808
<< obsm4 >>
rect 2083 22024 4214 22269
rect 4434 22024 4766 22269
rect 4986 22024 5318 22269
rect 5538 22024 5870 22269
rect 6090 22024 6422 22269
rect 6642 22024 6974 22269
rect 7194 22024 7526 22269
rect 7746 22024 8078 22269
rect 8298 22024 8630 22269
rect 8850 22024 9182 22269
rect 9402 22024 9734 22269
rect 9954 22024 10286 22269
rect 10506 22024 10838 22269
rect 11058 22024 11390 22269
rect 11610 22024 11942 22269
rect 12162 22024 12494 22269
rect 12714 22024 13046 22269
rect 13266 22024 13598 22269
rect 13818 22024 14150 22269
rect 14370 22024 14702 22269
rect 14922 22024 15254 22269
rect 15474 22024 15806 22269
rect 16026 22024 16358 22269
rect 16578 22024 16910 22269
rect 17130 22024 17462 22269
rect 17682 22024 18014 22269
rect 18234 22024 18566 22269
rect 18786 22024 19118 22269
rect 19338 22024 19670 22269
rect 19890 22024 20222 22269
rect 20442 22024 20774 22269
rect 20994 22024 21326 22269
rect 21546 22024 21878 22269
rect 22098 22024 22430 22269
rect 22650 22024 22982 22269
rect 23202 22024 23534 22269
rect 23754 22024 24086 22269
rect 24306 22024 24638 22269
rect 24858 22024 25190 22269
rect 25410 22024 25742 22269
rect 25962 22024 26294 22269
rect 26514 22024 26846 22269
rect 27066 22024 27398 22269
rect 27618 22024 27725 22269
rect 2083 21888 27725 22024
rect 2083 2075 4107 21888
rect 4587 2075 7902 21888
rect 8382 2075 11697 21888
rect 12177 2075 15492 21888
rect 15972 2075 19287 21888
rect 19767 2075 23082 21888
rect 23562 2075 26877 21888
rect 27357 2075 27725 21888
<< labels >>
rlabel metal4 s 7982 496 8302 21808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 15572 496 15892 21808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 23162 496 23482 21808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 30752 496 31072 21808 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4187 496 4507 21808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 11777 496 12097 21808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 19367 496 19687 21808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 26957 496 27277 21808 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 26926 22104 26986 22304 6 clk
port 3 nsew signal input
rlabel metal4 s 27478 22104 27538 22304 6 ena
port 4 nsew signal input
rlabel metal4 s 26374 22104 26434 22304 6 rst_n
port 5 nsew signal input
rlabel metal4 s 25822 22104 25882 22304 6 ui_in[0]
port 6 nsew signal input
rlabel metal4 s 25270 22104 25330 22304 6 ui_in[1]
port 7 nsew signal input
rlabel metal4 s 24718 22104 24778 22304 6 ui_in[2]
port 8 nsew signal input
rlabel metal4 s 24166 22104 24226 22304 6 ui_in[3]
port 9 nsew signal input
rlabel metal4 s 23614 22104 23674 22304 6 ui_in[4]
port 10 nsew signal input
rlabel metal4 s 23062 22104 23122 22304 6 ui_in[5]
port 11 nsew signal input
rlabel metal4 s 22510 22104 22570 22304 6 ui_in[6]
port 12 nsew signal input
rlabel metal4 s 21958 22104 22018 22304 6 ui_in[7]
port 13 nsew signal input
rlabel metal4 s 21406 22104 21466 22304 6 uio_in[0]
port 14 nsew signal input
rlabel metal4 s 20854 22104 20914 22304 6 uio_in[1]
port 15 nsew signal input
rlabel metal4 s 20302 22104 20362 22304 6 uio_in[2]
port 16 nsew signal input
rlabel metal4 s 19750 22104 19810 22304 6 uio_in[3]
port 17 nsew signal input
rlabel metal4 s 19198 22104 19258 22304 6 uio_in[4]
port 18 nsew signal input
rlabel metal4 s 18646 22104 18706 22304 6 uio_in[5]
port 19 nsew signal input
rlabel metal4 s 18094 22104 18154 22304 6 uio_in[6]
port 20 nsew signal input
rlabel metal4 s 17542 22104 17602 22304 6 uio_in[7]
port 21 nsew signal input
rlabel metal4 s 8158 22104 8218 22304 6 uio_oe[0]
port 22 nsew signal output
rlabel metal4 s 7606 22104 7666 22304 6 uio_oe[1]
port 23 nsew signal output
rlabel metal4 s 7054 22104 7114 22304 6 uio_oe[2]
port 24 nsew signal output
rlabel metal4 s 6502 22104 6562 22304 6 uio_oe[3]
port 25 nsew signal output
rlabel metal4 s 5950 22104 6010 22304 6 uio_oe[4]
port 26 nsew signal output
rlabel metal4 s 5398 22104 5458 22304 6 uio_oe[5]
port 27 nsew signal output
rlabel metal4 s 4846 22104 4906 22304 6 uio_oe[6]
port 28 nsew signal output
rlabel metal4 s 4294 22104 4354 22304 6 uio_oe[7]
port 29 nsew signal output
rlabel metal4 s 12574 22104 12634 22304 6 uio_out[0]
port 30 nsew signal output
rlabel metal4 s 12022 22104 12082 22304 6 uio_out[1]
port 31 nsew signal output
rlabel metal4 s 11470 22104 11530 22304 6 uio_out[2]
port 32 nsew signal output
rlabel metal4 s 10918 22104 10978 22304 6 uio_out[3]
port 33 nsew signal output
rlabel metal4 s 10366 22104 10426 22304 6 uio_out[4]
port 34 nsew signal output
rlabel metal4 s 9814 22104 9874 22304 6 uio_out[5]
port 35 nsew signal output
rlabel metal4 s 9262 22104 9322 22304 6 uio_out[6]
port 36 nsew signal output
rlabel metal4 s 8710 22104 8770 22304 6 uio_out[7]
port 37 nsew signal output
rlabel metal4 s 16990 22104 17050 22304 6 uo_out[0]
port 38 nsew signal output
rlabel metal4 s 16438 22104 16498 22304 6 uo_out[1]
port 39 nsew signal output
rlabel metal4 s 15886 22104 15946 22304 6 uo_out[2]
port 40 nsew signal output
rlabel metal4 s 15334 22104 15394 22304 6 uo_out[3]
port 41 nsew signal output
rlabel metal4 s 14782 22104 14842 22304 6 uo_out[4]
port 42 nsew signal output
rlabel metal4 s 14230 22104 14290 22304 6 uo_out[5]
port 43 nsew signal output
rlabel metal4 s 13678 22104 13738 22304 6 uo_out[6]
port 44 nsew signal output
rlabel metal4 s 13126 22104 13186 22304 6 uo_out[7]
port 45 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 31464 22304
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2907524
string GDS_FILE /work/runs/wokwi/results/signoff/tt_um_htfab_cell_tester.magic.gds
string GDS_START 252564
<< end >>

