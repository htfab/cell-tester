magic
tech sky130A
magscale 1 2
timestamp 1699029708
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 1 21 1931 203
rect 29 -17 63 21
<< scnmos >>
rect 81 47 111 177
rect 165 47 195 177
rect 353 47 383 177
rect 545 47 575 177
rect 629 47 659 177
rect 793 47 823 177
rect 877 47 907 177
rect 1629 47 1659 177
rect 1713 47 1743 177
rect 1797 47 1827 177
rect 1065 47 1095 177
rect 1161 47 1191 177
rect 1245 47 1275 177
rect 1425 47 1455 177
<< scpmoshvt >>
rect 81 297 111 497
rect 165 297 195 497
rect 353 297 383 497
rect 449 297 479 497
rect 545 297 575 497
rect 793 297 823 497
rect 877 297 907 497
rect 1629 297 1659 497
rect 1713 297 1743 497
rect 1797 297 1827 497
rect 1065 297 1095 497
rect 1245 297 1275 497
rect 1341 297 1371 497
rect 1425 297 1455 497
<< ndiff >>
rect 1577 47 1629 59
rect 1577 59 1585 93
rect 1619 59 1629 93
rect 1577 93 1629 177
rect 1275 47 1425 177
rect 301 47 353 59
rect 301 59 309 93
rect 343 59 353 93
rect 301 93 353 177
rect 29 47 81 67
rect 29 67 37 101
rect 71 67 81 101
rect 29 101 81 177
rect 111 47 165 59
rect 111 59 121 93
rect 155 59 165 93
rect 111 93 165 177
rect 195 47 247 67
rect 195 67 205 101
rect 239 67 247 101
rect 195 101 247 177
rect 383 47 545 59
rect 383 59 405 93
rect 439 59 545 93
rect 383 93 545 127
rect 383 127 405 161
rect 439 127 545 161
rect 383 161 545 177
rect 575 47 629 59
rect 575 59 585 93
rect 619 59 629 93
rect 575 93 629 177
rect 659 47 793 177
rect 823 47 877 177
rect 907 47 959 59
rect 907 59 917 93
rect 951 59 959 93
rect 907 93 959 177
rect 1659 47 1713 177
rect 1743 47 1797 59
rect 1743 59 1753 93
rect 1787 59 1797 93
rect 1743 93 1797 177
rect 1827 47 1879 59
rect 1827 59 1837 93
rect 1871 59 1879 93
rect 1827 93 1879 177
rect 1095 47 1161 67
rect 1095 67 1105 101
rect 1139 67 1161 101
rect 1095 101 1161 177
rect 1191 47 1245 59
rect 1191 59 1201 93
rect 1235 59 1245 93
rect 1191 93 1245 127
rect 1191 127 1201 161
rect 1235 127 1245 161
rect 1191 161 1245 177
rect 1455 47 1523 59
rect 1455 59 1481 93
rect 1515 59 1523 93
rect 1455 93 1523 177
rect 1013 47 1065 59
rect 1013 59 1021 93
rect 1055 59 1065 93
rect 1013 93 1065 177
<< pdiff >>
rect 1371 297 1425 497
rect 1455 297 1523 451
rect 1455 451 1481 485
rect 1515 451 1523 485
rect 1455 485 1523 497
rect 1013 297 1065 443
rect 1013 443 1021 477
rect 1055 443 1065 477
rect 1013 477 1065 497
rect 1577 297 1629 451
rect 1577 451 1585 485
rect 1619 451 1629 485
rect 1577 485 1629 497
rect 301 297 353 383
rect 301 383 309 417
rect 343 383 353 417
rect 301 417 353 451
rect 301 451 309 485
rect 343 451 353 485
rect 301 485 353 497
rect 29 297 81 375
rect 29 375 37 409
rect 71 375 81 409
rect 29 409 81 443
rect 29 443 37 477
rect 71 443 81 477
rect 29 477 81 497
rect 111 297 165 451
rect 111 451 121 485
rect 155 451 165 485
rect 111 485 165 497
rect 195 297 247 443
rect 195 443 205 477
rect 239 443 247 477
rect 195 477 247 497
rect 383 297 449 383
rect 383 383 405 417
rect 439 383 449 417
rect 383 417 449 451
rect 383 451 405 485
rect 439 451 449 485
rect 383 485 449 497
rect 479 297 545 443
rect 479 443 501 477
rect 535 443 545 477
rect 479 477 545 497
rect 823 297 877 451
rect 823 451 833 485
rect 867 451 877 485
rect 823 485 877 497
rect 907 297 959 443
rect 907 443 917 477
rect 951 443 959 477
rect 907 477 959 497
rect 1659 297 1713 443
rect 1659 443 1669 477
rect 1703 443 1713 477
rect 1659 477 1713 497
rect 1743 297 1797 451
rect 1743 451 1753 485
rect 1787 451 1797 485
rect 1743 485 1797 497
rect 1827 297 1879 451
rect 1827 451 1837 485
rect 1871 451 1879 485
rect 1827 485 1879 497
rect 1095 297 1245 443
rect 1095 443 1117 477
rect 1151 443 1201 477
rect 1235 443 1245 477
rect 1095 477 1245 497
rect 1275 297 1341 451
rect 1275 451 1297 485
rect 1331 451 1341 485
rect 1275 485 1341 497
rect 575 297 793 443
rect 575 443 749 477
rect 783 443 793 477
rect 575 477 793 497
<< ndiffc >>
rect 1201 127 1235 161
rect 405 127 439 161
rect 1105 67 1139 101
rect 205 67 239 101
rect 37 67 71 101
rect 309 59 343 93
rect 1837 59 1871 93
rect 585 59 619 93
rect 1201 59 1235 93
rect 1753 59 1787 93
rect 121 59 155 93
rect 1021 59 1055 93
rect 405 59 439 93
rect 1585 59 1619 93
rect 917 59 951 93
rect 1481 59 1515 93
<< pdiffc >>
rect 1297 451 1331 485
rect 121 451 155 485
rect 309 451 343 485
rect 405 451 439 485
rect 833 451 867 485
rect 1481 451 1515 485
rect 1585 451 1619 485
rect 1753 451 1787 485
rect 1837 451 1871 485
rect 1021 443 1055 477
rect 1669 443 1703 477
rect 501 443 535 477
rect 37 443 71 477
rect 205 443 239 477
rect 749 443 783 477
rect 1201 443 1235 477
rect 1117 443 1151 477
rect 917 443 951 477
rect 405 383 439 417
rect 309 383 343 417
rect 37 375 71 409
<< poly >>
rect 1713 497 1743 523
rect 449 497 479 523
rect 1425 497 1455 523
rect 165 497 195 523
rect 793 497 823 523
rect 1245 497 1275 523
rect 1341 497 1371 523
rect 545 497 575 523
rect 877 497 907 523
rect 1629 497 1659 523
rect 81 497 111 523
rect 353 497 383 523
rect 1797 497 1827 523
rect 1065 497 1095 523
rect 165 177 195 199
rect 153 199 207 215
rect 153 215 163 249
rect 197 215 207 249
rect 153 249 207 265
rect 165 265 195 297
rect 1629 177 1659 199
rect 1521 199 1659 215
rect 1521 215 1531 249
rect 1565 215 1659 249
rect 1521 249 1659 265
rect 1629 265 1659 297
rect 81 177 111 199
rect 57 199 111 215
rect 57 215 67 249
rect 101 215 111 249
rect 57 249 111 265
rect 81 265 111 297
rect 877 177 907 199
rect 865 199 919 215
rect 865 215 875 249
rect 909 215 919 249
rect 865 249 919 265
rect 877 265 907 297
rect 793 177 823 199
rect 769 199 823 215
rect 769 215 779 249
rect 813 215 823 249
rect 769 249 823 265
rect 793 265 823 297
rect 545 177 575 199
rect 533 199 587 215
rect 533 215 543 249
rect 577 215 587 249
rect 533 249 587 265
rect 545 265 575 297
rect 437 199 491 215
rect 437 215 447 249
rect 481 215 491 249
rect 437 249 491 265
rect 449 265 479 297
rect 353 177 383 199
rect 297 199 383 215
rect 297 215 307 249
rect 341 215 383 249
rect 297 249 383 265
rect 353 265 383 297
rect 1425 177 1455 199
rect 1425 199 1479 215
rect 1425 215 1435 249
rect 1469 215 1479 249
rect 1425 249 1479 265
rect 1425 265 1455 297
rect 1329 199 1383 215
rect 1329 215 1339 249
rect 1373 215 1383 249
rect 1329 249 1383 265
rect 1341 265 1371 297
rect 1245 177 1275 199
rect 1233 199 1287 215
rect 1233 215 1243 249
rect 1277 215 1287 249
rect 1233 249 1287 265
rect 1245 265 1275 297
rect 1065 177 1095 199
rect 961 199 1095 215
rect 961 215 971 249
rect 1005 215 1095 249
rect 961 249 1095 265
rect 1065 265 1095 297
rect 1797 177 1827 199
rect 1797 199 1851 215
rect 1797 215 1807 249
rect 1841 215 1851 249
rect 1797 249 1851 265
rect 1797 265 1827 297
rect 1713 177 1743 199
rect 1701 199 1755 215
rect 1701 215 1711 249
rect 1745 215 1755 249
rect 1701 249 1755 265
rect 1713 265 1743 297
rect 1161 177 1191 199
rect 1137 199 1191 215
rect 1137 215 1147 249
rect 1181 215 1191 249
rect 1137 249 1191 265
rect 629 177 659 199
rect 629 199 683 215
rect 629 215 639 249
rect 673 215 683 249
rect 629 249 683 265
rect 81 21 111 47
rect 877 21 907 47
rect 793 21 823 47
rect 629 21 659 47
rect 545 21 575 47
rect 353 21 383 47
rect 1425 21 1455 47
rect 1245 21 1275 47
rect 1161 21 1191 47
rect 1065 21 1095 47
rect 1797 21 1827 47
rect 1713 21 1743 47
rect 1629 21 1659 47
rect 165 21 195 47
<< polycont >>
rect 543 215 577 249
rect 307 215 341 249
rect 1243 215 1277 249
rect 1435 215 1469 249
rect 67 215 101 249
rect 1711 215 1745 249
rect 779 215 813 249
rect 1807 215 1841 249
rect 875 215 909 249
rect 971 215 1005 249
rect 639 215 673 249
rect 1339 215 1373 249
rect 447 215 481 249
rect 1531 215 1565 249
rect 1147 215 1181 249
rect 163 215 197 249
<< locali >>
rect 121 485 155 527
rect 63 527 121 561
rect 155 527 213 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 205 477 239 493
rect 619 59 743 93
rect 709 93 743 127
rect 709 127 1003 161
rect 709 161 743 199
rect 969 161 1003 199
rect 709 199 743 215
rect 969 199 1005 215
rect 709 215 743 249
rect 969 215 971 249
rect 709 249 743 265
rect 971 249 1005 265
rect 709 265 743 299
rect 681 299 743 333
rect 681 333 715 427
rect 501 427 535 443
rect 681 427 715 443
rect 535 443 715 477
rect 501 477 535 493
rect 1105 101 1139 127
rect 1041 127 1139 161
rect 1041 161 1075 215
rect 813 215 815 249
rect 1041 215 1075 249
rect 779 249 815 265
rect 1041 249 1075 265
rect 781 265 815 299
rect 1041 265 1075 299
rect 781 299 1075 333
rect 1041 333 1075 357
rect 1041 357 1123 391
rect 1089 391 1123 427
rect 1089 427 1235 443
rect 1089 443 1117 477
rect 1151 443 1201 477
rect 1117 477 1235 493
rect 917 477 951 493
rect 749 477 783 493
rect 37 477 71 493
rect 1669 477 1703 493
rect 1185 59 1201 93
rect 1235 59 1251 93
rect 1185 93 1251 127
rect 1185 127 1201 161
rect 1235 127 1547 161
rect 1513 161 1547 199
rect 1513 199 1565 215
rect 1513 215 1531 249
rect 1513 249 1565 265
rect 1513 265 1547 357
rect 1405 357 1547 391
rect 1405 391 1439 451
rect 1331 451 1439 485
rect 1871 59 1903 93
rect 1869 93 1903 127
rect 1869 127 1915 161
rect 1881 161 1915 315
rect 1869 315 1915 349
rect 1869 349 1903 451
rect 1871 451 1903 485
rect 389 59 405 93
rect 439 59 455 93
rect 389 93 455 127
rect 377 127 405 161
rect 439 127 455 161
rect 377 161 411 383
rect 377 383 405 417
rect 439 383 455 417
rect 389 417 455 451
rect 389 451 405 485
rect 439 451 455 485
rect 1821 451 1837 485
rect 1281 451 1297 485
rect 309 417 343 451
rect 121 435 155 451
rect 1753 435 1787 451
rect 749 375 951 409
rect 749 409 783 443
rect 917 409 951 443
rect 239 67 267 101
rect 233 101 267 357
rect 247 357 267 391
rect 37 409 71 443
rect 1021 427 1055 443
rect 1605 215 1711 221
rect 1605 221 1685 249
rect 1605 249 1639 299
rect 1593 299 1639 333
rect 1593 333 1627 391
rect 639 199 673 215
rect 481 215 483 249
rect 613 215 639 249
rect 447 249 483 265
rect 613 249 673 265
rect 449 265 483 299
rect 613 265 647 299
rect 449 299 647 333
rect 581 333 615 357
rect 1181 215 1191 249
rect 1147 249 1191 265
rect 1157 265 1191 357
rect 1157 357 1317 391
rect 309 367 343 383
rect 1619 59 1719 93
rect 1685 93 1719 143
rect 1685 143 1831 177
rect 1797 177 1831 199
rect 1797 199 1841 215
rect 1797 215 1807 249
rect 1797 249 1841 265
rect 1797 265 1831 289
rect 1811 289 1831 323
rect 1797 323 1831 357
rect 1669 357 1831 391
rect 1669 391 1703 443
rect 29 215 67 249
rect 29 249 63 323
rect 1435 199 1469 215
rect 1409 215 1435 249
rect 1409 249 1469 265
rect 1409 265 1443 289
rect 63 101 71 119
rect 29 119 71 125
rect 37 125 71 143
rect 37 143 195 177
rect 161 177 195 199
rect 161 199 197 215
rect 161 215 163 249
rect 161 249 197 265
rect 161 265 195 289
rect 155 289 195 323
rect 121 323 155 359
rect 37 359 71 367
rect 121 359 155 367
rect 37 367 155 375
rect 71 375 155 401
rect 1243 199 1277 215
rect 1225 215 1243 249
rect 1225 249 1277 265
rect 1225 265 1259 289
rect 891 249 909 255
rect 875 255 909 265
rect 307 199 341 215
rect 305 215 307 249
rect 305 249 341 255
rect 307 255 341 265
rect 489 119 523 127
rect 489 127 575 161
rect 541 161 575 199
rect 541 199 577 215
rect 541 215 543 249
rect 543 249 577 265
rect 1745 215 1761 249
rect 101 215 117 249
rect 779 199 813 215
rect 447 199 481 215
rect 1147 199 1181 215
rect 875 199 909 215
rect 121 93 155 109
rect 309 93 343 109
rect 1753 93 1787 109
rect 189 67 205 101
rect 1569 59 1585 93
rect 1903 -17 1932 17
rect 1821 59 1837 93
rect 569 59 585 93
rect 1105 51 1139 67
rect 0 527 29 561
rect 1481 435 1619 451
rect 1515 451 1585 485
rect 1481 485 1619 527
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1351 527 1409 561
rect 1259 527 1317 561
rect 1167 527 1225 561
rect 1075 527 1133 561
rect 1021 477 1055 527
rect 983 527 1041 561
rect 891 527 949 561
rect 309 485 343 527
rect 339 527 397 561
rect 247 527 305 561
rect 817 451 833 485
rect 867 451 883 485
rect 817 485 883 527
rect 799 527 857 561
rect 707 527 765 561
rect 615 527 673 561
rect 523 527 581 561
rect 431 527 489 561
rect 1753 485 1787 527
rect 1719 527 1777 561
rect 1627 527 1685 561
rect 205 357 213 391
rect 205 391 239 443
rect 1339 199 1373 215
rect 1329 215 1339 249
rect 1329 249 1373 265
rect 1329 265 1363 357
rect 1351 357 1363 391
rect 29 51 71 67
rect 29 67 37 85
rect 1811 -17 1869 17
rect 1719 -17 1777 17
rect 1753 17 1787 59
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1465 17 1531 59
rect 1465 59 1481 93
rect 1515 59 1531 93
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 901 17 1071 59
rect 901 59 917 93
rect 951 59 1021 93
rect 1055 59 1071 93
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 309 17 343 59
rect 247 -17 305 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 121 17 155 59
rect 0 -17 29 17
<< viali >>
rect 1869 527 1903 561
rect 673 527 707 561
rect 29 527 63 561
rect 1041 527 1075 561
rect 1501 527 1535 561
rect 213 527 247 561
rect 1225 527 1259 561
rect 1777 527 1811 561
rect 1409 527 1443 561
rect 949 527 983 561
rect 581 527 615 561
rect 305 527 339 561
rect 857 527 891 561
rect 397 527 431 561
rect 1593 527 1627 561
rect 1133 527 1167 561
rect 1317 527 1351 561
rect 489 527 523 561
rect 1685 527 1719 561
rect 121 527 155 561
rect 765 527 799 561
rect 581 357 615 391
rect 1317 357 1351 391
rect 213 357 247 391
rect 1777 289 1811 323
rect 1409 289 1443 323
rect 1225 289 1259 323
rect 121 289 155 323
rect 857 221 891 255
rect 1685 221 1719 255
rect 489 85 523 119
rect 29 85 63 119
rect 1317 -17 1351 17
rect 1685 -17 1719 17
rect 857 -17 891 17
rect 489 -17 523 17
rect 397 -17 431 17
rect 305 -17 339 17
rect 121 -17 155 17
rect 949 -17 983 17
rect 1593 -17 1627 17
rect 29 -17 63 17
rect 213 -17 247 17
rect 673 -17 707 17
rect 1225 -17 1259 17
rect 1041 -17 1075 17
rect 581 -17 615 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1133 -17 1167 17
rect 765 -17 799 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 496 1932 527
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 561 1932 592
rect 201 351 259 357
rect 569 351 627 357
rect 1305 351 1363 357
rect 201 357 213 360
rect 247 357 259 360
rect 569 357 581 360
rect 615 357 627 360
rect 1305 357 1317 360
rect 1351 357 1363 360
rect 201 360 213 388
rect 247 360 581 388
rect 615 360 1317 388
rect 1351 360 1363 388
rect 201 388 213 391
rect 247 388 259 391
rect 569 388 581 391
rect 615 388 627 391
rect 1305 388 1317 391
rect 1351 388 1363 391
rect 201 391 259 397
rect 569 391 627 397
rect 1305 391 1363 397
rect 109 283 167 289
rect 1213 283 1271 289
rect 109 289 121 292
rect 155 289 167 292
rect 1213 289 1225 292
rect 1259 289 1271 292
rect 109 292 121 320
rect 155 292 1225 320
rect 1259 292 1271 320
rect 109 320 121 323
rect 155 320 167 323
rect 1213 320 1225 323
rect 1259 320 1271 323
rect 109 323 167 329
rect 1213 323 1271 329
rect 1397 283 1455 289
rect 1765 283 1823 289
rect 1397 289 1409 292
rect 1443 289 1455 292
rect 1765 289 1777 292
rect 1811 289 1823 292
rect 1397 292 1409 320
rect 1443 292 1777 320
rect 1811 292 1823 320
rect 1397 320 1409 323
rect 1443 320 1455 323
rect 1765 320 1777 323
rect 1811 320 1823 323
rect 1397 323 1455 329
rect 1765 323 1823 329
rect 845 215 903 221
rect 1673 215 1731 221
rect 845 221 857 224
rect 891 221 903 224
rect 1673 221 1685 224
rect 1719 221 1731 224
rect 845 224 857 252
rect 891 224 1685 252
rect 1719 224 1731 252
rect 845 252 857 255
rect 891 252 903 255
rect 1673 252 1685 255
rect 1719 252 1731 255
rect 845 255 903 261
rect 1673 255 1731 261
rect 17 79 75 85
rect 477 79 535 85
rect 17 85 29 88
rect 63 85 75 88
rect 477 85 489 88
rect 523 85 535 88
rect 17 88 29 116
rect 63 88 489 116
rect 523 88 535 116
rect 17 116 29 119
rect 63 116 75 119
rect 477 116 489 119
rect 523 116 535 119
rect 17 119 75 125
rect 477 119 535 125
rect 0 -48 1932 -17
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 17 1932 48
<< labels >>
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 CLK
port 1 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 1593 357 1627 391 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1869 85 1903 119 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1869 357 1903 391 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1869 425 1903 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 -48 1932 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 1 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 dfrtp_1
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ht_sc_tt05.gds
string GDS_START 23748
string GDS_END 37828
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
