magic
tech sky130A
magscale 1 2
timestamp 1698891296
<< viali >>
rect 2421 21641 2455 21675
rect 6377 21641 6411 21675
rect 6929 21641 6963 21675
rect 9965 21641 9999 21675
rect 12817 21641 12851 21675
rect 19165 21641 19199 21675
rect 21005 21641 21039 21675
rect 5457 21573 5491 21607
rect 8217 21573 8251 21607
rect 10333 21573 10367 21607
rect 13185 21573 13219 21607
rect 18429 21573 18463 21607
rect 25697 21573 25731 21607
rect 30021 21573 30055 21607
rect 3712 21505 3746 21539
rect 7113 21505 7147 21539
rect 8677 21505 8711 21539
rect 11440 21505 11474 21539
rect 16865 21505 16899 21539
rect 17141 21505 17175 21539
rect 19441 21505 19475 21539
rect 19717 21505 19751 21539
rect 21465 21505 21499 21539
rect 21925 21505 21959 21539
rect 22477 21505 22511 21539
rect 23857 21505 23891 21539
rect 24501 21505 24535 21539
rect 24894 21505 24928 21539
rect 25053 21505 25087 21539
rect 949 21437 983 21471
rect 2145 21437 2179 21471
rect 2697 21437 2731 21471
rect 3249 21437 3283 21471
rect 3985 21437 4019 21471
rect 5641 21437 5675 21471
rect 6101 21437 6135 21471
rect 7389 21437 7423 21471
rect 8585 21437 8619 21471
rect 8953 21437 8987 21471
rect 10517 21437 10551 21471
rect 10793 21437 10827 21471
rect 10977 21437 11011 21471
rect 11304 21437 11338 21471
rect 11713 21437 11747 21471
rect 13369 21437 13403 21471
rect 13645 21437 13679 21471
rect 14289 21437 14323 21471
rect 14565 21437 14599 21471
rect 16313 21437 16347 21471
rect 16681 21437 16715 21471
rect 18705 21437 18739 21471
rect 18889 21437 18923 21471
rect 19073 21437 19107 21471
rect 19349 21437 19383 21471
rect 21281 21437 21315 21471
rect 22201 21437 22235 21471
rect 22318 21437 22352 21471
rect 23213 21437 23247 21471
rect 23397 21437 23431 21471
rect 23581 21437 23615 21471
rect 23673 21437 23707 21471
rect 24041 21437 24075 21471
rect 24777 21437 24811 21471
rect 26433 21437 26467 21471
rect 26709 21437 26743 21471
rect 28273 21437 28307 21471
rect 29469 21437 29503 21471
rect 29929 21437 29963 21471
rect 30205 21437 30239 21471
rect 30573 21437 30607 21471
rect 1225 21369 1259 21403
rect 1593 21369 1627 21403
rect 3065 21369 3099 21403
rect 6653 21369 6687 21403
rect 8033 21369 8067 21403
rect 9781 21369 9815 21403
rect 15945 21369 15979 21403
rect 16773 21369 16807 21403
rect 25881 21369 25915 21403
rect 29101 21369 29135 21403
rect 1869 21301 1903 21335
rect 3715 21301 3749 21335
rect 5089 21301 5123 21335
rect 8401 21301 8435 21335
rect 10609 21301 10643 21335
rect 13737 21301 13771 21335
rect 16129 21301 16163 21335
rect 23121 21301 23155 21335
rect 25973 21301 26007 21335
rect 27813 21301 27847 21335
rect 28365 21301 28399 21335
rect 29745 21301 29779 21335
rect 30389 21301 30423 21335
rect 857 21097 891 21131
rect 1599 21097 1633 21131
rect 6291 21097 6325 21131
rect 9873 21097 9907 21131
rect 13001 21097 13035 21131
rect 18797 21097 18831 21131
rect 20821 21097 20855 21131
rect 23121 21097 23155 21131
rect 27813 21097 27847 21131
rect 10425 21029 10459 21063
rect 10793 21029 10827 21063
rect 15669 21029 15703 21063
rect 25308 21029 25342 21063
rect 26157 21029 26191 21063
rect 1041 20961 1075 20995
rect 5457 20961 5491 20995
rect 8033 20961 8067 20995
rect 11897 20961 11931 20995
rect 13461 20961 13495 20995
rect 14381 20961 14415 20995
rect 16129 20961 16163 20995
rect 17969 20961 18003 20995
rect 18337 20961 18371 20995
rect 21005 20961 21039 20995
rect 23305 20961 23339 20995
rect 25513 20961 25547 20995
rect 25789 20961 25823 20995
rect 26433 20961 26467 20995
rect 28600 20961 28634 20995
rect 1133 20893 1167 20927
rect 1639 20893 1673 20927
rect 1869 20893 1903 20927
rect 3341 20893 3375 20927
rect 3668 20893 3702 20927
rect 3804 20893 3838 20927
rect 4077 20893 4111 20927
rect 5825 20893 5859 20927
rect 6288 20893 6322 20927
rect 6561 20893 6595 20927
rect 8360 20893 8394 20927
rect 8512 20911 8546 20945
rect 8769 20893 8803 20927
rect 11161 20893 11195 20927
rect 11488 20893 11522 20927
rect 11624 20895 11658 20929
rect 14105 20893 14139 20927
rect 16405 20893 16439 20927
rect 18705 20893 18739 20927
rect 18981 20893 19015 20927
rect 19257 20893 19291 20927
rect 21281 20893 21315 20927
rect 21557 20893 21591 20927
rect 23489 20893 23523 20927
rect 23765 20893 23799 20927
rect 26709 20893 26743 20927
rect 28273 20893 28307 20927
rect 28779 20893 28813 20927
rect 29009 20893 29043 20927
rect 3157 20757 3191 20791
rect 7849 20757 7883 20791
rect 13553 20757 13587 20791
rect 15945 20757 15979 20791
rect 17509 20757 17543 20791
rect 30113 20757 30147 20791
rect 2789 20553 2823 20587
rect 7941 20553 7975 20587
rect 10425 20553 10459 20587
rect 13001 20553 13035 20587
rect 14105 20553 14139 20587
rect 14546 20553 14580 20587
rect 16037 20553 16071 20587
rect 5917 20485 5951 20519
rect 1455 20417 1489 20451
rect 4399 20417 4433 20451
rect 6428 20417 6462 20451
rect 6607 20417 6641 20451
rect 8907 20417 8941 20451
rect 11105 20417 11139 20451
rect 16129 20417 16163 20451
rect 18245 20417 18279 20451
rect 19257 20417 19291 20451
rect 19533 20417 19567 20451
rect 21278 20417 21312 20451
rect 21833 20417 21867 20451
rect 23857 20417 23891 20451
rect 24133 20417 24167 20451
rect 26709 20417 26743 20451
rect 27215 20417 27249 20451
rect 30297 20417 30331 20451
rect 949 20349 983 20383
rect 1685 20349 1719 20383
rect 3433 20349 3467 20383
rect 3893 20349 3927 20383
rect 4629 20349 4663 20383
rect 6101 20349 6135 20383
rect 6837 20349 6871 20383
rect 8401 20349 8435 20383
rect 9137 20349 9171 20383
rect 10609 20349 10643 20383
rect 11345 20349 11379 20383
rect 12909 20349 12943 20383
rect 14296 20349 14330 20383
rect 16405 20349 16439 20383
rect 21557 20349 21591 20383
rect 23581 20349 23615 20383
rect 25881 20349 25915 20383
rect 27036 20349 27070 20383
rect 27445 20349 27479 20383
rect 29101 20349 29135 20383
rect 29285 20349 29319 20383
rect 29377 20349 29411 20383
rect 30021 20349 30055 20383
rect 30205 20349 30239 20383
rect 13829 20281 13863 20315
rect 17969 20281 18003 20315
rect 18797 20281 18831 20315
rect 26157 20281 26191 20315
rect 1415 20213 1449 20247
rect 3709 20213 3743 20247
rect 4359 20213 4393 20247
rect 8867 20213 8901 20247
rect 11075 20213 11109 20247
rect 12633 20213 12667 20247
rect 17509 20213 17543 20247
rect 18889 20213 18923 20247
rect 21097 20213 21131 20247
rect 23397 20213 23431 20247
rect 25697 20213 25731 20247
rect 26249 20213 26283 20247
rect 28549 20213 28583 20247
rect 29653 20213 29687 20247
rect 30481 20213 30515 20247
rect 1599 20009 1633 20043
rect 3157 20009 3191 20043
rect 7849 20009 7883 20043
rect 12547 20009 12581 20043
rect 13921 20009 13955 20043
rect 16773 20009 16807 20043
rect 24041 20009 24075 20043
rect 27813 20009 27847 20043
rect 30205 20009 30239 20043
rect 1041 19873 1075 19907
rect 1133 19873 1167 19907
rect 5641 19873 5675 19907
rect 8217 19873 8251 19907
rect 12817 19873 12851 19907
rect 16313 19873 16347 19907
rect 16497 19873 16531 19907
rect 17233 19873 17267 19907
rect 18705 19873 18739 19907
rect 20545 19873 20579 19907
rect 21557 19873 21591 19907
rect 21925 19873 21959 19907
rect 22201 19873 22235 19907
rect 24225 19873 24259 19907
rect 24409 19873 24443 19907
rect 26065 19873 26099 19907
rect 26709 19873 26743 19907
rect 1629 19823 1663 19857
rect 1869 19805 1903 19839
rect 3525 19805 3559 19839
rect 3852 19805 3886 19839
rect 4031 19805 4065 19839
rect 4261 19805 4295 19839
rect 5825 19805 5859 19839
rect 6152 19805 6186 19839
rect 6288 19805 6322 19839
rect 6561 19805 6595 19839
rect 8401 19805 8435 19839
rect 8493 19805 8527 19839
rect 8820 19805 8854 19839
rect 8956 19805 8990 19839
rect 9229 19805 9263 19839
rect 10977 19805 11011 19839
rect 11253 19805 11287 19839
rect 12081 19805 12115 19839
rect 12544 19805 12578 19839
rect 14289 19805 14323 19839
rect 14565 19805 14599 19839
rect 16221 19805 16255 19839
rect 16957 19805 16991 19839
rect 18981 19805 19015 19839
rect 22477 19805 22511 19839
rect 24685 19805 24719 19839
rect 26433 19805 26467 19839
rect 28365 19805 28399 19839
rect 28692 19805 28726 19839
rect 28871 19805 28905 19839
rect 29101 19805 29135 19839
rect 10517 19737 10551 19771
rect 21373 19737 21407 19771
rect 857 19669 891 19703
rect 15853 19669 15887 19703
rect 18521 19669 18555 19703
rect 20085 19669 20119 19703
rect 20821 19669 20855 19703
rect 7113 19465 7147 19499
rect 10241 19465 10275 19499
rect 15393 19465 15427 19499
rect 20085 19465 20119 19499
rect 22017 19465 22051 19499
rect 28549 19465 28583 19499
rect 29929 19465 29963 19499
rect 4997 19397 5031 19431
rect 18061 19397 18095 19431
rect 23581 19397 23615 19431
rect 1455 19329 1489 19363
rect 5273 19329 5307 19363
rect 5736 19329 5770 19363
rect 8125 19329 8159 19363
rect 8864 19329 8898 19363
rect 11716 19329 11750 19363
rect 14016 19329 14050 19363
rect 16221 19329 16255 19363
rect 18705 19329 18739 19363
rect 20729 19329 20763 19363
rect 25007 19329 25041 19363
rect 27215 19329 27249 19363
rect 949 19261 983 19295
rect 1685 19261 1719 19295
rect 3065 19261 3099 19295
rect 3525 19261 3559 19295
rect 3617 19261 3651 19295
rect 3893 19261 3927 19295
rect 6009 19261 6043 19295
rect 7665 19261 7699 19295
rect 8401 19261 8435 19295
rect 9137 19261 9171 19295
rect 10701 19261 10735 19295
rect 11253 19261 11287 19295
rect 11989 19261 12023 19295
rect 13553 19261 13587 19295
rect 13880 19261 13914 19295
rect 14289 19261 14323 19295
rect 15945 19261 15979 19295
rect 17601 19261 17635 19295
rect 18245 19261 18279 19295
rect 18521 19261 18555 19295
rect 18981 19261 19015 19295
rect 20453 19261 20487 19295
rect 24501 19261 24535 19295
rect 25237 19261 25271 19295
rect 26709 19261 26743 19295
rect 27445 19261 27479 19295
rect 29469 19261 29503 19295
rect 29837 19261 29871 19295
rect 4261 19193 4295 19227
rect 4813 19193 4847 19227
rect 7849 19193 7883 19227
rect 10977 19193 11011 19227
rect 17785 19193 17819 19227
rect 17969 19193 18003 19227
rect 22477 19193 22511 19227
rect 24041 19193 24075 19227
rect 29101 19193 29135 19227
rect 30205 19193 30239 19227
rect 1415 19125 1449 19159
rect 3341 19125 3375 19159
rect 4353 19125 4387 19159
rect 5739 19125 5773 19159
rect 7481 19125 7515 19159
rect 8867 19125 8901 19159
rect 11719 19125 11753 19159
rect 13093 19125 13127 19159
rect 18337 19125 18371 19159
rect 24133 19125 24167 19159
rect 24967 19125 25001 19159
rect 26341 19125 26375 19159
rect 27175 19125 27209 19159
rect 30297 19125 30331 19159
rect 1783 18921 1817 18955
rect 4997 18921 5031 18955
rect 11529 18921 11563 18955
rect 15853 18921 15887 18955
rect 16773 18921 16807 18955
rect 20269 18921 20303 18955
rect 23397 18921 23431 18955
rect 24599 18921 24633 18955
rect 5641 18853 5675 18887
rect 8033 18853 8067 18887
rect 10793 18853 10827 18887
rect 11253 18853 11287 18887
rect 1225 18785 1259 18819
rect 4077 18785 4111 18819
rect 4361 18789 4395 18823
rect 4629 18785 4663 18819
rect 4905 18785 4939 18819
rect 5181 18785 5215 18819
rect 5457 18785 5491 18819
rect 5917 18785 5951 18819
rect 6653 18785 6687 18819
rect 8217 18785 8251 18819
rect 9004 18785 9038 18819
rect 10977 18785 11011 18819
rect 11713 18785 11747 18819
rect 14197 18785 14231 18819
rect 14289 18785 14323 18819
rect 16313 18785 16347 18819
rect 16497 18785 16531 18819
rect 16957 18785 16991 18819
rect 18613 18785 18647 18819
rect 18981 18785 19015 18819
rect 20545 18785 20579 18819
rect 21557 18785 21591 18819
rect 23489 18785 23523 18819
rect 24041 18785 24075 18819
rect 24869 18785 24903 18819
rect 26617 18785 26651 18819
rect 27128 18785 27162 18819
rect 29009 18785 29043 18819
rect 29285 18785 29319 18819
rect 30113 18785 30147 18819
rect 30573 18785 30607 18819
rect 1317 18717 1351 18751
rect 1823 18717 1857 18751
rect 2053 18717 2087 18751
rect 6244 18717 6278 18751
rect 6380 18719 6414 18753
rect 8677 18717 8711 18751
rect 9140 18735 9174 18769
rect 9413 18717 9447 18751
rect 11805 18717 11839 18751
rect 12132 18717 12166 18751
rect 12311 18717 12345 18751
rect 12541 18717 12575 18751
rect 14565 18717 14599 18751
rect 16589 18717 16623 18751
rect 17233 18717 17267 18751
rect 18705 18717 18739 18751
rect 21281 18717 21315 18751
rect 23673 18717 23707 18751
rect 24133 18717 24167 18751
rect 24596 18717 24630 18751
rect 26801 18717 26835 18751
rect 27307 18717 27341 18751
rect 27537 18717 27571 18751
rect 3893 18649 3927 18683
rect 4445 18649 4479 18683
rect 4721 18649 4755 18683
rect 14013 18649 14047 18683
rect 23029 18649 23063 18683
rect 1041 18581 1075 18615
rect 3341 18581 3375 18615
rect 3709 18581 3743 18615
rect 4169 18581 4203 18615
rect 8493 18581 8527 18615
rect 13829 18581 13863 18615
rect 20637 18581 20671 18615
rect 22661 18581 22695 18615
rect 23857 18581 23891 18615
rect 25973 18581 26007 18615
rect 26433 18581 26467 18615
rect 28641 18581 28675 18615
rect 30297 18581 30331 18615
rect 30389 18581 30423 18615
rect 2789 18377 2823 18411
rect 5089 18377 5123 18411
rect 5549 18377 5583 18411
rect 5825 18377 5859 18411
rect 12541 18377 12575 18411
rect 13093 18377 13127 18411
rect 13829 18377 13863 18411
rect 17969 18377 18003 18411
rect 23397 18377 23431 18411
rect 24593 18377 24627 18411
rect 20269 18309 20303 18343
rect 23029 18309 23063 18343
rect 24225 18309 24259 18343
rect 26617 18309 26651 18343
rect 1455 18241 1489 18275
rect 3249 18241 3283 18275
rect 3712 18241 3746 18275
rect 6564 18241 6598 18275
rect 8956 18241 8990 18275
rect 10609 18241 10643 18275
rect 11164 18241 11198 18275
rect 14887 18241 14921 18275
rect 16865 18241 16899 18275
rect 18981 18241 19015 18275
rect 21051 18241 21085 18275
rect 21281 18241 21315 18275
rect 25283 18241 25317 18275
rect 949 18173 983 18207
rect 1685 18173 1719 18207
rect 3985 18173 4019 18207
rect 5733 18173 5767 18207
rect 6009 18173 6043 18207
rect 6101 18173 6135 18207
rect 6837 18173 6871 18207
rect 8493 18173 8527 18207
rect 8820 18173 8854 18207
rect 9229 18173 9263 18207
rect 10701 18173 10735 18207
rect 11437 18173 11471 18207
rect 14381 18173 14415 18207
rect 15117 18173 15151 18207
rect 16589 18173 16623 18207
rect 18521 18173 18555 18207
rect 18705 18173 18739 18207
rect 20545 18173 20579 18207
rect 20872 18173 20906 18207
rect 22845 18173 22879 18207
rect 23581 18173 23615 18207
rect 23949 18173 23983 18207
rect 24409 18173 24443 18207
rect 24777 18173 24811 18207
rect 25513 18173 25547 18207
rect 27077 18173 27111 18207
rect 29009 18173 29043 18207
rect 29285 18173 29319 18207
rect 30573 18173 30607 18207
rect 8217 18105 8251 18139
rect 13001 18105 13035 18139
rect 13737 18105 13771 18139
rect 27353 18105 27387 18139
rect 1415 18037 1449 18071
rect 3715 18037 3749 18071
rect 6567 18037 6601 18071
rect 11167 18037 11201 18071
rect 14847 18037 14881 18071
rect 16221 18037 16255 18071
rect 18337 18037 18371 18071
rect 22385 18037 22419 18071
rect 25243 18037 25277 18071
rect 28825 18037 28859 18071
rect 29929 18037 29963 18071
rect 30113 18037 30147 18071
rect 30389 18037 30423 18071
rect 5549 17833 5583 17867
rect 6935 17833 6969 17867
rect 8493 17833 8527 17867
rect 10701 17833 10735 17867
rect 11995 17833 12029 17867
rect 17049 17833 17083 17867
rect 25973 17833 26007 17867
rect 26899 17833 26933 17867
rect 28273 17833 28307 17867
rect 3433 17765 3467 17799
rect 30205 17765 30239 17799
rect 1225 17697 1259 17731
rect 5917 17697 5951 17731
rect 7205 17697 7239 17731
rect 9413 17697 9447 17731
rect 11069 17697 11103 17731
rect 12265 17697 12299 17731
rect 14013 17697 14047 17731
rect 14289 17697 14323 17731
rect 16221 17697 16255 17731
rect 16681 17697 16715 17731
rect 17877 17697 17911 17731
rect 19717 17697 19751 17731
rect 21608 17697 21642 17731
rect 23489 17697 23523 17731
rect 24869 17697 24903 17731
rect 28641 17697 28675 17731
rect 28917 17697 28951 17731
rect 1317 17629 1351 17663
rect 1644 17629 1678 17663
rect 1813 17647 1847 17681
rect 2053 17629 2087 17663
rect 3525 17629 3559 17663
rect 3852 17629 3886 17663
rect 4031 17629 4065 17663
rect 4261 17629 4295 17663
rect 6469 17629 6503 17663
rect 6932 17631 6966 17665
rect 8677 17629 8711 17663
rect 9004 17629 9038 17663
rect 9140 17631 9174 17665
rect 11529 17629 11563 17663
rect 12035 17629 12069 17663
rect 14565 17629 14599 17663
rect 15945 17629 15979 17663
rect 16957 17629 16991 17663
rect 17141 17629 17175 17663
rect 17468 17629 17502 17663
rect 17647 17629 17681 17663
rect 19441 17629 19475 17663
rect 21281 17629 21315 17663
rect 21777 17647 21811 17681
rect 22017 17629 22051 17663
rect 24133 17629 24167 17663
rect 24460 17629 24494 17663
rect 24639 17629 24673 17663
rect 26433 17629 26467 17663
rect 26896 17629 26930 17663
rect 27169 17629 27203 17663
rect 30481 17629 30515 17663
rect 23581 17561 23615 17595
rect 1041 17493 1075 17527
rect 6009 17493 6043 17527
rect 11161 17493 11195 17527
rect 13369 17493 13403 17527
rect 18981 17493 19015 17527
rect 20821 17493 20855 17527
rect 23121 17493 23155 17527
rect 2973 17289 3007 17323
rect 8401 17289 8435 17323
rect 10517 17289 10551 17323
rect 11069 17289 11103 17323
rect 16037 17289 16071 17323
rect 30389 17289 30423 17323
rect 13829 17221 13863 17255
rect 20361 17221 20395 17255
rect 23305 17221 23339 17255
rect 1455 17153 1489 17187
rect 4399 17153 4433 17187
rect 4583 17153 4617 17187
rect 6009 17153 6043 17187
rect 6564 17153 6598 17187
rect 6837 17153 6871 17187
rect 8217 17153 8251 17187
rect 9140 17153 9174 17187
rect 11759 17153 11793 17187
rect 14197 17153 14231 17187
rect 14703 17153 14737 17187
rect 16732 17153 16766 17187
rect 16911 17153 16945 17187
rect 21051 17153 21085 17187
rect 21281 17153 21315 17187
rect 25104 17153 25138 17187
rect 25240 17151 25274 17185
rect 25513 17153 25547 17187
rect 29837 17153 29871 17187
rect 949 17085 983 17119
rect 1685 17085 1719 17119
rect 3249 17085 3283 17119
rect 3893 17085 3927 17119
rect 6101 17085 6135 17119
rect 8585 17085 8619 17119
rect 8677 17085 8711 17119
rect 9413 17085 9447 17119
rect 10885 17085 10919 17119
rect 11253 17085 11287 17119
rect 11989 17085 12023 17119
rect 13645 17085 13679 17119
rect 14524 17085 14558 17119
rect 14933 17085 14967 17119
rect 16405 17085 16439 17119
rect 17141 17085 17175 17119
rect 18797 17085 18831 17119
rect 19073 17085 19107 17119
rect 20545 17085 20579 17119
rect 22845 17085 22879 17119
rect 23489 17085 23523 17119
rect 24041 17085 24075 17119
rect 24225 17085 24259 17119
rect 24777 17085 24811 17119
rect 26985 17085 27019 17119
rect 27261 17085 27295 17119
rect 29101 17085 29135 17119
rect 29653 17085 29687 17119
rect 3525 17017 3559 17051
rect 24501 17017 24535 17051
rect 30113 17017 30147 17051
rect 1415 16949 1449 16983
rect 4359 16949 4393 16983
rect 6567 16949 6601 16983
rect 9143 16949 9177 16983
rect 11719 16949 11753 16983
rect 13093 16949 13127 16983
rect 18245 16949 18279 16983
rect 21011 16949 21045 16983
rect 22385 16949 22419 16983
rect 23121 16949 23155 16983
rect 23857 16949 23891 16983
rect 26617 16949 26651 16983
rect 28365 16949 28399 16983
rect 29929 16949 29963 16983
rect 3157 16745 3191 16779
rect 3991 16745 4025 16779
rect 6291 16745 6325 16779
rect 7665 16745 7699 16779
rect 8033 16745 8067 16779
rect 10425 16745 10459 16779
rect 13461 16745 13495 16779
rect 14295 16745 14329 16779
rect 15669 16745 15703 16779
rect 17515 16745 17549 16779
rect 21005 16745 21039 16779
rect 23955 16745 23989 16779
rect 26065 16745 26099 16779
rect 26801 16745 26835 16779
rect 28279 16745 28313 16779
rect 29653 16745 29687 16779
rect 30389 16745 30423 16779
rect 5641 16677 5675 16711
rect 23397 16677 23431 16711
rect 30113 16677 30147 16711
rect 1225 16609 1259 16643
rect 1317 16609 1351 16643
rect 1644 16609 1678 16643
rect 3525 16609 3559 16643
rect 4261 16609 4295 16643
rect 5825 16609 5859 16643
rect 6561 16609 6595 16643
rect 8217 16609 8251 16643
rect 8493 16609 8527 16643
rect 9321 16609 9355 16643
rect 11161 16609 11195 16643
rect 11621 16609 11655 16643
rect 11948 16609 11982 16643
rect 13829 16609 13863 16643
rect 16405 16609 16439 16643
rect 16681 16609 16715 16643
rect 19717 16609 19751 16643
rect 21608 16609 21642 16643
rect 22017 16609 22051 16643
rect 23489 16609 23523 16643
rect 25789 16609 25823 16643
rect 26709 16609 26743 16643
rect 27261 16609 27295 16643
rect 27813 16609 27847 16643
rect 28549 16609 28583 16643
rect 1813 16559 1847 16593
rect 2053 16541 2087 16575
rect 3988 16543 4022 16577
rect 6331 16543 6365 16577
rect 8585 16541 8619 16575
rect 8912 16541 8946 16575
rect 9091 16543 9125 16577
rect 12117 16543 12151 16577
rect 12357 16541 12391 16575
rect 14292 16543 14326 16577
rect 14565 16541 14599 16575
rect 17049 16541 17083 16575
rect 17545 16559 17579 16593
rect 17785 16541 17819 16575
rect 19441 16541 19475 16575
rect 21281 16541 21315 16575
rect 21787 16541 21821 16575
rect 23968 16541 24002 16575
rect 24225 16541 24259 16575
rect 28319 16541 28353 16575
rect 8309 16473 8343 16507
rect 11437 16473 11471 16507
rect 1041 16405 1075 16439
rect 16221 16405 16255 16439
rect 18889 16405 18923 16439
rect 25329 16405 25363 16439
rect 27537 16405 27571 16439
rect 2973 16201 3007 16235
rect 5641 16201 5675 16235
rect 7941 16201 7975 16235
rect 10977 16201 11011 16235
rect 23581 16201 23615 16235
rect 30297 16201 30331 16235
rect 16497 16133 16531 16167
rect 18429 16133 18463 16167
rect 20729 16133 20763 16167
rect 949 16065 983 16099
rect 1455 16065 1489 16099
rect 4307 16065 4341 16099
rect 6607 16063 6641 16097
rect 8585 16065 8619 16099
rect 9091 16065 9125 16099
rect 11759 16065 11793 16099
rect 14984 16065 15018 16099
rect 15120 16063 15154 16097
rect 19032 16065 19066 16099
rect 19211 16065 19245 16099
rect 21884 16065 21918 16099
rect 22053 16047 22087 16081
rect 23857 16065 23891 16099
rect 24184 16065 24218 16099
rect 24363 16063 24397 16097
rect 24593 16065 24627 16099
rect 26065 16065 26099 16099
rect 26528 16065 26562 16099
rect 26801 16065 26835 16099
rect 1685 15997 1719 16031
rect 3801 15997 3835 16031
rect 4128 15997 4162 16031
rect 4537 15997 4571 16031
rect 6101 15997 6135 16031
rect 6428 15997 6462 16031
rect 6837 15997 6871 16031
rect 9321 15997 9355 16031
rect 11161 15997 11195 16031
rect 11253 15997 11287 16031
rect 11989 15997 12023 16031
rect 14565 15997 14599 16031
rect 14657 15997 14691 16031
rect 15393 15997 15427 16031
rect 16865 15997 16899 16031
rect 17141 15997 17175 16031
rect 18705 15997 18739 16031
rect 19441 15997 19475 16031
rect 20913 15997 20947 16031
rect 21557 15997 21591 16031
rect 22293 15997 22327 16031
rect 28273 15997 28307 16031
rect 29285 15997 29319 16031
rect 29377 15997 29411 16031
rect 29745 15997 29779 16031
rect 30205 15997 30239 16031
rect 3341 15929 3375 15963
rect 13829 15929 13863 15963
rect 21189 15929 21223 15963
rect 28549 15929 28583 15963
rect 29101 15929 29135 15963
rect 1415 15861 1449 15895
rect 3617 15861 3651 15895
rect 9051 15861 9085 15895
rect 10425 15861 10459 15895
rect 11719 15861 11753 15895
rect 13093 15861 13127 15895
rect 14105 15861 14139 15895
rect 14381 15861 14415 15895
rect 25697 15861 25731 15895
rect 26531 15861 26565 15895
rect 27905 15861 27939 15895
rect 29561 15861 29595 15895
rect 29929 15861 29963 15895
rect 3157 15657 3191 15691
rect 5365 15657 5399 15691
rect 14295 15657 14329 15691
rect 18981 15657 19015 15691
rect 23121 15657 23155 15691
rect 23955 15657 23989 15691
rect 28273 15657 28307 15691
rect 30389 15657 30423 15691
rect 11069 15589 11103 15623
rect 11437 15589 11471 15623
rect 16221 15589 16255 15623
rect 16589 15589 16623 15623
rect 25881 15589 25915 15623
rect 1133 15521 1167 15555
rect 1644 15521 1678 15555
rect 5917 15521 5951 15555
rect 8585 15521 8619 15555
rect 11621 15521 11655 15555
rect 11948 15521 11982 15555
rect 13829 15521 13863 15555
rect 14565 15521 14599 15555
rect 15945 15521 15979 15555
rect 17049 15521 17083 15555
rect 17141 15521 17175 15555
rect 19441 15521 19475 15555
rect 21281 15521 21315 15555
rect 22017 15521 22051 15555
rect 26760 15521 26794 15555
rect 28917 15521 28951 15555
rect 30573 15521 30607 15555
rect 1317 15453 1351 15487
rect 1813 15471 1847 15505
rect 2053 15453 2087 15487
rect 3525 15453 3559 15487
rect 3852 15453 3886 15487
rect 4031 15453 4065 15487
rect 4261 15453 4295 15487
rect 6193 15453 6227 15487
rect 6377 15453 6411 15487
rect 6704 15453 6738 15487
rect 6883 15453 6917 15487
rect 7113 15453 7147 15487
rect 8912 15453 8946 15487
rect 9081 15471 9115 15505
rect 9321 15453 9355 15487
rect 12127 15453 12161 15487
rect 12357 15453 12391 15487
rect 14335 15453 14369 15487
rect 17468 15453 17502 15487
rect 17647 15453 17681 15487
rect 17877 15453 17911 15487
rect 19717 15453 19751 15487
rect 21608 15453 21642 15487
rect 21787 15453 21821 15487
rect 23489 15453 23523 15487
rect 23952 15455 23986 15489
rect 24225 15453 24259 15487
rect 26433 15453 26467 15487
rect 26939 15453 26973 15487
rect 27169 15453 27203 15487
rect 28641 15453 28675 15487
rect 16865 15385 16899 15419
rect 949 15317 983 15351
rect 8217 15317 8251 15351
rect 10425 15317 10459 15351
rect 13461 15317 13495 15351
rect 21005 15317 21039 15351
rect 25329 15317 25363 15351
rect 26157 15317 26191 15351
rect 30021 15317 30055 15351
rect 2789 15113 2823 15147
rect 5825 15113 5859 15147
rect 10977 15113 11011 15147
rect 13921 15113 13955 15147
rect 16037 15113 16071 15147
rect 18245 15113 18279 15147
rect 21649 15113 21683 15147
rect 28457 15113 28491 15147
rect 30113 15113 30147 15147
rect 30389 15113 30423 15147
rect 13093 15045 13127 15079
rect 23581 15045 23615 15079
rect 28089 15045 28123 15079
rect 949 14977 983 15011
rect 1455 14977 1489 15011
rect 4307 14977 4341 15011
rect 6607 14977 6641 15011
rect 8912 14977 8946 15011
rect 9091 14977 9125 15011
rect 11759 14977 11793 15011
rect 14703 14977 14737 15011
rect 16405 14977 16439 15011
rect 16911 14977 16945 15011
rect 20305 14959 20339 14993
rect 22293 14977 22327 15011
rect 23857 14977 23891 15011
rect 24184 14977 24218 15011
rect 24363 14977 24397 15011
rect 26528 14959 26562 14993
rect 1685 14909 1719 14943
rect 3249 14909 3283 14943
rect 3801 14909 3835 14943
rect 4537 14909 4571 14943
rect 6101 14909 6135 14943
rect 6837 14909 6871 14943
rect 8585 14909 8619 14943
rect 9321 14909 9355 14943
rect 11161 14909 11195 14943
rect 11253 14909 11287 14943
rect 11989 14909 12023 14943
rect 14197 14909 14231 14943
rect 14933 14909 14967 14943
rect 17141 14909 17175 14943
rect 18705 14909 18739 14943
rect 19349 14909 19383 14943
rect 19717 14909 19751 14943
rect 19809 14909 19843 14943
rect 20545 14909 20579 14943
rect 22017 14909 22051 14943
rect 24593 14909 24627 14943
rect 26065 14909 26099 14943
rect 26801 14909 26835 14943
rect 29469 14909 29503 14943
rect 30297 14909 30331 14943
rect 30573 14909 30607 14943
rect 3525 14841 3559 14875
rect 13645 14841 13679 14875
rect 18981 14841 19015 14875
rect 28365 14841 28399 14875
rect 29101 14841 29135 14875
rect 29653 14841 29687 14875
rect 1415 14773 1449 14807
rect 4267 14773 4301 14807
rect 6567 14773 6601 14807
rect 7941 14773 7975 14807
rect 10425 14773 10459 14807
rect 11719 14773 11753 14807
rect 14663 14773 14697 14807
rect 16871 14773 16905 14807
rect 20275 14773 20309 14807
rect 25697 14773 25731 14807
rect 26531 14773 26565 14807
rect 29929 14773 29963 14807
rect 3065 14569 3099 14603
rect 3991 14569 4025 14603
rect 5549 14569 5583 14603
rect 6101 14569 6135 14603
rect 9413 14569 9447 14603
rect 9689 14569 9723 14603
rect 9965 14569 9999 14603
rect 11069 14569 11103 14603
rect 11345 14569 11379 14603
rect 13461 14569 13495 14603
rect 14295 14569 14329 14603
rect 15669 14569 15703 14603
rect 19717 14569 19751 14603
rect 19993 14569 20027 14603
rect 20269 14569 20303 14603
rect 20545 14569 20579 14603
rect 21747 14569 21781 14603
rect 23121 14569 23155 14603
rect 23581 14569 23615 14603
rect 24599 14569 24633 14603
rect 26157 14569 26191 14603
rect 30389 14569 30423 14603
rect 9137 14501 9171 14535
rect 10517 14501 10551 14535
rect 1133 14433 1167 14467
rect 1225 14433 1259 14467
rect 3525 14433 3559 14467
rect 6009 14433 6043 14467
rect 6285 14433 6319 14467
rect 6561 14433 6595 14467
rect 8861 14433 8895 14467
rect 9597 14433 9631 14467
rect 9873 14433 9907 14467
rect 10149 14433 10183 14467
rect 10425 14433 10459 14467
rect 11253 14433 11287 14467
rect 11529 14433 11563 14467
rect 11948 14433 11982 14467
rect 16221 14433 16255 14467
rect 16865 14433 16899 14467
rect 17049 14433 17083 14467
rect 19441 14433 19475 14467
rect 19901 14433 19935 14467
rect 20177 14433 20211 14467
rect 20453 14433 20487 14467
rect 20729 14433 20763 14467
rect 21005 14433 21039 14467
rect 22017 14433 22051 14467
rect 23765 14433 23799 14467
rect 24041 14433 24075 14467
rect 24869 14433 24903 14467
rect 26433 14433 26467 14467
rect 26709 14433 26743 14467
rect 28508 14433 28542 14467
rect 30573 14433 30607 14467
rect 1552 14365 1586 14399
rect 1721 14383 1755 14417
rect 1961 14365 1995 14399
rect 4031 14365 4065 14399
rect 4261 14365 4295 14399
rect 6653 14365 6687 14399
rect 6980 14365 7014 14399
rect 7116 14365 7150 14399
rect 7389 14365 7423 14399
rect 11621 14365 11655 14399
rect 12127 14365 12161 14399
rect 12357 14365 12391 14399
rect 13829 14365 13863 14399
rect 14335 14365 14369 14399
rect 14565 14365 14599 14399
rect 17376 14365 17410 14399
rect 17545 14383 17579 14417
rect 17785 14365 17819 14399
rect 21281 14365 21315 14399
rect 21787 14365 21821 14399
rect 24133 14365 24167 14399
rect 24639 14365 24673 14399
rect 28181 14365 28215 14399
rect 28687 14365 28721 14399
rect 28917 14365 28951 14399
rect 6377 14297 6411 14331
rect 10241 14297 10275 14331
rect 16681 14297 16715 14331
rect 19257 14297 19291 14331
rect 30021 14297 30055 14331
rect 949 14229 983 14263
rect 5825 14229 5859 14263
rect 8677 14229 8711 14263
rect 16313 14229 16347 14263
rect 18889 14229 18923 14263
rect 20821 14229 20855 14263
rect 23857 14229 23891 14263
rect 27997 14229 28031 14263
rect 8401 14025 8435 14059
rect 8677 14025 8711 14059
rect 9045 14025 9079 14059
rect 9321 14025 9355 14059
rect 12633 14025 12667 14059
rect 13737 14025 13771 14059
rect 18705 14025 18739 14059
rect 21649 14025 21683 14059
rect 23397 14025 23431 14059
rect 28549 14025 28583 14059
rect 29285 14025 29319 14059
rect 29561 14025 29595 14059
rect 29837 14025 29871 14059
rect 30113 14025 30147 14059
rect 3341 13957 3375 13991
rect 7941 13957 7975 13991
rect 12357 13957 12391 13991
rect 13369 13957 13403 13991
rect 18245 13957 18279 13991
rect 19533 13957 19567 13991
rect 26249 13957 26283 13991
rect 949 13889 983 13923
rect 1455 13889 1489 13923
rect 3709 13889 3743 13923
rect 4215 13889 4249 13923
rect 6101 13889 6135 13923
rect 6607 13889 6641 13923
rect 10060 13889 10094 13923
rect 11713 13889 11747 13923
rect 14197 13889 14231 13923
rect 14524 13889 14558 13923
rect 14703 13889 14737 13923
rect 14933 13889 14967 13923
rect 16732 13889 16766 13923
rect 16911 13889 16945 13923
rect 20315 13889 20349 13923
rect 20545 13889 20579 13923
rect 22293 13889 22327 13923
rect 24504 13889 24538 13923
rect 24777 13889 24811 13923
rect 26709 13889 26743 13923
rect 27205 13871 27239 13905
rect 1685 13821 1719 13855
rect 3525 13821 3559 13855
rect 4445 13821 4479 13855
rect 6428 13821 6462 13855
rect 6837 13821 6871 13855
rect 8585 13821 8619 13855
rect 8861 13821 8895 13855
rect 9229 13821 9263 13855
rect 9505 13821 9539 13855
rect 9623 13821 9657 13855
rect 10333 13821 10367 13855
rect 11805 13821 11839 13855
rect 12081 13821 12115 13855
rect 12541 13821 12575 13855
rect 12817 13821 12851 13855
rect 12909 13821 12943 13855
rect 13185 13821 13219 13855
rect 13553 13821 13587 13855
rect 16313 13821 16347 13855
rect 16405 13821 16439 13855
rect 17141 13821 17175 13855
rect 18889 13821 18923 13855
rect 19165 13821 19199 13855
rect 19717 13821 19751 13855
rect 19809 13821 19843 13855
rect 22006 13821 22040 13855
rect 24041 13821 24075 13855
rect 24368 13821 24402 13855
rect 26425 13821 26459 13855
rect 27445 13821 27479 13855
rect 29193 13821 29227 13855
rect 29469 13821 29503 13855
rect 29745 13821 29779 13855
rect 30021 13821 30055 13855
rect 30297 13821 30331 13855
rect 30573 13821 30607 13855
rect 5825 13753 5859 13787
rect 26157 13753 26191 13787
rect 1415 13685 1449 13719
rect 2789 13685 2823 13719
rect 4175 13685 4209 13719
rect 10063 13685 10097 13719
rect 13829 13685 13863 13719
rect 20275 13685 20309 13719
rect 27175 13685 27209 13719
rect 29009 13685 29043 13719
rect 30389 13685 30423 13719
rect 3991 13481 4025 13515
rect 5825 13481 5859 13515
rect 6193 13481 6227 13515
rect 8953 13481 8987 13515
rect 9413 13481 9447 13515
rect 9965 13481 9999 13515
rect 10977 13481 11011 13515
rect 13007 13481 13041 13515
rect 15485 13481 15519 13515
rect 15761 13481 15795 13515
rect 16589 13481 16623 13515
rect 16773 13481 16807 13515
rect 17877 13481 17911 13515
rect 20637 13481 20671 13515
rect 20913 13481 20947 13515
rect 21649 13481 21683 13515
rect 22391 13481 22425 13515
rect 24599 13481 24633 13515
rect 26899 13481 26933 13515
rect 30389 13481 30423 13515
rect 8861 13413 8895 13447
rect 24041 13413 24075 13447
rect 26249 13413 26283 13447
rect 1225 13345 1259 13379
rect 2053 13345 2087 13379
rect 3433 13345 3467 13379
rect 6009 13345 6043 13379
rect 6377 13345 6411 13379
rect 6653 13345 6687 13379
rect 9137 13345 9171 13379
rect 9229 13345 9263 13379
rect 9781 13345 9815 13379
rect 10333 13345 10367 13379
rect 10609 13345 10643 13379
rect 11161 13345 11195 13379
rect 11253 13345 11287 13379
rect 11805 13345 11839 13379
rect 12081 13345 12115 13379
rect 14933 13345 14967 13379
rect 15669 13345 15703 13379
rect 15945 13345 15979 13379
rect 16957 13345 16991 13379
rect 17233 13345 17267 13379
rect 17785 13345 17819 13379
rect 18061 13345 18095 13379
rect 20813 13345 20847 13379
rect 21097 13345 21131 13379
rect 21557 13345 21591 13379
rect 21833 13345 21867 13379
rect 22661 13345 22695 13379
rect 24133 13345 24167 13379
rect 24869 13345 24903 13379
rect 27169 13345 27203 13379
rect 28917 13345 28951 13379
rect 30573 13345 30607 13379
rect 1317 13277 1351 13311
rect 1644 13277 1678 13311
rect 1823 13279 1857 13313
rect 3525 13277 3559 13311
rect 3988 13279 4022 13313
rect 4261 13277 4295 13311
rect 6745 13277 6779 13311
rect 7072 13277 7106 13311
rect 7208 13277 7242 13311
rect 7481 13277 7515 13311
rect 9505 13277 9539 13311
rect 11529 13277 11563 13311
rect 12541 13277 12575 13311
rect 13004 13277 13038 13311
rect 13277 13277 13311 13311
rect 15117 13277 15151 13311
rect 18337 13277 18371 13311
rect 18664 13277 18698 13311
rect 18800 13277 18834 13311
rect 19073 13277 19107 13311
rect 21925 13277 21959 13311
rect 22431 13277 22465 13311
rect 24639 13277 24673 13311
rect 26433 13277 26467 13311
rect 26896 13295 26930 13329
rect 28641 13277 28675 13311
rect 10425 13209 10459 13243
rect 17601 13209 17635 13243
rect 28273 13209 28307 13243
rect 1041 13141 1075 13175
rect 5549 13141 5583 13175
rect 6469 13141 6503 13175
rect 10149 13141 10183 13175
rect 11437 13141 11471 13175
rect 11989 13141 12023 13175
rect 14381 13141 14415 13175
rect 20361 13141 20395 13175
rect 21373 13141 21407 13175
rect 30021 13141 30055 13175
rect 2973 12937 3007 12971
rect 5917 12937 5951 12971
rect 8769 12937 8803 12971
rect 9229 12937 9263 12971
rect 12909 12937 12943 12971
rect 17601 12937 17635 12971
rect 22937 12937 22971 12971
rect 25697 12937 25731 12971
rect 28457 12937 28491 12971
rect 30297 12937 30331 12971
rect 30481 12937 30515 12971
rect 3617 12869 3651 12903
rect 8585 12869 8619 12903
rect 9321 12869 9355 12903
rect 11989 12869 12023 12903
rect 18245 12869 18279 12903
rect 23121 12869 23155 12903
rect 29561 12869 29595 12903
rect 1445 12783 1479 12817
rect 3433 12801 3467 12835
rect 4356 12801 4390 12835
rect 6564 12801 6598 12835
rect 6837 12801 6871 12835
rect 9597 12801 9631 12835
rect 9924 12801 9958 12835
rect 10103 12799 10137 12833
rect 10333 12801 10367 12835
rect 11713 12801 11747 12835
rect 14016 12801 14050 12835
rect 16240 12799 16274 12833
rect 18705 12801 18739 12835
rect 19168 12801 19202 12835
rect 21376 12801 21410 12835
rect 24320 12801 24354 12835
rect 26341 12801 26375 12835
rect 26944 12801 26978 12835
rect 27123 12801 27157 12835
rect 27353 12801 27387 12835
rect 949 12733 983 12767
rect 1685 12733 1719 12767
rect 3801 12733 3835 12767
rect 3893 12733 3927 12767
rect 4629 12733 4663 12767
rect 6101 12733 6135 12767
rect 8401 12733 8435 12767
rect 8953 12733 8987 12767
rect 9045 12733 9079 12767
rect 9505 12733 9539 12767
rect 11805 12733 11839 12767
rect 12265 12733 12299 12767
rect 12817 12733 12851 12767
rect 13093 12733 13127 12767
rect 13369 12733 13403 12767
rect 13553 12733 13587 12767
rect 14289 12733 14323 12767
rect 15761 12733 15795 12767
rect 16088 12733 16122 12767
rect 16497 12733 16531 12767
rect 18429 12733 18463 12767
rect 19441 12733 19475 12767
rect 20913 12733 20947 12767
rect 21649 12733 21683 12767
rect 23305 12733 23339 12767
rect 23581 12733 23615 12767
rect 23857 12733 23891 12767
rect 24593 12733 24627 12767
rect 26065 12733 26099 12767
rect 26617 12733 26651 12767
rect 29745 12733 29779 12767
rect 29837 12733 29871 12767
rect 30113 12733 30147 12767
rect 30389 12733 30423 12767
rect 12357 12665 12391 12699
rect 29101 12665 29135 12699
rect 1415 12597 1449 12631
rect 4359 12597 4393 12631
rect 6567 12597 6601 12631
rect 8125 12597 8159 12631
rect 12081 12597 12115 12631
rect 12633 12597 12667 12631
rect 13185 12597 13219 12631
rect 14019 12597 14053 12631
rect 15393 12597 15427 12631
rect 19171 12597 19205 12631
rect 20729 12597 20763 12631
rect 21379 12597 21413 12631
rect 23397 12597 23431 12631
rect 24323 12597 24357 12631
rect 29193 12597 29227 12631
rect 30021 12597 30055 12631
rect 1783 12393 1817 12427
rect 5549 12393 5583 12427
rect 5825 12393 5859 12427
rect 8493 12393 8527 12427
rect 10977 12393 11011 12427
rect 11253 12393 11287 12427
rect 12081 12393 12115 12427
rect 16681 12393 16715 12427
rect 18981 12393 19015 12427
rect 19717 12393 19751 12427
rect 19993 12393 20027 12427
rect 20637 12393 20671 12427
rect 23121 12393 23155 12427
rect 25329 12393 25363 12427
rect 28555 12393 28589 12427
rect 29929 12393 29963 12427
rect 25973 12325 26007 12359
rect 26893 12325 26927 12359
rect 1225 12257 1259 12291
rect 3433 12257 3467 12291
rect 3852 12257 3886 12291
rect 4261 12257 4295 12291
rect 6009 12257 6043 12291
rect 6377 12257 6411 12291
rect 6469 12257 6503 12291
rect 6796 12257 6830 12291
rect 9004 12257 9038 12291
rect 9413 12257 9447 12291
rect 11161 12257 11195 12291
rect 11437 12257 11471 12291
rect 11713 12257 11747 12291
rect 11989 12257 12023 12291
rect 12265 12257 12299 12291
rect 12541 12257 12575 12291
rect 13369 12257 13403 12291
rect 14841 12257 14875 12291
rect 16865 12257 16899 12291
rect 17693 12257 17727 12291
rect 19165 12257 19199 12291
rect 19901 12257 19935 12291
rect 20177 12257 20211 12291
rect 20545 12257 20579 12291
rect 20821 12257 20855 12291
rect 21097 12257 21131 12291
rect 21281 12257 21315 12291
rect 22017 12257 22051 12291
rect 24225 12257 24259 12291
rect 25697 12257 25731 12291
rect 26525 12257 26559 12291
rect 27077 12257 27111 12291
rect 27537 12257 27571 12291
rect 28089 12257 28123 12291
rect 30389 12257 30423 12291
rect 1317 12189 1351 12223
rect 1823 12191 1857 12225
rect 2053 12189 2087 12223
rect 3525 12189 3559 12223
rect 3988 12191 4022 12225
rect 6932 12189 6966 12223
rect 7205 12189 7239 12223
rect 8677 12189 8711 12223
rect 9140 12189 9174 12223
rect 12633 12189 12667 12223
rect 12960 12189 12994 12223
rect 13112 12191 13146 12225
rect 15025 12189 15059 12223
rect 15669 12189 15703 12223
rect 16313 12189 16347 12223
rect 16957 12189 16991 12223
rect 17284 12189 17318 12223
rect 17463 12189 17497 12223
rect 19349 12189 19383 12223
rect 21608 12189 21642 12223
rect 21787 12189 21821 12223
rect 23489 12189 23523 12223
rect 23816 12189 23850 12223
rect 23952 12189 23986 12223
rect 28595 12189 28629 12223
rect 28825 12189 28859 12223
rect 10701 12121 10735 12155
rect 20361 12121 20395 12155
rect 27721 12121 27755 12155
rect 1041 12053 1075 12087
rect 6193 12053 6227 12087
rect 11529 12053 11563 12087
rect 11805 12053 11839 12087
rect 12357 12053 12391 12087
rect 14473 12053 14507 12087
rect 20913 12053 20947 12087
rect 27169 12053 27203 12087
rect 30573 12053 30607 12087
rect 2973 11849 3007 11883
rect 5365 11849 5399 11883
rect 7757 11849 7791 11883
rect 8861 11849 8895 11883
rect 12173 11849 12207 11883
rect 13277 11849 13311 11883
rect 22937 11849 22971 11883
rect 25973 11849 26007 11883
rect 27997 11849 28031 11883
rect 28641 11849 28675 11883
rect 29561 11849 29595 11883
rect 8585 11781 8619 11815
rect 11529 11781 11563 11815
rect 23489 11781 23523 11815
rect 28365 11781 28399 11815
rect 949 11713 983 11747
rect 1276 11713 1310 11747
rect 1455 11713 1489 11747
rect 3804 11713 3838 11747
rect 6012 11713 6046 11747
rect 9689 11713 9723 11747
rect 10152 11713 10186 11747
rect 10425 11713 10459 11747
rect 14016 11713 14050 11747
rect 16868 11713 16902 11747
rect 19168 11711 19202 11745
rect 19441 11713 19475 11747
rect 21376 11713 21410 11747
rect 21649 11713 21683 11747
rect 24455 11711 24489 11745
rect 26663 11711 26697 11745
rect 1685 11645 1719 11679
rect 3341 11645 3375 11679
rect 4077 11645 4111 11679
rect 5549 11645 5583 11679
rect 6285 11645 6319 11679
rect 7941 11645 7975 11679
rect 8217 11645 8251 11679
rect 8401 11645 8435 11679
rect 8677 11645 8711 11679
rect 9229 11645 9263 11679
rect 12081 11645 12115 11679
rect 12357 11645 12391 11679
rect 12541 11645 12575 11679
rect 13001 11645 13035 11679
rect 13553 11645 13587 11679
rect 14289 11645 14323 11679
rect 16405 11645 16439 11679
rect 17141 11645 17175 11679
rect 18705 11645 18739 11679
rect 20913 11645 20947 11679
rect 23397 11645 23431 11679
rect 23673 11645 23707 11679
rect 23949 11645 23983 11679
rect 24276 11645 24310 11679
rect 24685 11645 24719 11679
rect 26157 11645 26191 11679
rect 26893 11645 26927 11679
rect 28549 11645 28583 11679
rect 28825 11645 28859 11679
rect 29745 11645 29779 11679
rect 13185 11577 13219 11611
rect 20821 11577 20855 11611
rect 29101 11577 29135 11611
rect 3807 11509 3841 11543
rect 6015 11509 6049 11543
rect 7389 11509 7423 11543
rect 8033 11509 8067 11543
rect 9321 11509 9355 11543
rect 10155 11509 10189 11543
rect 11897 11509 11931 11543
rect 12633 11509 12667 11543
rect 12817 11509 12851 11543
rect 14019 11509 14053 11543
rect 15393 11509 15427 11543
rect 16037 11509 16071 11543
rect 16871 11509 16905 11543
rect 18429 11509 18463 11543
rect 19171 11509 19205 11543
rect 21379 11509 21413 11543
rect 23213 11509 23247 11543
rect 26623 11509 26657 11543
rect 29193 11509 29227 11543
rect 1133 11305 1167 11339
rect 3525 11305 3559 11339
rect 4261 11305 4295 11339
rect 5089 11305 5123 11339
rect 5365 11305 5399 11339
rect 6009 11305 6043 11339
rect 9413 11305 9447 11339
rect 9689 11305 9723 11339
rect 10977 11305 11011 11339
rect 16681 11305 16715 11339
rect 18797 11305 18831 11339
rect 22851 11305 22885 11339
rect 24409 11305 24443 11339
rect 1041 11237 1075 11271
rect 12265 11237 12299 11271
rect 14841 11237 14875 11271
rect 2237 11169 2271 11203
rect 3709 11169 3743 11203
rect 3985 11169 4019 11203
rect 4421 11169 4455 11203
rect 4629 11169 4663 11203
rect 5273 11169 5307 11203
rect 5549 11169 5583 11203
rect 6469 11169 6503 11203
rect 6653 11169 6687 11203
rect 6980 11169 7014 11203
rect 7389 11169 7423 11203
rect 8861 11169 8895 11203
rect 9229 11169 9263 11203
rect 9505 11169 9539 11203
rect 9781 11169 9815 11203
rect 10333 11169 10367 11203
rect 10609 11169 10643 11203
rect 11161 11169 11195 11203
rect 11437 11169 11471 11203
rect 11713 11169 11747 11203
rect 11805 11169 11839 11203
rect 12868 11169 12902 11203
rect 15485 11169 15519 11203
rect 16589 11169 16623 11203
rect 16865 11169 16899 11203
rect 16957 11169 16991 11203
rect 17693 11169 17727 11203
rect 19257 11169 19291 11203
rect 19993 11169 20027 11203
rect 21465 11169 21499 11203
rect 22385 11169 22419 11203
rect 23121 11169 23155 11203
rect 24685 11169 24719 11203
rect 25237 11169 25271 11203
rect 25789 11169 25823 11203
rect 26433 11169 26467 11203
rect 28641 11169 28675 11203
rect 28917 11169 28951 11203
rect 1501 11101 1535 11135
rect 1828 11101 1862 11135
rect 2007 11103 2041 11137
rect 4905 11101 4939 11135
rect 7116 11101 7150 11135
rect 8769 11101 8803 11135
rect 12449 11101 12483 11135
rect 12541 11101 12575 11135
rect 13004 11101 13038 11135
rect 13277 11101 13311 11135
rect 15117 11101 15151 11135
rect 17284 11101 17318 11135
rect 17463 11101 17497 11135
rect 22848 11103 22882 11137
rect 26065 11101 26099 11135
rect 26760 11101 26794 11135
rect 26929 11119 26963 11153
rect 27169 11101 27203 11135
rect 6285 11033 6319 11067
rect 10425 11033 10459 11067
rect 11253 11033 11287 11067
rect 11529 11033 11563 11067
rect 11989 11033 12023 11067
rect 15301 11033 15335 11067
rect 15761 11033 15795 11067
rect 16405 11033 16439 11067
rect 28273 11033 28307 11067
rect 30021 11033 30055 11067
rect 9045 10965 9079 10999
rect 9965 10965 9999 10999
rect 10149 10965 10183 10999
rect 14381 10965 14415 10999
rect 19533 10965 19567 10999
rect 21281 10965 21315 10999
rect 24869 10965 24903 10999
rect 25329 10965 25363 10999
rect 5273 10761 5307 10795
rect 7941 10761 7975 10795
rect 11621 10761 11655 10795
rect 13553 10761 13587 10795
rect 22753 10761 22787 10795
rect 23489 10761 23523 10795
rect 19625 10693 19659 10727
rect 29009 10693 29043 10727
rect 949 10625 983 10659
rect 1455 10625 1489 10659
rect 3065 10625 3099 10659
rect 3712 10625 3746 10659
rect 6012 10625 6046 10659
rect 8677 10625 8711 10659
rect 10060 10625 10094 10659
rect 10333 10625 10367 10659
rect 13829 10625 13863 10659
rect 14292 10623 14326 10657
rect 16868 10625 16902 10659
rect 20499 10625 20533 10659
rect 24320 10625 24354 10659
rect 26484 10625 26518 10659
rect 26663 10625 26697 10659
rect 26893 10625 26927 10659
rect 1685 10557 1719 10591
rect 3249 10557 3283 10591
rect 3985 10557 4019 10591
rect 5549 10557 5583 10591
rect 5876 10557 5910 10591
rect 6285 10557 6319 10591
rect 8401 10557 8435 10591
rect 8953 10557 8987 10591
rect 9505 10557 9539 10591
rect 9597 10557 9631 10591
rect 11897 10557 11931 10591
rect 12909 10557 12943 10591
rect 13737 10557 13771 10591
rect 14156 10557 14190 10591
rect 14565 10557 14599 10591
rect 16221 10557 16255 10591
rect 16405 10557 16439 10591
rect 17141 10557 17175 10591
rect 18889 10557 18923 10591
rect 19993 10557 20027 10591
rect 20320 10557 20354 10591
rect 20729 10557 20763 10591
rect 22477 10557 22511 10591
rect 22937 10557 22971 10591
rect 23673 10557 23707 10591
rect 23857 10557 23891 10591
rect 24184 10557 24218 10591
rect 24593 10557 24627 10591
rect 26157 10557 26191 10591
rect 29193 10557 29227 10591
rect 29469 10557 29503 10591
rect 29745 10557 29779 10591
rect 30021 10557 30055 10591
rect 7665 10489 7699 10523
rect 7849 10489 7883 10523
rect 12265 10489 12299 10523
rect 12449 10489 12483 10523
rect 13185 10489 13219 10523
rect 15945 10489 15979 10523
rect 18521 10489 18555 10523
rect 28457 10489 28491 10523
rect 1415 10421 1449 10455
rect 3715 10421 3749 10455
rect 9137 10421 9171 10455
rect 9321 10421 9355 10455
rect 10063 10421 10097 10455
rect 12725 10421 12759 10455
rect 16037 10421 16071 10455
rect 16871 10421 16905 10455
rect 18705 10421 18739 10455
rect 19165 10421 19199 10455
rect 21833 10421 21867 10455
rect 22293 10421 22327 10455
rect 25697 10421 25731 10455
rect 28181 10421 28215 10455
rect 28549 10421 28583 10455
rect 29285 10421 29319 10455
rect 29561 10421 29595 10455
rect 29837 10421 29871 10455
rect 1599 10217 1633 10251
rect 3807 10217 3841 10251
rect 6935 10217 6969 10251
rect 9143 10217 9177 10251
rect 11627 10217 11661 10251
rect 14295 10217 14329 10251
rect 17239 10217 17273 10251
rect 20361 10217 20395 10251
rect 21747 10217 21781 10251
rect 23121 10217 23155 10251
rect 30021 10217 30055 10251
rect 5457 10149 5491 10183
rect 6193 10149 6227 10183
rect 16497 10149 16531 10183
rect 18889 10149 18923 10183
rect 1041 10081 1075 10115
rect 1133 10081 1167 10115
rect 3249 10081 3283 10115
rect 5917 10081 5951 10115
rect 8585 10081 8619 10115
rect 9413 10081 9447 10115
rect 13553 10081 13587 10115
rect 13829 10081 13863 10115
rect 14565 10081 14599 10115
rect 16221 10081 16255 10115
rect 17509 10081 17543 10115
rect 19349 10081 19383 10115
rect 19809 10081 19843 10115
rect 20085 10081 20119 10115
rect 20545 10081 20579 10115
rect 20729 10081 20763 10115
rect 21281 10081 21315 10115
rect 22017 10081 22051 10115
rect 23908 10081 23942 10115
rect 25973 10081 26007 10115
rect 26433 10081 26467 10115
rect 27169 10081 27203 10115
rect 28641 10081 28675 10115
rect 28917 10081 28951 10115
rect 1629 10031 1663 10065
rect 1869 10013 1903 10047
rect 3341 10013 3375 10047
rect 3804 10013 3838 10047
rect 4077 10013 4111 10047
rect 6469 10013 6503 10047
rect 6932 10015 6966 10049
rect 7205 10013 7239 10047
rect 8677 10013 8711 10047
rect 9140 10015 9174 10049
rect 11161 10013 11195 10047
rect 11624 10031 11658 10065
rect 11897 10013 11931 10047
rect 14335 10013 14369 10047
rect 16773 10013 16807 10047
rect 17279 10013 17313 10047
rect 21744 10013 21778 10047
rect 23581 10013 23615 10047
rect 24087 10013 24121 10047
rect 24317 10013 24351 10047
rect 26760 10013 26794 10047
rect 26896 10013 26930 10047
rect 19625 9945 19659 9979
rect 25605 9945 25639 9979
rect 857 9877 891 9911
rect 10701 9877 10735 9911
rect 13001 9877 13035 9911
rect 15669 9877 15703 9911
rect 19165 9877 19199 9911
rect 19901 9877 19935 9911
rect 20821 9877 20855 9911
rect 26157 9877 26191 9911
rect 28273 9877 28307 9911
rect 5825 9673 5859 9707
rect 10977 9673 11011 9707
rect 16129 9673 16163 9707
rect 22753 9673 22787 9707
rect 26433 9673 26467 9707
rect 28457 9673 28491 9707
rect 29009 9673 29043 9707
rect 3433 9605 3467 9639
rect 8585 9605 8619 9639
rect 18245 9605 18279 9639
rect 20545 9605 20579 9639
rect 949 9537 983 9571
rect 1455 9537 1489 9571
rect 3065 9537 3099 9571
rect 4080 9537 4114 9571
rect 6101 9537 6135 9571
rect 6607 9537 6641 9571
rect 9280 9537 9314 9571
rect 9416 9535 9450 9569
rect 9689 9537 9723 9571
rect 11624 9537 11658 9571
rect 14064 9537 14098 9571
rect 14243 9537 14277 9571
rect 16911 9537 16945 9571
rect 19168 9537 19202 9571
rect 21376 9537 21410 9571
rect 24409 9537 24443 9571
rect 24872 9537 24906 9571
rect 27080 9537 27114 9571
rect 1685 9469 1719 9503
rect 3617 9469 3651 9503
rect 3944 9469 3978 9503
rect 4353 9469 4387 9503
rect 6009 9469 6043 9503
rect 6837 9469 6871 9503
rect 8401 9469 8435 9503
rect 8953 9469 8987 9503
rect 11161 9469 11195 9503
rect 11897 9469 11931 9503
rect 13737 9469 13771 9503
rect 14473 9469 14507 9503
rect 16313 9469 16347 9503
rect 16405 9469 16439 9503
rect 17141 9469 17175 9503
rect 18705 9469 18739 9503
rect 19441 9469 19475 9503
rect 20913 9469 20947 9503
rect 21649 9469 21683 9503
rect 23489 9469 23523 9503
rect 24041 9469 24075 9503
rect 24317 9445 24351 9479
rect 25145 9469 25179 9503
rect 26617 9469 26651 9503
rect 27353 9469 27387 9503
rect 29193 9469 29227 9503
rect 29469 9469 29503 9503
rect 5733 9401 5767 9435
rect 8217 9401 8251 9435
rect 1415 9333 1449 9367
rect 6567 9333 6601 9367
rect 11627 9333 11661 9367
rect 13001 9333 13035 9367
rect 15577 9333 15611 9367
rect 16871 9333 16905 9367
rect 19171 9333 19205 9367
rect 21379 9333 21413 9367
rect 23305 9333 23339 9367
rect 23857 9333 23891 9367
rect 24133 9333 24167 9367
rect 24875 9333 24909 9367
rect 27083 9333 27117 9367
rect 29285 9333 29319 9367
rect 857 9129 891 9163
rect 4629 9129 4663 9163
rect 4905 9129 4939 9163
rect 5181 9129 5215 9163
rect 5457 9129 5491 9163
rect 7389 9129 7423 9163
rect 9505 9129 9539 9163
rect 9873 9129 9907 9163
rect 10609 9129 10643 9163
rect 14295 9129 14329 9163
rect 16129 9129 16163 9163
rect 17883 9129 17917 9163
rect 21747 9129 21781 9163
rect 23121 9129 23155 9163
rect 25329 9129 25363 9163
rect 25697 9129 25731 9163
rect 25973 9129 26007 9163
rect 26899 9129 26933 9163
rect 28273 9129 28307 9163
rect 30205 9129 30239 9163
rect 1961 9061 1995 9095
rect 13461 9061 13495 9095
rect 17141 9061 17175 9095
rect 19717 9061 19751 9095
rect 1041 8993 1075 9027
rect 1133 8993 1167 9027
rect 1685 8993 1719 9027
rect 2564 8993 2598 9027
rect 4813 8993 4847 9027
rect 5089 8993 5123 9027
rect 5365 8993 5399 9027
rect 5641 8993 5675 9027
rect 6009 8993 6043 9027
rect 6377 8993 6411 9027
rect 6653 8993 6687 9027
rect 6929 8993 6963 9027
rect 7205 8993 7239 9027
rect 7573 8993 7607 9027
rect 7665 8993 7699 9027
rect 7992 8993 8026 9027
rect 8401 8993 8435 9027
rect 10057 8993 10091 9027
rect 10517 8993 10551 9027
rect 10793 8993 10827 9027
rect 11897 8993 11931 9027
rect 13829 8993 13863 9027
rect 14565 8993 14599 9027
rect 16313 8993 16347 9027
rect 16589 8993 16623 9027
rect 16865 8993 16899 9027
rect 17417 8993 17451 9027
rect 18153 8993 18187 9027
rect 21281 8993 21315 9027
rect 24225 8993 24259 9027
rect 25881 8993 25915 9027
rect 26157 8993 26191 9027
rect 26433 8993 26467 9027
rect 27169 8993 27203 9027
rect 28641 8993 28675 9027
rect 28917 8993 28951 9027
rect 1409 8925 1443 8959
rect 2237 8925 2271 8959
rect 2743 8925 2777 8959
rect 2973 8925 3007 8959
rect 8128 8925 8162 8959
rect 11161 8925 11195 8959
rect 11488 8925 11522 8959
rect 11624 8927 11658 8961
rect 14325 8943 14359 8977
rect 17923 8925 17957 8959
rect 21787 8927 21821 8961
rect 22017 8925 22051 8959
rect 23479 8925 23513 8959
rect 23816 8925 23850 8959
rect 23995 8925 24029 8959
rect 26896 8925 26930 8959
rect 10333 8857 10367 8891
rect 19993 8857 20027 8891
rect 4077 8789 4111 8823
rect 5825 8789 5859 8823
rect 6193 8789 6227 8823
rect 6469 8789 6503 8823
rect 6745 8789 6779 8823
rect 7021 8789 7055 8823
rect 13001 8789 13035 8823
rect 13553 8789 13587 8823
rect 15669 8789 15703 8823
rect 16405 8789 16439 8823
rect 19257 8789 19291 8823
rect 20453 8789 20487 8823
rect 5089 8585 5123 8619
rect 7389 8585 7423 8619
rect 8033 8585 8067 8619
rect 11713 8585 11747 8619
rect 20545 8585 20579 8619
rect 25881 8585 25915 8619
rect 26065 8585 26099 8619
rect 28549 8585 28583 8619
rect 8401 8517 8435 8551
rect 8861 8517 8895 8551
rect 9413 8517 9447 8551
rect 21281 8517 21315 8551
rect 1455 8449 1489 8483
rect 3712 8449 3746 8483
rect 6012 8449 6046 8483
rect 10152 8449 10186 8483
rect 14064 8449 14098 8483
rect 14200 8449 14234 8483
rect 14473 8449 14507 8483
rect 15853 8449 15887 8483
rect 16408 8449 16442 8483
rect 19201 8431 19235 8465
rect 22063 8449 22097 8483
rect 23673 8449 23707 8483
rect 24320 8449 24354 8483
rect 27036 8449 27070 8483
rect 27215 8449 27249 8483
rect 949 8381 983 8415
rect 1685 8381 1719 8415
rect 3249 8381 3283 8415
rect 3985 8381 4019 8415
rect 5549 8381 5583 8415
rect 5876 8381 5910 8415
rect 6285 8381 6319 8415
rect 7941 8381 7975 8415
rect 8217 8381 8251 8415
rect 8585 8381 8619 8415
rect 8677 8381 8711 8415
rect 9321 8381 9355 8415
rect 9597 8381 9631 8415
rect 9689 8381 9723 8415
rect 10425 8381 10459 8415
rect 12541 8381 12575 8415
rect 12817 8381 12851 8415
rect 13093 8381 13127 8415
rect 13369 8381 13403 8415
rect 13737 8381 13771 8415
rect 15945 8381 15979 8415
rect 16681 8381 16715 8415
rect 18337 8381 18371 8415
rect 18705 8381 18739 8415
rect 19441 8381 19475 8415
rect 21465 8381 21499 8415
rect 21557 8381 21591 8415
rect 22293 8381 22327 8415
rect 23857 8381 23891 8415
rect 24593 8381 24627 8415
rect 26249 8381 26283 8415
rect 26709 8381 26743 8415
rect 27445 8381 27479 8415
rect 29101 8381 29135 8415
rect 3065 8313 3099 8347
rect 12173 8313 12207 8347
rect 18061 8313 18095 8347
rect 29653 8313 29687 8347
rect 1415 8245 1449 8279
rect 3715 8245 3749 8279
rect 7757 8245 7791 8279
rect 9137 8245 9171 8279
rect 10155 8245 10189 8279
rect 12633 8245 12667 8279
rect 12909 8245 12943 8279
rect 13185 8245 13219 8279
rect 16411 8245 16445 8279
rect 18153 8245 18187 8279
rect 19171 8245 19205 8279
rect 21097 8245 21131 8279
rect 22023 8245 22057 8279
rect 24323 8245 24357 8279
rect 29193 8245 29227 8279
rect 29929 8245 29963 8279
rect 857 8041 891 8075
rect 10517 8041 10551 8075
rect 12087 8041 12121 8075
rect 18803 8041 18837 8075
rect 20177 8041 20211 8075
rect 20821 8041 20855 8075
rect 23121 8041 23155 8075
rect 23955 8041 23989 8075
rect 28095 8041 28129 8075
rect 29469 8041 29503 8075
rect 1041 7905 1075 7939
rect 3341 7905 3375 7939
rect 3525 7905 3559 7939
rect 5917 7905 5951 7939
rect 6796 7905 6830 7939
rect 7205 7905 7239 7939
rect 8677 7905 8711 7939
rect 11069 7905 11103 7939
rect 11437 7905 11471 7939
rect 11621 7905 11655 7939
rect 12357 7905 12391 7939
rect 13829 7905 13863 7939
rect 14156 7905 14190 7939
rect 14565 7905 14599 7939
rect 20729 7905 20763 7939
rect 21005 7905 21039 7939
rect 21608 7905 21642 7939
rect 23489 7905 23523 7939
rect 25697 7905 25731 7939
rect 26617 7905 26651 7939
rect 27261 7905 27295 7939
rect 27537 7905 27571 7939
rect 28365 7905 28399 7939
rect 30021 7905 30055 7939
rect 1225 7837 1259 7871
rect 1552 7837 1586 7871
rect 1721 7855 1755 7889
rect 1961 7837 1995 7871
rect 3852 7837 3886 7871
rect 4031 7837 4065 7871
rect 4261 7837 4295 7871
rect 6193 7837 6227 7871
rect 6469 7837 6503 7871
rect 6975 7837 7009 7871
rect 9004 7837 9038 7871
rect 9183 7837 9217 7871
rect 9413 7837 9447 7871
rect 12127 7837 12161 7871
rect 14335 7837 14369 7871
rect 16129 7837 16163 7871
rect 16456 7837 16490 7871
rect 16592 7837 16626 7871
rect 16865 7837 16899 7871
rect 18337 7837 18371 7871
rect 18843 7837 18877 7871
rect 19073 7837 19107 7871
rect 21281 7837 21315 7871
rect 21777 7839 21811 7873
rect 22017 7837 22051 7871
rect 23952 7837 23986 7871
rect 24225 7837 24259 7871
rect 25881 7837 25915 7871
rect 27629 7837 27663 7871
rect 28125 7855 28159 7889
rect 27077 7769 27111 7803
rect 5549 7701 5583 7735
rect 8309 7701 8343 7735
rect 13461 7701 13495 7735
rect 15669 7701 15703 7735
rect 17969 7701 18003 7735
rect 20545 7701 20579 7735
rect 25329 7701 25363 7735
rect 26433 7701 26467 7735
rect 27353 7701 27387 7735
rect 29837 7701 29871 7735
rect 5365 7497 5399 7531
rect 5733 7497 5767 7531
rect 18337 7497 18371 7531
rect 23489 7497 23523 7531
rect 25881 7497 25915 7531
rect 3249 7429 3283 7463
rect 17969 7429 18003 7463
rect 29285 7429 29319 7463
rect 1455 7361 1489 7395
rect 4031 7361 4065 7395
rect 6607 7361 6641 7395
rect 6837 7361 6871 7395
rect 9045 7361 9079 7395
rect 9551 7361 9585 7395
rect 11253 7361 11287 7395
rect 11759 7361 11793 7395
rect 14384 7361 14418 7395
rect 14657 7361 14691 7395
rect 16592 7359 16626 7393
rect 18705 7361 18739 7395
rect 19211 7361 19245 7395
rect 19441 7361 19475 7395
rect 21792 7361 21826 7395
rect 21971 7361 22005 7395
rect 23857 7361 23891 7395
rect 24363 7361 24397 7395
rect 26561 7343 26595 7377
rect 949 7293 983 7327
rect 1685 7293 1719 7327
rect 3433 7293 3467 7327
rect 3525 7293 3559 7327
rect 4261 7293 4295 7327
rect 5917 7293 5951 7327
rect 6101 7293 6135 7327
rect 8217 7293 8251 7327
rect 8401 7293 8435 7327
rect 9372 7293 9406 7327
rect 9781 7293 9815 7327
rect 11989 7293 12023 7327
rect 13829 7293 13863 7327
rect 13921 7293 13955 7327
rect 16129 7293 16163 7327
rect 16865 7293 16899 7327
rect 18521 7293 18555 7327
rect 21097 7293 21131 7327
rect 21465 7293 21499 7327
rect 22201 7293 22235 7327
rect 24593 7293 24627 7327
rect 26065 7293 26099 7327
rect 26801 7293 26835 7327
rect 29193 7293 29227 7327
rect 29469 7293 29503 7327
rect 29745 7293 29779 7327
rect 8677 7225 8711 7259
rect 28365 7225 28399 7259
rect 1415 7157 1449 7191
rect 2789 7157 2823 7191
rect 3991 7157 4025 7191
rect 6567 7157 6601 7191
rect 10885 7157 10919 7191
rect 11719 7157 11753 7191
rect 13093 7157 13127 7191
rect 13645 7157 13679 7191
rect 14387 7157 14421 7191
rect 15761 7157 15795 7191
rect 16595 7157 16629 7191
rect 19171 7157 19205 7191
rect 20545 7157 20579 7191
rect 24323 7157 24357 7191
rect 26531 7157 26565 7191
rect 27905 7157 27939 7191
rect 28457 7157 28491 7191
rect 29009 7157 29043 7191
rect 29561 7157 29595 7191
rect 1599 6953 1633 6987
rect 5825 6953 5859 6987
rect 6101 6953 6135 6987
rect 6935 6953 6969 6987
rect 9143 6953 9177 6987
rect 10517 6953 10551 6987
rect 11253 6953 11287 6987
rect 15025 6953 15059 6987
rect 20637 6953 20671 6987
rect 21281 6953 21315 6987
rect 23949 6953 23983 6987
rect 26433 6953 26467 6987
rect 28095 6953 28129 6987
rect 3249 6885 3283 6919
rect 14565 6885 14599 6919
rect 1041 6817 1075 6851
rect 1133 6817 1167 6851
rect 3668 6817 3702 6851
rect 4077 6817 4111 6851
rect 5457 6817 5491 6851
rect 6009 6817 6043 6851
rect 6285 6817 6319 6851
rect 6469 6817 6503 6851
rect 7205 6817 7239 6851
rect 8677 6817 8711 6851
rect 9413 6817 9447 6851
rect 11161 6817 11195 6851
rect 11437 6817 11471 6851
rect 11529 6817 11563 6851
rect 11989 6817 12023 6851
rect 12081 6817 12115 6851
rect 12408 6817 12442 6851
rect 12817 6817 12851 6851
rect 14289 6817 14323 6851
rect 15209 6817 15243 6851
rect 15301 6817 15335 6851
rect 15761 6817 15795 6851
rect 16313 6817 16347 6851
rect 18613 6817 18647 6851
rect 21097 6817 21131 6851
rect 21465 6817 21499 6851
rect 21741 6817 21775 6851
rect 22252 6817 22286 6851
rect 22661 6817 22695 6851
rect 24133 6817 24167 6851
rect 24460 6817 24494 6851
rect 24869 6817 24903 6851
rect 26617 6817 26651 6851
rect 27169 6817 27203 6851
rect 28365 6817 28399 6851
rect 29745 6817 29779 6851
rect 1639 6749 1673 6783
rect 1869 6749 1903 6783
rect 3341 6749 3375 6783
rect 3847 6749 3881 6783
rect 6975 6751 7009 6785
rect 9183 6749 9217 6783
rect 12544 6751 12578 6785
rect 16405 6749 16439 6783
rect 16732 6749 16766 6783
rect 16911 6749 16945 6783
rect 17141 6749 17175 6783
rect 18940 6749 18974 6783
rect 19119 6751 19153 6785
rect 19349 6749 19383 6783
rect 21925 6749 21959 6783
rect 22388 6749 22422 6783
rect 24639 6749 24673 6783
rect 27629 6749 27663 6783
rect 28092 6749 28126 6783
rect 8309 6681 8343 6715
rect 10977 6681 11011 6715
rect 11805 6681 11839 6715
rect 15485 6681 15519 6715
rect 857 6613 891 6647
rect 11713 6613 11747 6647
rect 13921 6613 13955 6647
rect 15945 6613 15979 6647
rect 16129 6613 16163 6647
rect 18429 6613 18463 6647
rect 20913 6613 20947 6647
rect 21557 6613 21591 6647
rect 25973 6613 26007 6647
rect 27261 6613 27295 6647
rect 7941 6409 7975 6443
rect 8953 6409 8987 6443
rect 11069 6409 11103 6443
rect 12633 6409 12667 6443
rect 13093 6409 13127 6443
rect 13185 6409 13219 6443
rect 13737 6409 13771 6443
rect 16405 6409 16439 6443
rect 18337 6409 18371 6443
rect 28549 6409 28583 6443
rect 5825 6341 5859 6375
rect 11805 6341 11839 6375
rect 1455 6273 1489 6307
rect 3065 6273 3099 6307
rect 3847 6273 3881 6307
rect 4077 6273 4111 6307
rect 6101 6273 6135 6307
rect 6428 6273 6462 6307
rect 6607 6271 6641 6305
rect 6837 6273 6871 6307
rect 9229 6273 9263 6307
rect 9556 6273 9590 6307
rect 9735 6273 9769 6307
rect 9965 6273 9999 6307
rect 14892 6273 14926 6307
rect 15071 6273 15105 6307
rect 17877 6273 17911 6307
rect 19901 6273 19935 6307
rect 20407 6273 20441 6307
rect 23029 6273 23063 6307
rect 23397 6273 23431 6307
rect 24547 6273 24581 6307
rect 27172 6271 27206 6305
rect 27445 6273 27479 6307
rect 949 6205 983 6239
rect 1685 6205 1719 6239
rect 3341 6205 3375 6239
rect 5733 6205 5767 6239
rect 6009 6205 6043 6239
rect 8401 6205 8435 6239
rect 8861 6205 8895 6239
rect 9137 6205 9171 6239
rect 11713 6205 11747 6239
rect 11989 6205 12023 6239
rect 12265 6205 12299 6239
rect 12541 6205 12575 6239
rect 12809 6205 12843 6239
rect 12909 6205 12943 6239
rect 13369 6205 13403 6239
rect 13921 6205 13955 6239
rect 14105 6205 14139 6239
rect 14565 6205 14599 6239
rect 15301 6205 15335 6239
rect 16773 6205 16807 6239
rect 17509 6205 17543 6239
rect 17601 6205 17635 6239
rect 18521 6205 18555 6239
rect 18889 6205 18923 6239
rect 19165 6205 19199 6239
rect 19441 6205 19475 6239
rect 19717 6205 19751 6239
rect 20228 6205 20262 6239
rect 20637 6205 20671 6239
rect 22293 6205 22327 6239
rect 22569 6205 22603 6239
rect 22753 6205 22787 6239
rect 24041 6205 24075 6239
rect 24777 6205 24811 6239
rect 26709 6205 26743 6239
rect 29193 6205 29227 6239
rect 17049 6137 17083 6171
rect 26157 6137 26191 6171
rect 1415 6069 1449 6103
rect 3807 6069 3841 6103
rect 5181 6069 5215 6103
rect 5549 6069 5583 6103
rect 8585 6069 8619 6103
rect 8677 6069 8711 6103
rect 11529 6069 11563 6103
rect 12081 6069 12115 6103
rect 12357 6069 12391 6103
rect 14197 6069 14231 6103
rect 17325 6069 17359 6103
rect 18705 6069 18739 6103
rect 18981 6069 19015 6103
rect 19257 6069 19291 6103
rect 19533 6069 19567 6103
rect 21925 6069 21959 6103
rect 22109 6069 22143 6103
rect 22385 6069 22419 6103
rect 24507 6069 24541 6103
rect 27175 6069 27209 6103
rect 29009 6069 29043 6103
rect 857 5865 891 5899
rect 7205 5865 7239 5899
rect 8315 5865 8349 5899
rect 10793 5865 10827 5899
rect 11069 5865 11103 5899
rect 12087 5865 12121 5899
rect 20545 5865 20579 5899
rect 20821 5865 20855 5899
rect 24599 5865 24633 5899
rect 28003 5865 28037 5899
rect 29377 5865 29411 5899
rect 6101 5797 6135 5831
rect 1041 5729 1075 5763
rect 1644 5729 1678 5763
rect 3852 5729 3886 5763
rect 5825 5729 5859 5763
rect 6561 5729 6595 5763
rect 6837 5729 6871 5763
rect 7113 5729 7147 5763
rect 7389 5729 7423 5763
rect 7665 5729 7699 5763
rect 8585 5729 8619 5763
rect 10241 5729 10275 5763
rect 10517 5729 10551 5763
rect 10609 5729 10643 5763
rect 11253 5729 11287 5763
rect 11529 5729 11563 5763
rect 11621 5729 11655 5763
rect 12357 5729 12391 5763
rect 13737 5729 13771 5763
rect 14565 5729 14599 5763
rect 16456 5729 16490 5763
rect 16865 5729 16899 5763
rect 19073 5729 19107 5763
rect 20729 5729 20763 5763
rect 21005 5729 21039 5763
rect 21465 5729 21499 5763
rect 21741 5729 21775 5763
rect 22661 5729 22695 5763
rect 24041 5729 24075 5763
rect 26617 5729 26651 5763
rect 26893 5729 26927 5763
rect 27169 5729 27203 5763
rect 27445 5729 27479 5763
rect 27545 5729 27579 5763
rect 28273 5729 28307 5763
rect 1317 5661 1351 5695
rect 1813 5679 1847 5713
rect 2053 5661 2087 5695
rect 3525 5661 3559 5695
rect 4031 5661 4065 5695
rect 4261 5661 4295 5695
rect 7849 5661 7883 5695
rect 8355 5661 8389 5695
rect 9965 5661 9999 5695
rect 12084 5661 12118 5695
rect 13829 5661 13863 5695
rect 14156 5661 14190 5695
rect 14292 5663 14326 5697
rect 16129 5661 16163 5695
rect 16592 5661 16626 5695
rect 18337 5661 18371 5695
rect 18664 5661 18698 5695
rect 18800 5661 18834 5695
rect 21925 5661 21959 5695
rect 22252 5661 22286 5695
rect 22388 5663 22422 5697
rect 24133 5661 24167 5695
rect 24596 5661 24630 5695
rect 24869 5661 24903 5695
rect 28043 5661 28077 5695
rect 6653 5593 6687 5627
rect 21281 5593 21315 5627
rect 26433 5593 26467 5627
rect 3341 5525 3375 5559
rect 5549 5525 5583 5559
rect 6377 5525 6411 5559
rect 6929 5525 6963 5559
rect 7481 5525 7515 5559
rect 10057 5525 10091 5559
rect 10333 5525 10367 5559
rect 11345 5525 11379 5559
rect 15853 5525 15887 5559
rect 18153 5525 18187 5559
rect 20361 5525 20395 5559
rect 21557 5525 21591 5559
rect 26157 5525 26191 5559
rect 26709 5525 26743 5559
rect 26985 5525 27019 5559
rect 27261 5525 27295 5559
rect 2973 5321 3007 5355
rect 13277 5321 13311 5355
rect 15761 5321 15795 5355
rect 20729 5321 20763 5355
rect 25697 5321 25731 5355
rect 29469 5321 29503 5355
rect 3525 5253 3559 5287
rect 8677 5253 8711 5287
rect 23121 5253 23155 5287
rect 1445 5167 1479 5201
rect 1685 5185 1719 5219
rect 4399 5185 4433 5219
rect 6009 5185 6043 5219
rect 6564 5185 6598 5219
rect 6837 5185 6871 5219
rect 9508 5185 9542 5219
rect 9781 5185 9815 5219
rect 11161 5185 11195 5219
rect 11716 5185 11750 5219
rect 14200 5185 14234 5219
rect 16408 5185 16442 5219
rect 19168 5185 19202 5219
rect 21240 5185 21274 5219
rect 21392 5167 21426 5201
rect 21649 5185 21683 5219
rect 24320 5185 24354 5219
rect 26709 5185 26743 5219
rect 27205 5167 27239 5201
rect 949 5117 983 5151
rect 3893 5117 3927 5151
rect 4220 5117 4254 5151
rect 4629 5117 4663 5151
rect 6101 5117 6135 5151
rect 6428 5117 6462 5151
rect 8585 5117 8619 5151
rect 8861 5117 8895 5151
rect 9045 5117 9079 5151
rect 9372 5117 9406 5151
rect 11253 5117 11287 5151
rect 11989 5117 12023 5151
rect 13737 5117 13771 5151
rect 14473 5117 14507 5151
rect 15945 5117 15979 5151
rect 16681 5117 16715 5151
rect 18521 5117 18555 5151
rect 18705 5117 18739 5151
rect 19441 5117 19475 5151
rect 20913 5117 20947 5151
rect 23305 5117 23339 5151
rect 23857 5117 23891 5151
rect 24593 5117 24627 5151
rect 27445 5117 27479 5151
rect 29193 5117 29227 5151
rect 29285 5117 29319 5151
rect 3341 5049 3375 5083
rect 8217 5049 8251 5083
rect 18061 5049 18095 5083
rect 1415 4981 1449 5015
rect 8401 4981 8435 5015
rect 11719 4981 11753 5015
rect 14203 4981 14237 5015
rect 16411 4981 16445 5015
rect 18337 4981 18371 5015
rect 19171 4981 19205 5015
rect 22753 4981 22787 5015
rect 24323 4981 24357 5015
rect 27175 4981 27209 5015
rect 28549 4981 28583 5015
rect 29009 4981 29043 5015
rect 857 4777 891 4811
rect 3157 4777 3191 4811
rect 3991 4777 4025 4811
rect 7941 4777 7975 4811
rect 9143 4777 9177 4811
rect 10701 4777 10735 4811
rect 12087 4777 12121 4811
rect 14295 4777 14329 4811
rect 18153 4777 18187 4811
rect 20361 4777 20395 4811
rect 22483 4777 22517 4811
rect 24225 4777 24259 4811
rect 24777 4777 24811 4811
rect 26617 4777 26651 4811
rect 27261 4777 27295 4811
rect 28279 4777 28313 4811
rect 15945 4709 15979 4743
rect 1041 4641 1075 4675
rect 1460 4641 1494 4675
rect 1869 4641 1903 4675
rect 6244 4641 6278 4675
rect 6653 4641 6687 4675
rect 8309 4641 8343 4675
rect 8585 4641 8619 4675
rect 11161 4641 11195 4675
rect 11529 4641 11563 4675
rect 12357 4641 12391 4675
rect 13737 4641 13771 4675
rect 19073 4641 19107 4675
rect 20729 4641 20763 4675
rect 21005 4641 21039 4675
rect 21465 4641 21499 4675
rect 21741 4641 21775 4675
rect 22017 4641 22051 4675
rect 24409 4641 24443 4675
rect 24685 4641 24719 4675
rect 24961 4641 24995 4675
rect 25237 4641 25271 4675
rect 25513 4641 25547 4675
rect 26433 4641 26467 4675
rect 27077 4641 27111 4675
rect 27813 4641 27847 4675
rect 28549 4641 28583 4675
rect 1133 4573 1167 4607
rect 1639 4573 1673 4607
rect 3525 4573 3559 4607
rect 3988 4573 4022 4607
rect 4261 4573 4295 4607
rect 5917 4573 5951 4607
rect 6423 4573 6457 4607
rect 8677 4573 8711 4607
rect 9183 4573 9217 4607
rect 9413 4573 9447 4607
rect 11621 4573 11655 4607
rect 12127 4573 12161 4607
rect 13829 4573 13863 4607
rect 14292 4575 14326 4609
rect 14565 4573 14599 4607
rect 16129 4573 16163 4607
rect 16456 4573 16490 4607
rect 16635 4573 16669 4607
rect 16865 4573 16899 4607
rect 18337 4573 18371 4607
rect 18664 4573 18698 4607
rect 18816 4591 18850 4625
rect 22523 4573 22557 4607
rect 22753 4573 22787 4607
rect 28276 4573 28310 4607
rect 8125 4505 8159 4539
rect 10977 4505 11011 4539
rect 20545 4505 20579 4539
rect 21281 4505 21315 4539
rect 29653 4505 29687 4539
rect 5549 4437 5583 4471
rect 8401 4437 8435 4471
rect 11345 4437 11379 4471
rect 20821 4437 20855 4471
rect 21557 4437 21591 4471
rect 24041 4437 24075 4471
rect 24501 4437 24535 4471
rect 25053 4437 25087 4471
rect 25329 4437 25363 4471
rect 5733 4233 5767 4267
rect 11897 4233 11931 4267
rect 13277 4233 13311 4267
rect 16221 4233 16255 4267
rect 18245 4165 18279 4199
rect 1445 4079 1479 4113
rect 4215 4097 4249 4131
rect 6380 4097 6414 4131
rect 6653 4097 6687 4131
rect 10336 4097 10370 4131
rect 12265 4097 12299 4131
rect 13921 4097 13955 4131
rect 14693 4079 14727 4113
rect 16901 4079 16935 4113
rect 17141 4097 17175 4131
rect 19441 4097 19475 4131
rect 20456 4097 20490 4131
rect 20729 4097 20763 4131
rect 24041 4097 24075 4131
rect 24504 4097 24538 4131
rect 24777 4097 24811 4131
rect 26712 4097 26746 4131
rect 26985 4097 27019 4131
rect 949 4029 983 4063
rect 1685 4029 1719 4063
rect 3617 4029 3651 4063
rect 3709 4029 3743 4063
rect 4036 4029 4070 4063
rect 4445 4029 4479 4063
rect 5917 4029 5951 4063
rect 6244 4029 6278 4063
rect 8493 4029 8527 4063
rect 9229 4029 9263 4063
rect 9505 4029 9539 4063
rect 9781 4029 9815 4063
rect 9873 4029 9907 4063
rect 10609 4029 10643 4063
rect 12081 4029 12115 4063
rect 12817 4029 12851 4063
rect 13645 4029 13679 4063
rect 14197 4029 14231 4063
rect 14933 4029 14967 4063
rect 16405 4029 16439 4063
rect 19257 4029 19291 4063
rect 19993 4029 20027 4063
rect 22385 4029 22419 4063
rect 23121 4029 23155 4063
rect 23397 4029 23431 4063
rect 26249 4029 26283 4063
rect 13001 3961 13035 3995
rect 18797 3961 18831 3995
rect 22109 3961 22143 3995
rect 22661 3961 22695 3995
rect 1415 3893 1449 3927
rect 2789 3893 2823 3927
rect 3433 3893 3467 3927
rect 7757 3893 7791 3927
rect 8585 3893 8619 3927
rect 9045 3893 9079 3927
rect 9321 3893 9355 3927
rect 9597 3893 9631 3927
rect 10339 3893 10373 3927
rect 12633 3893 12667 3927
rect 14663 3893 14697 3927
rect 16871 3893 16905 3927
rect 18889 3893 18923 3927
rect 20459 3893 20493 3927
rect 22937 3893 22971 3927
rect 23213 3893 23247 3927
rect 24507 3893 24541 3927
rect 26065 3893 26099 3927
rect 26715 3893 26749 3927
rect 28089 3893 28123 3927
rect 857 3689 891 3723
rect 1783 3689 1817 3723
rect 3991 3689 4025 3723
rect 5825 3689 5859 3723
rect 6653 3689 6687 3723
rect 8315 3689 8349 3723
rect 9689 3689 9723 3723
rect 11161 3689 11195 3723
rect 12087 3689 12121 3723
rect 14295 3689 14329 3723
rect 16595 3689 16629 3723
rect 21747 3689 21781 3723
rect 27353 3689 27387 3723
rect 28371 3689 28405 3723
rect 7573 3621 7607 3655
rect 26893 3621 26927 3655
rect 27261 3621 27295 3655
rect 1041 3553 1075 3587
rect 1317 3553 1351 3587
rect 3525 3553 3559 3587
rect 4261 3553 4295 3587
rect 6009 3553 6043 3587
rect 6377 3553 6411 3587
rect 7205 3553 7239 3587
rect 7297 3553 7331 3587
rect 10057 3553 10091 3587
rect 10793 3553 10827 3587
rect 11069 3553 11103 3587
rect 12357 3553 12391 3587
rect 13737 3553 13771 3587
rect 14565 3553 14599 3587
rect 15945 3553 15979 3587
rect 18245 3553 18279 3587
rect 19073 3553 19107 3587
rect 20637 3553 20671 3587
rect 21281 3553 21315 3587
rect 22017 3553 22051 3587
rect 23397 3553 23431 3587
rect 24225 3553 24259 3587
rect 25697 3553 25731 3587
rect 26617 3553 26651 3587
rect 27905 3553 27939 3587
rect 28641 3553 28675 3587
rect 1813 3503 1847 3537
rect 2053 3485 2087 3519
rect 3433 3485 3467 3519
rect 3988 3487 4022 3521
rect 5641 3485 5675 3519
rect 7849 3485 7883 3519
rect 8312 3485 8346 3519
rect 8585 3485 8619 3519
rect 10241 3485 10275 3519
rect 11621 3485 11655 3519
rect 12127 3485 12161 3519
rect 13829 3485 13863 3519
rect 14292 3487 14326 3521
rect 16129 3485 16163 3519
rect 16592 3487 16626 3521
rect 16865 3485 16899 3519
rect 18337 3485 18371 3519
rect 18664 3485 18698 3519
rect 18800 3487 18834 3521
rect 20453 3485 20487 3519
rect 21744 3503 21778 3537
rect 23489 3485 23523 3519
rect 23816 3485 23850 3519
rect 23952 3487 23986 3521
rect 25881 3485 25915 3519
rect 28368 3485 28402 3519
rect 29745 3417 29779 3451
rect 7021 3349 7055 3383
rect 10609 3349 10643 3383
rect 20729 3349 20763 3383
rect 25329 3349 25363 3383
rect 3433 3145 3467 3179
rect 3617 3145 3651 3179
rect 18153 3145 18187 3179
rect 28641 3145 28675 3179
rect 2973 3077 3007 3111
rect 8677 3077 8711 3111
rect 25697 3077 25731 3111
rect 1455 3009 1489 3043
rect 3893 3009 3927 3043
rect 4399 3007 4433 3041
rect 4629 3009 4663 3043
rect 6101 3009 6135 3043
rect 6607 3007 6641 3041
rect 8217 3009 8251 3043
rect 9508 3009 9542 3043
rect 11161 3009 11195 3043
rect 11716 3009 11750 3043
rect 11989 3009 12023 3043
rect 13369 3009 13403 3043
rect 14200 3009 14234 3043
rect 14473 3009 14507 3043
rect 15853 3009 15887 3043
rect 16408 3009 16442 3043
rect 18061 3009 18095 3043
rect 19168 3009 19202 3043
rect 19441 3009 19475 3043
rect 20821 3009 20855 3043
rect 21376 3009 21410 3043
rect 21649 3009 21683 3043
rect 23029 3009 23063 3043
rect 24320 3009 24354 3043
rect 24593 3009 24627 3043
rect 26712 3009 26746 3043
rect 26985 3009 27019 3043
rect 29193 3009 29227 3043
rect 949 2941 983 2975
rect 1685 2941 1719 2975
rect 3801 2941 3835 2975
rect 6837 2941 6871 2975
rect 8493 2941 8527 2975
rect 9045 2941 9079 2975
rect 9781 2941 9815 2975
rect 11253 2941 11287 2975
rect 13737 2941 13771 2975
rect 15945 2941 15979 2975
rect 16681 2941 16715 2975
rect 18337 2941 18371 2975
rect 18705 2941 18739 2975
rect 20913 2941 20947 2975
rect 23213 2941 23247 2975
rect 23857 2941 23891 2975
rect 26249 2941 26283 2975
rect 28457 2941 28491 2975
rect 29009 2941 29043 2975
rect 6009 2873 6043 2907
rect 1415 2805 1449 2839
rect 4359 2805 4393 2839
rect 6567 2805 6601 2839
rect 9511 2805 9545 2839
rect 11719 2805 11753 2839
rect 14203 2805 14237 2839
rect 16411 2805 16445 2839
rect 19171 2805 19205 2839
rect 21379 2805 21413 2839
rect 23305 2805 23339 2839
rect 24323 2805 24357 2839
rect 26715 2805 26749 2839
rect 28089 2805 28123 2839
rect 857 2601 891 2635
rect 1783 2601 1817 2635
rect 3157 2601 3191 2635
rect 6935 2601 6969 2635
rect 9143 2601 9177 2635
rect 11253 2601 11287 2635
rect 12087 2601 12121 2635
rect 14295 2601 14329 2635
rect 16595 2601 16629 2635
rect 21747 2601 21781 2635
rect 26899 2601 26933 2635
rect 28825 2601 28859 2635
rect 29377 2601 29411 2635
rect 6101 2533 6135 2567
rect 20453 2533 20487 2567
rect 23949 2533 23983 2567
rect 1041 2465 1075 2499
rect 1317 2465 1351 2499
rect 3525 2465 3559 2499
rect 4261 2465 4295 2499
rect 5825 2465 5859 2499
rect 6469 2465 6503 2499
rect 7205 2465 7239 2499
rect 8585 2465 8619 2499
rect 9413 2465 9447 2499
rect 11161 2465 11195 2499
rect 15945 2465 15979 2499
rect 18245 2465 18279 2499
rect 20545 2465 20579 2499
rect 21281 2465 21315 2499
rect 23581 2465 23615 2499
rect 24133 2465 24167 2499
rect 24869 2465 24903 2499
rect 27169 2465 27203 2499
rect 28641 2465 28675 2499
rect 28917 2465 28951 2499
rect 29193 2465 29227 2499
rect 1823 2399 1857 2433
rect 2053 2397 2087 2431
rect 3852 2397 3886 2431
rect 3988 2397 4022 2431
rect 6932 2399 6966 2433
rect 8677 2397 8711 2431
rect 9140 2397 9174 2431
rect 11621 2397 11655 2431
rect 12127 2397 12161 2431
rect 12357 2397 12391 2431
rect 13829 2397 13863 2431
rect 14292 2397 14326 2431
rect 14565 2397 14599 2431
rect 16129 2397 16163 2431
rect 16592 2397 16626 2431
rect 16865 2397 16899 2431
rect 18337 2397 18371 2431
rect 18664 2397 18698 2431
rect 18800 2397 18834 2431
rect 19073 2397 19107 2431
rect 20729 2397 20763 2431
rect 21744 2397 21778 2431
rect 22017 2397 22051 2431
rect 24460 2397 24494 2431
rect 24629 2415 24663 2449
rect 26433 2397 26467 2431
rect 26896 2397 26930 2431
rect 29101 2329 29135 2363
rect 5549 2261 5583 2295
rect 10701 2261 10735 2295
rect 13645 2261 13679 2295
rect 23121 2261 23155 2295
rect 25973 2261 26007 2295
rect 28273 2261 28307 2295
rect 2973 2057 3007 2091
rect 5365 2057 5399 2091
rect 7757 2057 7791 2091
rect 8769 2057 8803 2091
rect 13277 2057 13311 2091
rect 18061 2057 18095 2091
rect 23857 2057 23891 2091
rect 26341 2057 26375 2091
rect 28733 2057 28767 2091
rect 3249 1989 3283 2023
rect 18337 1989 18371 2023
rect 23121 1989 23155 2023
rect 29193 1989 29227 2023
rect 949 1921 983 1955
rect 1455 1921 1489 1955
rect 1685 1921 1719 1955
rect 4031 1919 4065 1953
rect 4261 1921 4295 1955
rect 5917 1921 5951 1955
rect 6380 1921 6414 1955
rect 9045 1921 9079 1955
rect 9372 1921 9406 1955
rect 9508 1921 9542 1955
rect 11161 1921 11195 1955
rect 11716 1921 11750 1955
rect 11989 1921 12023 1955
rect 13645 1921 13679 1955
rect 13972 1921 14006 1955
rect 14124 1921 14158 1955
rect 15761 1921 15795 1955
rect 16316 1921 16350 1955
rect 16589 1921 16623 1955
rect 18705 1921 18739 1955
rect 19168 1921 19202 1955
rect 20821 1921 20855 1955
rect 21376 1921 21410 1955
rect 21649 1921 21683 1955
rect 24780 1921 24814 1955
rect 25053 1921 25087 1955
rect 26709 1921 26743 1955
rect 27215 1921 27249 1955
rect 27445 1921 27479 1955
rect 3433 1853 3467 1887
rect 3525 1853 3559 1887
rect 3852 1853 3886 1887
rect 6653 1853 6687 1887
rect 8493 1853 8527 1887
rect 9781 1853 9815 1887
rect 11253 1853 11287 1887
rect 11580 1853 11614 1887
rect 14381 1853 14415 1887
rect 15853 1853 15887 1887
rect 18245 1853 18279 1887
rect 18521 1853 18555 1887
rect 19032 1853 19066 1887
rect 19441 1853 19475 1887
rect 20913 1853 20947 1887
rect 23305 1853 23339 1887
rect 23581 1853 23615 1887
rect 24041 1853 24075 1887
rect 24317 1853 24351 1887
rect 29009 1853 29043 1887
rect 17969 1785 18003 1819
rect 23029 1785 23063 1819
rect 1415 1717 1449 1751
rect 6383 1717 6417 1751
rect 16319 1717 16353 1751
rect 21379 1717 21413 1751
rect 23397 1717 23431 1751
rect 24783 1717 24817 1751
rect 27175 1717 27209 1751
rect 1783 1513 1817 1547
rect 3991 1513 4025 1547
rect 5549 1513 5583 1547
rect 6935 1513 6969 1547
rect 11345 1513 11379 1547
rect 12087 1513 12121 1547
rect 13645 1513 13679 1547
rect 14295 1513 14329 1547
rect 16595 1513 16629 1547
rect 18803 1513 18837 1547
rect 20545 1513 20579 1547
rect 21747 1513 21781 1547
rect 26433 1513 26467 1547
rect 27169 1513 27203 1547
rect 27445 1513 27479 1547
rect 28003 1513 28037 1547
rect 29377 1513 29411 1547
rect 6101 1445 6135 1479
rect 20453 1445 20487 1479
rect 1225 1377 1259 1411
rect 1317 1377 1351 1411
rect 3433 1377 3467 1411
rect 5825 1377 5859 1411
rect 6469 1377 6503 1411
rect 8677 1377 8711 1411
rect 11253 1377 11287 1411
rect 11529 1377 11563 1411
rect 11621 1377 11655 1411
rect 15945 1377 15979 1411
rect 18245 1377 18279 1411
rect 20729 1377 20763 1411
rect 21005 1377 21039 1411
rect 23397 1377 23431 1411
rect 23816 1377 23850 1411
rect 25605 1377 25639 1411
rect 25789 1377 25823 1411
rect 26617 1377 26651 1411
rect 26893 1377 26927 1411
rect 26985 1377 27019 1411
rect 27261 1377 27295 1411
rect 27537 1377 27571 1411
rect 29745 1377 29779 1411
rect 1823 1311 1857 1345
rect 2053 1309 2087 1343
rect 3525 1309 3559 1343
rect 4031 1309 4065 1343
rect 4261 1309 4295 1343
rect 6932 1327 6966 1361
rect 7205 1309 7239 1343
rect 8585 1309 8619 1343
rect 9004 1309 9038 1343
rect 9183 1309 9217 1343
rect 9413 1309 9447 1343
rect 10793 1309 10827 1343
rect 12084 1309 12118 1343
rect 12357 1309 12391 1343
rect 13829 1309 13863 1343
rect 14292 1309 14326 1343
rect 14565 1309 14599 1343
rect 16129 1309 16163 1343
rect 16592 1309 16626 1343
rect 16865 1309 16899 1343
rect 18337 1309 18371 1343
rect 18800 1309 18834 1343
rect 19073 1309 19107 1343
rect 21281 1309 21315 1343
rect 21744 1309 21778 1343
rect 22017 1309 22051 1343
rect 23489 1309 23523 1343
rect 23952 1309 23986 1343
rect 24225 1309 24259 1343
rect 28033 1327 28067 1361
rect 28273 1309 28307 1343
rect 20821 1241 20855 1275
rect 1041 1173 1075 1207
rect 11069 1173 11103 1207
rect 25881 1173 25915 1207
rect 26709 1173 26743 1207
rect 29929 1173 29963 1207
rect 3525 969 3559 1003
rect 3893 969 3927 1003
rect 5181 969 5215 1003
rect 5457 969 5491 1003
rect 8125 969 8159 1003
rect 10977 969 11011 1003
rect 13553 969 13587 1003
rect 16129 969 16163 1003
rect 18705 969 18739 1003
rect 23581 969 23615 1003
rect 25697 969 25731 1003
rect 28549 969 28583 1003
rect 29193 969 29227 1003
rect 29469 969 29503 1003
rect 18245 901 18279 935
rect 21281 901 21315 935
rect 26065 901 26099 935
rect 949 833 983 867
rect 1455 831 1489 865
rect 3065 833 3099 867
rect 6101 833 6135 867
rect 6607 833 6641 867
rect 6837 833 6871 867
rect 8677 833 8711 867
rect 9004 833 9038 867
rect 9140 833 9174 867
rect 9413 833 9447 867
rect 11253 833 11287 867
rect 11759 833 11793 867
rect 14335 833 14369 867
rect 16911 833 16945 867
rect 18981 833 19015 867
rect 19308 833 19342 867
rect 19487 831 19521 865
rect 19717 833 19751 867
rect 21557 833 21591 867
rect 22063 833 22097 867
rect 24320 833 24354 867
rect 24593 833 24627 867
rect 27215 833 27249 867
rect 1685 765 1719 799
rect 5365 765 5399 799
rect 5641 765 5675 799
rect 6009 765 6043 799
rect 8585 765 8619 799
rect 11161 765 11195 799
rect 11989 765 12023 799
rect 13737 765 13771 799
rect 13829 765 13863 799
rect 14156 765 14190 799
rect 14565 765 14599 799
rect 16313 765 16347 799
rect 16405 765 16439 799
rect 16732 765 16766 799
rect 17141 765 17175 799
rect 18889 765 18923 799
rect 21465 765 21499 799
rect 22293 765 22327 799
rect 23857 765 23891 799
rect 26249 765 26283 799
rect 26433 765 26467 799
rect 26709 765 26743 799
rect 27445 765 27479 799
rect 29009 765 29043 799
rect 1415 629 1449 663
rect 4261 629 4295 663
rect 5825 629 5859 663
rect 6567 629 6601 663
rect 8401 629 8435 663
rect 10701 629 10735 663
rect 11719 629 11753 663
rect 13093 629 13127 663
rect 15669 629 15703 663
rect 20821 629 20855 663
rect 22023 629 22057 663
rect 24323 629 24357 663
rect 26617 629 26651 663
rect 27175 629 27209 663
<< metal1 >>
rect 8202 22244 8208 22296
rect 8260 22284 8266 22296
rect 8260 22256 11008 22284
rect 8260 22244 8266 22256
rect 10980 22228 11008 22256
rect 11146 22244 11152 22296
rect 11204 22284 11210 22296
rect 12250 22284 12256 22296
rect 11204 22256 12256 22284
rect 11204 22244 11210 22256
rect 12250 22244 12256 22256
rect 12308 22244 12314 22296
rect 24118 22284 24124 22296
rect 19720 22256 24124 22284
rect 6454 22176 6460 22228
rect 6512 22216 6518 22228
rect 10042 22216 10048 22228
rect 6512 22188 10048 22216
rect 6512 22176 6518 22188
rect 10042 22176 10048 22188
rect 10100 22176 10106 22228
rect 10962 22176 10968 22228
rect 11020 22176 11026 22228
rect 11054 22176 11060 22228
rect 11112 22216 11118 22228
rect 14458 22216 14464 22228
rect 11112 22188 14464 22216
rect 11112 22176 11118 22188
rect 14458 22176 14464 22188
rect 14516 22176 14522 22228
rect 6086 22108 6092 22160
rect 6144 22148 6150 22160
rect 6144 22120 8432 22148
rect 6144 22108 6150 22120
rect 8404 22080 8432 22120
rect 9398 22108 9404 22160
rect 9456 22148 9462 22160
rect 9456 22120 14228 22148
rect 9456 22108 9462 22120
rect 9950 22080 9956 22092
rect 8404 22052 9956 22080
rect 9950 22040 9956 22052
rect 10008 22040 10014 22092
rect 10410 22040 10416 22092
rect 10468 22080 10474 22092
rect 13998 22080 14004 22092
rect 10468 22052 14004 22080
rect 10468 22040 10474 22052
rect 13998 22040 14004 22052
rect 14056 22040 14062 22092
rect 2746 21984 12848 22012
rect 2130 21836 2136 21888
rect 2188 21876 2194 21888
rect 2746 21876 2774 21984
rect 6638 21904 6644 21956
rect 6696 21944 6702 21956
rect 12066 21944 12072 21956
rect 6696 21916 12072 21944
rect 6696 21904 6702 21916
rect 12066 21904 12072 21916
rect 12124 21904 12130 21956
rect 12250 21904 12256 21956
rect 12308 21944 12314 21956
rect 12710 21944 12716 21956
rect 12308 21916 12716 21944
rect 12308 21904 12314 21916
rect 12710 21904 12716 21916
rect 12768 21904 12774 21956
rect 12820 21888 12848 21984
rect 14200 21888 14228 22120
rect 19720 22092 19748 22256
rect 24118 22244 24124 22256
rect 24176 22244 24182 22296
rect 22462 22176 22468 22228
rect 22520 22216 22526 22228
rect 25590 22216 25596 22228
rect 22520 22188 25596 22216
rect 22520 22176 22526 22188
rect 25590 22176 25596 22188
rect 25648 22176 25654 22228
rect 23750 22148 23756 22160
rect 20548 22120 23756 22148
rect 14274 22040 14280 22092
rect 14332 22080 14338 22092
rect 19334 22080 19340 22092
rect 14332 22052 19340 22080
rect 14332 22040 14338 22052
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 19702 22040 19708 22092
rect 19760 22040 19766 22092
rect 19886 22012 19892 22024
rect 16868 21984 19892 22012
rect 16868 21888 16896 21984
rect 19886 21972 19892 21984
rect 19944 21972 19950 22024
rect 20548 22012 20576 22120
rect 23750 22108 23756 22120
rect 23808 22108 23814 22160
rect 21082 22040 21088 22092
rect 21140 22080 21146 22092
rect 27982 22080 27988 22092
rect 21140 22052 27988 22080
rect 21140 22040 21146 22052
rect 27982 22040 27988 22052
rect 28040 22040 28046 22092
rect 20456 21984 20576 22012
rect 20346 21944 20352 21956
rect 18892 21916 20352 21944
rect 18892 21888 18920 21916
rect 20346 21904 20352 21916
rect 20404 21904 20410 21956
rect 2188 21848 2774 21876
rect 2188 21836 2194 21848
rect 6914 21836 6920 21888
rect 6972 21876 6978 21888
rect 10226 21876 10232 21888
rect 6972 21848 10232 21876
rect 6972 21836 6978 21848
rect 10226 21836 10232 21848
rect 10284 21836 10290 21888
rect 10318 21836 10324 21888
rect 10376 21876 10382 21888
rect 12618 21876 12624 21888
rect 10376 21848 12624 21876
rect 10376 21836 10382 21848
rect 12618 21836 12624 21848
rect 12676 21836 12682 21888
rect 12802 21836 12808 21888
rect 12860 21836 12866 21888
rect 14182 21836 14188 21888
rect 14240 21836 14246 21888
rect 16850 21836 16856 21888
rect 16908 21836 16914 21888
rect 18874 21836 18880 21888
rect 18932 21836 18938 21888
rect 19242 21836 19248 21888
rect 19300 21876 19306 21888
rect 20456 21876 20484 21984
rect 22462 21972 22468 22024
rect 22520 22012 22526 22024
rect 25406 22012 25412 22024
rect 22520 21984 25412 22012
rect 22520 21972 22526 21984
rect 25406 21972 25412 21984
rect 25464 21972 25470 22024
rect 21450 21904 21456 21956
rect 21508 21944 21514 21956
rect 23658 21944 23664 21956
rect 21508 21916 23664 21944
rect 21508 21904 21514 21916
rect 23658 21904 23664 21916
rect 23716 21904 23722 21956
rect 23934 21904 23940 21956
rect 23992 21944 23998 21956
rect 31294 21944 31300 21956
rect 23992 21916 31300 21944
rect 23992 21904 23998 21916
rect 31294 21904 31300 21916
rect 31352 21904 31358 21956
rect 19300 21848 20484 21876
rect 19300 21836 19306 21848
rect 20530 21836 20536 21888
rect 20588 21876 20594 21888
rect 23566 21876 23572 21888
rect 20588 21848 23572 21876
rect 20588 21836 20594 21848
rect 23566 21836 23572 21848
rect 23624 21836 23630 21888
rect 24118 21836 24124 21888
rect 24176 21876 24182 21888
rect 25682 21876 25688 21888
rect 24176 21848 25688 21876
rect 24176 21836 24182 21848
rect 25682 21836 25688 21848
rect 25740 21836 25746 21888
rect 552 21786 30912 21808
rect 552 21734 4193 21786
rect 4245 21734 4257 21786
rect 4309 21734 4321 21786
rect 4373 21734 4385 21786
rect 4437 21734 4449 21786
rect 4501 21734 11783 21786
rect 11835 21734 11847 21786
rect 11899 21734 11911 21786
rect 11963 21734 11975 21786
rect 12027 21734 12039 21786
rect 12091 21734 19373 21786
rect 19425 21734 19437 21786
rect 19489 21734 19501 21786
rect 19553 21734 19565 21786
rect 19617 21734 19629 21786
rect 19681 21734 26963 21786
rect 27015 21734 27027 21786
rect 27079 21734 27091 21786
rect 27143 21734 27155 21786
rect 27207 21734 27219 21786
rect 27271 21734 30912 21786
rect 552 21712 30912 21734
rect 2409 21675 2467 21681
rect 2409 21641 2421 21675
rect 2455 21672 2467 21675
rect 2498 21672 2504 21684
rect 2455 21644 2504 21672
rect 2455 21641 2467 21644
rect 2409 21635 2467 21641
rect 2498 21632 2504 21644
rect 2556 21632 2562 21684
rect 2866 21672 2872 21684
rect 2746 21644 2872 21672
rect 2746 21604 2774 21644
rect 2866 21632 2872 21644
rect 2924 21632 2930 21684
rect 6365 21675 6423 21681
rect 2976 21644 6224 21672
rect 952 21576 2774 21604
rect 952 21477 980 21576
rect 2976 21536 3004 21644
rect 5445 21607 5503 21613
rect 5445 21573 5457 21607
rect 5491 21604 5503 21607
rect 5491 21576 6040 21604
rect 5491 21573 5503 21576
rect 5445 21567 5503 21573
rect 2700 21508 3004 21536
rect 937 21471 995 21477
rect 937 21437 949 21471
rect 983 21437 995 21471
rect 937 21431 995 21437
rect 2130 21428 2136 21480
rect 2188 21428 2194 21480
rect 2700 21477 2728 21508
rect 3050 21496 3056 21548
rect 3108 21536 3114 21548
rect 3700 21539 3758 21545
rect 3700 21536 3712 21539
rect 3108 21508 3712 21536
rect 3108 21496 3114 21508
rect 3700 21505 3712 21508
rect 3746 21505 3758 21539
rect 3700 21499 3758 21505
rect 3896 21508 5948 21536
rect 2685 21471 2743 21477
rect 2685 21437 2697 21471
rect 2731 21437 2743 21471
rect 3234 21468 3240 21480
rect 2685 21431 2743 21437
rect 2884 21440 3240 21468
rect 1213 21403 1271 21409
rect 1213 21369 1225 21403
rect 1259 21400 1271 21403
rect 1394 21400 1400 21412
rect 1259 21372 1400 21400
rect 1259 21369 1271 21372
rect 1213 21363 1271 21369
rect 1394 21360 1400 21372
rect 1452 21360 1458 21412
rect 1581 21403 1639 21409
rect 1581 21369 1593 21403
rect 1627 21400 1639 21403
rect 2774 21400 2780 21412
rect 1627 21372 2780 21400
rect 1627 21369 1639 21372
rect 1581 21363 1639 21369
rect 2774 21360 2780 21372
rect 2832 21360 2838 21412
rect 1486 21292 1492 21344
rect 1544 21332 1550 21344
rect 1857 21335 1915 21341
rect 1857 21332 1869 21335
rect 1544 21304 1869 21332
rect 1544 21292 1550 21304
rect 1857 21301 1869 21304
rect 1903 21332 1915 21335
rect 2884 21332 2912 21440
rect 3234 21428 3240 21440
rect 3292 21428 3298 21480
rect 3896 21468 3924 21508
rect 3344 21440 3924 21468
rect 3053 21403 3111 21409
rect 3053 21369 3065 21403
rect 3099 21400 3111 21403
rect 3344 21400 3372 21440
rect 3970 21428 3976 21480
rect 4028 21428 4034 21480
rect 5626 21428 5632 21480
rect 5684 21428 5690 21480
rect 3099 21372 3372 21400
rect 3099 21369 3111 21372
rect 3053 21363 3111 21369
rect 1903 21304 2912 21332
rect 1903 21301 1915 21304
rect 1857 21295 1915 21301
rect 3694 21292 3700 21344
rect 3752 21341 3758 21344
rect 3752 21332 3761 21341
rect 3752 21304 3797 21332
rect 3752 21295 3761 21304
rect 3752 21292 3758 21295
rect 5074 21292 5080 21344
rect 5132 21292 5138 21344
rect 5920 21332 5948 21508
rect 6012 21400 6040 21576
rect 6086 21564 6092 21616
rect 6144 21564 6150 21616
rect 6104 21477 6132 21564
rect 6196 21536 6224 21644
rect 6365 21641 6377 21675
rect 6411 21672 6423 21675
rect 6454 21672 6460 21684
rect 6411 21644 6460 21672
rect 6411 21641 6423 21644
rect 6365 21635 6423 21641
rect 6454 21632 6460 21644
rect 6512 21632 6518 21684
rect 6914 21632 6920 21684
rect 6972 21632 6978 21684
rect 9398 21672 9404 21684
rect 7116 21644 9404 21672
rect 6914 21536 6920 21548
rect 6196 21508 6920 21536
rect 6914 21496 6920 21508
rect 6972 21496 6978 21548
rect 7116 21545 7144 21644
rect 8202 21564 8208 21616
rect 8260 21564 8266 21616
rect 8570 21604 8576 21616
rect 8312 21576 8576 21604
rect 7101 21539 7159 21545
rect 7101 21505 7113 21539
rect 7147 21505 7159 21539
rect 8312 21536 8340 21576
rect 8570 21564 8576 21576
rect 8628 21564 8634 21616
rect 8680 21545 8708 21644
rect 9398 21632 9404 21644
rect 9456 21632 9462 21684
rect 9953 21675 10011 21681
rect 9953 21641 9965 21675
rect 9999 21672 10011 21675
rect 9999 21644 12664 21672
rect 9999 21641 10011 21644
rect 9953 21635 10011 21641
rect 10318 21564 10324 21616
rect 10376 21564 10382 21616
rect 7101 21499 7159 21505
rect 7944 21508 8340 21536
rect 8665 21539 8723 21545
rect 6089 21471 6147 21477
rect 6089 21437 6101 21471
rect 6135 21437 6147 21471
rect 7282 21468 7288 21480
rect 6089 21431 6147 21437
rect 6564 21440 7288 21468
rect 6564 21400 6592 21440
rect 7282 21428 7288 21440
rect 7340 21428 7346 21480
rect 7377 21471 7435 21477
rect 7377 21437 7389 21471
rect 7423 21468 7435 21471
rect 7944 21468 7972 21508
rect 8665 21505 8677 21539
rect 8711 21505 8723 21539
rect 8665 21499 8723 21505
rect 11422 21496 11428 21548
rect 11480 21536 11486 21548
rect 12636 21536 12664 21644
rect 12710 21632 12716 21684
rect 12768 21632 12774 21684
rect 12802 21632 12808 21684
rect 12860 21632 12866 21684
rect 14550 21632 14556 21684
rect 14608 21672 14614 21684
rect 17126 21672 17132 21684
rect 14608 21644 17132 21672
rect 14608 21632 14614 21644
rect 17126 21632 17132 21644
rect 17184 21632 17190 21684
rect 19153 21675 19211 21681
rect 19153 21641 19165 21675
rect 19199 21672 19211 21675
rect 20993 21675 21051 21681
rect 19199 21644 20668 21672
rect 19199 21641 19211 21644
rect 19153 21635 19211 21641
rect 12728 21604 12756 21632
rect 13173 21607 13231 21613
rect 13173 21604 13185 21607
rect 12728 21576 13185 21604
rect 13173 21573 13185 21576
rect 13219 21573 13231 21607
rect 13173 21567 13231 21573
rect 18417 21607 18475 21613
rect 18417 21573 18429 21607
rect 18463 21604 18475 21607
rect 19058 21604 19064 21616
rect 18463 21576 19064 21604
rect 18463 21573 18475 21576
rect 18417 21567 18475 21573
rect 19058 21564 19064 21576
rect 19116 21564 19122 21616
rect 20640 21604 20668 21644
rect 20993 21641 21005 21675
rect 21039 21672 21051 21675
rect 21082 21672 21088 21684
rect 21039 21644 21088 21672
rect 21039 21641 21051 21644
rect 20993 21635 21051 21641
rect 21082 21632 21088 21644
rect 21140 21632 21146 21684
rect 22370 21672 22376 21684
rect 21192 21644 22376 21672
rect 21192 21604 21220 21644
rect 22370 21632 22376 21644
rect 22428 21632 22434 21684
rect 24504 21644 28396 21672
rect 23934 21604 23940 21616
rect 20640 21576 21220 21604
rect 23676 21576 23940 21604
rect 13814 21536 13820 21548
rect 11480 21508 11525 21536
rect 12636 21508 13820 21536
rect 11480 21496 11486 21508
rect 13814 21496 13820 21508
rect 13872 21496 13878 21548
rect 14200 21508 16804 21536
rect 7423 21440 7972 21468
rect 7423 21437 7435 21440
rect 7377 21431 7435 21437
rect 8570 21428 8576 21480
rect 8628 21428 8634 21480
rect 8846 21428 8852 21480
rect 8904 21468 8910 21480
rect 8941 21471 8999 21477
rect 8941 21468 8953 21471
rect 8904 21440 8953 21468
rect 8904 21428 8910 21440
rect 8941 21437 8953 21440
rect 8987 21468 8999 21471
rect 10410 21468 10416 21480
rect 8987 21440 10416 21468
rect 8987 21437 8999 21440
rect 8941 21431 8999 21437
rect 10410 21428 10416 21440
rect 10468 21428 10474 21480
rect 10505 21471 10563 21477
rect 10505 21437 10517 21471
rect 10551 21468 10563 21471
rect 10686 21468 10692 21480
rect 10551 21440 10692 21468
rect 10551 21437 10563 21440
rect 10505 21431 10563 21437
rect 10686 21428 10692 21440
rect 10744 21428 10750 21480
rect 10778 21428 10784 21480
rect 10836 21428 10842 21480
rect 10870 21428 10876 21480
rect 10928 21468 10934 21480
rect 10965 21471 11023 21477
rect 10965 21468 10977 21471
rect 10928 21440 10977 21468
rect 10928 21428 10934 21440
rect 10965 21437 10977 21440
rect 11011 21437 11023 21471
rect 10965 21431 11023 21437
rect 11054 21428 11060 21480
rect 11112 21428 11118 21480
rect 11238 21428 11244 21480
rect 11296 21477 11302 21480
rect 11296 21471 11350 21477
rect 11296 21437 11304 21471
rect 11338 21437 11350 21471
rect 11296 21431 11350 21437
rect 11296 21428 11302 21431
rect 11698 21428 11704 21480
rect 11756 21428 11762 21480
rect 13354 21428 13360 21480
rect 13412 21428 13418 21480
rect 13633 21471 13691 21477
rect 13633 21437 13645 21471
rect 13679 21468 13691 21471
rect 14200 21468 14228 21508
rect 13679 21440 14228 21468
rect 13679 21437 13691 21440
rect 13633 21431 13691 21437
rect 14274 21428 14280 21480
rect 14332 21428 14338 21480
rect 14550 21428 14556 21480
rect 14608 21428 14614 21480
rect 14642 21428 14648 21480
rect 14700 21468 14706 21480
rect 16301 21471 16359 21477
rect 16301 21468 16313 21471
rect 14700 21440 16313 21468
rect 14700 21428 14706 21440
rect 16301 21437 16313 21440
rect 16347 21437 16359 21471
rect 16301 21431 16359 21437
rect 16669 21471 16727 21477
rect 16669 21437 16681 21471
rect 16715 21437 16727 21471
rect 16776 21468 16804 21508
rect 16850 21496 16856 21548
rect 16908 21496 16914 21548
rect 17129 21539 17187 21545
rect 17129 21505 17141 21539
rect 17175 21536 17187 21539
rect 19242 21536 19248 21548
rect 17175 21508 19248 21536
rect 17175 21505 17187 21508
rect 17129 21499 17187 21505
rect 19242 21496 19248 21508
rect 19300 21496 19306 21548
rect 19429 21539 19487 21545
rect 19429 21505 19441 21539
rect 19475 21536 19487 21539
rect 19610 21536 19616 21548
rect 19475 21508 19616 21536
rect 19475 21505 19487 21508
rect 19429 21499 19487 21505
rect 19610 21496 19616 21508
rect 19668 21496 19674 21548
rect 19705 21539 19763 21545
rect 19705 21505 19717 21539
rect 19751 21536 19763 21539
rect 19751 21508 21404 21536
rect 19751 21505 19763 21508
rect 19705 21499 19763 21505
rect 18693 21471 18751 21477
rect 18693 21468 18705 21471
rect 16776 21440 18705 21468
rect 16669 21431 16727 21437
rect 18693 21437 18705 21440
rect 18739 21468 18751 21471
rect 18782 21468 18788 21480
rect 18739 21440 18788 21468
rect 18739 21437 18751 21440
rect 18693 21431 18751 21437
rect 6012 21372 6592 21400
rect 6638 21360 6644 21412
rect 6696 21360 6702 21412
rect 8021 21403 8079 21409
rect 8021 21369 8033 21403
rect 8067 21400 8079 21403
rect 8478 21400 8484 21412
rect 8067 21372 8484 21400
rect 8067 21369 8079 21372
rect 8021 21363 8079 21369
rect 8478 21360 8484 21372
rect 8536 21360 8542 21412
rect 9306 21360 9312 21412
rect 9364 21400 9370 21412
rect 9769 21403 9827 21409
rect 9769 21400 9781 21403
rect 9364 21372 9781 21400
rect 9364 21360 9370 21372
rect 9769 21369 9781 21372
rect 9815 21400 9827 21403
rect 11072 21400 11100 21428
rect 9815 21372 11100 21400
rect 15933 21403 15991 21409
rect 9815 21369 9827 21372
rect 9769 21363 9827 21369
rect 15933 21369 15945 21403
rect 15979 21400 15991 21403
rect 16390 21400 16396 21412
rect 15979 21372 16396 21400
rect 15979 21369 15991 21372
rect 15933 21363 15991 21369
rect 16390 21360 16396 21372
rect 16448 21360 16454 21412
rect 8294 21332 8300 21344
rect 5920 21304 8300 21332
rect 8294 21292 8300 21304
rect 8352 21292 8358 21344
rect 8389 21335 8447 21341
rect 8389 21301 8401 21335
rect 8435 21332 8447 21335
rect 8662 21332 8668 21344
rect 8435 21304 8668 21332
rect 8435 21301 8447 21304
rect 8389 21295 8447 21301
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 10597 21335 10655 21341
rect 10597 21301 10609 21335
rect 10643 21332 10655 21335
rect 11330 21332 11336 21344
rect 10643 21304 11336 21332
rect 10643 21301 10655 21304
rect 10597 21295 10655 21301
rect 11330 21292 11336 21304
rect 11388 21292 11394 21344
rect 11606 21292 11612 21344
rect 11664 21332 11670 21344
rect 12342 21332 12348 21344
rect 11664 21304 12348 21332
rect 11664 21292 11670 21304
rect 12342 21292 12348 21304
rect 12400 21292 12406 21344
rect 13722 21292 13728 21344
rect 13780 21292 13786 21344
rect 16114 21292 16120 21344
rect 16172 21292 16178 21344
rect 16684 21332 16712 21431
rect 18782 21428 18788 21440
rect 18840 21428 18846 21480
rect 18874 21428 18880 21480
rect 18932 21428 18938 21480
rect 19061 21471 19119 21477
rect 19061 21437 19073 21471
rect 19107 21468 19119 21471
rect 19337 21471 19395 21477
rect 19337 21468 19349 21471
rect 19107 21440 19349 21468
rect 19107 21437 19119 21440
rect 19061 21431 19119 21437
rect 19337 21437 19349 21440
rect 19383 21437 19395 21471
rect 20714 21468 20720 21480
rect 19337 21431 19395 21437
rect 19444 21440 20720 21468
rect 16758 21360 16764 21412
rect 16816 21360 16822 21412
rect 19444 21400 19472 21440
rect 20714 21428 20720 21440
rect 20772 21428 20778 21480
rect 21269 21471 21327 21477
rect 21269 21437 21281 21471
rect 21315 21437 21327 21471
rect 21269 21431 21327 21437
rect 18892 21372 19472 21400
rect 18892 21332 18920 21372
rect 21284 21344 21312 21431
rect 16684 21304 18920 21332
rect 18966 21292 18972 21344
rect 19024 21332 19030 21344
rect 20530 21332 20536 21344
rect 19024 21304 20536 21332
rect 19024 21292 19030 21304
rect 20530 21292 20536 21304
rect 20588 21292 20594 21344
rect 21266 21292 21272 21344
rect 21324 21292 21330 21344
rect 21376 21332 21404 21508
rect 21450 21496 21456 21548
rect 21508 21496 21514 21548
rect 21913 21539 21971 21545
rect 21913 21505 21925 21539
rect 21959 21536 21971 21539
rect 22002 21536 22008 21548
rect 21959 21508 22008 21536
rect 21959 21505 21971 21508
rect 21913 21499 21971 21505
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 22462 21496 22468 21548
rect 22520 21496 22526 21548
rect 22186 21428 22192 21480
rect 22244 21428 22250 21480
rect 22278 21428 22284 21480
rect 22336 21477 22342 21480
rect 22336 21471 22364 21477
rect 22352 21437 22364 21471
rect 22336 21431 22364 21437
rect 22336 21428 22342 21431
rect 23198 21428 23204 21480
rect 23256 21428 23262 21480
rect 23385 21471 23443 21477
rect 23385 21437 23397 21471
rect 23431 21437 23443 21471
rect 23385 21431 23443 21437
rect 23400 21400 23428 21431
rect 23566 21428 23572 21480
rect 23624 21428 23630 21480
rect 23676 21477 23704 21576
rect 23934 21564 23940 21576
rect 23992 21564 23998 21616
rect 24504 21548 24532 21644
rect 25498 21564 25504 21616
rect 25556 21604 25562 21616
rect 25685 21607 25743 21613
rect 25685 21604 25697 21607
rect 25556 21576 25697 21604
rect 25556 21564 25562 21576
rect 25685 21573 25697 21576
rect 25731 21573 25743 21607
rect 25685 21567 25743 21573
rect 28368 21548 28396 21644
rect 28994 21564 29000 21616
rect 29052 21604 29058 21616
rect 30009 21607 30067 21613
rect 30009 21604 30021 21607
rect 29052 21576 30021 21604
rect 29052 21564 29058 21576
rect 30009 21573 30021 21576
rect 30055 21573 30067 21607
rect 30009 21567 30067 21573
rect 23845 21539 23903 21545
rect 23845 21505 23857 21539
rect 23891 21536 23903 21539
rect 23891 21508 23983 21536
rect 23891 21505 23903 21508
rect 23845 21499 23903 21505
rect 23955 21480 23983 21508
rect 24486 21496 24492 21548
rect 24544 21496 24550 21548
rect 24578 21496 24584 21548
rect 24636 21536 24642 21548
rect 24882 21539 24940 21545
rect 24882 21536 24894 21539
rect 24636 21508 24894 21536
rect 24636 21496 24642 21508
rect 24882 21505 24894 21508
rect 24928 21505 24940 21539
rect 24882 21499 24940 21505
rect 25041 21539 25099 21545
rect 25041 21505 25053 21539
rect 25087 21536 25099 21539
rect 25406 21536 25412 21548
rect 25087 21508 25412 21536
rect 25087 21505 25099 21508
rect 25041 21499 25099 21505
rect 25406 21496 25412 21508
rect 25464 21496 25470 21548
rect 25774 21496 25780 21548
rect 25832 21536 25838 21548
rect 25832 21508 28304 21536
rect 25832 21496 25838 21508
rect 23661 21471 23719 21477
rect 23661 21437 23673 21471
rect 23707 21437 23719 21471
rect 23661 21431 23719 21437
rect 23934 21428 23940 21480
rect 23992 21428 23998 21480
rect 24029 21471 24087 21477
rect 24029 21437 24041 21471
rect 24075 21437 24087 21471
rect 24029 21431 24087 21437
rect 22940 21372 23428 21400
rect 22940 21344 22968 21372
rect 22738 21332 22744 21344
rect 21376 21304 22744 21332
rect 22738 21292 22744 21304
rect 22796 21292 22802 21344
rect 22922 21292 22928 21344
rect 22980 21292 22986 21344
rect 23014 21292 23020 21344
rect 23072 21332 23078 21344
rect 23109 21335 23167 21341
rect 23109 21332 23121 21335
rect 23072 21304 23121 21332
rect 23072 21292 23078 21304
rect 23109 21301 23121 21304
rect 23155 21301 23167 21335
rect 24044 21332 24072 21431
rect 24762 21428 24768 21480
rect 24820 21428 24826 21480
rect 25682 21428 25688 21480
rect 25740 21468 25746 21480
rect 26421 21471 26479 21477
rect 26421 21468 26433 21471
rect 25740 21440 26433 21468
rect 25740 21428 25746 21440
rect 26421 21437 26433 21440
rect 26467 21437 26479 21471
rect 26421 21431 26479 21437
rect 26697 21471 26755 21477
rect 26697 21437 26709 21471
rect 26743 21468 26755 21471
rect 27798 21468 27804 21480
rect 26743 21440 27804 21468
rect 26743 21437 26755 21440
rect 26697 21431 26755 21437
rect 27798 21428 27804 21440
rect 27856 21428 27862 21480
rect 28276 21477 28304 21508
rect 28350 21496 28356 21548
rect 28408 21496 28414 21548
rect 28261 21471 28319 21477
rect 28261 21437 28273 21471
rect 28307 21437 28319 21471
rect 29457 21471 29515 21477
rect 29457 21468 29469 21471
rect 28261 21431 28319 21437
rect 28368 21440 29469 21468
rect 25869 21403 25927 21409
rect 25869 21369 25881 21403
rect 25915 21400 25927 21403
rect 28074 21400 28080 21412
rect 25915 21372 26464 21400
rect 25915 21369 25927 21372
rect 25869 21363 25927 21369
rect 25038 21332 25044 21344
rect 24044 21304 25044 21332
rect 23109 21295 23167 21301
rect 25038 21292 25044 21304
rect 25096 21292 25102 21344
rect 25682 21292 25688 21344
rect 25740 21332 25746 21344
rect 25961 21335 26019 21341
rect 25961 21332 25973 21335
rect 25740 21304 25973 21332
rect 25740 21292 25746 21304
rect 25961 21301 25973 21304
rect 26007 21301 26019 21335
rect 26436 21332 26464 21372
rect 27356 21372 28080 21400
rect 27356 21332 27384 21372
rect 28074 21360 28080 21372
rect 28132 21400 28138 21412
rect 28368 21400 28396 21440
rect 29457 21437 29469 21440
rect 29503 21437 29515 21471
rect 29457 21431 29515 21437
rect 29917 21471 29975 21477
rect 29917 21437 29929 21471
rect 29963 21437 29975 21471
rect 29917 21431 29975 21437
rect 30193 21471 30251 21477
rect 30193 21437 30205 21471
rect 30239 21468 30251 21471
rect 30374 21468 30380 21480
rect 30239 21440 30380 21468
rect 30239 21437 30251 21440
rect 30193 21431 30251 21437
rect 28132 21372 28396 21400
rect 29089 21403 29147 21409
rect 28132 21360 28138 21372
rect 29089 21369 29101 21403
rect 29135 21369 29147 21403
rect 29932 21400 29960 21431
rect 30374 21428 30380 21440
rect 30432 21428 30438 21480
rect 30558 21428 30564 21480
rect 30616 21428 30622 21480
rect 30282 21400 30288 21412
rect 29932 21372 30288 21400
rect 29089 21363 29147 21369
rect 26436 21304 27384 21332
rect 25961 21295 26019 21301
rect 27430 21292 27436 21344
rect 27488 21332 27494 21344
rect 27801 21335 27859 21341
rect 27801 21332 27813 21335
rect 27488 21304 27813 21332
rect 27488 21292 27494 21304
rect 27801 21301 27813 21304
rect 27847 21301 27859 21335
rect 27801 21295 27859 21301
rect 28353 21335 28411 21341
rect 28353 21301 28365 21335
rect 28399 21332 28411 21335
rect 28442 21332 28448 21344
rect 28399 21304 28448 21332
rect 28399 21301 28411 21304
rect 28353 21295 28411 21301
rect 28442 21292 28448 21304
rect 28500 21332 28506 21344
rect 29104 21332 29132 21363
rect 30282 21360 30288 21372
rect 30340 21360 30346 21412
rect 28500 21304 29132 21332
rect 28500 21292 28506 21304
rect 29730 21292 29736 21344
rect 29788 21292 29794 21344
rect 30098 21292 30104 21344
rect 30156 21332 30162 21344
rect 30377 21335 30435 21341
rect 30377 21332 30389 21335
rect 30156 21304 30389 21332
rect 30156 21292 30162 21304
rect 30377 21301 30389 21304
rect 30423 21301 30435 21335
rect 30377 21295 30435 21301
rect 552 21242 31072 21264
rect 552 21190 7988 21242
rect 8040 21190 8052 21242
rect 8104 21190 8116 21242
rect 8168 21190 8180 21242
rect 8232 21190 8244 21242
rect 8296 21190 15578 21242
rect 15630 21190 15642 21242
rect 15694 21190 15706 21242
rect 15758 21190 15770 21242
rect 15822 21190 15834 21242
rect 15886 21190 23168 21242
rect 23220 21190 23232 21242
rect 23284 21190 23296 21242
rect 23348 21190 23360 21242
rect 23412 21190 23424 21242
rect 23476 21190 30758 21242
rect 30810 21190 30822 21242
rect 30874 21190 30886 21242
rect 30938 21190 30950 21242
rect 31002 21190 31014 21242
rect 31066 21190 31072 21242
rect 552 21168 31072 21190
rect 842 21088 848 21140
rect 900 21088 906 21140
rect 1587 21131 1645 21137
rect 1587 21097 1599 21131
rect 1633 21128 1645 21131
rect 3694 21128 3700 21140
rect 1633 21100 3700 21128
rect 1633 21097 1645 21100
rect 1587 21091 1645 21097
rect 3694 21088 3700 21100
rect 3752 21088 3758 21140
rect 6086 21088 6092 21140
rect 6144 21128 6150 21140
rect 6279 21131 6337 21137
rect 6279 21128 6291 21131
rect 6144 21100 6291 21128
rect 6144 21088 6150 21100
rect 6279 21097 6291 21100
rect 6325 21097 6337 21131
rect 6279 21091 6337 21097
rect 6638 21088 6644 21140
rect 6696 21128 6702 21140
rect 9861 21131 9919 21137
rect 9861 21128 9873 21131
rect 6696 21100 9873 21128
rect 6696 21088 6702 21100
rect 9861 21097 9873 21100
rect 9907 21097 9919 21131
rect 12989 21131 13047 21137
rect 12989 21128 13001 21131
rect 9861 21091 9919 21097
rect 10428 21100 13001 21128
rect 5902 21060 5908 21072
rect 5276 21032 5908 21060
rect 1029 20995 1087 21001
rect 1029 20961 1041 20995
rect 1075 20992 1087 20995
rect 5276 20992 5304 21032
rect 5902 21020 5908 21032
rect 5960 21020 5966 21072
rect 7834 21020 7840 21072
rect 7892 21060 7898 21072
rect 10428 21069 10456 21100
rect 12989 21097 13001 21100
rect 13035 21097 13047 21131
rect 16114 21128 16120 21140
rect 12989 21091 13047 21097
rect 13372 21100 16120 21128
rect 10413 21063 10471 21069
rect 7892 21032 8156 21060
rect 7892 21020 7898 21032
rect 1075 20964 5304 20992
rect 5445 20995 5503 21001
rect 1075 20961 1087 20964
rect 1029 20955 1087 20961
rect 5445 20961 5457 20995
rect 5491 20992 5503 20995
rect 5491 20964 6316 20992
rect 5491 20961 5503 20964
rect 5445 20955 5503 20961
rect 1121 20927 1179 20933
rect 1121 20893 1133 20927
rect 1167 20924 1179 20927
rect 1486 20924 1492 20936
rect 1167 20896 1492 20924
rect 1167 20893 1179 20896
rect 1121 20887 1179 20893
rect 1486 20884 1492 20896
rect 1544 20884 1550 20936
rect 1627 20927 1685 20933
rect 1627 20893 1639 20927
rect 1673 20924 1685 20927
rect 1762 20924 1768 20936
rect 1673 20896 1768 20924
rect 1673 20893 1685 20896
rect 1627 20887 1685 20893
rect 1762 20884 1768 20896
rect 1820 20884 1826 20936
rect 1854 20884 1860 20936
rect 1912 20884 1918 20936
rect 3234 20884 3240 20936
rect 3292 20924 3298 20936
rect 3329 20927 3387 20933
rect 3329 20924 3341 20927
rect 3292 20896 3341 20924
rect 3292 20884 3298 20896
rect 3329 20893 3341 20896
rect 3375 20924 3387 20927
rect 3510 20924 3516 20936
rect 3375 20896 3516 20924
rect 3375 20893 3387 20896
rect 3329 20887 3387 20893
rect 3510 20884 3516 20896
rect 3568 20884 3574 20936
rect 3694 20933 3700 20936
rect 3656 20927 3700 20933
rect 3656 20893 3668 20927
rect 3656 20887 3700 20893
rect 3694 20884 3700 20887
rect 3752 20884 3758 20936
rect 3786 20884 3792 20936
rect 3844 20884 3850 20936
rect 4062 20884 4068 20936
rect 4120 20884 4126 20936
rect 5810 20884 5816 20936
rect 5868 20884 5874 20936
rect 6288 20933 6316 20964
rect 7742 20952 7748 21004
rect 7800 20992 7806 21004
rect 8021 20995 8079 21001
rect 8021 20992 8033 20995
rect 7800 20964 8033 20992
rect 7800 20952 7806 20964
rect 8021 20961 8033 20964
rect 8067 20961 8079 20995
rect 8128 20992 8156 21032
rect 10413 21029 10425 21063
rect 10459 21029 10471 21063
rect 10413 21023 10471 21029
rect 10781 21063 10839 21069
rect 10781 21029 10793 21063
rect 10827 21060 10839 21063
rect 10962 21060 10968 21072
rect 10827 21032 10968 21060
rect 10827 21029 10839 21032
rect 10781 21023 10839 21029
rect 10962 21020 10968 21032
rect 11020 21020 11026 21072
rect 8404 20992 8527 20996
rect 8128 20968 8527 20992
rect 8128 20964 8432 20968
rect 8021 20955 8079 20961
rect 8499 20951 8527 20968
rect 8662 20952 8668 21004
rect 8720 20992 8726 21004
rect 8720 20964 10456 20992
rect 8720 20952 8726 20964
rect 8499 20945 8558 20951
rect 6276 20927 6334 20933
rect 6276 20893 6288 20927
rect 6322 20893 6334 20927
rect 6276 20887 6334 20893
rect 6546 20884 6552 20936
rect 6604 20884 6610 20936
rect 8348 20927 8406 20933
rect 8348 20924 8360 20927
rect 7760 20896 8360 20924
rect 3145 20791 3203 20797
rect 3145 20757 3157 20791
rect 3191 20788 3203 20791
rect 5534 20788 5540 20800
rect 3191 20760 5540 20788
rect 3191 20757 3203 20760
rect 3145 20751 3203 20757
rect 5534 20748 5540 20760
rect 5592 20748 5598 20800
rect 6454 20748 6460 20800
rect 6512 20788 6518 20800
rect 7650 20788 7656 20800
rect 6512 20760 7656 20788
rect 6512 20748 6518 20760
rect 7650 20748 7656 20760
rect 7708 20788 7714 20800
rect 7760 20788 7788 20896
rect 8348 20893 8360 20896
rect 8394 20893 8406 20927
rect 8499 20914 8512 20945
rect 8500 20911 8512 20914
rect 8546 20911 8558 20945
rect 8500 20905 8558 20911
rect 8348 20887 8406 20893
rect 8754 20884 8760 20936
rect 8812 20884 8818 20936
rect 8846 20884 8852 20936
rect 8904 20924 8910 20936
rect 10428 20924 10456 20964
rect 10502 20952 10508 21004
rect 10560 20992 10566 21004
rect 11885 20995 11943 21001
rect 11491 20992 11655 20995
rect 10560 20967 11655 20992
rect 10560 20964 11519 20967
rect 10560 20952 10566 20964
rect 11054 20924 11060 20936
rect 8904 20896 10364 20924
rect 10428 20896 11060 20924
rect 8904 20884 8910 20896
rect 7708 20760 7788 20788
rect 7837 20791 7895 20797
rect 7708 20748 7714 20760
rect 7837 20757 7849 20791
rect 7883 20788 7895 20791
rect 8938 20788 8944 20800
rect 7883 20760 8944 20788
rect 7883 20757 7895 20760
rect 7837 20751 7895 20757
rect 8938 20748 8944 20760
rect 8996 20748 9002 20800
rect 10336 20788 10364 20896
rect 11054 20884 11060 20896
rect 11112 20884 11118 20936
rect 11514 20933 11520 20936
rect 11149 20927 11207 20933
rect 11149 20893 11161 20927
rect 11195 20893 11207 20927
rect 11149 20887 11207 20893
rect 11476 20927 11520 20933
rect 11476 20893 11488 20927
rect 11476 20887 11520 20893
rect 10870 20816 10876 20868
rect 10928 20856 10934 20868
rect 11164 20856 11192 20887
rect 11514 20884 11520 20887
rect 11572 20884 11578 20936
rect 11627 20935 11655 20967
rect 11885 20961 11897 20995
rect 11931 20992 11943 20995
rect 13372 20992 13400 21100
rect 16114 21088 16120 21100
rect 16172 21088 16178 21140
rect 17954 21088 17960 21140
rect 18012 21128 18018 21140
rect 18785 21131 18843 21137
rect 18785 21128 18797 21131
rect 18012 21100 18797 21128
rect 18012 21088 18018 21100
rect 18785 21097 18797 21100
rect 18831 21097 18843 21131
rect 18785 21091 18843 21097
rect 20809 21131 20867 21137
rect 20809 21097 20821 21131
rect 20855 21128 20867 21131
rect 21266 21128 21272 21140
rect 20855 21100 21272 21128
rect 20855 21097 20867 21100
rect 20809 21091 20867 21097
rect 21266 21088 21272 21100
rect 21324 21088 21330 21140
rect 22186 21088 22192 21140
rect 22244 21128 22250 21140
rect 23109 21131 23167 21137
rect 23109 21128 23121 21131
rect 22244 21100 23121 21128
rect 22244 21088 22250 21100
rect 23109 21097 23121 21100
rect 23155 21097 23167 21131
rect 27801 21131 27859 21137
rect 27801 21128 27813 21131
rect 23109 21091 23167 21097
rect 23216 21100 27813 21128
rect 13998 21020 14004 21072
rect 14056 21020 14062 21072
rect 14182 21020 14188 21072
rect 14240 21060 14246 21072
rect 15562 21060 15568 21072
rect 14240 21032 15568 21060
rect 14240 21020 14246 21032
rect 15562 21020 15568 21032
rect 15620 21020 15626 21072
rect 15657 21063 15715 21069
rect 15657 21029 15669 21063
rect 15703 21060 15715 21063
rect 15703 21032 15884 21060
rect 15703 21029 15715 21032
rect 15657 21023 15715 21029
rect 11931 20964 13400 20992
rect 13449 20995 13507 21001
rect 11931 20961 11943 20964
rect 11885 20955 11943 20961
rect 13449 20961 13461 20995
rect 13495 20992 13507 20995
rect 13906 20992 13912 21004
rect 13495 20964 13912 20992
rect 13495 20961 13507 20964
rect 13449 20955 13507 20961
rect 13906 20952 13912 20964
rect 13964 20952 13970 21004
rect 14016 20992 14044 21020
rect 14366 20992 14372 21004
rect 14016 20964 14372 20992
rect 14366 20952 14372 20964
rect 14424 20952 14430 21004
rect 15856 20992 15884 21032
rect 15930 21020 15936 21072
rect 15988 21060 15994 21072
rect 15988 21032 16160 21060
rect 15988 21020 15994 21032
rect 16132 21001 16160 21032
rect 22830 21020 22836 21072
rect 22888 21060 22894 21072
rect 23216 21060 23244 21100
rect 27801 21097 27813 21100
rect 27847 21097 27859 21131
rect 27801 21091 27859 21097
rect 22888 21032 23244 21060
rect 22888 21020 22894 21032
rect 25038 21020 25044 21072
rect 25096 21060 25102 21072
rect 25296 21063 25354 21069
rect 25296 21060 25308 21063
rect 25096 21032 25308 21060
rect 25096 21020 25102 21032
rect 25296 21029 25308 21032
rect 25342 21029 25354 21063
rect 25296 21023 25354 21029
rect 25866 21020 25872 21072
rect 25924 21060 25930 21072
rect 26145 21063 26203 21069
rect 26145 21060 26157 21063
rect 25924 21032 26157 21060
rect 25924 21020 25930 21032
rect 26145 21029 26157 21032
rect 26191 21029 26203 21063
rect 26145 21023 26203 21029
rect 16117 20995 16175 21001
rect 15856 20964 15976 20992
rect 11612 20929 11670 20935
rect 11612 20895 11624 20929
rect 11658 20895 11670 20929
rect 11612 20889 11670 20895
rect 13814 20884 13820 20936
rect 13872 20884 13878 20936
rect 14093 20927 14151 20933
rect 14093 20893 14105 20927
rect 14139 20893 14151 20927
rect 15948 20924 15976 20964
rect 16117 20961 16129 20995
rect 16163 20961 16175 20995
rect 16117 20955 16175 20961
rect 16206 20952 16212 21004
rect 16264 20992 16270 21004
rect 17957 20995 18015 21001
rect 17957 20992 17969 20995
rect 16264 20964 17969 20992
rect 16264 20952 16270 20964
rect 17957 20961 17969 20964
rect 18003 20961 18015 20995
rect 17957 20955 18015 20961
rect 18325 20995 18383 21001
rect 18325 20961 18337 20995
rect 18371 20961 18383 20995
rect 20622 20992 20628 21004
rect 20378 20964 20628 20992
rect 18325 20955 18383 20961
rect 16224 20924 16252 20952
rect 15948 20896 16252 20924
rect 14093 20887 14151 20893
rect 10928 20828 11192 20856
rect 12912 20828 13584 20856
rect 10928 20816 10934 20828
rect 11422 20788 11428 20800
rect 10336 20760 11428 20788
rect 11422 20748 11428 20760
rect 11480 20748 11486 20800
rect 12250 20748 12256 20800
rect 12308 20788 12314 20800
rect 12912 20788 12940 20828
rect 13556 20797 13584 20828
rect 12308 20760 12940 20788
rect 13541 20791 13599 20797
rect 12308 20748 12314 20760
rect 13541 20757 13553 20791
rect 13587 20757 13599 20791
rect 13832 20788 13860 20884
rect 14108 20856 14136 20887
rect 16298 20884 16304 20936
rect 16356 20924 16362 20936
rect 16393 20927 16451 20933
rect 16393 20924 16405 20927
rect 16356 20896 16405 20924
rect 16356 20884 16362 20896
rect 16393 20893 16405 20896
rect 16439 20924 16451 20927
rect 18340 20924 18368 20955
rect 20622 20952 20628 20964
rect 20680 20952 20686 21004
rect 20993 20995 21051 21001
rect 20993 20961 21005 20995
rect 21039 20961 21051 20995
rect 23106 20992 23112 21004
rect 22678 20964 23112 20992
rect 20993 20955 21051 20961
rect 16439 20896 18368 20924
rect 18693 20927 18751 20933
rect 16439 20893 16451 20896
rect 16393 20887 16451 20893
rect 18693 20893 18705 20927
rect 18739 20924 18751 20927
rect 18874 20924 18880 20936
rect 18739 20896 18880 20924
rect 18739 20893 18751 20896
rect 18693 20887 18751 20893
rect 14274 20856 14280 20868
rect 14108 20828 14280 20856
rect 14274 20816 14280 20828
rect 14332 20816 14338 20868
rect 18708 20856 18736 20887
rect 18874 20884 18880 20896
rect 18932 20884 18938 20936
rect 18969 20927 19027 20933
rect 18969 20893 18981 20927
rect 19015 20893 19027 20927
rect 18969 20887 19027 20893
rect 17144 20828 18736 20856
rect 15933 20791 15991 20797
rect 15933 20788 15945 20791
rect 13832 20760 15945 20788
rect 13541 20751 13599 20757
rect 15933 20757 15945 20760
rect 15979 20757 15991 20791
rect 15933 20751 15991 20757
rect 16758 20748 16764 20800
rect 16816 20788 16822 20800
rect 17144 20788 17172 20828
rect 16816 20760 17172 20788
rect 16816 20748 16822 20760
rect 17218 20748 17224 20800
rect 17276 20788 17282 20800
rect 17497 20791 17555 20797
rect 17497 20788 17509 20791
rect 17276 20760 17509 20788
rect 17276 20748 17282 20760
rect 17497 20757 17509 20760
rect 17543 20757 17555 20791
rect 18984 20788 19012 20887
rect 19242 20884 19248 20936
rect 19300 20924 19306 20936
rect 21008 20924 21036 20955
rect 23106 20952 23112 20964
rect 23164 20952 23170 21004
rect 23293 20995 23351 21001
rect 23293 20961 23305 20995
rect 23339 20961 23351 20995
rect 25130 20992 25136 21004
rect 24886 20964 25136 20992
rect 23293 20955 23351 20961
rect 19300 20896 21036 20924
rect 19300 20884 19306 20896
rect 21174 20884 21180 20936
rect 21232 20924 21238 20936
rect 21269 20927 21327 20933
rect 21269 20924 21281 20927
rect 21232 20896 21281 20924
rect 21232 20884 21238 20896
rect 21269 20893 21281 20896
rect 21315 20893 21327 20927
rect 21269 20887 21327 20893
rect 21545 20927 21603 20933
rect 21545 20893 21557 20927
rect 21591 20924 21603 20927
rect 23308 20924 23336 20955
rect 25130 20952 25136 20964
rect 25188 20952 25194 21004
rect 25501 20995 25559 21001
rect 25501 20961 25513 20995
rect 25547 20961 25559 20995
rect 25501 20955 25559 20961
rect 25777 20995 25835 21001
rect 25777 20961 25789 20995
rect 25823 20961 25835 20995
rect 25777 20955 25835 20961
rect 26421 20995 26479 21001
rect 26421 20961 26433 20995
rect 26467 20992 26479 20995
rect 26467 20964 26832 20992
rect 26467 20961 26479 20964
rect 26421 20955 26479 20961
rect 23477 20927 23535 20933
rect 23477 20924 23489 20927
rect 21591 20896 23489 20924
rect 21591 20893 21603 20896
rect 21545 20887 21603 20893
rect 23477 20893 23489 20896
rect 23523 20893 23535 20927
rect 23753 20927 23811 20933
rect 23753 20924 23765 20927
rect 23477 20887 23535 20893
rect 23584 20896 23765 20924
rect 23584 20856 23612 20896
rect 23753 20893 23765 20896
rect 23799 20924 23811 20927
rect 25516 20924 25544 20955
rect 23799 20896 25544 20924
rect 23799 20893 23811 20896
rect 23753 20887 23811 20893
rect 22756 20828 23612 20856
rect 22756 20800 22784 20828
rect 22646 20788 22652 20800
rect 18984 20760 22652 20788
rect 17497 20751 17555 20757
rect 22646 20748 22652 20760
rect 22704 20748 22710 20800
rect 22738 20748 22744 20800
rect 22796 20748 22802 20800
rect 24486 20748 24492 20800
rect 24544 20788 24550 20800
rect 25792 20788 25820 20955
rect 26804 20936 26832 20964
rect 27430 20952 27436 21004
rect 27488 20992 27494 21004
rect 28588 20995 28646 21001
rect 28588 20992 28600 20995
rect 27488 20964 28600 20992
rect 27488 20952 27494 20964
rect 28588 20961 28600 20964
rect 28634 20961 28646 20995
rect 28588 20955 28646 20961
rect 28920 20964 29684 20992
rect 26694 20884 26700 20936
rect 26752 20884 26758 20936
rect 26786 20884 26792 20936
rect 26844 20884 26850 20936
rect 26878 20884 26884 20936
rect 26936 20924 26942 20936
rect 28261 20927 28319 20933
rect 28261 20924 28273 20927
rect 26936 20896 28273 20924
rect 26936 20884 26942 20896
rect 28261 20893 28273 20896
rect 28307 20893 28319 20927
rect 28261 20887 28319 20893
rect 28767 20927 28825 20933
rect 28767 20893 28779 20927
rect 28813 20924 28825 20927
rect 28920 20924 28948 20964
rect 29656 20936 29684 20964
rect 28813 20896 28948 20924
rect 28997 20927 29055 20933
rect 28813 20893 28825 20896
rect 28767 20887 28825 20893
rect 28997 20893 29009 20927
rect 29043 20924 29055 20927
rect 29454 20924 29460 20936
rect 29043 20896 29460 20924
rect 29043 20893 29055 20896
rect 28997 20887 29055 20893
rect 29454 20884 29460 20896
rect 29512 20884 29518 20936
rect 29638 20884 29644 20936
rect 29696 20884 29702 20936
rect 24544 20760 25820 20788
rect 24544 20748 24550 20760
rect 26878 20748 26884 20800
rect 26936 20788 26942 20800
rect 30101 20791 30159 20797
rect 30101 20788 30113 20791
rect 26936 20760 30113 20788
rect 26936 20748 26942 20760
rect 30101 20757 30113 20760
rect 30147 20757 30159 20791
rect 30101 20751 30159 20757
rect 552 20698 30912 20720
rect 552 20646 4193 20698
rect 4245 20646 4257 20698
rect 4309 20646 4321 20698
rect 4373 20646 4385 20698
rect 4437 20646 4449 20698
rect 4501 20646 11783 20698
rect 11835 20646 11847 20698
rect 11899 20646 11911 20698
rect 11963 20646 11975 20698
rect 12027 20646 12039 20698
rect 12091 20646 19373 20698
rect 19425 20646 19437 20698
rect 19489 20646 19501 20698
rect 19553 20646 19565 20698
rect 19617 20646 19629 20698
rect 19681 20646 26963 20698
rect 27015 20646 27027 20698
rect 27079 20646 27091 20698
rect 27143 20646 27155 20698
rect 27207 20646 27219 20698
rect 27271 20646 30912 20698
rect 552 20624 30912 20646
rect 1762 20544 1768 20596
rect 1820 20584 1826 20596
rect 2777 20587 2835 20593
rect 2777 20584 2789 20587
rect 1820 20556 2789 20584
rect 1820 20544 1826 20556
rect 2777 20553 2789 20556
rect 2823 20553 2835 20587
rect 6638 20584 6644 20596
rect 2777 20547 2835 20553
rect 3804 20556 6644 20584
rect 1443 20451 1501 20457
rect 1443 20417 1455 20451
rect 1489 20448 1501 20451
rect 3234 20448 3240 20460
rect 1489 20420 3240 20448
rect 1489 20417 1501 20420
rect 1443 20411 1501 20417
rect 3234 20408 3240 20420
rect 3292 20408 3298 20460
rect 937 20383 995 20389
rect 937 20349 949 20383
rect 983 20380 995 20383
rect 1210 20380 1216 20392
rect 983 20352 1216 20380
rect 983 20349 995 20352
rect 937 20343 995 20349
rect 1210 20340 1216 20352
rect 1268 20340 1274 20392
rect 1670 20340 1676 20392
rect 1728 20340 1734 20392
rect 2774 20340 2780 20392
rect 2832 20340 2838 20392
rect 3421 20383 3479 20389
rect 3421 20349 3433 20383
rect 3467 20380 3479 20383
rect 3804 20380 3832 20556
rect 6638 20544 6644 20556
rect 6696 20544 6702 20596
rect 6914 20544 6920 20596
rect 6972 20584 6978 20596
rect 7929 20587 7987 20593
rect 7929 20584 7941 20587
rect 6972 20556 7941 20584
rect 6972 20544 6978 20556
rect 7929 20553 7941 20556
rect 7975 20553 7987 20587
rect 10413 20587 10471 20593
rect 7929 20547 7987 20553
rect 8404 20556 10364 20584
rect 5905 20519 5963 20525
rect 5905 20485 5917 20519
rect 5951 20516 5963 20519
rect 5994 20516 6000 20528
rect 5951 20488 6000 20516
rect 5951 20485 5963 20488
rect 5905 20479 5963 20485
rect 5994 20476 6000 20488
rect 6052 20476 6058 20528
rect 7742 20476 7748 20528
rect 7800 20516 7806 20528
rect 8404 20516 8432 20556
rect 7800 20488 8432 20516
rect 10336 20516 10364 20556
rect 10413 20553 10425 20587
rect 10459 20584 10471 20587
rect 10502 20584 10508 20596
rect 10459 20556 10508 20584
rect 10459 20553 10471 20556
rect 10413 20547 10471 20553
rect 10502 20544 10508 20556
rect 10560 20544 10566 20596
rect 10870 20584 10876 20596
rect 10612 20556 10876 20584
rect 10612 20516 10640 20556
rect 10870 20544 10876 20556
rect 10928 20544 10934 20596
rect 10962 20544 10968 20596
rect 11020 20584 11026 20596
rect 12989 20587 13047 20593
rect 12989 20584 13001 20587
rect 11020 20556 13001 20584
rect 11020 20544 11026 20556
rect 12989 20553 13001 20556
rect 13035 20553 13047 20587
rect 12989 20547 13047 20553
rect 14093 20587 14151 20593
rect 14093 20553 14105 20587
rect 14139 20584 14151 20587
rect 14182 20584 14188 20596
rect 14139 20556 14188 20584
rect 14139 20553 14151 20556
rect 14093 20547 14151 20553
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 14366 20544 14372 20596
rect 14424 20584 14430 20596
rect 14534 20587 14592 20593
rect 14534 20584 14546 20587
rect 14424 20556 14546 20584
rect 14424 20544 14430 20556
rect 14534 20553 14546 20556
rect 14580 20584 14592 20587
rect 15102 20584 15108 20596
rect 14580 20556 15108 20584
rect 14580 20553 14592 20556
rect 14534 20547 14592 20553
rect 15102 20544 15108 20556
rect 15160 20544 15166 20596
rect 15194 20544 15200 20596
rect 15252 20584 15258 20596
rect 16025 20587 16083 20593
rect 16025 20584 16037 20587
rect 15252 20556 16037 20584
rect 15252 20544 15258 20556
rect 16025 20553 16037 20556
rect 16071 20553 16083 20587
rect 16025 20547 16083 20553
rect 16390 20544 16396 20596
rect 16448 20584 16454 20596
rect 21358 20584 21364 20596
rect 16448 20556 21364 20584
rect 16448 20544 16454 20556
rect 21358 20544 21364 20556
rect 21416 20544 21422 20596
rect 21542 20544 21548 20596
rect 21600 20584 21606 20596
rect 21600 20556 23152 20584
rect 21600 20544 21606 20556
rect 10336 20488 10640 20516
rect 7800 20476 7806 20488
rect 4387 20451 4445 20457
rect 4387 20417 4399 20451
rect 4433 20448 4445 20451
rect 5074 20448 5080 20460
rect 4433 20420 5080 20448
rect 4433 20417 4445 20420
rect 4387 20411 4445 20417
rect 5074 20408 5080 20420
rect 5132 20408 5138 20460
rect 6454 20457 6460 20460
rect 6416 20451 6460 20457
rect 6416 20417 6428 20451
rect 6416 20411 6460 20417
rect 6454 20408 6460 20411
rect 6512 20408 6518 20460
rect 6595 20451 6653 20457
rect 6595 20417 6607 20451
rect 6641 20448 6653 20451
rect 8895 20451 8953 20457
rect 6641 20420 7144 20448
rect 6641 20417 6653 20420
rect 6595 20411 6653 20417
rect 7116 20392 7144 20420
rect 8895 20417 8907 20451
rect 8941 20448 8953 20451
rect 11093 20451 11151 20457
rect 11093 20448 11105 20451
rect 8941 20420 10272 20448
rect 8941 20417 8953 20420
rect 8895 20411 8953 20417
rect 10244 20392 10272 20420
rect 10980 20420 11105 20448
rect 10980 20392 11008 20420
rect 11093 20417 11105 20420
rect 11139 20417 11151 20451
rect 15930 20448 15936 20460
rect 11093 20411 11151 20417
rect 13832 20420 15936 20448
rect 3467 20352 3832 20380
rect 3881 20383 3939 20389
rect 3467 20349 3479 20352
rect 3421 20343 3479 20349
rect 3881 20349 3893 20383
rect 3927 20349 3939 20383
rect 3881 20343 3939 20349
rect 4617 20383 4675 20389
rect 4617 20349 4629 20383
rect 4663 20380 4675 20383
rect 4706 20380 4712 20392
rect 4663 20352 4712 20380
rect 4663 20349 4675 20352
rect 4617 20343 4675 20349
rect 2792 20312 2820 20340
rect 3896 20312 3924 20343
rect 4706 20340 4712 20352
rect 4764 20340 4770 20392
rect 4890 20340 4896 20392
rect 4948 20380 4954 20392
rect 5442 20380 5448 20392
rect 4948 20352 5448 20380
rect 4948 20340 4954 20352
rect 5442 20340 5448 20352
rect 5500 20380 5506 20392
rect 6089 20383 6147 20389
rect 6089 20380 6101 20383
rect 5500 20352 6101 20380
rect 5500 20340 5506 20352
rect 6089 20349 6101 20352
rect 6135 20349 6147 20383
rect 6089 20343 6147 20349
rect 6822 20340 6828 20392
rect 6880 20340 6886 20392
rect 7098 20340 7104 20392
rect 7156 20340 7162 20392
rect 8386 20340 8392 20392
rect 8444 20340 8450 20392
rect 9125 20383 9183 20389
rect 9125 20380 9137 20383
rect 8496 20352 9137 20380
rect 3970 20312 3976 20324
rect 2792 20284 3976 20312
rect 3970 20272 3976 20284
rect 4028 20272 4034 20324
rect 1394 20204 1400 20256
rect 1452 20253 1458 20256
rect 1452 20244 1461 20253
rect 1762 20244 1768 20256
rect 1452 20216 1768 20244
rect 1452 20207 1461 20216
rect 1452 20204 1458 20207
rect 1762 20204 1768 20216
rect 1820 20204 1826 20256
rect 3697 20247 3755 20253
rect 3697 20213 3709 20247
rect 3743 20244 3755 20247
rect 4246 20244 4252 20256
rect 3743 20216 4252 20244
rect 3743 20213 3755 20216
rect 3697 20207 3755 20213
rect 4246 20204 4252 20216
rect 4304 20204 4310 20256
rect 4347 20247 4405 20253
rect 4347 20213 4359 20247
rect 4393 20244 4405 20247
rect 4614 20244 4620 20256
rect 4393 20216 4620 20244
rect 4393 20213 4405 20216
rect 4347 20207 4405 20213
rect 4614 20204 4620 20216
rect 4672 20204 4678 20256
rect 4890 20204 4896 20256
rect 4948 20244 4954 20256
rect 8496 20244 8524 20352
rect 9125 20349 9137 20352
rect 9171 20349 9183 20383
rect 9125 20343 9183 20349
rect 9490 20340 9496 20392
rect 9548 20380 9554 20392
rect 9548 20352 10180 20380
rect 9548 20340 9554 20352
rect 10152 20312 10180 20352
rect 10226 20340 10232 20392
rect 10284 20340 10290 20392
rect 10597 20383 10655 20389
rect 10597 20349 10609 20383
rect 10643 20349 10655 20383
rect 10597 20343 10655 20349
rect 10612 20312 10640 20343
rect 10962 20340 10968 20392
rect 11020 20340 11026 20392
rect 11238 20340 11244 20392
rect 11296 20380 11302 20392
rect 11333 20383 11391 20389
rect 11333 20380 11345 20383
rect 11296 20352 11345 20380
rect 11296 20340 11302 20352
rect 11333 20349 11345 20352
rect 11379 20349 11391 20383
rect 11333 20343 11391 20349
rect 12897 20383 12955 20389
rect 12897 20349 12909 20383
rect 12943 20380 12955 20383
rect 12943 20352 13768 20380
rect 12943 20349 12955 20352
rect 12897 20343 12955 20349
rect 10152 20284 10640 20312
rect 4948 20216 8524 20244
rect 4948 20204 4954 20216
rect 8662 20204 8668 20256
rect 8720 20244 8726 20256
rect 8855 20247 8913 20253
rect 8855 20244 8867 20247
rect 8720 20216 8867 20244
rect 8720 20204 8726 20216
rect 8855 20213 8867 20216
rect 8901 20244 8913 20247
rect 11063 20247 11121 20253
rect 11063 20244 11075 20247
rect 8901 20216 11075 20244
rect 8901 20213 8913 20216
rect 8855 20207 8913 20213
rect 11063 20213 11075 20216
rect 11109 20244 11121 20247
rect 11606 20244 11612 20256
rect 11109 20216 11612 20244
rect 11109 20213 11121 20216
rect 11063 20207 11121 20213
rect 11606 20204 11612 20216
rect 11664 20204 11670 20256
rect 12621 20247 12679 20253
rect 12621 20213 12633 20247
rect 12667 20244 12679 20247
rect 13262 20244 13268 20256
rect 12667 20216 13268 20244
rect 12667 20213 12679 20216
rect 12621 20207 12679 20213
rect 13262 20204 13268 20216
rect 13320 20204 13326 20256
rect 13740 20244 13768 20352
rect 13832 20321 13860 20420
rect 15930 20408 15936 20420
rect 15988 20448 15994 20460
rect 16117 20451 16175 20457
rect 16117 20448 16129 20451
rect 15988 20420 16129 20448
rect 15988 20408 15994 20420
rect 16117 20417 16129 20420
rect 16163 20448 16175 20451
rect 18233 20451 18291 20457
rect 18233 20448 18245 20451
rect 16163 20420 18245 20448
rect 16163 20417 16175 20420
rect 16117 20411 16175 20417
rect 18233 20417 18245 20420
rect 18279 20417 18291 20451
rect 18233 20411 18291 20417
rect 19242 20408 19248 20460
rect 19300 20408 19306 20460
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20448 19579 20451
rect 21174 20448 21180 20460
rect 19567 20420 21180 20448
rect 19567 20417 19579 20420
rect 19521 20411 19579 20417
rect 21174 20408 21180 20420
rect 21232 20448 21238 20460
rect 21266 20451 21324 20457
rect 21266 20448 21278 20451
rect 21232 20420 21278 20448
rect 21232 20408 21238 20420
rect 21266 20417 21278 20420
rect 21312 20417 21324 20451
rect 21560 20448 21588 20544
rect 23124 20528 23152 20556
rect 27062 20544 27068 20596
rect 27120 20584 27126 20596
rect 27430 20584 27436 20596
rect 27120 20556 27436 20584
rect 27120 20544 27126 20556
rect 27430 20544 27436 20556
rect 27488 20544 27494 20596
rect 29362 20544 29368 20596
rect 29420 20584 29426 20596
rect 29420 20556 30420 20584
rect 29420 20544 29426 20556
rect 23106 20476 23112 20528
rect 23164 20476 23170 20528
rect 29104 20488 30328 20516
rect 21266 20411 21324 20417
rect 21468 20420 21588 20448
rect 21821 20451 21879 20457
rect 14274 20340 14280 20392
rect 14332 20389 14338 20392
rect 14332 20343 14342 20389
rect 14332 20340 14338 20343
rect 16390 20340 16396 20392
rect 16448 20340 16454 20392
rect 20622 20340 20628 20392
rect 20680 20380 20686 20392
rect 21468 20380 21496 20420
rect 21821 20417 21833 20451
rect 21867 20448 21879 20451
rect 23845 20451 23903 20457
rect 23845 20448 23857 20451
rect 21867 20420 23857 20448
rect 21867 20417 21879 20420
rect 21821 20411 21879 20417
rect 23584 20389 23612 20420
rect 23845 20417 23857 20420
rect 23891 20417 23903 20451
rect 23845 20411 23903 20417
rect 24121 20451 24179 20457
rect 24121 20417 24133 20451
rect 24167 20448 24179 20451
rect 24167 20420 25912 20448
rect 24167 20417 24179 20420
rect 24121 20411 24179 20417
rect 20680 20352 21496 20380
rect 21545 20383 21603 20389
rect 20680 20340 20686 20352
rect 21545 20349 21557 20383
rect 21591 20349 21603 20383
rect 21545 20343 21603 20349
rect 23569 20383 23627 20389
rect 23569 20349 23581 20383
rect 23615 20349 23627 20383
rect 23569 20343 23627 20349
rect 13817 20315 13875 20321
rect 13817 20281 13829 20315
rect 13863 20281 13875 20315
rect 14292 20312 14320 20340
rect 14826 20312 14832 20324
rect 14292 20284 14832 20312
rect 13817 20275 13875 20281
rect 14826 20272 14832 20284
rect 14884 20272 14890 20324
rect 16206 20312 16212 20324
rect 15778 20284 16212 20312
rect 16206 20272 16212 20284
rect 16264 20272 16270 20324
rect 17954 20272 17960 20324
rect 18012 20312 18018 20324
rect 18012 20284 18184 20312
rect 18012 20272 18018 20284
rect 15378 20244 15384 20256
rect 13740 20216 15384 20244
rect 15378 20204 15384 20216
rect 15436 20204 15442 20256
rect 17494 20204 17500 20256
rect 17552 20204 17558 20256
rect 18156 20244 18184 20284
rect 18782 20272 18788 20324
rect 18840 20272 18846 20324
rect 21560 20312 21588 20343
rect 25130 20340 25136 20392
rect 25188 20380 25194 20392
rect 25188 20352 25254 20380
rect 25188 20340 25194 20352
rect 25682 20340 25688 20392
rect 25740 20340 25746 20392
rect 25884 20389 25912 20420
rect 26418 20408 26424 20460
rect 26476 20448 26482 20460
rect 26602 20448 26608 20460
rect 26476 20420 26608 20448
rect 26476 20408 26482 20420
rect 26602 20408 26608 20420
rect 26660 20448 26666 20460
rect 26697 20451 26755 20457
rect 26697 20448 26709 20451
rect 26660 20420 26709 20448
rect 26660 20408 26666 20420
rect 26697 20417 26709 20420
rect 26743 20417 26755 20451
rect 26697 20411 26755 20417
rect 27203 20451 27261 20457
rect 27203 20417 27215 20451
rect 27249 20448 27261 20451
rect 27249 20420 28764 20448
rect 27249 20417 27261 20420
rect 27203 20411 27261 20417
rect 27062 20389 27068 20392
rect 25869 20383 25927 20389
rect 25869 20349 25881 20383
rect 25915 20349 25927 20383
rect 27024 20383 27068 20389
rect 27024 20380 27036 20383
rect 25869 20343 25927 20349
rect 26620 20352 27036 20380
rect 23106 20312 23112 20324
rect 21560 20284 22140 20312
rect 23046 20284 23112 20312
rect 18690 20244 18696 20256
rect 18156 20216 18696 20244
rect 18690 20204 18696 20216
rect 18748 20244 18754 20256
rect 18877 20247 18935 20253
rect 18877 20244 18889 20247
rect 18748 20216 18889 20244
rect 18748 20204 18754 20216
rect 18877 20213 18889 20216
rect 18923 20213 18935 20247
rect 18877 20207 18935 20213
rect 21085 20247 21143 20253
rect 21085 20213 21097 20247
rect 21131 20244 21143 20247
rect 22002 20244 22008 20256
rect 21131 20216 22008 20244
rect 21131 20213 21143 20216
rect 21085 20207 21143 20213
rect 22002 20204 22008 20216
rect 22060 20204 22066 20256
rect 22112 20244 22140 20284
rect 23106 20272 23112 20284
rect 23164 20312 23170 20324
rect 23474 20312 23480 20324
rect 23164 20284 23480 20312
rect 23164 20272 23170 20284
rect 23474 20272 23480 20284
rect 23532 20272 23538 20324
rect 24394 20272 24400 20324
rect 24452 20272 24458 20324
rect 25700 20312 25728 20340
rect 26620 20324 26648 20352
rect 27024 20349 27036 20352
rect 27024 20343 27068 20349
rect 27062 20340 27068 20343
rect 27120 20340 27126 20392
rect 27433 20383 27491 20389
rect 27433 20349 27445 20383
rect 27479 20380 27491 20383
rect 27479 20352 28672 20380
rect 27479 20349 27491 20352
rect 27433 20343 27491 20349
rect 26145 20315 26203 20321
rect 26145 20312 26157 20315
rect 25700 20284 26157 20312
rect 26145 20281 26157 20284
rect 26191 20281 26203 20315
rect 26145 20275 26203 20281
rect 26602 20272 26608 20324
rect 26660 20272 26666 20324
rect 22462 20244 22468 20256
rect 22112 20216 22468 20244
rect 22462 20204 22468 20216
rect 22520 20204 22526 20256
rect 23385 20247 23443 20253
rect 23385 20213 23397 20247
rect 23431 20244 23443 20247
rect 24412 20244 24440 20272
rect 23431 20216 24440 20244
rect 23431 20213 23443 20216
rect 23385 20207 23443 20213
rect 24762 20204 24768 20256
rect 24820 20244 24826 20256
rect 25685 20247 25743 20253
rect 25685 20244 25697 20247
rect 24820 20216 25697 20244
rect 24820 20204 24826 20216
rect 25685 20213 25697 20216
rect 25731 20213 25743 20247
rect 25685 20207 25743 20213
rect 26234 20204 26240 20256
rect 26292 20204 26298 20256
rect 26510 20204 26516 20256
rect 26568 20244 26574 20256
rect 28537 20247 28595 20253
rect 28537 20244 28549 20247
rect 26568 20216 28549 20244
rect 26568 20204 26574 20216
rect 28537 20213 28549 20216
rect 28583 20213 28595 20247
rect 28644 20244 28672 20352
rect 28736 20312 28764 20420
rect 29104 20392 29132 20488
rect 30300 20457 30328 20488
rect 30285 20451 30343 20457
rect 29288 20420 30052 20448
rect 29288 20392 29316 20420
rect 29086 20340 29092 20392
rect 29144 20340 29150 20392
rect 29270 20340 29276 20392
rect 29328 20340 29334 20392
rect 29362 20340 29368 20392
rect 29420 20340 29426 20392
rect 30024 20389 30052 20420
rect 30285 20417 30297 20451
rect 30331 20417 30343 20451
rect 30285 20411 30343 20417
rect 30009 20383 30067 20389
rect 30009 20349 30021 20383
rect 30055 20349 30067 20383
rect 30009 20343 30067 20349
rect 30193 20383 30251 20389
rect 30193 20349 30205 20383
rect 30239 20380 30251 20383
rect 30392 20380 30420 20556
rect 30239 20352 30420 20380
rect 30239 20349 30251 20352
rect 30193 20343 30251 20349
rect 28736 20284 30236 20312
rect 30208 20256 30236 20284
rect 28994 20244 29000 20256
rect 28644 20216 29000 20244
rect 28537 20207 28595 20213
rect 28994 20204 29000 20216
rect 29052 20204 29058 20256
rect 29641 20247 29699 20253
rect 29641 20213 29653 20247
rect 29687 20244 29699 20247
rect 29822 20244 29828 20256
rect 29687 20216 29828 20244
rect 29687 20213 29699 20216
rect 29641 20207 29699 20213
rect 29822 20204 29828 20216
rect 29880 20204 29886 20256
rect 30190 20204 30196 20256
rect 30248 20204 30254 20256
rect 30469 20247 30527 20253
rect 30469 20213 30481 20247
rect 30515 20244 30527 20247
rect 31202 20244 31208 20256
rect 30515 20216 31208 20244
rect 30515 20213 30527 20216
rect 30469 20207 30527 20213
rect 31202 20204 31208 20216
rect 31260 20204 31266 20256
rect 552 20154 31072 20176
rect 552 20102 7988 20154
rect 8040 20102 8052 20154
rect 8104 20102 8116 20154
rect 8168 20102 8180 20154
rect 8232 20102 8244 20154
rect 8296 20102 15578 20154
rect 15630 20102 15642 20154
rect 15694 20102 15706 20154
rect 15758 20102 15770 20154
rect 15822 20102 15834 20154
rect 15886 20102 23168 20154
rect 23220 20102 23232 20154
rect 23284 20102 23296 20154
rect 23348 20102 23360 20154
rect 23412 20102 23424 20154
rect 23476 20102 30758 20154
rect 30810 20102 30822 20154
rect 30874 20102 30886 20154
rect 30938 20102 30950 20154
rect 31002 20102 31014 20154
rect 31066 20102 31072 20154
rect 552 20080 31072 20102
rect 1587 20043 1645 20049
rect 1587 20009 1599 20043
rect 1633 20040 1645 20043
rect 1762 20040 1768 20052
rect 1633 20012 1768 20040
rect 1633 20009 1645 20012
rect 1587 20003 1645 20009
rect 1762 20000 1768 20012
rect 1820 20000 1826 20052
rect 3145 20043 3203 20049
rect 3145 20009 3157 20043
rect 3191 20040 3203 20043
rect 3786 20040 3792 20052
rect 3191 20012 3792 20040
rect 3191 20009 3203 20012
rect 3145 20003 3203 20009
rect 3786 20000 3792 20012
rect 3844 20000 3850 20052
rect 4246 20000 4252 20052
rect 4304 20040 4310 20052
rect 4304 20012 7236 20040
rect 4304 20000 4310 20012
rect 7208 19972 7236 20012
rect 7834 20000 7840 20052
rect 7892 20000 7898 20052
rect 9582 20040 9588 20052
rect 7944 20012 9588 20040
rect 7944 19972 7972 20012
rect 9582 20000 9588 20012
rect 9640 20000 9646 20052
rect 11238 20040 11244 20052
rect 10336 20012 11244 20040
rect 8386 19972 8392 19984
rect 7208 19944 7972 19972
rect 8036 19944 8392 19972
rect 658 19864 664 19916
rect 716 19904 722 19916
rect 1029 19907 1087 19913
rect 1029 19904 1041 19907
rect 716 19876 1041 19904
rect 716 19864 722 19876
rect 1029 19873 1041 19876
rect 1075 19873 1087 19907
rect 1029 19867 1087 19873
rect 1121 19907 1179 19913
rect 1121 19873 1133 19907
rect 1167 19904 1179 19907
rect 1210 19904 1216 19916
rect 1167 19876 1216 19904
rect 1167 19873 1179 19876
rect 1121 19867 1179 19873
rect 1210 19864 1216 19876
rect 1268 19864 1274 19916
rect 2866 19904 2872 19916
rect 1786 19876 2872 19904
rect 1617 19857 1675 19863
rect 1617 19854 1629 19857
rect 1596 19823 1629 19854
rect 1663 19836 1675 19857
rect 1786 19836 1814 19876
rect 2866 19864 2872 19876
rect 2924 19864 2930 19916
rect 5629 19907 5687 19913
rect 4178 19876 5212 19904
rect 1663 19823 1814 19836
rect 1596 19808 1814 19823
rect 1854 19796 1860 19848
rect 1912 19796 1918 19848
rect 3510 19796 3516 19848
rect 3568 19836 3574 19848
rect 3694 19836 3700 19848
rect 3568 19808 3700 19836
rect 3568 19796 3574 19808
rect 3694 19796 3700 19808
rect 3752 19796 3758 19848
rect 3878 19845 3884 19848
rect 3840 19839 3884 19845
rect 3840 19805 3852 19839
rect 3840 19799 3884 19805
rect 3878 19796 3884 19799
rect 3936 19796 3942 19848
rect 4019 19839 4077 19845
rect 4019 19805 4031 19839
rect 4065 19836 4077 19839
rect 4178 19836 4206 19876
rect 5184 19848 5212 19876
rect 5629 19873 5641 19907
rect 5675 19904 5687 19907
rect 5675 19876 6316 19904
rect 5675 19873 5687 19876
rect 5629 19867 5687 19873
rect 4065 19808 4206 19836
rect 4249 19839 4307 19845
rect 4065 19805 4077 19808
rect 4019 19799 4077 19805
rect 4249 19805 4261 19839
rect 4295 19836 4307 19839
rect 4706 19836 4712 19848
rect 4295 19808 4712 19836
rect 4295 19805 4307 19808
rect 4249 19799 4307 19805
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 5074 19796 5080 19848
rect 5132 19796 5138 19848
rect 5166 19796 5172 19848
rect 5224 19796 5230 19848
rect 5810 19796 5816 19848
rect 5868 19796 5874 19848
rect 6178 19845 6184 19848
rect 6140 19839 6184 19845
rect 6140 19805 6152 19839
rect 6140 19799 6184 19805
rect 6178 19796 6184 19799
rect 6236 19796 6242 19848
rect 6288 19845 6316 19876
rect 6914 19864 6920 19916
rect 6972 19904 6978 19916
rect 8036 19904 8064 19944
rect 8386 19932 8392 19944
rect 8444 19932 8450 19984
rect 6972 19876 8064 19904
rect 6972 19864 6978 19876
rect 8202 19864 8208 19916
rect 8260 19864 8266 19916
rect 8312 19876 8616 19904
rect 6276 19839 6334 19845
rect 6276 19805 6288 19839
rect 6322 19805 6334 19839
rect 6276 19799 6334 19805
rect 6546 19796 6552 19848
rect 6604 19796 6610 19848
rect 7650 19796 7656 19848
rect 7708 19836 7714 19848
rect 8312 19836 8340 19876
rect 7708 19808 8340 19836
rect 7708 19796 7714 19808
rect 8386 19796 8392 19848
rect 8444 19796 8450 19848
rect 8481 19839 8539 19845
rect 8481 19805 8493 19839
rect 8527 19805 8539 19839
rect 8588 19836 8616 19876
rect 9030 19864 9036 19916
rect 9088 19904 9094 19916
rect 10336 19904 10364 20012
rect 11238 20000 11244 20012
rect 11296 20000 11302 20052
rect 11514 20000 11520 20052
rect 11572 20040 11578 20052
rect 12535 20043 12593 20049
rect 12535 20040 12547 20043
rect 11572 20012 12547 20040
rect 11572 20000 11578 20012
rect 12535 20009 12547 20012
rect 12581 20040 12593 20043
rect 13630 20040 13636 20052
rect 12581 20012 13636 20040
rect 12581 20009 12593 20012
rect 12535 20003 12593 20009
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 13906 20000 13912 20052
rect 13964 20000 13970 20052
rect 14826 20000 14832 20052
rect 14884 20040 14890 20052
rect 14884 20012 16344 20040
rect 14884 20000 14890 20012
rect 9088 19876 10364 19904
rect 9088 19864 9094 19876
rect 10870 19864 10876 19916
rect 10928 19904 10934 19916
rect 11238 19904 11244 19938
rect 10928 19886 11244 19904
rect 11296 19904 11302 19938
rect 16316 19916 16344 20012
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 16761 20043 16819 20049
rect 16761 20040 16773 20043
rect 16632 20012 16773 20040
rect 16632 20000 16638 20012
rect 16761 20009 16773 20012
rect 16807 20009 16819 20043
rect 16761 20003 16819 20009
rect 22186 20000 22192 20052
rect 22244 20040 22250 20052
rect 22830 20040 22836 20052
rect 22244 20012 22836 20040
rect 22244 20000 22250 20012
rect 22830 20000 22836 20012
rect 22888 20040 22894 20052
rect 22888 20012 23796 20040
rect 22888 20000 22894 20012
rect 22738 19972 22744 19984
rect 22204 19944 22744 19972
rect 12805 19907 12863 19913
rect 11296 19886 12112 19904
rect 10928 19876 12112 19886
rect 10928 19864 10934 19876
rect 8846 19845 8852 19848
rect 8808 19839 8852 19845
rect 8808 19836 8820 19839
rect 8588 19808 8820 19836
rect 8481 19799 8539 19805
rect 8808 19805 8820 19808
rect 8808 19799 8852 19805
rect 5092 19768 5120 19796
rect 5828 19768 5856 19796
rect 8496 19768 8524 19799
rect 8846 19796 8852 19799
rect 8904 19796 8910 19848
rect 8938 19796 8944 19848
rect 8996 19836 9002 19848
rect 8996 19808 9041 19836
rect 8996 19796 9002 19808
rect 9214 19796 9220 19848
rect 9272 19796 9278 19848
rect 10965 19839 11023 19845
rect 10965 19805 10977 19839
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 11241 19839 11299 19845
rect 11241 19805 11253 19839
rect 11287 19836 11299 19839
rect 11422 19836 11428 19848
rect 11287 19808 11428 19836
rect 11287 19805 11299 19808
rect 11241 19799 11299 19805
rect 5092 19740 5856 19768
rect 8404 19740 8524 19768
rect 842 19660 848 19712
rect 900 19660 906 19712
rect 5442 19660 5448 19712
rect 5500 19700 5506 19712
rect 7742 19700 7748 19712
rect 5500 19672 7748 19700
rect 5500 19660 5506 19672
rect 7742 19660 7748 19672
rect 7800 19700 7806 19712
rect 8404 19700 8432 19740
rect 9950 19728 9956 19780
rect 10008 19768 10014 19780
rect 10505 19771 10563 19777
rect 10505 19768 10517 19771
rect 10008 19740 10517 19768
rect 10008 19728 10014 19740
rect 10505 19737 10517 19740
rect 10551 19737 10563 19771
rect 10505 19731 10563 19737
rect 7800 19672 8432 19700
rect 7800 19660 7806 19672
rect 8478 19660 8484 19712
rect 8536 19700 8542 19712
rect 10318 19700 10324 19712
rect 8536 19672 10324 19700
rect 8536 19660 8542 19672
rect 10318 19660 10324 19672
rect 10376 19660 10382 19712
rect 10980 19700 11008 19799
rect 11422 19796 11428 19808
rect 11480 19796 11486 19848
rect 12084 19845 12112 19876
rect 12805 19873 12817 19907
rect 12851 19904 12863 19907
rect 16022 19904 16028 19916
rect 12851 19876 16028 19904
rect 12851 19873 12863 19876
rect 12805 19867 12863 19873
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 16298 19864 16304 19916
rect 16356 19864 16362 19916
rect 16485 19907 16543 19913
rect 16485 19873 16497 19907
rect 16531 19873 16543 19907
rect 16485 19867 16543 19873
rect 17221 19907 17279 19913
rect 17221 19873 17233 19907
rect 17267 19904 17279 19907
rect 17494 19904 17500 19916
rect 17267 19876 17500 19904
rect 17267 19873 17279 19876
rect 17221 19867 17279 19873
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19836 12127 19839
rect 12250 19836 12256 19848
rect 12115 19808 12256 19836
rect 12115 19805 12127 19808
rect 12069 19799 12127 19805
rect 12250 19796 12256 19808
rect 12308 19796 12314 19848
rect 12526 19796 12532 19848
rect 12584 19836 12590 19848
rect 12584 19808 12629 19836
rect 12584 19796 12590 19808
rect 14182 19796 14188 19848
rect 14240 19836 14246 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 14240 19808 14289 19836
rect 14240 19796 14246 19808
rect 14277 19805 14289 19808
rect 14323 19805 14335 19839
rect 14277 19799 14335 19805
rect 14458 19796 14464 19848
rect 14516 19836 14522 19848
rect 14553 19839 14611 19845
rect 14553 19836 14565 19839
rect 14516 19808 14565 19836
rect 14516 19796 14522 19808
rect 14553 19805 14565 19808
rect 14599 19836 14611 19839
rect 16206 19836 16212 19848
rect 14599 19808 16212 19836
rect 14599 19805 14611 19808
rect 14553 19799 14611 19805
rect 16206 19796 16212 19808
rect 16264 19796 16270 19848
rect 16500 19768 16528 19867
rect 17494 19864 17500 19876
rect 17552 19864 17558 19916
rect 17954 19864 17960 19916
rect 18012 19864 18018 19916
rect 18693 19907 18751 19913
rect 18693 19873 18705 19907
rect 18739 19904 18751 19907
rect 18782 19904 18788 19916
rect 18739 19876 18788 19904
rect 18739 19873 18751 19876
rect 18693 19867 18751 19873
rect 18782 19864 18788 19876
rect 18840 19864 18846 19916
rect 20533 19907 20591 19913
rect 20533 19873 20545 19907
rect 20579 19904 20591 19907
rect 20622 19904 20628 19916
rect 20579 19876 20628 19904
rect 20579 19873 20591 19876
rect 20533 19867 20591 19873
rect 20622 19864 20628 19876
rect 20680 19864 20686 19916
rect 21542 19864 21548 19916
rect 21600 19864 21606 19916
rect 22204 19913 22232 19944
rect 22738 19932 22744 19944
rect 22796 19932 22802 19984
rect 23768 19972 23796 20012
rect 23934 20000 23940 20052
rect 23992 20040 23998 20052
rect 24029 20043 24087 20049
rect 24029 20040 24041 20043
rect 23992 20012 24041 20040
rect 23992 20000 23998 20012
rect 24029 20009 24041 20012
rect 24075 20009 24087 20043
rect 24029 20003 24087 20009
rect 24762 20000 24768 20052
rect 24820 20040 24826 20052
rect 26510 20040 26516 20052
rect 24820 20012 26516 20040
rect 24820 20000 24826 20012
rect 26510 20000 26516 20012
rect 26568 20000 26574 20052
rect 27798 20000 27804 20052
rect 27856 20000 27862 20052
rect 30190 20000 30196 20052
rect 30248 20000 30254 20052
rect 23768 19944 24440 19972
rect 21913 19907 21971 19913
rect 21913 19873 21925 19907
rect 21959 19904 21971 19907
rect 22189 19907 22247 19913
rect 21959 19876 22140 19904
rect 21959 19873 21971 19876
rect 21913 19867 21971 19873
rect 16942 19796 16948 19848
rect 17000 19836 17006 19848
rect 17972 19836 18000 19864
rect 17000 19808 18000 19836
rect 18969 19839 19027 19845
rect 17000 19796 17006 19808
rect 18969 19805 18981 19839
rect 19015 19836 19027 19839
rect 20070 19836 20076 19848
rect 19015 19808 20076 19836
rect 19015 19805 19027 19808
rect 18969 19799 19027 19805
rect 20070 19796 20076 19808
rect 20128 19796 20134 19848
rect 16666 19768 16672 19780
rect 15212 19740 16672 19768
rect 15212 19712 15240 19740
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 20714 19728 20720 19780
rect 20772 19768 20778 19780
rect 21361 19771 21419 19777
rect 21361 19768 21373 19771
rect 20772 19740 21373 19768
rect 20772 19728 20778 19740
rect 21361 19737 21373 19740
rect 21407 19737 21419 19771
rect 21361 19731 21419 19737
rect 22112 19712 22140 19876
rect 22189 19873 22201 19907
rect 22235 19873 22247 19907
rect 22189 19867 22247 19873
rect 23566 19864 23572 19916
rect 23624 19904 23630 19916
rect 23624 19876 23704 19904
rect 23624 19864 23630 19876
rect 22462 19796 22468 19848
rect 22520 19836 22526 19848
rect 23106 19836 23112 19848
rect 22520 19808 23112 19836
rect 22520 19796 22526 19808
rect 23106 19796 23112 19808
rect 23164 19796 23170 19848
rect 23676 19836 23704 19876
rect 23934 19864 23940 19916
rect 23992 19904 23998 19916
rect 24412 19913 24440 19944
rect 24213 19907 24271 19913
rect 24213 19904 24225 19907
rect 23992 19876 24225 19904
rect 23992 19864 23998 19876
rect 24213 19873 24225 19876
rect 24259 19873 24271 19907
rect 24213 19867 24271 19873
rect 24397 19907 24455 19913
rect 24397 19873 24409 19907
rect 24443 19873 24455 19907
rect 25130 19904 25136 19916
rect 24397 19867 24455 19873
rect 24504 19876 25136 19904
rect 24504 19836 24532 19876
rect 25130 19864 25136 19876
rect 25188 19864 25194 19916
rect 26053 19907 26111 19913
rect 26053 19873 26065 19907
rect 26099 19904 26111 19907
rect 26697 19907 26755 19913
rect 26697 19904 26709 19907
rect 26099 19876 26709 19904
rect 26099 19873 26111 19876
rect 26053 19867 26111 19873
rect 26697 19873 26709 19876
rect 26743 19873 26755 19907
rect 26697 19867 26755 19873
rect 23676 19808 24532 19836
rect 24670 19796 24676 19848
rect 24728 19796 24734 19848
rect 26421 19839 26479 19845
rect 26421 19805 26433 19839
rect 26467 19836 26479 19839
rect 26786 19836 26792 19848
rect 26467 19808 26792 19836
rect 26467 19805 26479 19808
rect 26421 19799 26479 19805
rect 26786 19796 26792 19808
rect 26844 19796 26850 19848
rect 27614 19796 27620 19848
rect 27672 19836 27678 19848
rect 28353 19839 28411 19845
rect 28353 19836 28365 19839
rect 27672 19808 28365 19836
rect 27672 19796 27678 19808
rect 28353 19805 28365 19808
rect 28399 19805 28411 19839
rect 28353 19799 28411 19805
rect 28534 19796 28540 19848
rect 28592 19836 28598 19848
rect 28680 19839 28738 19845
rect 28680 19836 28692 19839
rect 28592 19808 28692 19836
rect 28592 19796 28598 19808
rect 28680 19805 28692 19808
rect 28726 19805 28738 19839
rect 28680 19799 28738 19805
rect 28859 19839 28917 19845
rect 28859 19805 28871 19839
rect 28905 19836 28917 19839
rect 28994 19836 29000 19848
rect 28905 19808 29000 19836
rect 28905 19805 28917 19808
rect 28859 19799 28917 19805
rect 28994 19796 29000 19808
rect 29052 19796 29058 19848
rect 29089 19839 29147 19845
rect 29089 19805 29101 19839
rect 29135 19836 29147 19839
rect 29546 19836 29552 19848
rect 29135 19808 29552 19836
rect 29135 19805 29147 19808
rect 29089 19799 29147 19805
rect 29546 19796 29552 19808
rect 29604 19796 29610 19848
rect 14734 19700 14740 19712
rect 10980 19672 14740 19700
rect 14734 19660 14740 19672
rect 14792 19660 14798 19712
rect 15194 19660 15200 19712
rect 15252 19660 15258 19712
rect 15838 19660 15844 19712
rect 15896 19660 15902 19712
rect 18509 19703 18567 19709
rect 18509 19669 18521 19703
rect 18555 19700 18567 19703
rect 18598 19700 18604 19712
rect 18555 19672 18604 19700
rect 18555 19669 18567 19672
rect 18509 19663 18567 19669
rect 18598 19660 18604 19672
rect 18656 19660 18662 19712
rect 19794 19660 19800 19712
rect 19852 19700 19858 19712
rect 20073 19703 20131 19709
rect 20073 19700 20085 19703
rect 19852 19672 20085 19700
rect 19852 19660 19858 19672
rect 20073 19669 20085 19672
rect 20119 19669 20131 19703
rect 20073 19663 20131 19669
rect 20438 19660 20444 19712
rect 20496 19700 20502 19712
rect 20809 19703 20867 19709
rect 20809 19700 20821 19703
rect 20496 19672 20821 19700
rect 20496 19660 20502 19672
rect 20809 19669 20821 19672
rect 20855 19669 20867 19703
rect 20809 19663 20867 19669
rect 22094 19660 22100 19712
rect 22152 19660 22158 19712
rect 22462 19660 22468 19712
rect 22520 19700 22526 19712
rect 26694 19700 26700 19712
rect 22520 19672 26700 19700
rect 22520 19660 22526 19672
rect 26694 19660 26700 19672
rect 26752 19660 26758 19712
rect 29178 19660 29184 19712
rect 29236 19700 29242 19712
rect 30282 19700 30288 19712
rect 29236 19672 30288 19700
rect 29236 19660 29242 19672
rect 30282 19660 30288 19672
rect 30340 19660 30346 19712
rect 552 19610 30912 19632
rect 552 19558 4193 19610
rect 4245 19558 4257 19610
rect 4309 19558 4321 19610
rect 4373 19558 4385 19610
rect 4437 19558 4449 19610
rect 4501 19558 11783 19610
rect 11835 19558 11847 19610
rect 11899 19558 11911 19610
rect 11963 19558 11975 19610
rect 12027 19558 12039 19610
rect 12091 19558 19373 19610
rect 19425 19558 19437 19610
rect 19489 19558 19501 19610
rect 19553 19558 19565 19610
rect 19617 19558 19629 19610
rect 19681 19558 26963 19610
rect 27015 19558 27027 19610
rect 27079 19558 27091 19610
rect 27143 19558 27155 19610
rect 27207 19558 27219 19610
rect 27271 19558 30912 19610
rect 552 19536 30912 19558
rect 842 19456 848 19508
rect 900 19496 906 19508
rect 900 19468 3648 19496
rect 900 19456 906 19468
rect 1443 19363 1501 19369
rect 1443 19329 1455 19363
rect 1489 19360 1501 19363
rect 2774 19360 2780 19372
rect 1489 19332 2780 19360
rect 1489 19329 1501 19332
rect 1443 19323 1501 19329
rect 2774 19320 2780 19332
rect 2832 19320 2838 19372
rect 3620 19360 3648 19468
rect 3970 19456 3976 19508
rect 4028 19496 4034 19508
rect 4028 19468 4568 19496
rect 4028 19456 4034 19468
rect 3694 19388 3700 19440
rect 3752 19428 3758 19440
rect 4246 19428 4252 19440
rect 3752 19400 4252 19428
rect 3752 19388 3758 19400
rect 4246 19388 4252 19400
rect 4304 19388 4310 19440
rect 4540 19428 4568 19468
rect 4614 19456 4620 19508
rect 4672 19496 4678 19508
rect 6178 19496 6184 19508
rect 4672 19468 6184 19496
rect 4672 19456 4678 19468
rect 6178 19456 6184 19468
rect 6236 19496 6242 19508
rect 6236 19468 6684 19496
rect 6236 19456 6242 19468
rect 4985 19431 5043 19437
rect 4985 19428 4997 19431
rect 4540 19400 4997 19428
rect 4985 19397 4997 19400
rect 5031 19397 5043 19431
rect 6656 19428 6684 19468
rect 7098 19456 7104 19508
rect 7156 19456 7162 19508
rect 7558 19456 7564 19508
rect 7616 19496 7622 19508
rect 8202 19496 8208 19508
rect 7616 19468 8208 19496
rect 7616 19456 7622 19468
rect 8202 19456 8208 19468
rect 8260 19456 8266 19508
rect 8662 19496 8668 19508
rect 8404 19468 8668 19496
rect 8404 19428 8432 19468
rect 8662 19456 8668 19468
rect 8720 19456 8726 19508
rect 8846 19456 8852 19508
rect 8904 19496 8910 19508
rect 8904 19468 10180 19496
rect 8904 19456 8910 19468
rect 6656 19400 8432 19428
rect 4985 19391 5043 19397
rect 5000 19360 5028 19391
rect 5074 19360 5080 19372
rect 3620 19332 4936 19360
rect 5000 19332 5080 19360
rect 937 19295 995 19301
rect 937 19261 949 19295
rect 983 19292 995 19295
rect 1210 19292 1216 19304
rect 983 19264 1216 19292
rect 983 19261 995 19264
rect 937 19255 995 19261
rect 1210 19252 1216 19264
rect 1268 19252 1274 19304
rect 1673 19295 1731 19301
rect 1673 19261 1685 19295
rect 1719 19292 1731 19295
rect 2498 19292 2504 19304
rect 1719 19264 2504 19292
rect 1719 19261 1731 19264
rect 1673 19255 1731 19261
rect 2498 19252 2504 19264
rect 2556 19252 2562 19304
rect 3050 19252 3056 19304
rect 3108 19252 3114 19304
rect 3142 19252 3148 19304
rect 3200 19292 3206 19304
rect 3513 19295 3571 19301
rect 3513 19292 3525 19295
rect 3200 19264 3525 19292
rect 3200 19252 3206 19264
rect 3513 19261 3525 19264
rect 3559 19261 3571 19295
rect 3513 19255 3571 19261
rect 3605 19295 3663 19301
rect 3605 19261 3617 19295
rect 3651 19292 3663 19295
rect 3786 19292 3792 19304
rect 3651 19264 3792 19292
rect 3651 19261 3663 19264
rect 3605 19255 3663 19261
rect 2958 19184 2964 19236
rect 3016 19224 3022 19236
rect 3620 19224 3648 19255
rect 3786 19252 3792 19264
rect 3844 19252 3850 19304
rect 3878 19252 3884 19304
rect 3936 19252 3942 19304
rect 4338 19252 4344 19304
rect 4396 19292 4402 19304
rect 4908 19292 4936 19332
rect 5074 19320 5080 19332
rect 5132 19360 5138 19372
rect 5261 19363 5319 19369
rect 5261 19360 5273 19363
rect 5132 19332 5273 19360
rect 5132 19320 5138 19332
rect 5261 19329 5273 19332
rect 5307 19329 5319 19363
rect 5261 19323 5319 19329
rect 5534 19320 5540 19372
rect 5592 19360 5598 19372
rect 5724 19363 5782 19369
rect 5724 19360 5736 19363
rect 5592 19332 5736 19360
rect 5592 19320 5598 19332
rect 5724 19329 5736 19332
rect 5770 19329 5782 19363
rect 6454 19360 6460 19372
rect 5724 19323 5782 19329
rect 5920 19332 6460 19360
rect 5920 19292 5948 19332
rect 6454 19320 6460 19332
rect 6512 19320 6518 19372
rect 6914 19320 6920 19372
rect 6972 19360 6978 19372
rect 8113 19363 8171 19369
rect 8113 19360 8125 19363
rect 6972 19332 8125 19360
rect 6972 19320 6978 19332
rect 8113 19329 8125 19332
rect 8159 19360 8171 19363
rect 8202 19360 8208 19372
rect 8159 19332 8208 19360
rect 8159 19329 8171 19332
rect 8113 19323 8171 19329
rect 8202 19320 8208 19332
rect 8260 19320 8266 19372
rect 8312 19332 8524 19360
rect 4396 19264 4752 19292
rect 4908 19264 5948 19292
rect 5997 19295 6055 19301
rect 4396 19252 4402 19264
rect 4724 19236 4752 19264
rect 5997 19261 6009 19295
rect 6043 19292 6055 19295
rect 6270 19292 6276 19304
rect 6043 19264 6276 19292
rect 6043 19261 6055 19264
rect 5997 19255 6055 19261
rect 6270 19252 6276 19264
rect 6328 19252 6334 19304
rect 7650 19252 7656 19304
rect 7708 19252 7714 19304
rect 7742 19252 7748 19304
rect 7800 19292 7806 19304
rect 8312 19292 8340 19332
rect 7800 19264 8340 19292
rect 8389 19295 8447 19301
rect 7800 19252 7806 19264
rect 8389 19261 8401 19295
rect 8435 19261 8447 19295
rect 8496 19292 8524 19332
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 8852 19363 8910 19369
rect 8852 19360 8864 19363
rect 8628 19332 8864 19360
rect 8628 19320 8634 19332
rect 8852 19329 8864 19332
rect 8898 19329 8910 19363
rect 8852 19323 8910 19329
rect 9125 19295 9183 19301
rect 9125 19292 9137 19295
rect 8496 19264 9137 19292
rect 8389 19255 8447 19261
rect 9125 19261 9137 19264
rect 9171 19261 9183 19295
rect 9125 19255 9183 19261
rect 3016 19196 3648 19224
rect 3016 19184 3022 19196
rect 4246 19184 4252 19236
rect 4304 19224 4310 19236
rect 4614 19224 4620 19236
rect 4304 19196 4620 19224
rect 4304 19184 4310 19196
rect 4614 19184 4620 19196
rect 4672 19184 4678 19236
rect 4706 19184 4712 19236
rect 4764 19184 4770 19236
rect 4798 19184 4804 19236
rect 4856 19184 4862 19236
rect 4982 19184 4988 19236
rect 5040 19224 5046 19236
rect 5350 19224 5356 19236
rect 5040 19196 5356 19224
rect 5040 19184 5046 19196
rect 5350 19184 5356 19196
rect 5408 19184 5414 19236
rect 6656 19196 7604 19224
rect 1403 19159 1461 19165
rect 1403 19125 1415 19159
rect 1449 19156 1461 19159
rect 1762 19156 1768 19168
rect 1449 19128 1768 19156
rect 1449 19125 1461 19128
rect 1403 19119 1461 19125
rect 1762 19116 1768 19128
rect 1820 19116 1826 19168
rect 3329 19159 3387 19165
rect 3329 19125 3341 19159
rect 3375 19156 3387 19159
rect 4062 19156 4068 19168
rect 3375 19128 4068 19156
rect 3375 19125 3387 19128
rect 3329 19119 3387 19125
rect 4062 19116 4068 19128
rect 4120 19116 4126 19168
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 4341 19159 4399 19165
rect 4341 19156 4353 19159
rect 4212 19128 4353 19156
rect 4212 19116 4218 19128
rect 4341 19125 4353 19128
rect 4387 19125 4399 19159
rect 4341 19119 4399 19125
rect 5727 19159 5785 19165
rect 5727 19125 5739 19159
rect 5773 19156 5785 19159
rect 5902 19156 5908 19168
rect 5773 19128 5908 19156
rect 5773 19125 5785 19128
rect 5727 19119 5785 19125
rect 5902 19116 5908 19128
rect 5960 19116 5966 19168
rect 5994 19116 6000 19168
rect 6052 19156 6058 19168
rect 6656 19156 6684 19196
rect 6052 19128 6684 19156
rect 6052 19116 6058 19128
rect 7466 19116 7472 19168
rect 7524 19116 7530 19168
rect 7576 19156 7604 19196
rect 7834 19184 7840 19236
rect 7892 19184 7898 19236
rect 8404 19156 8432 19255
rect 10152 19224 10180 19468
rect 10226 19456 10232 19508
rect 10284 19456 10290 19508
rect 10318 19456 10324 19508
rect 10376 19496 10382 19508
rect 14642 19496 14648 19508
rect 10376 19468 14648 19496
rect 10376 19456 10382 19468
rect 14642 19456 14648 19468
rect 14700 19456 14706 19508
rect 15378 19456 15384 19508
rect 15436 19456 15442 19508
rect 20070 19456 20076 19508
rect 20128 19456 20134 19508
rect 20622 19456 20628 19508
rect 20680 19496 20686 19508
rect 22005 19499 22063 19505
rect 20680 19468 21404 19496
rect 20680 19456 20686 19468
rect 13262 19388 13268 19440
rect 13320 19388 13326 19440
rect 18049 19431 18107 19437
rect 18049 19428 18061 19431
rect 17512 19400 18061 19428
rect 10778 19320 10784 19372
rect 10836 19360 10842 19372
rect 11704 19363 11762 19369
rect 11704 19360 11716 19363
rect 10836 19332 11716 19360
rect 10836 19320 10842 19332
rect 11704 19329 11716 19332
rect 11750 19329 11762 19363
rect 13280 19360 13308 19388
rect 14004 19363 14062 19369
rect 14004 19360 14016 19363
rect 13280 19332 14016 19360
rect 11704 19323 11762 19329
rect 14004 19329 14016 19332
rect 14050 19329 14062 19363
rect 14004 19323 14062 19329
rect 15838 19320 15844 19372
rect 15896 19360 15902 19372
rect 16209 19363 16267 19369
rect 16209 19360 16221 19363
rect 15896 19332 16221 19360
rect 15896 19320 15902 19332
rect 16209 19329 16221 19332
rect 16255 19329 16267 19363
rect 16209 19323 16267 19329
rect 10686 19252 10692 19304
rect 10744 19252 10750 19304
rect 11146 19252 11152 19304
rect 11204 19252 11210 19304
rect 11238 19252 11244 19304
rect 11296 19252 11302 19304
rect 11977 19295 12035 19301
rect 11977 19292 11989 19295
rect 11348 19264 11989 19292
rect 10965 19227 11023 19233
rect 10965 19224 10977 19227
rect 10152 19196 10977 19224
rect 10965 19193 10977 19196
rect 11011 19193 11023 19227
rect 11164 19224 11192 19252
rect 11348 19224 11376 19264
rect 11977 19261 11989 19264
rect 12023 19261 12035 19295
rect 11977 19255 12035 19261
rect 12250 19252 12256 19304
rect 12308 19292 12314 19304
rect 13538 19292 13544 19304
rect 12308 19264 13544 19292
rect 12308 19252 12314 19264
rect 13538 19252 13544 19264
rect 13596 19252 13602 19304
rect 13630 19252 13636 19304
rect 13688 19292 13694 19304
rect 13868 19295 13926 19301
rect 13868 19292 13880 19295
rect 13688 19264 13880 19292
rect 13688 19252 13694 19264
rect 13868 19261 13880 19264
rect 13914 19261 13926 19295
rect 13868 19255 13926 19261
rect 14090 19252 14096 19304
rect 14148 19292 14154 19304
rect 14277 19295 14335 19301
rect 14277 19292 14289 19295
rect 14148 19264 14289 19292
rect 14148 19252 14154 19264
rect 14277 19261 14289 19264
rect 14323 19261 14335 19295
rect 14277 19255 14335 19261
rect 15930 19252 15936 19304
rect 15988 19252 15994 19304
rect 16022 19252 16028 19304
rect 16080 19292 16086 19304
rect 17512 19292 17540 19400
rect 18049 19397 18061 19400
rect 18095 19397 18107 19431
rect 21376 19428 21404 19468
rect 22005 19465 22017 19499
rect 22051 19496 22063 19499
rect 24670 19496 24676 19508
rect 22051 19468 24676 19496
rect 22051 19465 22063 19468
rect 22005 19459 22063 19465
rect 24670 19456 24676 19468
rect 24728 19456 24734 19508
rect 28537 19499 28595 19505
rect 28537 19496 28549 19499
rect 26712 19468 28549 19496
rect 22186 19428 22192 19440
rect 21376 19400 22192 19428
rect 18049 19391 18107 19397
rect 22186 19388 22192 19400
rect 22244 19388 22250 19440
rect 23569 19431 23627 19437
rect 23569 19397 23581 19431
rect 23615 19428 23627 19431
rect 23658 19428 23664 19440
rect 23615 19400 23664 19428
rect 23615 19397 23627 19400
rect 23569 19391 23627 19397
rect 23658 19388 23664 19400
rect 23716 19388 23722 19440
rect 18690 19320 18696 19372
rect 18748 19320 18754 19372
rect 20364 19332 20668 19360
rect 16080 19264 17540 19292
rect 17589 19295 17647 19301
rect 16080 19252 16086 19264
rect 17589 19261 17601 19295
rect 17635 19292 17647 19295
rect 17635 19264 18184 19292
rect 17635 19261 17647 19264
rect 17589 19255 17647 19261
rect 11164 19196 11376 19224
rect 10965 19187 11023 19193
rect 8754 19156 8760 19168
rect 7576 19128 8760 19156
rect 8754 19116 8760 19128
rect 8812 19116 8818 19168
rect 8846 19116 8852 19168
rect 8904 19165 8910 19168
rect 8904 19156 8913 19165
rect 10980 19156 11008 19187
rect 17034 19184 17040 19236
rect 17092 19224 17098 19236
rect 17773 19227 17831 19233
rect 17773 19224 17785 19227
rect 17092 19196 17785 19224
rect 17092 19184 17098 19196
rect 17773 19193 17785 19196
rect 17819 19193 17831 19227
rect 17773 19187 17831 19193
rect 17954 19184 17960 19236
rect 18012 19184 18018 19236
rect 18156 19224 18184 19264
rect 18230 19252 18236 19304
rect 18288 19252 18294 19304
rect 18322 19252 18328 19304
rect 18380 19292 18386 19304
rect 18509 19295 18567 19301
rect 18509 19292 18521 19295
rect 18380 19264 18521 19292
rect 18380 19252 18386 19264
rect 18509 19261 18521 19264
rect 18555 19261 18567 19295
rect 18969 19295 19027 19301
rect 18969 19292 18981 19295
rect 18509 19255 18567 19261
rect 18800 19264 18981 19292
rect 18800 19224 18828 19264
rect 18969 19261 18981 19264
rect 19015 19261 19027 19295
rect 18969 19255 19027 19261
rect 19242 19252 19248 19304
rect 19300 19292 19306 19304
rect 20364 19292 20392 19332
rect 19300 19264 20392 19292
rect 19300 19252 19306 19264
rect 20438 19252 20444 19304
rect 20496 19252 20502 19304
rect 20640 19292 20668 19332
rect 20714 19320 20720 19372
rect 20772 19320 20778 19372
rect 21082 19320 21088 19372
rect 21140 19360 21146 19372
rect 21910 19360 21916 19372
rect 21140 19332 21916 19360
rect 21140 19320 21146 19332
rect 21910 19320 21916 19332
rect 21968 19320 21974 19372
rect 22094 19320 22100 19372
rect 22152 19360 22158 19372
rect 24995 19363 25053 19369
rect 22152 19332 23244 19360
rect 22152 19320 22158 19332
rect 23216 19292 23244 19332
rect 24995 19329 25007 19363
rect 25041 19360 25053 19363
rect 26712 19360 26740 19468
rect 28537 19465 28549 19468
rect 28583 19465 28595 19499
rect 28537 19459 28595 19465
rect 29917 19499 29975 19505
rect 29917 19465 29929 19499
rect 29963 19496 29975 19499
rect 29963 19468 30696 19496
rect 29963 19465 29975 19468
rect 29917 19459 29975 19465
rect 29362 19388 29368 19440
rect 29420 19428 29426 19440
rect 29420 19400 30052 19428
rect 29420 19388 29426 19400
rect 25041 19332 26740 19360
rect 27203 19363 27261 19369
rect 25041 19329 25053 19332
rect 24995 19323 25053 19329
rect 27203 19329 27215 19363
rect 27249 19360 27261 19363
rect 29914 19360 29920 19372
rect 27249 19332 29920 19360
rect 27249 19329 27261 19332
rect 27203 19323 27261 19329
rect 29914 19320 29920 19332
rect 29972 19320 29978 19372
rect 23566 19292 23572 19304
rect 20640 19264 22094 19292
rect 23216 19278 23572 19292
rect 23230 19264 23572 19278
rect 18156 19196 18828 19224
rect 11514 19156 11520 19168
rect 8904 19128 8949 19156
rect 10980 19128 11520 19156
rect 8904 19119 8913 19128
rect 8904 19116 8910 19119
rect 11514 19116 11520 19128
rect 11572 19156 11578 19168
rect 11707 19159 11765 19165
rect 11707 19156 11719 19159
rect 11572 19128 11719 19156
rect 11572 19116 11578 19128
rect 11707 19125 11719 19128
rect 11753 19125 11765 19159
rect 11707 19119 11765 19125
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 13081 19159 13139 19165
rect 13081 19156 13093 19159
rect 12492 19128 13093 19156
rect 12492 19116 12498 19128
rect 13081 19125 13093 19128
rect 13127 19125 13139 19159
rect 13081 19119 13139 19125
rect 13998 19116 14004 19168
rect 14056 19156 14062 19168
rect 18325 19159 18383 19165
rect 18325 19156 18337 19159
rect 14056 19128 18337 19156
rect 14056 19116 14062 19128
rect 18325 19125 18337 19128
rect 18371 19125 18383 19159
rect 18325 19119 18383 19125
rect 18506 19116 18512 19168
rect 18564 19156 18570 19168
rect 21634 19156 21640 19168
rect 18564 19128 21640 19156
rect 18564 19116 18570 19128
rect 21634 19116 21640 19128
rect 21692 19116 21698 19168
rect 22066 19156 22094 19264
rect 23566 19252 23572 19264
rect 23624 19252 23630 19304
rect 23676 19264 24164 19292
rect 22370 19184 22376 19236
rect 22428 19224 22434 19236
rect 22465 19227 22523 19233
rect 22465 19224 22477 19227
rect 22428 19196 22477 19224
rect 22428 19184 22434 19196
rect 22465 19193 22477 19196
rect 22511 19193 22523 19227
rect 22465 19187 22523 19193
rect 22738 19184 22744 19236
rect 22796 19224 22802 19236
rect 22922 19224 22928 19236
rect 22796 19196 22928 19224
rect 22796 19184 22802 19196
rect 22922 19184 22928 19196
rect 22980 19184 22986 19236
rect 23676 19156 23704 19264
rect 24026 19184 24032 19236
rect 24084 19184 24090 19236
rect 24136 19224 24164 19264
rect 24394 19252 24400 19304
rect 24452 19292 24458 19304
rect 24489 19295 24547 19301
rect 24489 19292 24501 19295
rect 24452 19264 24501 19292
rect 24452 19252 24458 19264
rect 24489 19261 24501 19264
rect 24535 19261 24547 19295
rect 24489 19255 24547 19261
rect 25225 19295 25283 19301
rect 25225 19261 25237 19295
rect 25271 19292 25283 19295
rect 25590 19292 25596 19304
rect 25271 19264 25596 19292
rect 25271 19261 25283 19264
rect 25225 19255 25283 19261
rect 25590 19252 25596 19264
rect 25648 19252 25654 19304
rect 26697 19295 26755 19301
rect 26697 19261 26709 19295
rect 26743 19292 26755 19295
rect 26970 19292 26976 19304
rect 26743 19264 26976 19292
rect 26743 19261 26755 19264
rect 26697 19255 26755 19261
rect 26970 19252 26976 19264
rect 27028 19252 27034 19304
rect 27433 19295 27491 19301
rect 27433 19261 27445 19295
rect 27479 19292 27491 19295
rect 27479 19264 29040 19292
rect 27479 19261 27491 19264
rect 27433 19255 27491 19261
rect 24136 19196 24532 19224
rect 24504 19168 24532 19196
rect 28534 19184 28540 19236
rect 28592 19184 28598 19236
rect 22066 19128 23704 19156
rect 24118 19116 24124 19168
rect 24176 19116 24182 19168
rect 24486 19116 24492 19168
rect 24544 19116 24550 19168
rect 24946 19116 24952 19168
rect 25004 19165 25010 19168
rect 25004 19119 25013 19165
rect 25004 19116 25010 19119
rect 25314 19116 25320 19168
rect 25372 19156 25378 19168
rect 26329 19159 26387 19165
rect 26329 19156 26341 19159
rect 25372 19128 26341 19156
rect 25372 19116 25378 19128
rect 26329 19125 26341 19128
rect 26375 19125 26387 19159
rect 26329 19119 26387 19125
rect 27163 19159 27221 19165
rect 27163 19125 27175 19159
rect 27209 19156 27221 19159
rect 28552 19156 28580 19184
rect 27209 19128 28580 19156
rect 29012 19156 29040 19264
rect 29270 19252 29276 19304
rect 29328 19292 29334 19304
rect 29457 19295 29515 19301
rect 29457 19292 29469 19295
rect 29328 19264 29469 19292
rect 29328 19252 29334 19264
rect 29457 19261 29469 19264
rect 29503 19261 29515 19295
rect 29457 19255 29515 19261
rect 29825 19295 29883 19301
rect 29825 19261 29837 19295
rect 29871 19292 29883 19295
rect 30024 19292 30052 19400
rect 30668 19372 30696 19468
rect 30650 19320 30656 19372
rect 30708 19320 30714 19372
rect 29871 19264 30052 19292
rect 29871 19261 29883 19264
rect 29825 19255 29883 19261
rect 29086 19184 29092 19236
rect 29144 19184 29150 19236
rect 30006 19224 30012 19236
rect 29840 19196 30012 19224
rect 29840 19156 29868 19196
rect 30006 19184 30012 19196
rect 30064 19184 30070 19236
rect 30193 19227 30251 19233
rect 30193 19193 30205 19227
rect 30239 19224 30251 19227
rect 30466 19224 30472 19236
rect 30239 19196 30472 19224
rect 30239 19193 30251 19196
rect 30193 19187 30251 19193
rect 30466 19184 30472 19196
rect 30524 19184 30530 19236
rect 29012 19128 29868 19156
rect 27209 19125 27221 19128
rect 27163 19119 27221 19125
rect 30282 19116 30288 19168
rect 30340 19116 30346 19168
rect 552 19066 31072 19088
rect 552 19014 7988 19066
rect 8040 19014 8052 19066
rect 8104 19014 8116 19066
rect 8168 19014 8180 19066
rect 8232 19014 8244 19066
rect 8296 19014 15578 19066
rect 15630 19014 15642 19066
rect 15694 19014 15706 19066
rect 15758 19014 15770 19066
rect 15822 19014 15834 19066
rect 15886 19014 23168 19066
rect 23220 19014 23232 19066
rect 23284 19014 23296 19066
rect 23348 19014 23360 19066
rect 23412 19014 23424 19066
rect 23476 19014 30758 19066
rect 30810 19014 30822 19066
rect 30874 19014 30886 19066
rect 30938 19014 30950 19066
rect 31002 19014 31014 19066
rect 31066 19014 31072 19066
rect 552 18992 31072 19014
rect 1578 18912 1584 18964
rect 1636 18952 1642 18964
rect 1771 18955 1829 18961
rect 1771 18952 1783 18955
rect 1636 18924 1783 18952
rect 1636 18912 1642 18924
rect 1771 18921 1783 18924
rect 1817 18921 1829 18955
rect 4985 18955 5043 18961
rect 1771 18915 1829 18921
rect 3068 18924 4936 18952
rect 1213 18819 1271 18825
rect 1213 18785 1225 18819
rect 1259 18816 1271 18819
rect 3068 18816 3096 18924
rect 3694 18816 3700 18828
rect 1259 18788 3096 18816
rect 3160 18788 3700 18816
rect 1259 18785 1271 18788
rect 1213 18779 1271 18785
rect 1302 18708 1308 18760
rect 1360 18708 1366 18760
rect 1811 18751 1869 18757
rect 1811 18717 1823 18751
rect 1857 18748 1869 18751
rect 1946 18748 1952 18760
rect 1857 18720 1952 18748
rect 1857 18717 1869 18720
rect 1811 18711 1869 18717
rect 1946 18708 1952 18720
rect 2004 18708 2010 18760
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18748 2099 18751
rect 3160 18748 3188 18788
rect 3694 18776 3700 18788
rect 3752 18776 3758 18828
rect 3970 18776 3976 18828
rect 4028 18816 4034 18828
rect 4065 18819 4123 18825
rect 4065 18816 4077 18819
rect 4028 18788 4077 18816
rect 4028 18776 4034 18788
rect 4065 18785 4077 18788
rect 4111 18785 4123 18819
rect 4065 18779 4123 18785
rect 4349 18823 4407 18829
rect 4349 18789 4361 18823
rect 4395 18820 4407 18823
rect 4448 18820 4476 18924
rect 4908 18884 4936 18924
rect 4985 18921 4997 18955
rect 5031 18952 5043 18955
rect 5534 18952 5540 18964
rect 5031 18924 5540 18952
rect 5031 18921 5043 18924
rect 4985 18915 5043 18921
rect 5534 18912 5540 18924
rect 5592 18912 5598 18964
rect 5902 18912 5908 18964
rect 5960 18952 5966 18964
rect 6178 18952 6184 18964
rect 5960 18924 6184 18952
rect 5960 18912 5966 18924
rect 6178 18912 6184 18924
rect 6236 18912 6242 18964
rect 7466 18912 7472 18964
rect 7524 18952 7530 18964
rect 9858 18952 9864 18964
rect 7524 18924 9864 18952
rect 7524 18912 7530 18924
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 11517 18955 11575 18961
rect 11517 18921 11529 18955
rect 11563 18952 11575 18955
rect 13906 18952 13912 18964
rect 11563 18924 13912 18952
rect 11563 18921 11575 18924
rect 11517 18915 11575 18921
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 15841 18955 15899 18961
rect 14016 18924 15332 18952
rect 5629 18887 5687 18893
rect 5629 18884 5641 18887
rect 4908 18856 5641 18884
rect 5629 18853 5641 18856
rect 5675 18853 5687 18887
rect 5629 18847 5687 18853
rect 8021 18887 8079 18893
rect 8021 18853 8033 18887
rect 8067 18884 8079 18887
rect 8570 18884 8576 18896
rect 8067 18856 8576 18884
rect 8067 18853 8079 18856
rect 8021 18847 8079 18853
rect 4395 18792 4476 18820
rect 4617 18819 4675 18825
rect 4617 18816 4629 18819
rect 4395 18789 4407 18792
rect 4349 18783 4407 18789
rect 4540 18788 4629 18816
rect 2087 18720 3188 18748
rect 2087 18717 2099 18720
rect 2041 18711 2099 18717
rect 3418 18708 3424 18760
rect 3476 18748 3482 18760
rect 4154 18748 4160 18760
rect 3476 18720 4160 18748
rect 3476 18708 3482 18720
rect 4154 18708 4160 18720
rect 4212 18708 4218 18760
rect 4540 18748 4568 18788
rect 4617 18785 4629 18788
rect 4663 18785 4675 18819
rect 4617 18779 4675 18785
rect 4890 18776 4896 18828
rect 4948 18776 4954 18828
rect 5169 18819 5227 18825
rect 5169 18785 5181 18819
rect 5215 18785 5227 18819
rect 5169 18779 5227 18785
rect 4356 18720 4568 18748
rect 4356 18692 4384 18720
rect 3510 18640 3516 18692
rect 3568 18680 3574 18692
rect 3881 18683 3939 18689
rect 3881 18680 3893 18683
rect 3568 18652 3893 18680
rect 3568 18640 3574 18652
rect 3881 18649 3893 18652
rect 3927 18649 3939 18683
rect 3881 18643 3939 18649
rect 4338 18640 4344 18692
rect 4396 18640 4402 18692
rect 4433 18683 4491 18689
rect 4433 18649 4445 18683
rect 4479 18680 4491 18683
rect 4522 18680 4528 18692
rect 4479 18652 4528 18680
rect 4479 18649 4491 18652
rect 4433 18643 4491 18649
rect 4522 18640 4528 18652
rect 4580 18640 4586 18692
rect 4614 18640 4620 18692
rect 4672 18640 4678 18692
rect 4706 18640 4712 18692
rect 4764 18640 4770 18692
rect 5184 18680 5212 18779
rect 5442 18776 5448 18828
rect 5500 18776 5506 18828
rect 4816 18652 5212 18680
rect 1026 18572 1032 18624
rect 1084 18572 1090 18624
rect 3326 18572 3332 18624
rect 3384 18572 3390 18624
rect 3694 18572 3700 18624
rect 3752 18572 3758 18624
rect 4157 18615 4215 18621
rect 4157 18581 4169 18615
rect 4203 18612 4215 18615
rect 4632 18612 4660 18640
rect 4816 18624 4844 18652
rect 4203 18584 4660 18612
rect 4203 18581 4215 18584
rect 4157 18575 4215 18581
rect 4798 18572 4804 18624
rect 4856 18572 4862 18624
rect 5644 18612 5672 18847
rect 8570 18844 8576 18856
rect 8628 18844 8634 18896
rect 8662 18844 8668 18896
rect 8720 18884 8726 18896
rect 8720 18856 8800 18884
rect 8720 18844 8726 18856
rect 5902 18776 5908 18828
rect 5960 18776 5966 18828
rect 6454 18776 6460 18828
rect 6512 18816 6518 18828
rect 6641 18819 6699 18825
rect 6641 18816 6653 18819
rect 6512 18788 6653 18816
rect 6512 18776 6518 18788
rect 6641 18785 6653 18788
rect 6687 18785 6699 18819
rect 6641 18779 6699 18785
rect 8205 18819 8263 18825
rect 8205 18785 8217 18819
rect 8251 18785 8263 18819
rect 8772 18816 8800 18856
rect 10778 18844 10784 18896
rect 10836 18844 10842 18896
rect 11241 18887 11299 18893
rect 11241 18853 11253 18887
rect 11287 18884 11299 18887
rect 11606 18884 11612 18896
rect 11287 18856 11612 18884
rect 11287 18853 11299 18856
rect 11241 18847 11299 18853
rect 11606 18844 11612 18856
rect 11664 18844 11670 18896
rect 14016 18884 14044 18924
rect 15304 18896 15332 18924
rect 15841 18921 15853 18955
rect 15887 18952 15899 18955
rect 16390 18952 16396 18964
rect 15887 18924 16396 18952
rect 15887 18921 15899 18924
rect 15841 18915 15899 18921
rect 16390 18912 16396 18924
rect 16448 18912 16454 18964
rect 16761 18955 16819 18961
rect 16761 18921 16773 18955
rect 16807 18921 16819 18955
rect 16761 18915 16819 18921
rect 13188 18856 14044 18884
rect 8992 18819 9050 18825
rect 8992 18816 9004 18819
rect 8772 18788 9004 18816
rect 8205 18779 8263 18785
rect 8992 18785 9004 18788
rect 9038 18785 9050 18819
rect 10965 18819 11023 18825
rect 8992 18779 9050 18785
rect 9324 18788 10548 18816
rect 6178 18708 6184 18760
rect 6236 18757 6242 18760
rect 6236 18751 6290 18757
rect 6236 18717 6244 18751
rect 6278 18717 6290 18751
rect 6236 18711 6290 18717
rect 6236 18708 6242 18711
rect 6362 18708 6368 18760
rect 6420 18708 6426 18760
rect 7466 18708 7472 18760
rect 7524 18748 7530 18760
rect 7742 18748 7748 18760
rect 7524 18720 7748 18748
rect 7524 18708 7530 18720
rect 7742 18708 7748 18720
rect 7800 18708 7806 18760
rect 8220 18624 8248 18779
rect 9128 18769 9186 18775
rect 8665 18751 8723 18757
rect 8665 18717 8677 18751
rect 8711 18717 8723 18751
rect 9128 18735 9140 18769
rect 9174 18748 9186 18769
rect 9324 18748 9352 18788
rect 10520 18760 10548 18788
rect 10965 18785 10977 18819
rect 11011 18785 11023 18819
rect 11701 18819 11759 18825
rect 11701 18816 11713 18819
rect 10965 18779 11023 18785
rect 11256 18788 11713 18816
rect 9174 18735 9352 18748
rect 9128 18729 9352 18735
rect 9143 18720 9352 18729
rect 8665 18711 8723 18717
rect 8294 18640 8300 18692
rect 8352 18680 8358 18692
rect 8352 18652 8616 18680
rect 8352 18640 8358 18652
rect 8588 18624 8616 18652
rect 8202 18612 8208 18624
rect 5644 18584 8208 18612
rect 8202 18572 8208 18584
rect 8260 18572 8266 18624
rect 8478 18572 8484 18624
rect 8536 18572 8542 18624
rect 8570 18572 8576 18624
rect 8628 18572 8634 18624
rect 8680 18612 8708 18711
rect 9398 18708 9404 18760
rect 9456 18708 9462 18760
rect 9582 18708 9588 18760
rect 9640 18748 9646 18760
rect 9640 18720 10186 18748
rect 9640 18708 9646 18720
rect 9490 18612 9496 18624
rect 8680 18584 9496 18612
rect 9490 18572 9496 18584
rect 9548 18572 9554 18624
rect 10158 18612 10186 18720
rect 10502 18708 10508 18760
rect 10560 18708 10566 18760
rect 10226 18640 10232 18692
rect 10284 18680 10290 18692
rect 10686 18680 10692 18692
rect 10284 18652 10692 18680
rect 10284 18640 10290 18652
rect 10686 18640 10692 18652
rect 10744 18680 10750 18692
rect 10980 18680 11008 18779
rect 11256 18760 11284 18788
rect 11701 18785 11713 18788
rect 11747 18785 11759 18819
rect 13188 18816 13216 18856
rect 15286 18844 15292 18896
rect 15344 18844 15350 18896
rect 16114 18844 16120 18896
rect 16172 18884 16178 18896
rect 16776 18884 16804 18915
rect 18414 18912 18420 18964
rect 18472 18952 18478 18964
rect 20257 18955 20315 18961
rect 18472 18924 19656 18952
rect 18472 18912 18478 18924
rect 16172 18856 16804 18884
rect 16172 18844 16178 18856
rect 18506 18844 18512 18896
rect 18564 18844 18570 18896
rect 19628 18884 19656 18924
rect 20257 18921 20269 18955
rect 20303 18952 20315 18955
rect 20714 18952 20720 18964
rect 20303 18924 20720 18952
rect 20303 18921 20315 18924
rect 20257 18915 20315 18921
rect 20714 18912 20720 18924
rect 20772 18912 20778 18964
rect 20824 18924 22968 18952
rect 20824 18884 20852 18924
rect 19628 18856 20852 18884
rect 22554 18844 22560 18896
rect 22612 18844 22618 18896
rect 22940 18884 22968 18924
rect 23014 18912 23020 18964
rect 23072 18952 23078 18964
rect 23385 18955 23443 18961
rect 23385 18952 23397 18955
rect 23072 18924 23397 18952
rect 23072 18912 23078 18924
rect 23385 18921 23397 18924
rect 23431 18921 23443 18955
rect 23385 18915 23443 18921
rect 24587 18955 24645 18961
rect 24587 18921 24599 18955
rect 24633 18952 24645 18955
rect 24946 18952 24952 18964
rect 24633 18924 24952 18952
rect 24633 18921 24645 18924
rect 24587 18915 24645 18921
rect 24946 18912 24952 18924
rect 25004 18912 25010 18964
rect 26436 18924 28994 18952
rect 22940 18856 24164 18884
rect 11701 18779 11759 18785
rect 12452 18788 13216 18816
rect 11238 18708 11244 18760
rect 11296 18708 11302 18760
rect 11514 18708 11520 18760
rect 11572 18748 11578 18760
rect 12158 18757 12164 18760
rect 11793 18751 11851 18757
rect 11793 18748 11805 18751
rect 11572 18720 11805 18748
rect 11572 18708 11578 18720
rect 11793 18717 11805 18720
rect 11839 18717 11851 18751
rect 11793 18711 11851 18717
rect 12120 18751 12164 18757
rect 12120 18717 12132 18751
rect 12120 18711 12164 18717
rect 12158 18708 12164 18711
rect 12216 18708 12222 18760
rect 12299 18751 12357 18757
rect 12299 18717 12311 18751
rect 12345 18748 12357 18751
rect 12452 18748 12480 18788
rect 14182 18776 14188 18828
rect 14240 18776 14246 18828
rect 14277 18819 14335 18825
rect 14277 18785 14289 18819
rect 14323 18816 14335 18819
rect 14366 18816 14372 18828
rect 14323 18788 14372 18816
rect 14323 18785 14335 18788
rect 14277 18779 14335 18785
rect 14366 18776 14372 18788
rect 14424 18776 14430 18828
rect 15930 18816 15936 18828
rect 14476 18788 15936 18816
rect 12345 18720 12480 18748
rect 12529 18751 12587 18757
rect 12345 18717 12357 18720
rect 12299 18711 12357 18717
rect 12529 18717 12541 18751
rect 12575 18748 12587 18751
rect 12894 18748 12900 18760
rect 12575 18720 12900 18748
rect 12575 18717 12587 18720
rect 12529 18711 12587 18717
rect 12894 18708 12900 18720
rect 12952 18708 12958 18760
rect 14476 18748 14504 18788
rect 15930 18776 15936 18788
rect 15988 18776 15994 18828
rect 16298 18776 16304 18828
rect 16356 18776 16362 18828
rect 16485 18819 16543 18825
rect 16485 18785 16497 18819
rect 16531 18816 16543 18819
rect 16666 18816 16672 18828
rect 16531 18788 16672 18816
rect 16531 18785 16543 18788
rect 16485 18779 16543 18785
rect 16666 18776 16672 18788
rect 16724 18776 16730 18828
rect 16942 18776 16948 18828
rect 17000 18776 17006 18828
rect 18524 18816 18552 18844
rect 17052 18788 18552 18816
rect 18601 18819 18659 18825
rect 14016 18720 14504 18748
rect 14553 18751 14611 18757
rect 14016 18689 14044 18720
rect 14553 18717 14565 18751
rect 14599 18748 14611 18751
rect 15010 18748 15016 18760
rect 14599 18720 15016 18748
rect 14599 18717 14611 18720
rect 14553 18711 14611 18717
rect 15010 18708 15016 18720
rect 15068 18708 15074 18760
rect 10744 18652 11008 18680
rect 14001 18683 14059 18689
rect 10744 18640 10750 18652
rect 14001 18649 14013 18683
rect 14047 18649 14059 18683
rect 16316 18680 16344 18776
rect 16390 18708 16396 18760
rect 16448 18748 16454 18760
rect 16577 18751 16635 18757
rect 16577 18748 16589 18751
rect 16448 18720 16589 18748
rect 16448 18708 16454 18720
rect 16577 18717 16589 18720
rect 16623 18748 16635 18751
rect 17052 18748 17080 18788
rect 18601 18785 18613 18819
rect 18647 18816 18659 18819
rect 18969 18819 19027 18825
rect 18969 18816 18981 18819
rect 18647 18788 18981 18816
rect 18647 18785 18659 18788
rect 18601 18779 18659 18785
rect 18969 18785 18981 18788
rect 19015 18785 19027 18819
rect 18969 18779 19027 18785
rect 20438 18776 20444 18828
rect 20496 18816 20502 18828
rect 20533 18819 20591 18825
rect 20533 18816 20545 18819
rect 20496 18788 20545 18816
rect 20496 18776 20502 18788
rect 20533 18785 20545 18788
rect 20579 18785 20591 18819
rect 21545 18819 21603 18825
rect 21545 18816 21557 18819
rect 20533 18779 20591 18785
rect 20640 18788 21557 18816
rect 16623 18720 17080 18748
rect 17221 18751 17279 18757
rect 16623 18717 16635 18720
rect 16577 18711 16635 18717
rect 17221 18717 17233 18751
rect 17267 18748 17279 18751
rect 17678 18748 17684 18760
rect 17267 18720 17684 18748
rect 17267 18717 17279 18720
rect 17221 18711 17279 18717
rect 17678 18708 17684 18720
rect 17736 18708 17742 18760
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18717 18751 18751
rect 18693 18711 18751 18717
rect 16666 18680 16672 18692
rect 16316 18652 16672 18680
rect 14001 18643 14059 18649
rect 16666 18640 16672 18652
rect 16724 18640 16730 18692
rect 18708 18624 18736 18711
rect 20346 18708 20352 18760
rect 20404 18748 20410 18760
rect 20640 18748 20668 18788
rect 21545 18785 21557 18788
rect 21591 18785 21603 18819
rect 21545 18779 21603 18785
rect 21634 18776 21640 18828
rect 21692 18816 21698 18828
rect 22572 18816 22600 18844
rect 23477 18819 23535 18825
rect 23477 18816 23489 18819
rect 21692 18788 22094 18816
rect 22572 18788 23489 18816
rect 21692 18776 21698 18788
rect 20404 18720 20668 18748
rect 21269 18751 21327 18757
rect 20404 18708 20410 18720
rect 21269 18717 21281 18751
rect 21315 18717 21327 18751
rect 22066 18748 22094 18788
rect 23477 18785 23489 18788
rect 23523 18785 23535 18819
rect 23477 18779 23535 18785
rect 23934 18776 23940 18828
rect 23992 18816 23998 18828
rect 24029 18819 24087 18825
rect 24029 18816 24041 18819
rect 23992 18788 24041 18816
rect 23992 18776 23998 18788
rect 24029 18785 24041 18788
rect 24075 18785 24087 18819
rect 24136 18816 24164 18856
rect 24857 18819 24915 18825
rect 24136 18788 24348 18816
rect 24029 18779 24087 18785
rect 24320 18760 24348 18788
rect 24857 18785 24869 18819
rect 24903 18816 24915 18819
rect 26436 18816 26464 18924
rect 28966 18884 28994 18924
rect 28966 18856 29776 18884
rect 29748 18828 29776 18856
rect 24903 18788 26464 18816
rect 24903 18785 24915 18788
rect 24857 18779 24915 18785
rect 26602 18776 26608 18828
rect 26660 18776 26666 18828
rect 26694 18776 26700 18828
rect 26752 18816 26758 18828
rect 27116 18819 27174 18825
rect 27116 18816 27128 18819
rect 26752 18788 27128 18816
rect 26752 18776 26758 18788
rect 27116 18785 27128 18788
rect 27162 18785 27174 18819
rect 28997 18819 29055 18825
rect 27116 18779 27174 18785
rect 27448 18788 28304 18816
rect 23661 18751 23719 18757
rect 22066 18720 23520 18748
rect 21269 18711 21327 18717
rect 20438 18640 20444 18692
rect 20496 18680 20502 18692
rect 21284 18680 21312 18711
rect 23492 18692 23520 18720
rect 23661 18717 23673 18751
rect 23707 18748 23719 18751
rect 23842 18748 23848 18760
rect 23707 18720 23848 18748
rect 23707 18717 23719 18720
rect 23661 18711 23719 18717
rect 23842 18708 23848 18720
rect 23900 18708 23906 18760
rect 24121 18751 24179 18757
rect 24121 18717 24133 18751
rect 24167 18717 24179 18751
rect 24121 18711 24179 18717
rect 20496 18652 21312 18680
rect 20496 18640 20502 18652
rect 22738 18640 22744 18692
rect 22796 18680 22802 18692
rect 23017 18683 23075 18689
rect 23017 18680 23029 18683
rect 22796 18652 23029 18680
rect 22796 18640 22802 18652
rect 23017 18649 23029 18652
rect 23063 18649 23075 18683
rect 23017 18643 23075 18649
rect 23474 18640 23480 18692
rect 23532 18640 23538 18692
rect 11146 18612 11152 18624
rect 10158 18584 11152 18612
rect 11146 18572 11152 18584
rect 11204 18572 11210 18624
rect 13814 18572 13820 18624
rect 13872 18572 13878 18624
rect 18690 18572 18696 18624
rect 18748 18612 18754 18624
rect 20625 18615 20683 18621
rect 20625 18612 20637 18615
rect 18748 18584 20637 18612
rect 18748 18572 18754 18584
rect 20625 18581 20637 18584
rect 20671 18581 20683 18615
rect 20625 18575 20683 18581
rect 20714 18572 20720 18624
rect 20772 18612 20778 18624
rect 22649 18615 22707 18621
rect 22649 18612 22661 18615
rect 20772 18584 22661 18612
rect 20772 18572 20778 18584
rect 22649 18581 22661 18584
rect 22695 18581 22707 18615
rect 22649 18575 22707 18581
rect 22922 18572 22928 18624
rect 22980 18612 22986 18624
rect 23845 18615 23903 18621
rect 23845 18612 23857 18615
rect 22980 18584 23857 18612
rect 22980 18572 22986 18584
rect 23845 18581 23857 18584
rect 23891 18581 23903 18615
rect 24136 18612 24164 18711
rect 24302 18708 24308 18760
rect 24360 18708 24366 18760
rect 24578 18708 24584 18760
rect 24636 18708 24642 18760
rect 26418 18708 26424 18760
rect 26476 18748 26482 18760
rect 26789 18751 26847 18757
rect 26789 18748 26801 18751
rect 26476 18720 26801 18748
rect 26476 18708 26482 18720
rect 26789 18717 26801 18720
rect 26835 18717 26847 18751
rect 26789 18711 26847 18717
rect 27295 18751 27353 18757
rect 27295 18717 27307 18751
rect 27341 18748 27353 18751
rect 27448 18748 27476 18788
rect 28276 18760 28304 18788
rect 28997 18785 29009 18819
rect 29043 18816 29055 18819
rect 29178 18816 29184 18828
rect 29043 18788 29184 18816
rect 29043 18785 29055 18788
rect 28997 18779 29055 18785
rect 29178 18776 29184 18788
rect 29236 18776 29242 18828
rect 29273 18819 29331 18825
rect 29273 18785 29285 18819
rect 29319 18816 29331 18819
rect 29362 18816 29368 18828
rect 29319 18788 29368 18816
rect 29319 18785 29331 18788
rect 29273 18779 29331 18785
rect 29362 18776 29368 18788
rect 29420 18776 29426 18828
rect 29730 18776 29736 18828
rect 29788 18776 29794 18828
rect 30101 18819 30159 18825
rect 30101 18785 30113 18819
rect 30147 18785 30159 18819
rect 30101 18779 30159 18785
rect 27341 18720 27476 18748
rect 27525 18751 27583 18757
rect 27341 18717 27353 18720
rect 27295 18711 27353 18717
rect 27525 18717 27537 18751
rect 27571 18748 27583 18751
rect 27571 18720 28212 18748
rect 27571 18717 27583 18720
rect 27525 18711 27583 18717
rect 26050 18680 26056 18692
rect 25516 18652 26056 18680
rect 24394 18612 24400 18624
rect 24136 18584 24400 18612
rect 23845 18575 23903 18581
rect 24394 18572 24400 18584
rect 24452 18612 24458 18624
rect 25516 18612 25544 18652
rect 26050 18640 26056 18652
rect 26108 18680 26114 18692
rect 26436 18680 26464 18708
rect 26108 18652 26464 18680
rect 28184 18680 28212 18720
rect 28258 18708 28264 18760
rect 28316 18708 28322 18760
rect 30116 18680 30144 18779
rect 30190 18776 30196 18828
rect 30248 18816 30254 18828
rect 30561 18819 30619 18825
rect 30561 18816 30573 18819
rect 30248 18788 30573 18816
rect 30248 18776 30254 18788
rect 30561 18785 30573 18788
rect 30607 18785 30619 18819
rect 30561 18779 30619 18785
rect 28184 18652 29132 18680
rect 26108 18640 26114 18652
rect 24452 18584 25544 18612
rect 24452 18572 24458 18584
rect 25958 18572 25964 18624
rect 26016 18572 26022 18624
rect 26418 18572 26424 18624
rect 26476 18572 26482 18624
rect 27706 18572 27712 18624
rect 27764 18612 27770 18624
rect 28629 18615 28687 18621
rect 28629 18612 28641 18615
rect 27764 18584 28641 18612
rect 27764 18572 27770 18584
rect 28629 18581 28641 18584
rect 28675 18581 28687 18615
rect 29104 18612 29132 18652
rect 29748 18652 30144 18680
rect 29748 18624 29776 18652
rect 29270 18612 29276 18624
rect 29104 18584 29276 18612
rect 28629 18575 28687 18581
rect 29270 18572 29276 18584
rect 29328 18572 29334 18624
rect 29730 18572 29736 18624
rect 29788 18572 29794 18624
rect 30282 18572 30288 18624
rect 30340 18572 30346 18624
rect 30377 18615 30435 18621
rect 30377 18581 30389 18615
rect 30423 18612 30435 18615
rect 30423 18584 30972 18612
rect 30423 18581 30435 18584
rect 30377 18575 30435 18581
rect 552 18522 30912 18544
rect 552 18470 4193 18522
rect 4245 18470 4257 18522
rect 4309 18470 4321 18522
rect 4373 18470 4385 18522
rect 4437 18470 4449 18522
rect 4501 18470 11783 18522
rect 11835 18470 11847 18522
rect 11899 18470 11911 18522
rect 11963 18470 11975 18522
rect 12027 18470 12039 18522
rect 12091 18470 19373 18522
rect 19425 18470 19437 18522
rect 19489 18470 19501 18522
rect 19553 18470 19565 18522
rect 19617 18470 19629 18522
rect 19681 18470 26963 18522
rect 27015 18470 27027 18522
rect 27079 18470 27091 18522
rect 27143 18470 27155 18522
rect 27207 18470 27219 18522
rect 27271 18470 30912 18522
rect 552 18448 30912 18470
rect 1210 18368 1216 18420
rect 1268 18408 1274 18420
rect 1268 18380 2360 18408
rect 1268 18368 1274 18380
rect 2332 18340 2360 18380
rect 2774 18368 2780 18420
rect 2832 18368 2838 18420
rect 3418 18408 3424 18420
rect 3252 18380 3424 18408
rect 3252 18340 3280 18380
rect 3418 18368 3424 18380
rect 3476 18368 3482 18420
rect 3970 18368 3976 18420
rect 4028 18408 4034 18420
rect 4798 18408 4804 18420
rect 4028 18380 4804 18408
rect 4028 18368 4034 18380
rect 4798 18368 4804 18380
rect 4856 18368 4862 18420
rect 5077 18411 5135 18417
rect 5077 18377 5089 18411
rect 5123 18408 5135 18411
rect 5166 18408 5172 18420
rect 5123 18380 5172 18408
rect 5123 18377 5135 18380
rect 5077 18371 5135 18377
rect 5166 18368 5172 18380
rect 5224 18368 5230 18420
rect 5258 18368 5264 18420
rect 5316 18408 5322 18420
rect 5537 18411 5595 18417
rect 5537 18408 5549 18411
rect 5316 18380 5549 18408
rect 5316 18368 5322 18380
rect 5537 18377 5549 18380
rect 5583 18377 5595 18411
rect 5537 18371 5595 18377
rect 5626 18368 5632 18420
rect 5684 18368 5690 18420
rect 5813 18411 5871 18417
rect 5813 18377 5825 18411
rect 5859 18408 5871 18411
rect 6730 18408 6736 18420
rect 5859 18380 6736 18408
rect 5859 18377 5871 18380
rect 5813 18371 5871 18377
rect 6730 18368 6736 18380
rect 6788 18368 6794 18420
rect 6914 18368 6920 18420
rect 6972 18408 6978 18420
rect 8846 18408 8852 18420
rect 6972 18380 8852 18408
rect 6972 18368 6978 18380
rect 8846 18368 8852 18380
rect 8904 18368 8910 18420
rect 9582 18368 9588 18420
rect 9640 18408 9646 18420
rect 9640 18380 10548 18408
rect 9640 18368 9646 18380
rect 2332 18312 3280 18340
rect 5644 18340 5672 18368
rect 5902 18340 5908 18352
rect 5644 18312 5908 18340
rect 1443 18275 1501 18281
rect 1443 18241 1455 18275
rect 1489 18272 1501 18275
rect 2958 18272 2964 18284
rect 1489 18244 2964 18272
rect 1489 18241 1501 18244
rect 1443 18235 1501 18241
rect 2958 18232 2964 18244
rect 3016 18232 3022 18284
rect 3252 18281 3280 18312
rect 5902 18300 5908 18312
rect 5960 18300 5966 18352
rect 8478 18300 8484 18352
rect 8536 18300 8542 18352
rect 3237 18275 3295 18281
rect 3237 18241 3249 18275
rect 3283 18241 3295 18275
rect 3700 18275 3758 18281
rect 3700 18272 3712 18275
rect 3237 18235 3295 18241
rect 3528 18244 3712 18272
rect 3528 18216 3556 18244
rect 3700 18241 3712 18244
rect 3746 18241 3758 18275
rect 3700 18235 3758 18241
rect 3878 18232 3884 18284
rect 3936 18272 3942 18284
rect 5534 18272 5540 18284
rect 3936 18244 5540 18272
rect 3936 18232 3942 18244
rect 5534 18232 5540 18244
rect 5592 18232 5598 18284
rect 5626 18232 5632 18284
rect 5684 18272 5690 18284
rect 6552 18275 6610 18281
rect 6552 18272 6564 18275
rect 5684 18244 6564 18272
rect 5684 18232 5690 18244
rect 6552 18241 6564 18244
rect 6598 18241 6610 18275
rect 6552 18235 6610 18241
rect 8294 18232 8300 18284
rect 8352 18232 8358 18284
rect 8496 18272 8524 18300
rect 8944 18275 9002 18281
rect 8944 18272 8956 18275
rect 8496 18244 8956 18272
rect 8944 18241 8956 18244
rect 8990 18241 9002 18275
rect 8944 18235 9002 18241
rect 9674 18232 9680 18284
rect 9732 18272 9738 18284
rect 9732 18244 10088 18272
rect 9732 18232 9738 18244
rect 937 18207 995 18213
rect 937 18173 949 18207
rect 983 18204 995 18207
rect 1210 18204 1216 18216
rect 983 18176 1216 18204
rect 983 18173 995 18176
rect 937 18167 995 18173
rect 1210 18164 1216 18176
rect 1268 18164 1274 18216
rect 1673 18207 1731 18213
rect 1673 18173 1685 18207
rect 1719 18204 1731 18207
rect 2682 18204 2688 18216
rect 1719 18176 2688 18204
rect 1719 18173 1731 18176
rect 1673 18167 1731 18173
rect 2682 18164 2688 18176
rect 2740 18164 2746 18216
rect 3510 18164 3516 18216
rect 3568 18164 3574 18216
rect 3970 18164 3976 18216
rect 4028 18164 4034 18216
rect 4062 18164 4068 18216
rect 4120 18204 4126 18216
rect 5721 18207 5779 18213
rect 4120 18176 5672 18204
rect 4120 18164 4126 18176
rect 5644 18136 5672 18176
rect 5721 18173 5733 18207
rect 5767 18204 5779 18207
rect 5994 18204 6000 18216
rect 5767 18176 6000 18204
rect 5767 18173 5779 18176
rect 5721 18167 5779 18173
rect 5994 18164 6000 18176
rect 6052 18164 6058 18216
rect 6086 18164 6092 18216
rect 6144 18164 6150 18216
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6196 18176 6837 18204
rect 6196 18136 6224 18176
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 8312 18204 8340 18232
rect 8846 18213 8852 18216
rect 8481 18207 8539 18213
rect 8481 18204 8493 18207
rect 8312 18176 8493 18204
rect 6825 18167 6883 18173
rect 8481 18173 8493 18176
rect 8527 18173 8539 18207
rect 8481 18167 8539 18173
rect 8808 18207 8852 18213
rect 8808 18173 8820 18207
rect 8808 18167 8852 18173
rect 8846 18164 8852 18167
rect 8904 18164 8910 18216
rect 9217 18207 9275 18213
rect 9217 18173 9229 18207
rect 9263 18204 9275 18207
rect 9950 18204 9956 18216
rect 9263 18176 9956 18204
rect 9263 18173 9275 18176
rect 9217 18167 9275 18173
rect 9950 18164 9956 18176
rect 10008 18164 10014 18216
rect 5644 18108 6224 18136
rect 8205 18139 8263 18145
rect 8205 18105 8217 18139
rect 8251 18136 8263 18139
rect 8570 18136 8576 18148
rect 8251 18108 8576 18136
rect 8251 18105 8263 18108
rect 8205 18099 8263 18105
rect 8570 18096 8576 18108
rect 8628 18096 8634 18148
rect 10060 18136 10088 18244
rect 10520 18204 10548 18380
rect 12526 18368 12532 18420
rect 12584 18368 12590 18420
rect 13078 18368 13084 18420
rect 13136 18368 13142 18420
rect 13446 18368 13452 18420
rect 13504 18408 13510 18420
rect 13817 18411 13875 18417
rect 13817 18408 13829 18411
rect 13504 18380 13829 18408
rect 13504 18368 13510 18380
rect 13817 18377 13829 18380
rect 13863 18377 13875 18411
rect 13817 18371 13875 18377
rect 14182 18368 14188 18420
rect 14240 18408 14246 18420
rect 16390 18408 16396 18420
rect 14240 18380 16396 18408
rect 14240 18368 14246 18380
rect 16390 18368 16396 18380
rect 16448 18368 16454 18420
rect 17678 18368 17684 18420
rect 17736 18408 17742 18420
rect 17957 18411 18015 18417
rect 17957 18408 17969 18411
rect 17736 18380 17969 18408
rect 17736 18368 17742 18380
rect 17957 18377 17969 18380
rect 18003 18377 18015 18411
rect 22554 18408 22560 18420
rect 17957 18371 18015 18377
rect 18524 18380 22560 18408
rect 10597 18275 10655 18281
rect 10597 18241 10609 18275
rect 10643 18272 10655 18275
rect 11152 18275 11210 18281
rect 11152 18272 11164 18275
rect 10643 18244 11164 18272
rect 10643 18241 10655 18244
rect 10597 18235 10655 18241
rect 11152 18241 11164 18244
rect 11198 18241 11210 18275
rect 11152 18235 11210 18241
rect 11606 18232 11612 18284
rect 11664 18232 11670 18284
rect 13722 18232 13728 18284
rect 13780 18272 13786 18284
rect 14875 18275 14933 18281
rect 13780 18244 14504 18272
rect 13780 18232 13786 18244
rect 10689 18207 10747 18213
rect 10689 18204 10701 18207
rect 10520 18176 10701 18204
rect 10689 18173 10701 18176
rect 10735 18173 10747 18207
rect 11425 18207 11483 18213
rect 11425 18204 11437 18207
rect 10689 18167 10747 18173
rect 10796 18176 11437 18204
rect 10796 18136 10824 18176
rect 11425 18173 11437 18176
rect 11471 18173 11483 18207
rect 11624 18204 11652 18232
rect 11624 18176 12112 18204
rect 11425 18167 11483 18173
rect 10060 18108 10824 18136
rect 1403 18071 1461 18077
rect 1403 18037 1415 18071
rect 1449 18068 1461 18071
rect 1670 18068 1676 18080
rect 1449 18040 1676 18068
rect 1449 18037 1461 18040
rect 1403 18031 1461 18037
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 1762 18028 1768 18080
rect 1820 18068 1826 18080
rect 3703 18071 3761 18077
rect 3703 18068 3715 18071
rect 1820 18040 3715 18068
rect 1820 18028 1826 18040
rect 3703 18037 3715 18040
rect 3749 18068 3761 18071
rect 6178 18068 6184 18080
rect 3749 18040 6184 18068
rect 3749 18037 3761 18040
rect 3703 18031 3761 18037
rect 6178 18028 6184 18040
rect 6236 18068 6242 18080
rect 6555 18071 6613 18077
rect 6555 18068 6567 18071
rect 6236 18040 6567 18068
rect 6236 18028 6242 18040
rect 6555 18037 6567 18040
rect 6601 18068 6613 18071
rect 6730 18068 6736 18080
rect 6601 18040 6736 18068
rect 6601 18037 6613 18040
rect 6555 18031 6613 18037
rect 6730 18028 6736 18040
rect 6788 18028 6794 18080
rect 7650 18028 7656 18080
rect 7708 18068 7714 18080
rect 10042 18068 10048 18080
rect 7708 18040 10048 18068
rect 7708 18028 7714 18040
rect 10042 18028 10048 18040
rect 10100 18068 10106 18080
rect 10686 18068 10692 18080
rect 10100 18040 10692 18068
rect 10100 18028 10106 18040
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 11155 18071 11213 18077
rect 11155 18037 11167 18071
rect 11201 18068 11213 18071
rect 12084 18068 12112 18176
rect 14366 18164 14372 18216
rect 14424 18164 14430 18216
rect 14476 18204 14504 18244
rect 14875 18241 14887 18275
rect 14921 18272 14933 18275
rect 16853 18275 16911 18281
rect 14921 18244 16804 18272
rect 14921 18241 14933 18244
rect 14875 18235 14933 18241
rect 15105 18207 15163 18213
rect 15105 18204 15117 18207
rect 14476 18176 15117 18204
rect 15105 18173 15117 18176
rect 15151 18173 15163 18207
rect 15105 18167 15163 18173
rect 16022 18164 16028 18216
rect 16080 18204 16086 18216
rect 16577 18207 16635 18213
rect 16577 18204 16589 18207
rect 16080 18176 16589 18204
rect 16080 18164 16086 18176
rect 16577 18173 16589 18176
rect 16623 18173 16635 18207
rect 16776 18204 16804 18244
rect 16853 18241 16865 18275
rect 16899 18272 16911 18275
rect 17218 18272 17224 18284
rect 16899 18244 17224 18272
rect 16899 18241 16911 18244
rect 16853 18235 16911 18241
rect 17218 18232 17224 18244
rect 17276 18232 17282 18284
rect 17954 18204 17960 18216
rect 16776 18176 17960 18204
rect 16577 18167 16635 18173
rect 17954 18164 17960 18176
rect 18012 18164 18018 18216
rect 18524 18213 18552 18380
rect 22554 18368 22560 18380
rect 22612 18368 22618 18420
rect 22646 18368 22652 18420
rect 22704 18408 22710 18420
rect 23385 18411 23443 18417
rect 23385 18408 23397 18411
rect 22704 18380 23397 18408
rect 22704 18368 22710 18380
rect 23385 18377 23397 18380
rect 23431 18377 23443 18411
rect 23385 18371 23443 18377
rect 24486 18368 24492 18420
rect 24544 18408 24550 18420
rect 24581 18411 24639 18417
rect 24581 18408 24593 18411
rect 24544 18380 24593 18408
rect 24544 18368 24550 18380
rect 24581 18377 24593 18380
rect 24627 18377 24639 18411
rect 26786 18408 26792 18420
rect 24581 18371 24639 18377
rect 24780 18380 26792 18408
rect 20257 18343 20315 18349
rect 20257 18309 20269 18343
rect 20303 18340 20315 18343
rect 20346 18340 20352 18352
rect 20303 18312 20352 18340
rect 20303 18309 20315 18312
rect 20257 18303 20315 18309
rect 20346 18300 20352 18312
rect 20404 18300 20410 18352
rect 22830 18300 22836 18352
rect 22888 18340 22894 18352
rect 23017 18343 23075 18349
rect 23017 18340 23029 18343
rect 22888 18312 23029 18340
rect 22888 18300 22894 18312
rect 23017 18309 23029 18312
rect 23063 18309 23075 18343
rect 23017 18303 23075 18309
rect 24213 18343 24271 18349
rect 24213 18309 24225 18343
rect 24259 18340 24271 18343
rect 24780 18340 24808 18380
rect 26786 18368 26792 18380
rect 26844 18368 26850 18420
rect 30944 18408 30972 18584
rect 28368 18380 30972 18408
rect 24259 18312 24808 18340
rect 24259 18309 24271 18312
rect 24213 18303 24271 18309
rect 18598 18232 18604 18284
rect 18656 18272 18662 18284
rect 18969 18275 19027 18281
rect 18969 18272 18981 18275
rect 18656 18244 18981 18272
rect 18656 18232 18662 18244
rect 18969 18241 18981 18244
rect 19015 18241 19027 18275
rect 18969 18235 19027 18241
rect 21039 18275 21097 18281
rect 21039 18241 21051 18275
rect 21085 18272 21097 18275
rect 21085 18244 21220 18272
rect 21085 18241 21097 18244
rect 21039 18235 21097 18241
rect 18509 18207 18567 18213
rect 18509 18173 18521 18207
rect 18555 18173 18567 18207
rect 18509 18167 18567 18173
rect 18690 18164 18696 18216
rect 18748 18164 18754 18216
rect 20346 18164 20352 18216
rect 20404 18204 20410 18216
rect 20898 18213 20904 18216
rect 20533 18207 20591 18213
rect 20533 18204 20545 18207
rect 20404 18176 20545 18204
rect 20404 18164 20410 18176
rect 20533 18173 20545 18176
rect 20579 18173 20591 18207
rect 20533 18167 20591 18173
rect 20860 18207 20904 18213
rect 20860 18173 20872 18207
rect 20860 18167 20904 18173
rect 20898 18164 20904 18167
rect 20956 18164 20962 18216
rect 21192 18204 21220 18244
rect 21266 18232 21272 18284
rect 21324 18232 21330 18284
rect 24228 18272 24256 18303
rect 26602 18300 26608 18352
rect 26660 18300 26666 18352
rect 22848 18244 24256 18272
rect 25271 18275 25329 18281
rect 22848 18213 22876 18244
rect 25271 18241 25283 18275
rect 25317 18272 25329 18275
rect 25958 18272 25964 18284
rect 25317 18244 25964 18272
rect 25317 18241 25329 18244
rect 25271 18235 25329 18241
rect 25958 18232 25964 18244
rect 26016 18232 26022 18284
rect 28368 18272 28396 18380
rect 26988 18244 28396 18272
rect 22833 18207 22891 18213
rect 21192 18176 21956 18204
rect 12618 18096 12624 18148
rect 12676 18136 12682 18148
rect 12989 18139 13047 18145
rect 12989 18136 13001 18139
rect 12676 18108 13001 18136
rect 12676 18096 12682 18108
rect 12989 18105 13001 18108
rect 13035 18105 13047 18139
rect 12989 18099 13047 18105
rect 13630 18096 13636 18148
rect 13688 18136 13694 18148
rect 13725 18139 13783 18145
rect 13725 18136 13737 18139
rect 13688 18108 13737 18136
rect 13688 18096 13694 18108
rect 13725 18105 13737 18108
rect 13771 18105 13783 18139
rect 21928 18136 21956 18176
rect 22833 18173 22845 18207
rect 22879 18173 22891 18207
rect 22833 18167 22891 18173
rect 23569 18207 23627 18213
rect 23569 18173 23581 18207
rect 23615 18204 23627 18207
rect 23658 18204 23664 18216
rect 23615 18176 23664 18204
rect 23615 18173 23627 18176
rect 23569 18167 23627 18173
rect 23658 18164 23664 18176
rect 23716 18164 23722 18216
rect 23842 18164 23848 18216
rect 23900 18204 23906 18216
rect 23937 18207 23995 18213
rect 23937 18204 23949 18207
rect 23900 18176 23949 18204
rect 23900 18164 23906 18176
rect 23937 18173 23949 18176
rect 23983 18204 23995 18207
rect 24118 18204 24124 18216
rect 23983 18176 24124 18204
rect 23983 18173 23995 18176
rect 23937 18167 23995 18173
rect 24118 18164 24124 18176
rect 24176 18164 24182 18216
rect 24302 18164 24308 18216
rect 24360 18204 24366 18216
rect 24397 18207 24455 18213
rect 24397 18204 24409 18207
rect 24360 18176 24409 18204
rect 24360 18164 24366 18176
rect 24397 18173 24409 18176
rect 24443 18173 24455 18207
rect 24397 18167 24455 18173
rect 24670 18164 24676 18216
rect 24728 18204 24734 18216
rect 24765 18207 24823 18213
rect 24765 18204 24777 18207
rect 24728 18176 24777 18204
rect 24728 18164 24734 18176
rect 24765 18173 24777 18176
rect 24811 18173 24823 18207
rect 24765 18167 24823 18173
rect 25501 18207 25559 18213
rect 25501 18173 25513 18207
rect 25547 18204 25559 18207
rect 26988 18204 27016 18244
rect 30374 18232 30380 18284
rect 30432 18232 30438 18284
rect 25547 18176 27016 18204
rect 27065 18207 27123 18213
rect 25547 18173 25559 18176
rect 25501 18167 25559 18173
rect 27065 18173 27077 18207
rect 27111 18173 27123 18207
rect 28997 18207 29055 18213
rect 28997 18204 29009 18207
rect 27065 18167 27123 18173
rect 28644 18176 29009 18204
rect 13725 18099 13783 18105
rect 17512 18108 18460 18136
rect 21928 18108 24532 18136
rect 11201 18040 12112 18068
rect 11201 18037 11213 18040
rect 11155 18031 11213 18037
rect 13906 18028 13912 18080
rect 13964 18068 13970 18080
rect 14642 18068 14648 18080
rect 13964 18040 14648 18068
rect 13964 18028 13970 18040
rect 14642 18028 14648 18040
rect 14700 18028 14706 18080
rect 14826 18028 14832 18080
rect 14884 18077 14890 18080
rect 14884 18031 14893 18077
rect 14884 18028 14890 18031
rect 16206 18028 16212 18080
rect 16264 18028 16270 18080
rect 16666 18028 16672 18080
rect 16724 18068 16730 18080
rect 17512 18068 17540 18108
rect 16724 18040 17540 18068
rect 16724 18028 16730 18040
rect 18322 18028 18328 18080
rect 18380 18028 18386 18080
rect 18432 18068 18460 18108
rect 24504 18080 24532 18108
rect 22186 18068 22192 18080
rect 18432 18040 22192 18068
rect 22186 18028 22192 18040
rect 22244 18028 22250 18080
rect 22370 18028 22376 18080
rect 22428 18028 22434 18080
rect 24486 18028 24492 18080
rect 24544 18028 24550 18080
rect 25130 18028 25136 18080
rect 25188 18068 25194 18080
rect 25231 18071 25289 18077
rect 25231 18068 25243 18071
rect 25188 18040 25243 18068
rect 25188 18028 25194 18040
rect 25231 18037 25243 18040
rect 25277 18068 25289 18071
rect 26142 18068 26148 18080
rect 25277 18040 26148 18068
rect 25277 18037 25289 18040
rect 25231 18031 25289 18037
rect 26142 18028 26148 18040
rect 26200 18028 26206 18080
rect 27086 18068 27114 18167
rect 27341 18139 27399 18145
rect 27341 18105 27353 18139
rect 27387 18136 27399 18139
rect 27430 18136 27436 18148
rect 27387 18108 27436 18136
rect 27387 18105 27399 18108
rect 27341 18099 27399 18105
rect 27430 18096 27436 18108
rect 27488 18096 27494 18148
rect 27798 18096 27804 18148
rect 27856 18096 27862 18148
rect 28644 18068 28672 18176
rect 28997 18173 29009 18176
rect 29043 18204 29055 18207
rect 29178 18204 29184 18216
rect 29043 18176 29184 18204
rect 29043 18173 29055 18176
rect 28997 18167 29055 18173
rect 29178 18164 29184 18176
rect 29236 18164 29242 18216
rect 29273 18207 29331 18213
rect 29273 18173 29285 18207
rect 29319 18204 29331 18207
rect 29362 18204 29368 18216
rect 29319 18176 29368 18204
rect 29319 18173 29331 18176
rect 29273 18167 29331 18173
rect 29362 18164 29368 18176
rect 29420 18164 29426 18216
rect 30392 18204 30420 18232
rect 30561 18207 30619 18213
rect 30561 18204 30573 18207
rect 30392 18176 30573 18204
rect 30561 18173 30573 18176
rect 30607 18173 30619 18207
rect 30561 18167 30619 18173
rect 28902 18096 28908 18148
rect 28960 18136 28966 18148
rect 28960 18108 30420 18136
rect 28960 18096 28966 18108
rect 27086 18040 28672 18068
rect 28810 18028 28816 18080
rect 28868 18028 28874 18080
rect 29086 18028 29092 18080
rect 29144 18068 29150 18080
rect 29730 18068 29736 18080
rect 29144 18040 29736 18068
rect 29144 18028 29150 18040
rect 29730 18028 29736 18040
rect 29788 18068 29794 18080
rect 29917 18071 29975 18077
rect 29917 18068 29929 18071
rect 29788 18040 29929 18068
rect 29788 18028 29794 18040
rect 29917 18037 29929 18040
rect 29963 18037 29975 18071
rect 29917 18031 29975 18037
rect 30101 18071 30159 18077
rect 30101 18037 30113 18071
rect 30147 18068 30159 18071
rect 30190 18068 30196 18080
rect 30147 18040 30196 18068
rect 30147 18037 30159 18040
rect 30101 18031 30159 18037
rect 30190 18028 30196 18040
rect 30248 18028 30254 18080
rect 30392 18077 30420 18108
rect 30377 18071 30435 18077
rect 30377 18037 30389 18071
rect 30423 18037 30435 18071
rect 30377 18031 30435 18037
rect 552 17978 31072 18000
rect 552 17926 7988 17978
rect 8040 17926 8052 17978
rect 8104 17926 8116 17978
rect 8168 17926 8180 17978
rect 8232 17926 8244 17978
rect 8296 17926 15578 17978
rect 15630 17926 15642 17978
rect 15694 17926 15706 17978
rect 15758 17926 15770 17978
rect 15822 17926 15834 17978
rect 15886 17926 23168 17978
rect 23220 17926 23232 17978
rect 23284 17926 23296 17978
rect 23348 17926 23360 17978
rect 23412 17926 23424 17978
rect 23476 17926 30758 17978
rect 30810 17926 30822 17978
rect 30874 17926 30886 17978
rect 30938 17926 30950 17978
rect 31002 17926 31014 17978
rect 31066 17926 31072 17978
rect 552 17904 31072 17926
rect 4522 17864 4528 17876
rect 3344 17836 4528 17864
rect 1118 17756 1124 17808
rect 1176 17756 1182 17808
rect 842 17688 848 17740
rect 900 17728 906 17740
rect 1136 17728 1164 17756
rect 1213 17731 1271 17737
rect 1213 17728 1225 17731
rect 900 17700 1225 17728
rect 900 17688 906 17700
rect 1213 17697 1225 17700
rect 1259 17697 1271 17731
rect 3142 17728 3148 17740
rect 1213 17691 1271 17697
rect 1964 17700 3148 17728
rect 1801 17681 1859 17687
rect 1670 17669 1676 17672
rect 1305 17663 1363 17669
rect 1305 17660 1317 17663
rect 1228 17632 1317 17660
rect 1228 17536 1256 17632
rect 1305 17629 1317 17632
rect 1351 17629 1363 17663
rect 1305 17623 1363 17629
rect 1632 17663 1676 17669
rect 1632 17629 1644 17663
rect 1632 17623 1676 17629
rect 1670 17620 1676 17623
rect 1728 17620 1734 17672
rect 1801 17647 1813 17681
rect 1847 17660 1859 17681
rect 1964 17660 1992 17700
rect 3142 17688 3148 17700
rect 3200 17688 3206 17740
rect 1847 17647 1992 17660
rect 1801 17641 1992 17647
rect 1826 17632 1992 17641
rect 2041 17663 2099 17669
rect 2041 17629 2053 17663
rect 2087 17660 2099 17663
rect 2406 17660 2412 17672
rect 2087 17632 2412 17660
rect 2087 17629 2099 17632
rect 2041 17623 2099 17629
rect 2406 17620 2412 17632
rect 2464 17620 2470 17672
rect 1029 17527 1087 17533
rect 1029 17524 1041 17527
rect 492 17496 1041 17524
rect 492 17320 520 17496
rect 1029 17493 1041 17496
rect 1075 17493 1087 17527
rect 1029 17487 1087 17493
rect 1210 17484 1216 17536
rect 1268 17484 1274 17536
rect 1946 17484 1952 17536
rect 2004 17524 2010 17536
rect 3344 17524 3372 17836
rect 4522 17824 4528 17836
rect 4580 17824 4586 17876
rect 4614 17824 4620 17876
rect 4672 17864 4678 17876
rect 5537 17867 5595 17873
rect 4672 17836 5488 17864
rect 4672 17824 4678 17836
rect 3421 17799 3479 17805
rect 3421 17765 3433 17799
rect 3467 17796 3479 17799
rect 3510 17796 3516 17808
rect 3467 17768 3516 17796
rect 3467 17765 3479 17768
rect 3421 17759 3479 17765
rect 3510 17756 3516 17768
rect 3568 17756 3574 17808
rect 5460 17796 5488 17836
rect 5537 17833 5549 17867
rect 5583 17864 5595 17867
rect 6362 17864 6368 17876
rect 5583 17836 6368 17864
rect 5583 17833 5595 17836
rect 5537 17827 5595 17833
rect 6362 17824 6368 17836
rect 6420 17824 6426 17876
rect 6730 17824 6736 17876
rect 6788 17864 6794 17876
rect 6923 17867 6981 17873
rect 6923 17864 6935 17867
rect 6788 17836 6935 17864
rect 6788 17824 6794 17836
rect 6923 17833 6935 17836
rect 6969 17833 6981 17867
rect 6923 17827 6981 17833
rect 7834 17824 7840 17876
rect 7892 17824 7898 17876
rect 8478 17824 8484 17876
rect 8536 17824 8542 17876
rect 10134 17864 10140 17876
rect 8772 17836 10140 17864
rect 7852 17796 7880 17824
rect 8772 17796 8800 17836
rect 10134 17824 10140 17836
rect 10192 17824 10198 17876
rect 10689 17867 10747 17873
rect 10689 17833 10701 17867
rect 10735 17864 10747 17867
rect 11054 17864 11060 17876
rect 10735 17836 11060 17864
rect 10735 17833 10747 17836
rect 10689 17827 10747 17833
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 11983 17867 12041 17873
rect 11983 17833 11995 17867
rect 12029 17864 12041 17867
rect 12158 17864 12164 17876
rect 12029 17836 12164 17864
rect 12029 17833 12041 17836
rect 11983 17827 12041 17833
rect 12158 17824 12164 17836
rect 12216 17824 12222 17876
rect 16206 17864 16212 17876
rect 13924 17836 16212 17864
rect 11422 17796 11428 17808
rect 5460 17768 6040 17796
rect 7852 17768 8800 17796
rect 11072 17768 11428 17796
rect 4178 17700 5580 17728
rect 3878 17669 3884 17672
rect 3513 17663 3571 17669
rect 3513 17629 3525 17663
rect 3559 17629 3571 17663
rect 3513 17623 3571 17629
rect 3840 17663 3884 17669
rect 3840 17629 3852 17663
rect 3840 17623 3884 17629
rect 2004 17496 3372 17524
rect 3528 17524 3556 17623
rect 3878 17620 3884 17623
rect 3936 17620 3942 17672
rect 4019 17663 4077 17669
rect 4019 17629 4031 17663
rect 4065 17660 4077 17663
rect 4178 17660 4206 17700
rect 5552 17672 5580 17700
rect 5810 17688 5816 17740
rect 5868 17728 5874 17740
rect 5905 17731 5963 17737
rect 5905 17728 5917 17731
rect 5868 17700 5917 17728
rect 5868 17688 5874 17700
rect 5905 17697 5917 17700
rect 5951 17697 5963 17731
rect 6012 17728 6040 17768
rect 7193 17731 7251 17737
rect 7193 17728 7205 17731
rect 6012 17700 7205 17728
rect 5905 17691 5963 17697
rect 7193 17697 7205 17700
rect 7239 17697 7251 17731
rect 7193 17691 7251 17697
rect 4065 17632 4206 17660
rect 4249 17663 4307 17669
rect 4065 17629 4077 17632
rect 4019 17623 4077 17629
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 5258 17660 5264 17672
rect 4295 17632 5264 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 5258 17620 5264 17632
rect 5316 17620 5322 17672
rect 5534 17620 5540 17672
rect 5592 17620 5598 17672
rect 5920 17660 5948 17691
rect 8570 17688 8576 17740
rect 8628 17728 8634 17740
rect 8628 17700 9171 17728
rect 8628 17688 8634 17700
rect 6086 17660 6092 17672
rect 5920 17632 6092 17660
rect 6086 17620 6092 17632
rect 6144 17660 6150 17672
rect 6457 17663 6515 17669
rect 6457 17660 6469 17663
rect 6144 17632 6469 17660
rect 6144 17620 6150 17632
rect 6457 17629 6469 17632
rect 6503 17629 6515 17663
rect 6457 17623 6515 17629
rect 6920 17665 6978 17671
rect 6920 17631 6932 17665
rect 6966 17660 6978 17665
rect 7006 17660 7012 17672
rect 6966 17632 7012 17660
rect 6966 17631 6978 17632
rect 6920 17625 6978 17631
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 8662 17620 8668 17672
rect 8720 17620 8726 17672
rect 9030 17669 9036 17672
rect 8992 17663 9036 17669
rect 8992 17629 9004 17663
rect 8992 17623 9036 17629
rect 9030 17620 9036 17623
rect 9088 17620 9094 17672
rect 9143 17671 9171 17700
rect 9214 17688 9220 17740
rect 9272 17728 9278 17740
rect 9401 17731 9459 17737
rect 9401 17728 9413 17731
rect 9272 17700 9413 17728
rect 9272 17688 9278 17700
rect 9401 17697 9413 17700
rect 9447 17697 9459 17731
rect 9401 17691 9459 17697
rect 9858 17688 9864 17740
rect 9916 17688 9922 17740
rect 11072 17737 11100 17768
rect 11422 17756 11428 17768
rect 11480 17756 11486 17808
rect 11057 17731 11115 17737
rect 11057 17697 11069 17731
rect 11103 17697 11115 17731
rect 12253 17731 12311 17737
rect 12253 17728 12265 17731
rect 11057 17691 11115 17697
rect 11164 17700 12265 17728
rect 9128 17665 9186 17671
rect 9128 17631 9140 17665
rect 9174 17631 9186 17665
rect 9876 17660 9904 17688
rect 11164 17660 11192 17700
rect 12253 17697 12265 17700
rect 12299 17697 12311 17731
rect 12253 17691 12311 17697
rect 9876 17632 11192 17660
rect 9128 17625 9186 17631
rect 11238 17620 11244 17672
rect 11296 17660 11302 17672
rect 11514 17660 11520 17672
rect 11296 17632 11520 17660
rect 11296 17620 11302 17632
rect 11514 17620 11520 17632
rect 11572 17620 11578 17672
rect 12023 17663 12081 17669
rect 12023 17629 12035 17663
rect 12069 17660 12081 17663
rect 13924 17660 13952 17836
rect 16206 17824 16212 17836
rect 16264 17824 16270 17876
rect 16482 17824 16488 17876
rect 16540 17864 16546 17876
rect 17037 17867 17095 17873
rect 17037 17864 17049 17867
rect 16540 17836 17049 17864
rect 16540 17824 16546 17836
rect 17037 17833 17049 17836
rect 17083 17833 17095 17867
rect 23290 17864 23296 17876
rect 17037 17827 17095 17833
rect 17236 17836 18920 17864
rect 16114 17756 16120 17808
rect 16172 17756 16178 17808
rect 14001 17731 14059 17737
rect 14001 17697 14013 17731
rect 14047 17728 14059 17731
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 14047 17700 14289 17728
rect 14047 17697 14059 17700
rect 14001 17691 14059 17697
rect 14277 17697 14289 17700
rect 14323 17728 14335 17731
rect 16132 17728 16160 17756
rect 16209 17731 16267 17737
rect 16209 17728 16221 17731
rect 14323 17700 15516 17728
rect 16132 17700 16221 17728
rect 14323 17697 14335 17700
rect 14277 17691 14335 17697
rect 15488 17672 15516 17700
rect 16209 17697 16221 17700
rect 16255 17697 16267 17731
rect 16209 17691 16267 17697
rect 16666 17688 16672 17740
rect 16724 17688 16730 17740
rect 17236 17728 17264 17836
rect 18892 17796 18920 17836
rect 19076 17836 23296 17864
rect 19076 17796 19104 17836
rect 23290 17824 23296 17836
rect 23348 17824 23354 17876
rect 25961 17867 26019 17873
rect 25961 17864 25973 17867
rect 23400 17836 25973 17864
rect 18892 17768 19104 17796
rect 20530 17756 20536 17808
rect 20588 17796 20594 17808
rect 21082 17796 21088 17808
rect 20588 17768 21088 17796
rect 20588 17756 20594 17768
rect 21082 17756 21088 17768
rect 21140 17756 21146 17808
rect 16868 17700 17264 17728
rect 17865 17731 17923 17737
rect 12069 17632 13952 17660
rect 14553 17663 14611 17669
rect 12069 17629 12081 17632
rect 12023 17623 12081 17629
rect 14553 17629 14565 17663
rect 14599 17660 14611 17663
rect 15010 17660 15016 17672
rect 14599 17632 15016 17660
rect 14599 17629 14611 17632
rect 14553 17623 14611 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 15470 17620 15476 17672
rect 15528 17620 15534 17672
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17660 15991 17663
rect 16868 17660 16896 17700
rect 17865 17697 17877 17731
rect 17911 17728 17923 17731
rect 18322 17728 18328 17740
rect 17911 17700 18328 17728
rect 17911 17697 17923 17700
rect 17865 17691 17923 17697
rect 18322 17688 18328 17700
rect 18380 17688 18386 17740
rect 19705 17731 19763 17737
rect 19705 17697 19717 17731
rect 19751 17728 19763 17731
rect 19794 17728 19800 17740
rect 19751 17700 19800 17728
rect 19751 17697 19763 17700
rect 19705 17691 19763 17697
rect 19794 17688 19800 17700
rect 19852 17688 19858 17740
rect 20898 17688 20904 17740
rect 20956 17728 20962 17740
rect 21596 17731 21654 17737
rect 21596 17728 21608 17731
rect 20956 17700 21608 17728
rect 20956 17688 20962 17700
rect 21100 17672 21128 17700
rect 21596 17697 21608 17700
rect 21642 17697 21654 17731
rect 23400 17728 23428 17836
rect 25961 17833 25973 17836
rect 26007 17833 26019 17867
rect 25961 17827 26019 17833
rect 26142 17824 26148 17876
rect 26200 17864 26206 17876
rect 26887 17867 26945 17873
rect 26887 17864 26899 17867
rect 26200 17836 26899 17864
rect 26200 17824 26206 17836
rect 26887 17833 26899 17836
rect 26933 17833 26945 17867
rect 26887 17827 26945 17833
rect 27062 17824 27068 17876
rect 27120 17864 27126 17876
rect 28261 17867 28319 17873
rect 28261 17864 28273 17867
rect 27120 17836 28273 17864
rect 27120 17824 27126 17836
rect 28261 17833 28273 17836
rect 28307 17833 28319 17867
rect 28902 17864 28908 17876
rect 28261 17827 28319 17833
rect 28558 17836 28908 17864
rect 21596 17691 21654 17697
rect 21828 17700 23428 17728
rect 21828 17694 21856 17700
rect 21780 17687 21856 17694
rect 23474 17688 23480 17740
rect 23532 17688 23538 17740
rect 24857 17731 24915 17737
rect 24857 17697 24869 17731
rect 24903 17697 24915 17731
rect 28558 17728 28586 17836
rect 28902 17824 28908 17836
rect 28960 17824 28966 17876
rect 28644 17768 29224 17796
rect 28644 17737 28672 17768
rect 29196 17740 29224 17768
rect 29730 17756 29736 17808
rect 29788 17796 29794 17808
rect 30193 17799 30251 17805
rect 30193 17796 30205 17799
rect 29788 17768 30205 17796
rect 29788 17756 29794 17768
rect 30193 17765 30205 17768
rect 30239 17765 30251 17799
rect 30193 17759 30251 17765
rect 24857 17691 24915 17697
rect 25700 17700 28586 17728
rect 28629 17731 28687 17737
rect 21765 17681 21856 17687
rect 15979 17632 16896 17660
rect 15979 17629 15991 17632
rect 15933 17623 15991 17629
rect 16942 17620 16948 17672
rect 17000 17620 17006 17672
rect 17494 17669 17500 17672
rect 17129 17663 17187 17669
rect 17129 17629 17141 17663
rect 17175 17629 17187 17663
rect 17129 17623 17187 17629
rect 17456 17663 17500 17669
rect 17456 17629 17468 17663
rect 17456 17623 17500 17629
rect 5828 17564 6500 17592
rect 3786 17524 3792 17536
rect 3528 17496 3792 17524
rect 2004 17484 2010 17496
rect 3786 17484 3792 17496
rect 3844 17484 3850 17536
rect 4062 17484 4068 17536
rect 4120 17524 4126 17536
rect 5828 17524 5856 17564
rect 4120 17496 5856 17524
rect 4120 17484 4126 17496
rect 5902 17484 5908 17536
rect 5960 17524 5966 17536
rect 5997 17527 6055 17533
rect 5997 17524 6009 17527
rect 5960 17496 6009 17524
rect 5960 17484 5966 17496
rect 5997 17493 6009 17496
rect 6043 17493 6055 17527
rect 6472 17524 6500 17564
rect 10704 17564 11284 17592
rect 10704 17536 10732 17564
rect 9490 17524 9496 17536
rect 6472 17496 9496 17524
rect 5997 17487 6055 17493
rect 9490 17484 9496 17496
rect 9548 17484 9554 17536
rect 10686 17484 10692 17536
rect 10744 17484 10750 17536
rect 10962 17484 10968 17536
rect 11020 17524 11026 17536
rect 11149 17527 11207 17533
rect 11149 17524 11161 17527
rect 11020 17496 11161 17524
rect 11020 17484 11026 17496
rect 11149 17493 11161 17496
rect 11195 17493 11207 17527
rect 11256 17524 11284 17564
rect 16390 17552 16396 17604
rect 16448 17592 16454 17604
rect 17144 17592 17172 17623
rect 17494 17620 17500 17623
rect 17552 17620 17558 17672
rect 17635 17663 17693 17669
rect 17635 17629 17647 17663
rect 17681 17660 17693 17663
rect 19429 17663 19487 17669
rect 17681 17632 19380 17660
rect 17681 17629 17693 17632
rect 17635 17623 17693 17629
rect 16448 17564 17172 17592
rect 16448 17552 16454 17564
rect 13357 17527 13415 17533
rect 13357 17524 13369 17527
rect 11256 17496 13369 17524
rect 11149 17487 11207 17493
rect 13357 17493 13369 17496
rect 13403 17493 13415 17527
rect 13357 17487 13415 17493
rect 15930 17484 15936 17536
rect 15988 17524 15994 17536
rect 17678 17524 17684 17536
rect 15988 17496 17684 17524
rect 15988 17484 15994 17496
rect 17678 17484 17684 17496
rect 17736 17484 17742 17536
rect 17954 17484 17960 17536
rect 18012 17524 18018 17536
rect 18969 17527 19027 17533
rect 18969 17524 18981 17527
rect 18012 17496 18981 17524
rect 18012 17484 18018 17496
rect 18969 17493 18981 17496
rect 19015 17493 19027 17527
rect 19352 17524 19380 17632
rect 19429 17629 19441 17663
rect 19475 17660 19487 17663
rect 20438 17660 20444 17672
rect 19475 17632 20444 17660
rect 19475 17629 19487 17632
rect 19429 17623 19487 17629
rect 20438 17620 20444 17632
rect 20496 17620 20502 17672
rect 21082 17620 21088 17672
rect 21140 17620 21146 17672
rect 21266 17620 21272 17672
rect 21324 17620 21330 17672
rect 21765 17647 21777 17681
rect 21811 17666 21856 17681
rect 21811 17647 21823 17666
rect 21765 17641 21823 17647
rect 22005 17663 22063 17669
rect 22005 17629 22017 17663
rect 22051 17660 22063 17663
rect 22922 17660 22928 17672
rect 22051 17632 22928 17660
rect 22051 17629 22063 17632
rect 22005 17623 22063 17629
rect 22922 17620 22928 17632
rect 22980 17620 22986 17672
rect 24486 17669 24492 17672
rect 24121 17663 24179 17669
rect 24121 17629 24133 17663
rect 24167 17629 24179 17663
rect 24121 17623 24179 17629
rect 24448 17663 24492 17669
rect 24448 17629 24460 17663
rect 24448 17623 24492 17629
rect 20732 17564 20944 17592
rect 20732 17524 20760 17564
rect 19352 17496 20760 17524
rect 18969 17487 19027 17493
rect 20806 17484 20812 17536
rect 20864 17484 20870 17536
rect 20916 17524 20944 17564
rect 23566 17552 23572 17604
rect 23624 17552 23630 17604
rect 23014 17524 23020 17536
rect 20916 17496 23020 17524
rect 23014 17484 23020 17496
rect 23072 17484 23078 17536
rect 23106 17484 23112 17536
rect 23164 17484 23170 17536
rect 23750 17484 23756 17536
rect 23808 17524 23814 17536
rect 24136 17524 24164 17623
rect 24486 17620 24492 17623
rect 24544 17620 24550 17672
rect 24627 17663 24685 17669
rect 24627 17629 24639 17663
rect 24673 17660 24685 17663
rect 24762 17660 24768 17672
rect 24673 17632 24768 17660
rect 24673 17629 24685 17632
rect 24627 17623 24685 17629
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 24872 17660 24900 17691
rect 25700 17660 25728 17700
rect 28629 17697 28641 17731
rect 28675 17697 28687 17731
rect 28629 17691 28687 17697
rect 28902 17688 28908 17740
rect 28960 17688 28966 17740
rect 29178 17688 29184 17740
rect 29236 17688 29242 17740
rect 24872 17632 25728 17660
rect 25774 17620 25780 17672
rect 25832 17660 25838 17672
rect 26421 17663 26479 17669
rect 26421 17660 26433 17663
rect 25832 17632 26433 17660
rect 25832 17620 25838 17632
rect 26421 17629 26433 17632
rect 26467 17629 26479 17663
rect 26421 17623 26479 17629
rect 26878 17620 26884 17672
rect 26936 17660 26942 17672
rect 27157 17663 27215 17669
rect 26936 17632 26981 17660
rect 26936 17620 26942 17632
rect 27157 17629 27169 17663
rect 27203 17660 27215 17663
rect 27203 17632 28586 17660
rect 27203 17629 27215 17632
rect 27157 17623 27215 17629
rect 24762 17524 24768 17536
rect 23808 17496 24768 17524
rect 23808 17484 23814 17496
rect 24762 17484 24768 17496
rect 24820 17524 24826 17536
rect 25774 17524 25780 17536
rect 24820 17496 25780 17524
rect 24820 17484 24826 17496
rect 25774 17484 25780 17496
rect 25832 17484 25838 17536
rect 25866 17484 25872 17536
rect 25924 17524 25930 17536
rect 27798 17524 27804 17536
rect 25924 17496 27804 17524
rect 25924 17484 25930 17496
rect 27798 17484 27804 17496
rect 27856 17484 27862 17536
rect 28558 17524 28586 17632
rect 30466 17620 30472 17672
rect 30524 17620 30530 17672
rect 30098 17552 30104 17604
rect 30156 17552 30162 17604
rect 30116 17524 30144 17552
rect 28558 17496 30144 17524
rect 552 17434 30912 17456
rect 552 17382 4193 17434
rect 4245 17382 4257 17434
rect 4309 17382 4321 17434
rect 4373 17382 4385 17434
rect 4437 17382 4449 17434
rect 4501 17382 11783 17434
rect 11835 17382 11847 17434
rect 11899 17382 11911 17434
rect 11963 17382 11975 17434
rect 12027 17382 12039 17434
rect 12091 17382 19373 17434
rect 19425 17382 19437 17434
rect 19489 17382 19501 17434
rect 19553 17382 19565 17434
rect 19617 17382 19629 17434
rect 19681 17382 26963 17434
rect 27015 17382 27027 17434
rect 27079 17382 27091 17434
rect 27143 17382 27155 17434
rect 27207 17382 27219 17434
rect 27271 17382 30912 17434
rect 552 17360 30912 17382
rect 492 17292 2774 17320
rect 2746 17252 2774 17292
rect 2866 17280 2872 17332
rect 2924 17320 2930 17332
rect 2961 17323 3019 17329
rect 2961 17320 2973 17323
rect 2924 17292 2973 17320
rect 2924 17280 2930 17292
rect 2961 17289 2973 17292
rect 3007 17289 3019 17323
rect 4522 17320 4528 17332
rect 2961 17283 3019 17289
rect 3896 17292 4528 17320
rect 3896 17252 3924 17292
rect 4522 17280 4528 17292
rect 4580 17280 4586 17332
rect 8389 17323 8447 17329
rect 8389 17289 8401 17323
rect 8435 17320 8447 17323
rect 9766 17320 9772 17332
rect 8435 17292 9772 17320
rect 8435 17289 8447 17292
rect 8389 17283 8447 17289
rect 9766 17280 9772 17292
rect 9824 17280 9830 17332
rect 10502 17280 10508 17332
rect 10560 17280 10566 17332
rect 11054 17280 11060 17332
rect 11112 17280 11118 17332
rect 16025 17323 16083 17329
rect 16025 17320 16037 17323
rect 11256 17292 16037 17320
rect 2746 17224 3924 17252
rect 1443 17187 1501 17193
rect 1443 17153 1455 17187
rect 1489 17184 1501 17187
rect 2774 17184 2780 17196
rect 1489 17156 2780 17184
rect 1489 17153 1501 17156
rect 1443 17147 1501 17153
rect 2774 17144 2780 17156
rect 2832 17144 2838 17196
rect 3510 17144 3516 17196
rect 3568 17184 3574 17196
rect 4062 17184 4068 17196
rect 3568 17156 4068 17184
rect 3568 17144 3574 17156
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 4430 17193 4436 17196
rect 4387 17187 4436 17193
rect 4387 17153 4399 17187
rect 4433 17153 4436 17187
rect 4387 17147 4436 17153
rect 4430 17144 4436 17147
rect 4488 17144 4494 17196
rect 4571 17187 4629 17193
rect 4571 17153 4583 17187
rect 4617 17184 4629 17187
rect 5350 17184 5356 17196
rect 4617 17156 5356 17184
rect 4617 17153 4629 17156
rect 4571 17147 4629 17153
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 5997 17187 6055 17193
rect 5997 17153 6009 17187
rect 6043 17184 6055 17187
rect 6552 17187 6610 17193
rect 6552 17184 6564 17187
rect 6043 17156 6564 17184
rect 6043 17153 6055 17156
rect 5997 17147 6055 17153
rect 6552 17153 6564 17156
rect 6598 17153 6610 17187
rect 6552 17147 6610 17153
rect 6638 17144 6644 17196
rect 6696 17184 6702 17196
rect 6825 17187 6883 17193
rect 6825 17184 6837 17187
rect 6696 17156 6837 17184
rect 6696 17144 6702 17156
rect 6825 17153 6837 17156
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17184 8263 17187
rect 9128 17187 9186 17193
rect 8251 17156 9082 17184
rect 8251 17153 8263 17156
rect 8205 17147 8263 17153
rect 937 17119 995 17125
rect 937 17085 949 17119
rect 983 17116 995 17119
rect 1210 17116 1216 17128
rect 983 17088 1216 17116
rect 983 17085 995 17088
rect 937 17079 995 17085
rect 1210 17076 1216 17088
rect 1268 17076 1274 17128
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17116 1731 17119
rect 1762 17116 1768 17128
rect 1719 17088 1768 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 1762 17076 1768 17088
rect 1820 17076 1826 17128
rect 3237 17119 3295 17125
rect 3237 17085 3249 17119
rect 3283 17116 3295 17119
rect 3418 17116 3424 17128
rect 3283 17088 3424 17116
rect 3283 17085 3295 17088
rect 3237 17079 3295 17085
rect 3418 17076 3424 17088
rect 3476 17076 3482 17128
rect 3786 17076 3792 17128
rect 3844 17116 3850 17128
rect 3881 17119 3939 17125
rect 3881 17116 3893 17119
rect 3844 17088 3893 17116
rect 3844 17076 3850 17088
rect 3881 17085 3893 17088
rect 3927 17116 3939 17119
rect 5902 17116 5908 17128
rect 3927 17112 4568 17116
rect 4724 17112 5908 17116
rect 3927 17088 5908 17112
rect 3927 17085 3939 17088
rect 3881 17079 3939 17085
rect 4540 17084 4752 17088
rect 5902 17076 5908 17088
rect 5960 17076 5966 17128
rect 6086 17076 6092 17128
rect 6144 17076 6150 17128
rect 8573 17119 8631 17125
rect 8573 17116 8585 17119
rect 8496 17088 8585 17116
rect 3513 17051 3571 17057
rect 3513 17017 3525 17051
rect 3559 17017 3571 17051
rect 3513 17011 3571 17017
rect 1403 16983 1461 16989
rect 1403 16949 1415 16983
rect 1449 16980 1461 16983
rect 1670 16980 1676 16992
rect 1449 16952 1676 16980
rect 1449 16949 1461 16952
rect 1403 16943 1461 16949
rect 1670 16940 1676 16952
rect 1728 16980 1734 16992
rect 3528 16980 3556 17011
rect 8496 16992 8524 17088
rect 8573 17085 8585 17088
rect 8619 17085 8631 17119
rect 8573 17079 8631 17085
rect 8662 17076 8668 17128
rect 8720 17076 8726 17128
rect 9054 17116 9082 17156
rect 9128 17153 9140 17187
rect 9174 17153 9186 17187
rect 9128 17147 9186 17153
rect 9143 17116 9171 17147
rect 9490 17144 9496 17196
rect 9548 17184 9554 17196
rect 11256 17184 11284 17292
rect 16025 17289 16037 17292
rect 16071 17289 16083 17323
rect 23106 17320 23112 17332
rect 16025 17283 16083 17289
rect 16408 17292 18092 17320
rect 12802 17212 12808 17264
rect 12860 17252 12866 17264
rect 13817 17255 13875 17261
rect 13817 17252 13829 17255
rect 12860 17224 13829 17252
rect 12860 17212 12866 17224
rect 13817 17221 13829 17224
rect 13863 17221 13875 17255
rect 13817 17215 13875 17221
rect 11747 17187 11805 17193
rect 11747 17184 11759 17187
rect 9548 17156 10456 17184
rect 11256 17156 11759 17184
rect 9548 17144 9554 17156
rect 9054 17088 9171 17116
rect 9398 17076 9404 17128
rect 9456 17076 9462 17128
rect 10428 16992 10456 17156
rect 11747 17153 11759 17156
rect 11793 17153 11805 17187
rect 11747 17147 11805 17153
rect 12710 17144 12716 17196
rect 12768 17144 12774 17196
rect 14182 17144 14188 17196
rect 14240 17184 14246 17196
rect 14366 17184 14372 17196
rect 14240 17156 14372 17184
rect 14240 17144 14246 17156
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 14691 17187 14749 17193
rect 14691 17153 14703 17187
rect 14737 17184 14749 17187
rect 16408 17184 16436 17292
rect 18064 17264 18092 17292
rect 19720 17292 23112 17320
rect 18046 17212 18052 17264
rect 18104 17212 18110 17264
rect 14737 17156 16436 17184
rect 14737 17153 14749 17156
rect 14691 17147 14749 17153
rect 16574 17144 16580 17196
rect 16632 17144 16638 17196
rect 16758 17193 16764 17196
rect 16720 17187 16764 17193
rect 16720 17153 16732 17187
rect 16720 17147 16764 17153
rect 16758 17144 16764 17147
rect 16816 17144 16822 17196
rect 16899 17187 16957 17193
rect 16899 17153 16911 17187
rect 16945 17184 16957 17187
rect 19720 17184 19748 17292
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 28810 17320 28816 17332
rect 23400 17292 28816 17320
rect 23400 17264 23428 17292
rect 28810 17280 28816 17292
rect 28868 17320 28874 17332
rect 29730 17320 29736 17332
rect 28868 17292 29736 17320
rect 28868 17280 28874 17292
rect 29730 17280 29736 17292
rect 29788 17280 29794 17332
rect 30377 17323 30435 17329
rect 30377 17289 30389 17323
rect 30423 17320 30435 17323
rect 30558 17320 30564 17332
rect 30423 17292 30564 17320
rect 30423 17289 30435 17292
rect 30377 17283 30435 17289
rect 30558 17280 30564 17292
rect 30616 17280 30622 17332
rect 20349 17255 20407 17261
rect 20349 17221 20361 17255
rect 20395 17252 20407 17255
rect 20530 17252 20536 17264
rect 20395 17224 20536 17252
rect 20395 17221 20407 17224
rect 20349 17215 20407 17221
rect 20530 17212 20536 17224
rect 20588 17212 20594 17264
rect 23293 17255 23351 17261
rect 23293 17252 23305 17255
rect 22066 17224 23305 17252
rect 20714 17184 20720 17196
rect 16945 17156 19748 17184
rect 20456 17156 20720 17184
rect 16945 17153 16957 17156
rect 16899 17147 16957 17153
rect 10870 17076 10876 17128
rect 10928 17076 10934 17128
rect 11238 17076 11244 17128
rect 11296 17076 11302 17128
rect 11330 17076 11336 17128
rect 11388 17116 11394 17128
rect 11977 17119 12035 17125
rect 11977 17116 11989 17119
rect 11388 17088 11989 17116
rect 11388 17076 11394 17088
rect 11977 17085 11989 17088
rect 12023 17085 12035 17119
rect 11977 17079 12035 17085
rect 12728 17048 12756 17144
rect 13630 17076 13636 17128
rect 13688 17076 13694 17128
rect 14512 17119 14570 17125
rect 14512 17085 14524 17119
rect 14558 17116 14570 17119
rect 14826 17116 14832 17128
rect 14558 17088 14832 17116
rect 14558 17085 14570 17088
rect 14512 17079 14570 17085
rect 14826 17076 14832 17088
rect 14884 17076 14890 17128
rect 14918 17076 14924 17128
rect 14976 17076 14982 17128
rect 16390 17076 16396 17128
rect 16448 17076 16454 17128
rect 16592 17116 16620 17144
rect 17129 17119 17187 17125
rect 17129 17116 17141 17119
rect 16592 17088 17141 17116
rect 17129 17085 17141 17088
rect 17175 17085 17187 17119
rect 17129 17079 17187 17085
rect 18785 17119 18843 17125
rect 18785 17085 18797 17119
rect 18831 17085 18843 17119
rect 18785 17079 18843 17085
rect 19061 17119 19119 17125
rect 19061 17085 19073 17119
rect 19107 17116 19119 17119
rect 20456 17116 20484 17156
rect 20714 17144 20720 17156
rect 20772 17144 20778 17196
rect 21039 17187 21097 17193
rect 21039 17153 21051 17187
rect 21085 17184 21097 17187
rect 21174 17184 21180 17196
rect 21085 17156 21180 17184
rect 21085 17153 21097 17156
rect 21039 17147 21097 17153
rect 21174 17144 21180 17156
rect 21232 17144 21238 17196
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17184 21327 17187
rect 22066 17184 22094 17224
rect 23293 17221 23305 17224
rect 23339 17221 23351 17255
rect 23293 17215 23351 17221
rect 23382 17212 23388 17264
rect 23440 17212 23446 17264
rect 23566 17212 23572 17264
rect 23624 17252 23630 17264
rect 23842 17252 23848 17264
rect 23624 17224 23848 17252
rect 23624 17212 23630 17224
rect 23842 17212 23848 17224
rect 23900 17212 23906 17264
rect 28442 17212 28448 17264
rect 28500 17252 28506 17264
rect 28626 17252 28632 17264
rect 28500 17224 28632 17252
rect 28500 17212 28506 17224
rect 28626 17212 28632 17224
rect 28684 17212 28690 17264
rect 28902 17212 28908 17264
rect 28960 17252 28966 17264
rect 29362 17252 29368 17264
rect 28960 17224 29368 17252
rect 28960 17212 28994 17224
rect 29362 17212 29368 17224
rect 29420 17252 29426 17264
rect 29420 17224 29868 17252
rect 29420 17212 29426 17224
rect 21315 17156 22094 17184
rect 21315 17153 21327 17156
rect 21269 17147 21327 17153
rect 22738 17144 22744 17196
rect 22796 17184 22802 17196
rect 25130 17193 25136 17196
rect 25092 17187 25136 17193
rect 22796 17156 24900 17184
rect 22796 17144 22802 17156
rect 19107 17088 20484 17116
rect 20533 17119 20591 17125
rect 19107 17085 19119 17088
rect 19061 17079 19119 17085
rect 20533 17085 20545 17119
rect 20579 17116 20591 17119
rect 21358 17116 21364 17128
rect 20579 17088 21364 17116
rect 20579 17085 20591 17088
rect 20533 17079 20591 17085
rect 12728 17020 14320 17048
rect 3878 16980 3884 16992
rect 1728 16952 3884 16980
rect 1728 16940 1734 16952
rect 3878 16940 3884 16952
rect 3936 16980 3942 16992
rect 4246 16980 4252 16992
rect 3936 16952 4252 16980
rect 3936 16940 3942 16952
rect 4246 16940 4252 16952
rect 4304 16980 4310 16992
rect 4347 16983 4405 16989
rect 4347 16980 4359 16983
rect 4304 16952 4359 16980
rect 4304 16940 4310 16952
rect 4347 16949 4359 16952
rect 4393 16949 4405 16983
rect 4347 16943 4405 16949
rect 4982 16940 4988 16992
rect 5040 16980 5046 16992
rect 5810 16980 5816 16992
rect 5040 16952 5816 16980
rect 5040 16940 5046 16952
rect 5810 16940 5816 16952
rect 5868 16940 5874 16992
rect 6555 16983 6613 16989
rect 6555 16949 6567 16983
rect 6601 16980 6613 16983
rect 6730 16980 6736 16992
rect 6601 16952 6736 16980
rect 6601 16949 6613 16952
rect 6555 16943 6613 16949
rect 6730 16940 6736 16952
rect 6788 16940 6794 16992
rect 8478 16940 8484 16992
rect 8536 16940 8542 16992
rect 9030 16940 9036 16992
rect 9088 16980 9094 16992
rect 9131 16983 9189 16989
rect 9131 16980 9143 16983
rect 9088 16952 9143 16980
rect 9088 16940 9094 16952
rect 9131 16949 9143 16952
rect 9177 16949 9189 16983
rect 9131 16943 9189 16949
rect 10410 16940 10416 16992
rect 10468 16940 10474 16992
rect 11707 16983 11765 16989
rect 11707 16949 11719 16983
rect 11753 16980 11765 16983
rect 11974 16980 11980 16992
rect 11753 16952 11980 16980
rect 11753 16949 11765 16952
rect 11707 16943 11765 16949
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 12066 16940 12072 16992
rect 12124 16980 12130 16992
rect 13081 16983 13139 16989
rect 13081 16980 13093 16983
rect 12124 16952 13093 16980
rect 12124 16940 12130 16952
rect 13081 16949 13093 16952
rect 13127 16949 13139 16983
rect 14292 16980 14320 17020
rect 14918 16980 14924 16992
rect 14292 16952 14924 16980
rect 13081 16943 13139 16949
rect 14918 16940 14924 16952
rect 14976 16940 14982 16992
rect 16114 16940 16120 16992
rect 16172 16980 16178 16992
rect 18233 16983 18291 16989
rect 18233 16980 18245 16983
rect 16172 16952 18245 16980
rect 16172 16940 16178 16952
rect 18233 16949 18245 16952
rect 18279 16949 18291 16983
rect 18800 16980 18828 17079
rect 20346 17008 20352 17060
rect 20404 17048 20410 17060
rect 20548 17048 20576 17079
rect 21358 17076 21364 17088
rect 21416 17116 21422 17128
rect 22833 17119 22891 17125
rect 22833 17116 22845 17119
rect 21416 17088 22845 17116
rect 21416 17076 21422 17088
rect 22833 17085 22845 17088
rect 22879 17085 22891 17119
rect 22833 17079 22891 17085
rect 23198 17076 23204 17128
rect 23256 17116 23262 17128
rect 23477 17119 23535 17125
rect 23477 17116 23489 17119
rect 23256 17088 23489 17116
rect 23256 17076 23262 17088
rect 23477 17085 23489 17088
rect 23523 17085 23535 17119
rect 23477 17079 23535 17085
rect 24029 17119 24087 17125
rect 24029 17085 24041 17119
rect 24075 17116 24087 17119
rect 24118 17116 24124 17128
rect 24075 17088 24124 17116
rect 24075 17085 24087 17088
rect 24029 17079 24087 17085
rect 20404 17020 20576 17048
rect 20404 17008 20410 17020
rect 22554 17008 22560 17060
rect 22612 17048 22618 17060
rect 24044 17048 24072 17079
rect 24118 17076 24124 17088
rect 24176 17076 24182 17128
rect 24210 17076 24216 17128
rect 24268 17116 24274 17128
rect 24670 17116 24676 17128
rect 24268 17088 24676 17116
rect 24268 17076 24274 17088
rect 24670 17076 24676 17088
rect 24728 17076 24734 17128
rect 24762 17076 24768 17128
rect 24820 17076 24826 17128
rect 24872 17116 24900 17156
rect 25092 17153 25104 17187
rect 25092 17147 25136 17153
rect 25130 17144 25136 17147
rect 25188 17144 25194 17196
rect 25228 17185 25286 17191
rect 25228 17151 25240 17185
rect 25274 17184 25286 17185
rect 25314 17184 25320 17196
rect 25274 17156 25320 17184
rect 25274 17151 25286 17156
rect 25228 17145 25286 17151
rect 25314 17144 25320 17156
rect 25372 17144 25378 17196
rect 25501 17187 25559 17193
rect 25501 17153 25513 17187
rect 25547 17184 25559 17187
rect 26418 17184 26424 17196
rect 25547 17156 26424 17184
rect 25547 17153 25559 17156
rect 25501 17147 25559 17153
rect 26418 17144 26424 17156
rect 26476 17144 26482 17196
rect 26528 17156 27292 17184
rect 26528 17116 26556 17156
rect 24872 17088 26556 17116
rect 26786 17076 26792 17128
rect 26844 17116 26850 17128
rect 27264 17125 27292 17156
rect 27430 17144 27436 17196
rect 27488 17184 27494 17196
rect 28966 17184 28994 17212
rect 27488 17156 28994 17184
rect 27488 17144 27494 17156
rect 29178 17144 29184 17196
rect 29236 17184 29242 17196
rect 29840 17193 29868 17224
rect 29825 17187 29883 17193
rect 29236 17156 29684 17184
rect 29236 17144 29242 17156
rect 26973 17119 27031 17125
rect 26973 17116 26985 17119
rect 26844 17088 26985 17116
rect 26844 17076 26850 17088
rect 26973 17085 26985 17088
rect 27019 17085 27031 17119
rect 26973 17079 27031 17085
rect 27249 17119 27307 17125
rect 27249 17085 27261 17119
rect 27295 17085 27307 17119
rect 27249 17079 27307 17085
rect 27706 17076 27712 17128
rect 27764 17116 27770 17128
rect 29086 17116 29092 17128
rect 27764 17088 29092 17116
rect 27764 17076 27770 17088
rect 29086 17076 29092 17088
rect 29144 17076 29150 17128
rect 29656 17125 29684 17156
rect 29825 17153 29837 17187
rect 29871 17153 29883 17187
rect 29825 17147 29883 17153
rect 29641 17119 29699 17125
rect 29641 17085 29653 17119
rect 29687 17116 29699 17119
rect 30466 17116 30472 17128
rect 29687 17088 30472 17116
rect 29687 17085 29699 17088
rect 29641 17079 29699 17085
rect 30466 17076 30472 17088
rect 30524 17076 30530 17128
rect 22612 17020 24072 17048
rect 22612 17008 22618 17020
rect 24486 17008 24492 17060
rect 24544 17008 24550 17060
rect 30101 17051 30159 17057
rect 30101 17017 30113 17051
rect 30147 17048 30159 17051
rect 30282 17048 30288 17060
rect 30147 17020 30288 17048
rect 30147 17017 30159 17020
rect 30101 17011 30159 17017
rect 30282 17008 30288 17020
rect 30340 17048 30346 17060
rect 31110 17048 31116 17060
rect 30340 17020 31116 17048
rect 30340 17008 30346 17020
rect 31110 17008 31116 17020
rect 31168 17008 31174 17060
rect 19426 16980 19432 16992
rect 18800 16952 19432 16980
rect 18233 16943 18291 16949
rect 19426 16940 19432 16952
rect 19484 16940 19490 16992
rect 20999 16983 21057 16989
rect 20999 16949 21011 16983
rect 21045 16980 21057 16983
rect 21174 16980 21180 16992
rect 21045 16952 21180 16980
rect 21045 16949 21057 16952
rect 20999 16943 21057 16949
rect 21174 16940 21180 16952
rect 21232 16940 21238 16992
rect 22094 16940 22100 16992
rect 22152 16980 22158 16992
rect 22373 16983 22431 16989
rect 22373 16980 22385 16983
rect 22152 16952 22385 16980
rect 22152 16940 22158 16952
rect 22373 16949 22385 16952
rect 22419 16949 22431 16983
rect 22373 16943 22431 16949
rect 23109 16983 23167 16989
rect 23109 16949 23121 16983
rect 23155 16980 23167 16983
rect 23750 16980 23756 16992
rect 23155 16952 23756 16980
rect 23155 16949 23167 16952
rect 23109 16943 23167 16949
rect 23750 16940 23756 16952
rect 23808 16940 23814 16992
rect 23842 16940 23848 16992
rect 23900 16940 23906 16992
rect 24504 16980 24532 17008
rect 25130 16980 25136 16992
rect 24504 16952 25136 16980
rect 25130 16940 25136 16952
rect 25188 16940 25194 16992
rect 25866 16940 25872 16992
rect 25924 16980 25930 16992
rect 26234 16980 26240 16992
rect 25924 16952 26240 16980
rect 25924 16940 25930 16952
rect 26234 16940 26240 16952
rect 26292 16940 26298 16992
rect 26602 16940 26608 16992
rect 26660 16940 26666 16992
rect 26694 16940 26700 16992
rect 26752 16980 26758 16992
rect 28353 16983 28411 16989
rect 28353 16980 28365 16983
rect 26752 16952 28365 16980
rect 26752 16940 26758 16952
rect 28353 16949 28365 16952
rect 28399 16949 28411 16983
rect 28353 16943 28411 16949
rect 29362 16940 29368 16992
rect 29420 16980 29426 16992
rect 29917 16983 29975 16989
rect 29917 16980 29929 16983
rect 29420 16952 29929 16980
rect 29420 16940 29426 16952
rect 29917 16949 29929 16952
rect 29963 16949 29975 16983
rect 29917 16943 29975 16949
rect 552 16890 31072 16912
rect 552 16838 7988 16890
rect 8040 16838 8052 16890
rect 8104 16838 8116 16890
rect 8168 16838 8180 16890
rect 8232 16838 8244 16890
rect 8296 16838 15578 16890
rect 15630 16838 15642 16890
rect 15694 16838 15706 16890
rect 15758 16838 15770 16890
rect 15822 16838 15834 16890
rect 15886 16838 23168 16890
rect 23220 16838 23232 16890
rect 23284 16838 23296 16890
rect 23348 16838 23360 16890
rect 23412 16838 23424 16890
rect 23476 16838 30758 16890
rect 30810 16838 30822 16890
rect 30874 16838 30886 16890
rect 30938 16838 30950 16890
rect 31002 16838 31014 16890
rect 31066 16838 31072 16890
rect 552 16816 31072 16838
rect 1210 16736 1216 16788
rect 1268 16776 1274 16788
rect 3145 16779 3203 16785
rect 1268 16748 2774 16776
rect 1268 16736 1274 16748
rect 658 16668 664 16720
rect 716 16668 722 16720
rect 676 16640 704 16668
rect 1320 16649 1348 16748
rect 2746 16708 2774 16748
rect 3145 16745 3157 16779
rect 3191 16776 3203 16779
rect 3234 16776 3240 16788
rect 3191 16748 3240 16776
rect 3191 16745 3203 16748
rect 3145 16739 3203 16745
rect 3234 16736 3240 16748
rect 3292 16736 3298 16788
rect 3979 16779 4037 16785
rect 3979 16745 3991 16779
rect 4025 16776 4037 16779
rect 4246 16776 4252 16788
rect 4025 16748 4252 16776
rect 4025 16745 4037 16748
rect 3979 16739 4037 16745
rect 4246 16736 4252 16748
rect 4304 16776 4310 16788
rect 6279 16779 6337 16785
rect 6279 16776 6291 16779
rect 4304 16748 6291 16776
rect 4304 16736 4310 16748
rect 6279 16745 6291 16748
rect 6325 16745 6337 16779
rect 6279 16739 6337 16745
rect 7006 16736 7012 16788
rect 7064 16776 7070 16788
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 7064 16748 7665 16776
rect 7064 16736 7070 16748
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 7653 16739 7711 16745
rect 8021 16779 8079 16785
rect 8021 16745 8033 16779
rect 8067 16776 8079 16779
rect 9306 16776 9312 16788
rect 8067 16748 9312 16776
rect 8067 16745 8079 16748
rect 8021 16739 8079 16745
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 9582 16736 9588 16788
rect 9640 16776 9646 16788
rect 9640 16748 10364 16776
rect 9640 16736 9646 16748
rect 3326 16708 3332 16720
rect 2746 16680 3332 16708
rect 3326 16668 3332 16680
rect 3384 16708 3390 16720
rect 3384 16680 3556 16708
rect 3384 16668 3390 16680
rect 1670 16649 1676 16652
rect 1213 16643 1271 16649
rect 1213 16640 1225 16643
rect 676 16612 1225 16640
rect 1213 16609 1225 16612
rect 1259 16609 1271 16643
rect 1213 16603 1271 16609
rect 1305 16643 1363 16649
rect 1305 16609 1317 16643
rect 1351 16609 1363 16643
rect 1305 16603 1363 16609
rect 1632 16643 1676 16649
rect 1632 16609 1644 16643
rect 1632 16603 1676 16609
rect 1670 16600 1676 16603
rect 1728 16600 1734 16652
rect 3050 16640 3056 16652
rect 1964 16612 3056 16640
rect 1801 16593 1859 16599
rect 1801 16559 1813 16593
rect 1847 16572 1859 16593
rect 1964 16572 1992 16612
rect 3050 16600 3056 16612
rect 3108 16600 3114 16652
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 3418 16640 3424 16652
rect 3292 16612 3424 16640
rect 3292 16600 3298 16612
rect 3418 16600 3424 16612
rect 3476 16600 3482 16652
rect 3528 16649 3556 16680
rect 5626 16668 5632 16720
rect 5684 16668 5690 16720
rect 5902 16668 5908 16720
rect 5960 16668 5966 16720
rect 10336 16708 10364 16748
rect 10410 16736 10416 16788
rect 10468 16736 10474 16788
rect 10870 16736 10876 16788
rect 10928 16776 10934 16788
rect 12618 16776 12624 16788
rect 10928 16748 12624 16776
rect 10928 16736 10934 16748
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 12802 16736 12808 16788
rect 12860 16776 12866 16788
rect 13449 16779 13507 16785
rect 13449 16776 13461 16779
rect 12860 16748 13461 16776
rect 12860 16736 12866 16748
rect 13449 16745 13461 16748
rect 13495 16745 13507 16779
rect 13449 16739 13507 16745
rect 14283 16779 14341 16785
rect 14283 16745 14295 16779
rect 14329 16776 14341 16779
rect 14458 16776 14464 16788
rect 14329 16748 14464 16776
rect 14329 16745 14341 16748
rect 14283 16739 14341 16745
rect 14458 16736 14464 16748
rect 14516 16776 14522 16788
rect 14826 16776 14832 16788
rect 14516 16748 14832 16776
rect 14516 16736 14522 16748
rect 14826 16736 14832 16748
rect 14884 16736 14890 16788
rect 15286 16736 15292 16788
rect 15344 16776 15350 16788
rect 15657 16779 15715 16785
rect 15657 16776 15669 16779
rect 15344 16748 15669 16776
rect 15344 16736 15350 16748
rect 15657 16745 15669 16748
rect 15703 16745 15715 16779
rect 15657 16739 15715 16745
rect 16114 16736 16120 16788
rect 16172 16736 16178 16788
rect 16758 16736 16764 16788
rect 16816 16776 16822 16788
rect 17494 16776 17500 16788
rect 17552 16785 17558 16788
rect 16816 16748 17500 16776
rect 16816 16736 16822 16748
rect 17494 16736 17500 16748
rect 17552 16776 17561 16785
rect 17552 16748 17597 16776
rect 17552 16739 17561 16748
rect 17552 16736 17558 16739
rect 18046 16736 18052 16788
rect 18104 16776 18110 16788
rect 18104 16748 20760 16776
rect 18104 16736 18110 16748
rect 8404 16680 8708 16708
rect 10336 16680 11284 16708
rect 3513 16643 3571 16649
rect 3513 16609 3525 16643
rect 3559 16640 3571 16643
rect 3786 16640 3792 16652
rect 3559 16612 3792 16640
rect 3559 16609 3571 16612
rect 3513 16603 3571 16609
rect 3786 16600 3792 16612
rect 3844 16600 3850 16652
rect 4249 16643 4307 16649
rect 4249 16609 4261 16643
rect 4295 16640 4307 16643
rect 5350 16640 5356 16652
rect 4295 16612 5356 16640
rect 4295 16609 4307 16612
rect 4249 16603 4307 16609
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 5813 16643 5871 16649
rect 5813 16609 5825 16643
rect 5859 16640 5871 16643
rect 5920 16640 5948 16668
rect 5859 16612 5948 16640
rect 6549 16643 6607 16649
rect 5859 16609 5871 16612
rect 5813 16603 5871 16609
rect 6549 16609 6561 16643
rect 6595 16640 6607 16643
rect 8110 16640 8116 16652
rect 6595 16612 8116 16640
rect 6595 16609 6607 16612
rect 6549 16603 6607 16609
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 8205 16643 8263 16649
rect 8205 16609 8217 16643
rect 8251 16609 8263 16643
rect 8205 16603 8263 16609
rect 1847 16559 1992 16572
rect 1801 16553 1992 16559
rect 1826 16544 1992 16553
rect 2038 16532 2044 16584
rect 2096 16532 2102 16584
rect 3976 16577 4034 16583
rect 3976 16543 3988 16577
rect 4022 16572 4034 16577
rect 4062 16572 4068 16584
rect 4022 16544 4068 16572
rect 4022 16543 4034 16544
rect 3976 16537 4034 16543
rect 4062 16532 4068 16544
rect 4120 16532 4126 16584
rect 4430 16532 4436 16584
rect 4488 16572 4494 16584
rect 6362 16583 6368 16584
rect 6319 16577 6368 16583
rect 4488 16544 5028 16572
rect 4488 16532 4494 16544
rect 5000 16516 5028 16544
rect 6319 16543 6331 16577
rect 6365 16543 6368 16577
rect 6319 16537 6368 16543
rect 6362 16532 6368 16537
rect 6420 16532 6426 16584
rect 8220 16516 8248 16603
rect 8404 16572 8432 16680
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16609 8539 16643
rect 8680 16640 8708 16680
rect 9309 16643 9367 16649
rect 9309 16640 9321 16643
rect 8680 16612 9321 16640
rect 8481 16603 8539 16609
rect 9309 16609 9321 16612
rect 9355 16609 9367 16643
rect 10778 16640 10784 16652
rect 9309 16603 9367 16609
rect 9416 16612 10784 16640
rect 8312 16544 8432 16572
rect 4982 16464 4988 16516
rect 5040 16464 5046 16516
rect 8202 16464 8208 16516
rect 8260 16464 8266 16516
rect 8312 16513 8340 16544
rect 8496 16516 8524 16603
rect 8570 16532 8576 16584
rect 8628 16532 8634 16584
rect 8938 16581 8944 16584
rect 8900 16575 8944 16581
rect 8900 16541 8912 16575
rect 8900 16535 8944 16541
rect 8938 16532 8944 16535
rect 8996 16532 9002 16584
rect 9079 16577 9137 16583
rect 9079 16543 9091 16577
rect 9125 16572 9137 16577
rect 9416 16572 9444 16612
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 11149 16643 11207 16649
rect 11149 16640 11161 16643
rect 11072 16612 11161 16640
rect 9125 16544 9444 16572
rect 9125 16543 9137 16544
rect 9079 16537 9137 16543
rect 9490 16532 9496 16584
rect 9548 16572 9554 16584
rect 11072 16572 11100 16612
rect 11149 16609 11161 16612
rect 11195 16609 11207 16643
rect 11149 16603 11207 16609
rect 9548 16544 11100 16572
rect 11256 16572 11284 16680
rect 11330 16600 11336 16652
rect 11388 16640 11394 16652
rect 11609 16643 11667 16649
rect 11609 16640 11621 16643
rect 11388 16612 11621 16640
rect 11388 16600 11394 16612
rect 11609 16609 11621 16612
rect 11655 16609 11667 16643
rect 11609 16603 11667 16609
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 11974 16649 11980 16652
rect 11936 16643 11980 16649
rect 11936 16640 11948 16643
rect 11756 16612 11948 16640
rect 11756 16600 11762 16612
rect 11936 16609 11948 16612
rect 11936 16603 11980 16609
rect 11974 16600 11980 16603
rect 12032 16600 12038 16652
rect 12360 16640 12480 16644
rect 12120 16616 12480 16640
rect 12120 16612 12388 16616
rect 12120 16583 12148 16612
rect 12105 16577 12163 16583
rect 11256 16544 11468 16572
rect 9548 16532 9554 16544
rect 8297 16507 8355 16513
rect 8297 16473 8309 16507
rect 8343 16473 8355 16507
rect 8297 16467 8355 16473
rect 8478 16464 8484 16516
rect 8536 16464 8542 16516
rect 11440 16513 11468 16544
rect 12105 16543 12117 16577
rect 12151 16543 12163 16577
rect 12105 16537 12163 16543
rect 12250 16532 12256 16584
rect 12308 16572 12314 16584
rect 12345 16575 12403 16581
rect 12345 16572 12357 16575
rect 12308 16544 12357 16572
rect 12308 16532 12314 16544
rect 12345 16541 12357 16544
rect 12391 16541 12403 16575
rect 12452 16572 12480 16616
rect 13817 16643 13875 16649
rect 13817 16609 13829 16643
rect 13863 16640 13875 16643
rect 14182 16640 14188 16652
rect 13863 16612 14188 16640
rect 13863 16609 13875 16612
rect 13817 16603 13875 16609
rect 14182 16600 14188 16612
rect 14240 16600 14246 16652
rect 16132 16640 16160 16736
rect 20732 16720 20760 16748
rect 20806 16736 20812 16788
rect 20864 16736 20870 16788
rect 20993 16779 21051 16785
rect 20993 16745 21005 16779
rect 21039 16776 21051 16779
rect 22738 16776 22744 16788
rect 21039 16748 22744 16776
rect 21039 16745 21051 16748
rect 20993 16739 21051 16745
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 23842 16776 23848 16788
rect 22940 16748 23848 16776
rect 20714 16668 20720 16720
rect 20772 16668 20778 16720
rect 14292 16612 16160 16640
rect 16393 16643 16451 16649
rect 14292 16583 14320 16612
rect 16393 16609 16405 16643
rect 16439 16640 16451 16643
rect 16574 16640 16580 16652
rect 16439 16612 16580 16640
rect 16439 16609 16451 16612
rect 16393 16603 16451 16609
rect 16574 16600 16580 16612
rect 16632 16640 16638 16652
rect 16669 16643 16727 16649
rect 16669 16640 16681 16643
rect 16632 16612 16681 16640
rect 16632 16600 16638 16612
rect 16669 16609 16681 16612
rect 16715 16609 16727 16643
rect 19518 16640 19524 16652
rect 17604 16624 19524 16640
rect 16669 16603 16727 16609
rect 17548 16612 19524 16624
rect 17548 16599 17632 16612
rect 19518 16600 19524 16612
rect 19576 16600 19582 16652
rect 19705 16643 19763 16649
rect 19705 16609 19717 16643
rect 19751 16640 19763 16643
rect 20824 16640 20852 16736
rect 21596 16643 21654 16649
rect 21596 16640 21608 16643
rect 19751 16612 20852 16640
rect 21192 16612 21608 16640
rect 19751 16609 19763 16612
rect 19705 16603 19763 16609
rect 17533 16596 17632 16599
rect 17533 16593 17591 16596
rect 14280 16577 14338 16583
rect 12452 16544 13768 16572
rect 12345 16535 12403 16541
rect 11425 16507 11483 16513
rect 11425 16473 11437 16507
rect 11471 16504 11483 16507
rect 11471 16476 11658 16504
rect 11471 16473 11483 16476
rect 11425 16467 11483 16473
rect 1026 16396 1032 16448
rect 1084 16396 1090 16448
rect 3970 16396 3976 16448
rect 4028 16436 4034 16448
rect 11054 16436 11060 16448
rect 4028 16408 11060 16436
rect 4028 16396 4034 16408
rect 11054 16396 11060 16408
rect 11112 16396 11118 16448
rect 11630 16436 11658 16476
rect 12158 16436 12164 16448
rect 11630 16408 12164 16436
rect 12158 16396 12164 16408
rect 12216 16396 12222 16448
rect 13740 16436 13768 16544
rect 14280 16543 14292 16577
rect 14326 16543 14338 16577
rect 14280 16537 14338 16543
rect 14553 16575 14611 16581
rect 14553 16541 14565 16575
rect 14599 16572 14611 16575
rect 14642 16572 14648 16584
rect 14599 16544 14648 16572
rect 14599 16541 14611 16544
rect 14553 16535 14611 16541
rect 14642 16532 14648 16544
rect 14700 16532 14706 16584
rect 17037 16575 17095 16581
rect 17037 16541 17049 16575
rect 17083 16572 17095 16575
rect 17218 16572 17224 16584
rect 17083 16544 17224 16572
rect 17083 16541 17095 16544
rect 17037 16535 17095 16541
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 17533 16559 17545 16593
rect 17579 16559 17591 16593
rect 21192 16584 21220 16612
rect 21596 16609 21608 16612
rect 21642 16609 21654 16643
rect 21596 16603 21654 16609
rect 22005 16643 22063 16649
rect 22005 16609 22017 16643
rect 22051 16640 22063 16643
rect 22940 16640 22968 16748
rect 23842 16736 23848 16748
rect 23900 16736 23906 16788
rect 23943 16779 24001 16785
rect 23943 16745 23955 16779
rect 23989 16776 24001 16779
rect 24302 16776 24308 16788
rect 23989 16748 24308 16776
rect 23989 16745 24001 16748
rect 23943 16739 24001 16745
rect 24302 16736 24308 16748
rect 24360 16776 24366 16788
rect 24486 16776 24492 16788
rect 24360 16748 24492 16776
rect 24360 16736 24366 16748
rect 24486 16736 24492 16748
rect 24544 16736 24550 16788
rect 26050 16736 26056 16788
rect 26108 16736 26114 16788
rect 26789 16779 26847 16785
rect 26789 16745 26801 16779
rect 26835 16776 26847 16779
rect 26878 16776 26884 16788
rect 26835 16748 26884 16776
rect 26835 16745 26847 16748
rect 26789 16739 26847 16745
rect 26878 16736 26884 16748
rect 26936 16736 26942 16788
rect 27798 16736 27804 16788
rect 27856 16776 27862 16788
rect 28267 16779 28325 16785
rect 28267 16776 28279 16779
rect 27856 16748 28279 16776
rect 27856 16736 27862 16748
rect 28267 16745 28279 16748
rect 28313 16776 28325 16779
rect 28534 16776 28540 16788
rect 28313 16748 28540 16776
rect 28313 16745 28325 16748
rect 28267 16739 28325 16745
rect 28534 16736 28540 16748
rect 28592 16736 28598 16788
rect 29638 16736 29644 16788
rect 29696 16736 29702 16788
rect 30374 16736 30380 16788
rect 30432 16736 30438 16788
rect 23014 16668 23020 16720
rect 23072 16708 23078 16720
rect 23385 16711 23443 16717
rect 23385 16708 23397 16711
rect 23072 16680 23397 16708
rect 23072 16668 23078 16680
rect 23385 16677 23397 16680
rect 23431 16677 23443 16711
rect 30101 16711 30159 16717
rect 23385 16671 23443 16677
rect 24872 16680 27476 16708
rect 22051 16612 22968 16640
rect 23477 16643 23535 16649
rect 22051 16609 22063 16612
rect 22005 16603 22063 16609
rect 23477 16609 23489 16643
rect 23523 16640 23535 16643
rect 23750 16640 23756 16652
rect 23523 16612 23756 16640
rect 23523 16609 23535 16612
rect 23477 16603 23535 16609
rect 23750 16600 23756 16612
rect 23808 16600 23814 16652
rect 23842 16600 23848 16652
rect 23900 16600 23906 16652
rect 24044 16612 24348 16640
rect 17533 16553 17591 16559
rect 17678 16532 17684 16584
rect 17736 16572 17742 16584
rect 17773 16575 17831 16581
rect 17773 16572 17785 16575
rect 17736 16544 17785 16572
rect 17736 16532 17742 16544
rect 17773 16541 17785 16544
rect 17819 16541 17831 16575
rect 17773 16535 17831 16541
rect 19426 16532 19432 16584
rect 19484 16572 19490 16584
rect 20622 16572 20628 16584
rect 19484 16544 20628 16572
rect 19484 16532 19490 16544
rect 20622 16532 20628 16544
rect 20680 16532 20686 16584
rect 21174 16532 21180 16584
rect 21232 16532 21238 16584
rect 21266 16532 21272 16584
rect 21324 16532 21330 16584
rect 21775 16575 21833 16581
rect 21775 16541 21787 16575
rect 21821 16572 21833 16575
rect 23860 16572 23888 16600
rect 21821 16544 23888 16572
rect 23956 16575 24014 16581
rect 21821 16541 21833 16544
rect 21775 16535 21833 16541
rect 23956 16541 23968 16575
rect 24002 16572 24014 16575
rect 24044 16572 24072 16612
rect 24002 16544 24072 16572
rect 24002 16541 24014 16544
rect 23956 16535 24014 16541
rect 24118 16532 24124 16584
rect 24176 16572 24182 16584
rect 24213 16575 24271 16581
rect 24213 16572 24225 16575
rect 24176 16544 24225 16572
rect 24176 16532 24182 16544
rect 24213 16541 24225 16544
rect 24259 16541 24271 16575
rect 24320 16572 24348 16612
rect 24486 16600 24492 16652
rect 24544 16640 24550 16652
rect 24872 16640 24900 16680
rect 27448 16652 27476 16680
rect 30101 16677 30113 16711
rect 30147 16708 30159 16711
rect 30190 16708 30196 16720
rect 30147 16680 30196 16708
rect 30147 16677 30159 16680
rect 30101 16671 30159 16677
rect 30190 16668 30196 16680
rect 30248 16668 30254 16720
rect 24544 16612 24900 16640
rect 24544 16600 24550 16612
rect 25774 16600 25780 16652
rect 25832 16600 25838 16652
rect 26234 16600 26240 16652
rect 26292 16640 26298 16652
rect 26697 16643 26755 16649
rect 26697 16640 26709 16643
rect 26292 16612 26709 16640
rect 26292 16600 26298 16612
rect 26697 16609 26709 16612
rect 26743 16609 26755 16643
rect 26697 16603 26755 16609
rect 26786 16600 26792 16652
rect 26844 16640 26850 16652
rect 27249 16643 27307 16649
rect 27249 16640 27261 16643
rect 26844 16612 27261 16640
rect 26844 16600 26850 16612
rect 27249 16609 27261 16612
rect 27295 16609 27307 16643
rect 27249 16603 27307 16609
rect 27430 16600 27436 16652
rect 27488 16600 27494 16652
rect 27614 16600 27620 16652
rect 27672 16640 27678 16652
rect 27801 16643 27859 16649
rect 27801 16640 27813 16643
rect 27672 16612 27813 16640
rect 27672 16600 27678 16612
rect 27801 16609 27813 16612
rect 27847 16640 27859 16643
rect 28166 16640 28172 16652
rect 27847 16612 28172 16640
rect 27847 16609 27859 16612
rect 27801 16603 27859 16609
rect 28166 16600 28172 16612
rect 28224 16600 28230 16652
rect 28537 16643 28595 16649
rect 28537 16609 28549 16643
rect 28583 16640 28595 16643
rect 28994 16640 29000 16652
rect 28583 16612 29000 16640
rect 28583 16609 28595 16612
rect 28537 16603 28595 16609
rect 28994 16600 29000 16612
rect 29052 16600 29058 16652
rect 27522 16572 27528 16584
rect 24320 16544 27528 16572
rect 24213 16535 24271 16541
rect 27522 16532 27528 16544
rect 27580 16532 27586 16584
rect 28307 16575 28365 16581
rect 28307 16541 28319 16575
rect 28353 16572 28365 16575
rect 28442 16572 28448 16584
rect 28353 16544 28448 16572
rect 28353 16541 28365 16544
rect 28307 16535 28365 16541
rect 28442 16532 28448 16544
rect 28500 16532 28506 16584
rect 15470 16464 15476 16516
rect 15528 16504 15534 16516
rect 16298 16504 16304 16516
rect 15528 16476 16304 16504
rect 15528 16464 15534 16476
rect 16298 16464 16304 16476
rect 16356 16504 16362 16516
rect 16850 16504 16856 16516
rect 16356 16476 16856 16504
rect 16356 16464 16362 16476
rect 16850 16464 16856 16476
rect 16908 16464 16914 16516
rect 18506 16464 18512 16516
rect 18564 16504 18570 16516
rect 18564 16476 19012 16504
rect 18564 16464 18570 16476
rect 15930 16436 15936 16448
rect 13740 16408 15936 16436
rect 15930 16396 15936 16408
rect 15988 16396 15994 16448
rect 16209 16439 16267 16445
rect 16209 16405 16221 16439
rect 16255 16436 16267 16439
rect 18782 16436 18788 16448
rect 16255 16408 18788 16436
rect 16255 16405 16267 16408
rect 16209 16399 16267 16405
rect 18782 16396 18788 16408
rect 18840 16396 18846 16448
rect 18874 16396 18880 16448
rect 18932 16396 18938 16448
rect 18984 16436 19012 16476
rect 23474 16436 23480 16448
rect 18984 16408 23480 16436
rect 23474 16396 23480 16408
rect 23532 16396 23538 16448
rect 23934 16396 23940 16448
rect 23992 16436 23998 16448
rect 25130 16436 25136 16448
rect 23992 16408 25136 16436
rect 23992 16396 23998 16408
rect 25130 16396 25136 16408
rect 25188 16396 25194 16448
rect 25314 16396 25320 16448
rect 25372 16396 25378 16448
rect 26418 16396 26424 16448
rect 26476 16436 26482 16448
rect 27525 16439 27583 16445
rect 27525 16436 27537 16439
rect 26476 16408 27537 16436
rect 26476 16396 26482 16408
rect 27525 16405 27537 16408
rect 27571 16436 27583 16439
rect 28902 16436 28908 16448
rect 27571 16408 28908 16436
rect 27571 16405 27583 16408
rect 27525 16399 27583 16405
rect 28902 16396 28908 16408
rect 28960 16396 28966 16448
rect 552 16346 30912 16368
rect 552 16294 4193 16346
rect 4245 16294 4257 16346
rect 4309 16294 4321 16346
rect 4373 16294 4385 16346
rect 4437 16294 4449 16346
rect 4501 16294 11783 16346
rect 11835 16294 11847 16346
rect 11899 16294 11911 16346
rect 11963 16294 11975 16346
rect 12027 16294 12039 16346
rect 12091 16294 19373 16346
rect 19425 16294 19437 16346
rect 19489 16294 19501 16346
rect 19553 16294 19565 16346
rect 19617 16294 19629 16346
rect 19681 16294 26963 16346
rect 27015 16294 27027 16346
rect 27079 16294 27091 16346
rect 27143 16294 27155 16346
rect 27207 16294 27219 16346
rect 27271 16294 30912 16346
rect 552 16272 30912 16294
rect 2958 16192 2964 16244
rect 3016 16192 3022 16244
rect 3970 16232 3976 16244
rect 3712 16204 3976 16232
rect 937 16099 995 16105
rect 937 16065 949 16099
rect 983 16096 995 16099
rect 1118 16096 1124 16108
rect 983 16068 1124 16096
rect 983 16065 995 16068
rect 937 16059 995 16065
rect 1118 16056 1124 16068
rect 1176 16056 1182 16108
rect 1443 16099 1501 16105
rect 1443 16065 1455 16099
rect 1489 16096 1501 16099
rect 3510 16096 3516 16108
rect 1489 16068 3516 16096
rect 1489 16065 1501 16068
rect 1443 16059 1501 16065
rect 3510 16056 3516 16068
rect 3568 16056 3574 16108
rect 1673 16031 1731 16037
rect 1673 15997 1685 16031
rect 1719 16028 1731 16031
rect 3712 16028 3740 16204
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 4062 16192 4068 16244
rect 4120 16232 4126 16244
rect 5629 16235 5687 16241
rect 5629 16232 5641 16235
rect 4120 16204 5641 16232
rect 4120 16192 4126 16204
rect 5629 16201 5641 16204
rect 5675 16201 5687 16235
rect 7929 16235 7987 16241
rect 7929 16232 7941 16235
rect 5629 16195 5687 16201
rect 6104 16204 7941 16232
rect 4295 16099 4353 16105
rect 4295 16065 4307 16099
rect 4341 16096 4353 16099
rect 6104 16096 6132 16204
rect 7929 16201 7941 16204
rect 7975 16201 7987 16235
rect 7929 16195 7987 16201
rect 8570 16192 8576 16244
rect 8628 16232 8634 16244
rect 10965 16235 11023 16241
rect 8628 16204 9996 16232
rect 8628 16192 8634 16204
rect 6638 16103 6644 16108
rect 4341 16068 6132 16096
rect 6595 16097 6644 16103
rect 4341 16065 4353 16068
rect 4295 16059 4353 16065
rect 6595 16063 6607 16097
rect 6641 16063 6644 16097
rect 6595 16057 6644 16063
rect 6638 16056 6644 16057
rect 6696 16056 6702 16108
rect 8588 16105 8616 16192
rect 9968 16164 9996 16204
rect 10965 16201 10977 16235
rect 11011 16232 11023 16235
rect 20530 16232 20536 16244
rect 11011 16204 12664 16232
rect 11011 16201 11023 16204
rect 10965 16195 11023 16201
rect 11054 16164 11060 16176
rect 9968 16136 11060 16164
rect 11054 16124 11060 16136
rect 11112 16124 11118 16176
rect 12636 16164 12664 16204
rect 14476 16204 16528 16232
rect 13722 16164 13728 16176
rect 12636 16136 13728 16164
rect 13722 16124 13728 16136
rect 13780 16124 13786 16176
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16065 8631 16099
rect 8573 16059 8631 16065
rect 8754 16056 8760 16108
rect 8812 16056 8818 16108
rect 9079 16099 9137 16105
rect 9079 16065 9091 16099
rect 9125 16096 9137 16099
rect 11514 16096 11520 16108
rect 9125 16068 11520 16096
rect 9125 16065 9137 16068
rect 9079 16059 9137 16065
rect 11514 16056 11520 16068
rect 11572 16056 11578 16108
rect 11747 16099 11805 16105
rect 11747 16065 11759 16099
rect 11793 16096 11805 16099
rect 14476 16096 14504 16204
rect 16500 16173 16528 16204
rect 16874 16204 20536 16232
rect 16485 16167 16543 16173
rect 16485 16133 16497 16167
rect 16531 16133 16543 16167
rect 16485 16127 16543 16133
rect 14826 16096 14832 16108
rect 11793 16068 14504 16096
rect 14568 16068 14832 16096
rect 11793 16065 11805 16068
rect 11747 16059 11805 16065
rect 1719 16000 3740 16028
rect 3789 16031 3847 16037
rect 1719 15997 1731 16000
rect 1673 15991 1731 15997
rect 3789 15997 3801 16031
rect 3835 15997 3847 16031
rect 3789 15991 3847 15997
rect 3326 15920 3332 15972
rect 3384 15920 3390 15972
rect 3804 15960 3832 15991
rect 3878 15988 3884 16040
rect 3936 16028 3942 16040
rect 4116 16031 4174 16037
rect 4116 16028 4128 16031
rect 3936 16000 4128 16028
rect 3936 15988 3942 16000
rect 4116 15997 4128 16000
rect 4162 15997 4174 16031
rect 4116 15991 4174 15997
rect 4522 15988 4528 16040
rect 4580 15988 4586 16040
rect 6086 15988 6092 16040
rect 6144 15988 6150 16040
rect 6454 16037 6460 16040
rect 6416 16031 6460 16037
rect 6416 15997 6428 16031
rect 6416 15991 6460 15997
rect 6454 15988 6460 15991
rect 6512 15988 6518 16040
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 7650 16028 7656 16040
rect 6871 16000 7656 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 7650 15988 7656 16000
rect 7708 15988 7714 16040
rect 8202 15988 8208 16040
rect 8260 16028 8266 16040
rect 8772 16028 8800 16056
rect 8260 16000 8800 16028
rect 8260 15988 8266 16000
rect 9214 15988 9220 16040
rect 9272 16028 9278 16040
rect 9309 16031 9367 16037
rect 9309 16028 9321 16031
rect 9272 16000 9321 16028
rect 9272 15988 9278 16000
rect 9309 15997 9321 16000
rect 9355 15997 9367 16031
rect 9309 15991 9367 15997
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 15997 11207 16031
rect 11149 15991 11207 15997
rect 11241 16031 11299 16037
rect 11241 15997 11253 16031
rect 11287 16028 11299 16031
rect 11330 16028 11336 16040
rect 11287 16000 11336 16028
rect 11287 15997 11299 16000
rect 11241 15991 11299 15997
rect 3620 15932 3832 15960
rect 1394 15852 1400 15904
rect 1452 15901 1458 15904
rect 1452 15855 1461 15901
rect 1452 15852 1458 15855
rect 3510 15852 3516 15904
rect 3568 15892 3574 15904
rect 3620 15901 3648 15932
rect 11164 15904 11192 15991
rect 11330 15988 11336 16000
rect 11388 15988 11394 16040
rect 11606 15988 11612 16040
rect 11664 16028 11670 16040
rect 11977 16031 12035 16037
rect 11977 16028 11989 16031
rect 11664 16000 11989 16028
rect 11664 15988 11670 16000
rect 11977 15997 11989 16000
rect 12023 15997 12035 16031
rect 11977 15991 12035 15997
rect 12342 15988 12348 16040
rect 12400 16028 12406 16040
rect 12400 16000 12664 16028
rect 12400 15988 12406 16000
rect 12636 15960 12664 16000
rect 14182 15988 14188 16040
rect 14240 16028 14246 16040
rect 14568 16037 14596 16068
rect 14826 16056 14832 16068
rect 14884 16056 14890 16108
rect 14918 16056 14924 16108
rect 14976 16105 14982 16108
rect 14976 16099 15030 16105
rect 14976 16065 14984 16099
rect 15018 16065 15030 16099
rect 14976 16059 15030 16065
rect 15108 16097 15166 16103
rect 15108 16063 15120 16097
rect 15154 16063 15166 16097
rect 14976 16056 14982 16059
rect 15108 16057 15166 16063
rect 14553 16031 14611 16037
rect 14240 16000 14504 16028
rect 14240 15988 14246 16000
rect 13817 15963 13875 15969
rect 12636 15932 13216 15960
rect 3605 15895 3663 15901
rect 3605 15892 3617 15895
rect 3568 15864 3617 15892
rect 3568 15852 3574 15864
rect 3605 15861 3617 15864
rect 3651 15861 3663 15895
rect 3605 15855 3663 15861
rect 4154 15852 4160 15904
rect 4212 15892 4218 15904
rect 7834 15892 7840 15904
rect 4212 15864 7840 15892
rect 4212 15852 4218 15864
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 8938 15852 8944 15904
rect 8996 15892 9002 15904
rect 9039 15895 9097 15901
rect 9039 15892 9051 15895
rect 8996 15864 9051 15892
rect 8996 15852 9002 15864
rect 9039 15861 9051 15864
rect 9085 15861 9097 15895
rect 9039 15855 9097 15861
rect 10410 15852 10416 15904
rect 10468 15852 10474 15904
rect 11146 15852 11152 15904
rect 11204 15852 11210 15904
rect 11698 15852 11704 15904
rect 11756 15901 11762 15904
rect 11756 15892 11765 15901
rect 11756 15864 11801 15892
rect 11756 15855 11765 15864
rect 11756 15852 11762 15855
rect 13078 15852 13084 15904
rect 13136 15852 13142 15904
rect 13188 15892 13216 15932
rect 13817 15929 13829 15963
rect 13863 15960 13875 15963
rect 13906 15960 13912 15972
rect 13863 15932 13912 15960
rect 13863 15929 13875 15932
rect 13817 15923 13875 15929
rect 13906 15920 13912 15932
rect 13964 15960 13970 15972
rect 14274 15960 14280 15972
rect 13964 15932 14280 15960
rect 13964 15920 13970 15932
rect 14274 15920 14280 15932
rect 14332 15920 14338 15972
rect 14476 15960 14504 16000
rect 14553 15997 14565 16031
rect 14599 15997 14611 16031
rect 14553 15991 14611 15997
rect 14642 15988 14648 16040
rect 14700 15988 14706 16040
rect 15123 16028 15151 16057
rect 15194 16056 15200 16108
rect 15252 16096 15258 16108
rect 16874 16096 16902 16204
rect 20530 16192 20536 16204
rect 20588 16192 20594 16244
rect 22370 16232 22376 16244
rect 20640 16204 22376 16232
rect 18417 16167 18475 16173
rect 18417 16133 18429 16167
rect 18463 16164 18475 16167
rect 18506 16164 18512 16176
rect 18463 16136 18512 16164
rect 18463 16133 18475 16136
rect 18417 16127 18475 16133
rect 18506 16124 18512 16136
rect 18564 16124 18570 16176
rect 15252 16068 16902 16096
rect 15252 16056 15258 16068
rect 17494 16056 17500 16108
rect 17552 16096 17558 16108
rect 19020 16099 19078 16105
rect 19020 16096 19032 16099
rect 17552 16068 19032 16096
rect 17552 16056 17558 16068
rect 19020 16065 19032 16068
rect 19066 16065 19078 16099
rect 19020 16059 19078 16065
rect 19199 16099 19257 16105
rect 19199 16065 19211 16099
rect 19245 16096 19257 16099
rect 20640 16096 20668 16204
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 23569 16235 23627 16241
rect 23569 16201 23581 16235
rect 23615 16232 23627 16235
rect 24578 16232 24584 16244
rect 23615 16204 24584 16232
rect 23615 16201 23627 16204
rect 23569 16195 23627 16201
rect 24578 16192 24584 16204
rect 24636 16192 24642 16244
rect 25958 16192 25964 16244
rect 26016 16232 26022 16244
rect 30285 16235 30343 16241
rect 30285 16232 30297 16235
rect 26016 16204 28488 16232
rect 26016 16192 26022 16204
rect 20714 16124 20720 16176
rect 20772 16124 20778 16176
rect 21910 16105 21916 16108
rect 19245 16068 20668 16096
rect 21872 16099 21916 16105
rect 19245 16065 19257 16068
rect 19199 16059 19257 16065
rect 21872 16065 21884 16099
rect 21872 16059 21916 16065
rect 21910 16056 21916 16059
rect 21968 16056 21974 16108
rect 22002 16056 22008 16108
rect 22060 16096 22066 16108
rect 22060 16087 22094 16096
rect 22060 16081 22099 16087
rect 22087 16078 22099 16081
rect 22041 16047 22053 16056
rect 22087 16050 22125 16078
rect 23750 16056 23756 16108
rect 23808 16096 23814 16108
rect 24210 16105 24216 16108
rect 23845 16099 23903 16105
rect 23845 16096 23857 16099
rect 23808 16068 23857 16096
rect 23808 16056 23814 16068
rect 23845 16065 23857 16068
rect 23891 16065 23903 16099
rect 23845 16059 23903 16065
rect 24172 16099 24216 16105
rect 24172 16065 24184 16099
rect 24172 16059 24216 16065
rect 24210 16056 24216 16059
rect 24268 16056 24274 16108
rect 24394 16103 24400 16108
rect 24351 16097 24400 16103
rect 24351 16063 24363 16097
rect 24397 16063 24400 16097
rect 24351 16057 24400 16063
rect 24394 16056 24400 16057
rect 24452 16056 24458 16108
rect 24581 16099 24639 16105
rect 24581 16065 24593 16099
rect 24627 16096 24639 16099
rect 24762 16096 24768 16108
rect 24627 16068 24768 16096
rect 24627 16065 24639 16068
rect 24581 16059 24639 16065
rect 24762 16056 24768 16068
rect 24820 16056 24826 16108
rect 26050 16056 26056 16108
rect 26108 16056 26114 16108
rect 26326 16056 26332 16108
rect 26384 16096 26390 16108
rect 26516 16099 26574 16105
rect 26516 16096 26528 16099
rect 26384 16068 26528 16096
rect 26384 16056 26390 16068
rect 26516 16065 26528 16068
rect 26562 16065 26574 16099
rect 26516 16059 26574 16065
rect 26789 16099 26847 16105
rect 26789 16065 26801 16099
rect 26835 16096 26847 16099
rect 27890 16096 27896 16108
rect 26835 16068 27896 16096
rect 26835 16065 26847 16068
rect 26789 16059 26847 16065
rect 27890 16056 27896 16068
rect 27948 16056 27954 16108
rect 22087 16047 22099 16050
rect 22041 16041 22099 16047
rect 15286 16028 15292 16040
rect 15123 16000 15292 16028
rect 15286 15988 15292 16000
rect 15344 15988 15350 16040
rect 15378 15988 15384 16040
rect 15436 15988 15442 16040
rect 16666 15988 16672 16040
rect 16724 15988 16730 16040
rect 16850 15988 16856 16040
rect 16908 15988 16914 16040
rect 17126 15988 17132 16040
rect 17184 15988 17190 16040
rect 17218 15988 17224 16040
rect 17276 16028 17282 16040
rect 18693 16031 18751 16037
rect 18693 16028 18705 16031
rect 17276 16000 18705 16028
rect 17276 15988 17282 16000
rect 18693 15997 18705 16000
rect 18739 15997 18751 16031
rect 18693 15991 18751 15997
rect 14666 15960 14694 15988
rect 14476 15932 14694 15960
rect 14093 15895 14151 15901
rect 14093 15892 14105 15895
rect 13188 15864 14105 15892
rect 14093 15861 14105 15864
rect 14139 15861 14151 15895
rect 14093 15855 14151 15861
rect 14369 15895 14427 15901
rect 14369 15861 14381 15895
rect 14415 15892 14427 15895
rect 16684 15892 16712 15988
rect 18414 15960 18420 15972
rect 17788 15932 18420 15960
rect 14415 15864 16712 15892
rect 14415 15861 14427 15864
rect 14369 15855 14427 15861
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 17788 15892 17816 15932
rect 18414 15920 18420 15932
rect 18472 15920 18478 15972
rect 18708 15960 18736 15991
rect 18782 15988 18788 16040
rect 18840 16028 18846 16040
rect 19429 16031 19487 16037
rect 19429 16028 19441 16031
rect 18840 16024 18971 16028
rect 19168 16024 19441 16028
rect 18840 16000 19441 16024
rect 18840 15988 18846 16000
rect 18943 15996 19196 16000
rect 19429 15997 19441 16000
rect 19475 15997 19487 16031
rect 19429 15991 19487 15997
rect 20901 16031 20959 16037
rect 20901 15997 20913 16031
rect 20947 15997 20959 16031
rect 20901 15991 20959 15997
rect 18708 15932 18828 15960
rect 18800 15904 18828 15932
rect 16908 15864 17816 15892
rect 16908 15852 16914 15864
rect 18782 15852 18788 15904
rect 18840 15852 18846 15904
rect 19150 15852 19156 15904
rect 19208 15892 19214 15904
rect 20806 15892 20812 15904
rect 19208 15864 20812 15892
rect 19208 15852 19214 15864
rect 20806 15852 20812 15864
rect 20864 15852 20870 15904
rect 20916 15892 20944 15991
rect 21450 15988 21456 16040
rect 21508 16028 21514 16040
rect 21545 16031 21603 16037
rect 21545 16028 21557 16031
rect 21508 16000 21557 16028
rect 21508 15988 21514 16000
rect 21545 15997 21557 16000
rect 21591 15997 21603 16031
rect 21545 15991 21603 15997
rect 22281 16031 22339 16037
rect 22281 15997 22293 16031
rect 22327 16028 22339 16031
rect 23014 16028 23020 16040
rect 22327 16000 23020 16028
rect 22327 15997 22339 16000
rect 22281 15991 22339 15997
rect 23014 15988 23020 16000
rect 23072 15988 23078 16040
rect 24670 15988 24676 16040
rect 24728 16028 24734 16040
rect 25406 16028 25412 16040
rect 24728 16000 25412 16028
rect 24728 15988 24734 16000
rect 25406 15988 25412 16000
rect 25464 16028 25470 16040
rect 28261 16031 28319 16037
rect 28261 16028 28273 16031
rect 25464 16000 28273 16028
rect 25464 15988 25470 16000
rect 28261 15997 28273 16000
rect 28307 15997 28319 16031
rect 28460 16028 28488 16204
rect 29104 16204 30297 16232
rect 29104 16176 29132 16204
rect 30285 16201 30297 16204
rect 30331 16201 30343 16235
rect 30285 16195 30343 16201
rect 31202 16192 31208 16244
rect 31260 16192 31266 16244
rect 29086 16124 29092 16176
rect 29144 16124 29150 16176
rect 30190 16164 30196 16176
rect 29748 16136 30196 16164
rect 28718 16056 28724 16108
rect 28776 16096 28782 16108
rect 28776 16094 28856 16096
rect 28920 16094 29592 16096
rect 28776 16068 29592 16094
rect 28776 16056 28782 16068
rect 28828 16066 28948 16068
rect 29273 16031 29331 16037
rect 29273 16028 29285 16031
rect 28460 16000 29285 16028
rect 28261 15991 28319 15997
rect 29273 15997 29285 16000
rect 29319 15997 29331 16031
rect 29273 15991 29331 15997
rect 29362 15988 29368 16040
rect 29420 15988 29426 16040
rect 29564 16028 29592 16068
rect 29638 16028 29644 16040
rect 29564 16000 29644 16028
rect 29638 15988 29644 16000
rect 29696 15988 29702 16040
rect 29748 16037 29776 16136
rect 30190 16124 30196 16136
rect 30248 16164 30254 16176
rect 31220 16164 31248 16192
rect 30248 16136 31248 16164
rect 30248 16124 30254 16136
rect 29733 16031 29791 16037
rect 29733 15997 29745 16031
rect 29779 15997 29791 16031
rect 29733 15991 29791 15997
rect 29822 15988 29828 16040
rect 29880 16028 29886 16040
rect 30193 16031 30251 16037
rect 30193 16028 30205 16031
rect 29880 16000 30205 16028
rect 29880 15988 29886 16000
rect 30193 15997 30205 16000
rect 30239 15997 30251 16031
rect 30193 15991 30251 15997
rect 21174 15920 21180 15972
rect 21232 15920 21238 15972
rect 23842 15960 23848 15972
rect 23124 15932 23848 15960
rect 23124 15892 23152 15932
rect 23842 15920 23848 15932
rect 23900 15920 23906 15972
rect 28537 15963 28595 15969
rect 28537 15960 28549 15963
rect 27816 15932 28549 15960
rect 20916 15864 23152 15892
rect 25682 15852 25688 15904
rect 25740 15852 25746 15904
rect 26510 15852 26516 15904
rect 26568 15901 26574 15904
rect 26568 15892 26577 15901
rect 27816 15892 27844 15932
rect 28537 15929 28549 15932
rect 28583 15929 28595 15963
rect 28537 15923 28595 15929
rect 28718 15920 28724 15972
rect 28776 15960 28782 15972
rect 29089 15963 29147 15969
rect 29089 15960 29101 15963
rect 28776 15932 29101 15960
rect 28776 15920 28782 15932
rect 29089 15929 29101 15932
rect 29135 15960 29147 15963
rect 30650 15960 30656 15972
rect 29135 15932 30656 15960
rect 29135 15929 29147 15932
rect 29089 15923 29147 15929
rect 30650 15920 30656 15932
rect 30708 15920 30714 15972
rect 26568 15864 27844 15892
rect 26568 15855 26577 15864
rect 26568 15852 26574 15855
rect 27890 15852 27896 15904
rect 27948 15852 27954 15904
rect 29362 15852 29368 15904
rect 29420 15892 29426 15904
rect 29549 15895 29607 15901
rect 29549 15892 29561 15895
rect 29420 15864 29561 15892
rect 29420 15852 29426 15864
rect 29549 15861 29561 15864
rect 29595 15861 29607 15895
rect 29549 15855 29607 15861
rect 29638 15852 29644 15904
rect 29696 15892 29702 15904
rect 29917 15895 29975 15901
rect 29917 15892 29929 15895
rect 29696 15864 29929 15892
rect 29696 15852 29702 15864
rect 29917 15861 29929 15864
rect 29963 15861 29975 15895
rect 29917 15855 29975 15861
rect 552 15802 31072 15824
rect 552 15750 7988 15802
rect 8040 15750 8052 15802
rect 8104 15750 8116 15802
rect 8168 15750 8180 15802
rect 8232 15750 8244 15802
rect 8296 15750 15578 15802
rect 15630 15750 15642 15802
rect 15694 15750 15706 15802
rect 15758 15750 15770 15802
rect 15822 15750 15834 15802
rect 15886 15750 23168 15802
rect 23220 15750 23232 15802
rect 23284 15750 23296 15802
rect 23348 15750 23360 15802
rect 23412 15750 23424 15802
rect 23476 15750 30758 15802
rect 30810 15750 30822 15802
rect 30874 15750 30886 15802
rect 30938 15750 30950 15802
rect 31002 15750 31014 15802
rect 31066 15750 31072 15802
rect 552 15728 31072 15750
rect 1136 15660 3096 15688
rect 1136 15561 1164 15660
rect 1394 15580 1400 15632
rect 1452 15580 1458 15632
rect 3068 15620 3096 15660
rect 3142 15648 3148 15700
rect 3200 15648 3206 15700
rect 4706 15688 4712 15700
rect 3620 15660 4712 15688
rect 3620 15620 3648 15660
rect 4706 15648 4712 15660
rect 4764 15648 4770 15700
rect 4982 15648 4988 15700
rect 5040 15688 5046 15700
rect 5353 15691 5411 15697
rect 5353 15688 5365 15691
rect 5040 15660 5365 15688
rect 5040 15648 5046 15660
rect 5353 15657 5365 15660
rect 5399 15657 5411 15691
rect 10410 15688 10416 15700
rect 5353 15651 5411 15657
rect 5828 15660 10416 15688
rect 3068 15592 3648 15620
rect 1121 15555 1179 15561
rect 1121 15521 1133 15555
rect 1167 15521 1179 15555
rect 1412 15552 1440 15580
rect 1632 15555 1690 15561
rect 1632 15552 1644 15555
rect 1412 15524 1644 15552
rect 1121 15515 1179 15521
rect 1632 15521 1644 15524
rect 1678 15521 1690 15555
rect 5828 15552 5856 15660
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 13078 15688 13084 15700
rect 10888 15660 13084 15688
rect 1632 15515 1690 15521
rect 1964 15524 5856 15552
rect 5905 15555 5963 15561
rect 1801 15505 1859 15511
rect 1305 15487 1363 15493
rect 1305 15453 1317 15487
rect 1351 15453 1363 15487
rect 1801 15471 1813 15505
rect 1847 15484 1859 15505
rect 1964 15484 1992 15524
rect 5905 15521 5917 15555
rect 5951 15521 5963 15555
rect 5905 15515 5963 15521
rect 1847 15471 1992 15484
rect 1801 15465 1992 15471
rect 1826 15456 1992 15465
rect 2041 15487 2099 15493
rect 1305 15447 1363 15453
rect 2041 15453 2053 15487
rect 2087 15484 2099 15487
rect 2866 15484 2872 15496
rect 2087 15456 2872 15484
rect 2087 15453 2099 15456
rect 2041 15447 2099 15453
rect 1118 15376 1124 15428
rect 1176 15416 1182 15428
rect 1320 15416 1348 15447
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 3510 15444 3516 15496
rect 3568 15444 3574 15496
rect 3878 15493 3884 15496
rect 3840 15487 3884 15493
rect 3840 15453 3852 15487
rect 3840 15447 3884 15453
rect 3878 15444 3884 15447
rect 3936 15444 3942 15496
rect 4019 15487 4077 15493
rect 4019 15453 4031 15487
rect 4065 15484 4077 15487
rect 4154 15484 4160 15496
rect 4065 15456 4160 15484
rect 4065 15453 4077 15456
rect 4019 15447 4077 15453
rect 4154 15444 4160 15456
rect 4212 15444 4218 15496
rect 4249 15487 4307 15493
rect 4249 15453 4261 15487
rect 4295 15484 4307 15487
rect 5442 15484 5448 15496
rect 4295 15456 5448 15484
rect 4295 15453 4307 15456
rect 4249 15447 4307 15453
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 1176 15388 1348 15416
rect 1176 15376 1182 15388
rect 937 15351 995 15357
rect 937 15317 949 15351
rect 983 15348 995 15351
rect 1210 15348 1216 15360
rect 983 15320 1216 15348
rect 983 15317 995 15320
rect 937 15311 995 15317
rect 1210 15308 1216 15320
rect 1268 15308 1274 15360
rect 1320 15348 1348 15388
rect 3528 15348 3556 15444
rect 3786 15348 3792 15360
rect 1320 15320 3792 15348
rect 3786 15308 3792 15320
rect 3844 15348 3850 15360
rect 5920 15348 5948 15515
rect 6454 15512 6460 15564
rect 6512 15512 6518 15564
rect 6876 15524 8340 15552
rect 6086 15444 6092 15496
rect 6144 15484 6150 15496
rect 6181 15487 6239 15493
rect 6181 15484 6193 15487
rect 6144 15456 6193 15484
rect 6144 15444 6150 15456
rect 6181 15453 6193 15456
rect 6227 15484 6239 15487
rect 6365 15487 6423 15493
rect 6365 15484 6377 15487
rect 6227 15456 6377 15484
rect 6227 15453 6239 15456
rect 6181 15447 6239 15453
rect 6365 15453 6377 15456
rect 6411 15453 6423 15487
rect 6472 15484 6500 15512
rect 6876 15493 6904 15524
rect 6692 15487 6750 15493
rect 6692 15484 6704 15487
rect 6472 15456 6704 15484
rect 6365 15447 6423 15453
rect 6692 15453 6704 15456
rect 6738 15453 6750 15487
rect 6692 15447 6750 15453
rect 6871 15487 6929 15493
rect 6871 15453 6883 15487
rect 6917 15453 6929 15487
rect 6871 15447 6929 15453
rect 7006 15444 7012 15496
rect 7064 15484 7070 15496
rect 7101 15487 7159 15493
rect 7101 15484 7113 15487
rect 7064 15456 7113 15484
rect 7064 15444 7070 15456
rect 7101 15453 7113 15456
rect 7147 15453 7159 15487
rect 7101 15447 7159 15453
rect 3844 15320 5948 15348
rect 3844 15308 3850 15320
rect 6270 15308 6276 15360
rect 6328 15348 6334 15360
rect 8205 15351 8263 15357
rect 8205 15348 8217 15351
rect 6328 15320 8217 15348
rect 6328 15308 6334 15320
rect 8205 15317 8217 15320
rect 8251 15317 8263 15351
rect 8312 15348 8340 15524
rect 8570 15512 8576 15564
rect 8628 15512 8634 15564
rect 10778 15552 10784 15564
rect 9232 15524 10784 15552
rect 9069 15505 9127 15511
rect 8938 15493 8944 15496
rect 8900 15487 8944 15493
rect 8900 15453 8912 15487
rect 8900 15447 8944 15453
rect 8938 15444 8944 15447
rect 8996 15444 9002 15496
rect 9069 15471 9081 15505
rect 9115 15484 9127 15505
rect 9232 15484 9260 15524
rect 10778 15512 10784 15524
rect 10836 15512 10842 15564
rect 9115 15471 9260 15484
rect 9069 15465 9260 15471
rect 9084 15456 9260 15465
rect 9306 15444 9312 15496
rect 9364 15444 9370 15496
rect 10888 15484 10916 15660
rect 13078 15648 13084 15660
rect 13136 15648 13142 15700
rect 14283 15691 14341 15697
rect 14283 15657 14295 15691
rect 14329 15688 14341 15691
rect 14458 15688 14464 15700
rect 14329 15660 14464 15688
rect 14329 15657 14341 15660
rect 14283 15651 14341 15657
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 14642 15648 14648 15700
rect 14700 15688 14706 15700
rect 17218 15688 17224 15700
rect 14700 15660 16252 15688
rect 14700 15648 14706 15660
rect 11054 15580 11060 15632
rect 11112 15580 11118 15632
rect 11330 15580 11336 15632
rect 11388 15620 11394 15632
rect 11425 15623 11483 15629
rect 11425 15620 11437 15623
rect 11388 15592 11437 15620
rect 11388 15580 11394 15592
rect 11425 15589 11437 15592
rect 11471 15589 11483 15623
rect 11425 15583 11483 15589
rect 11440 15552 11468 15583
rect 11698 15580 11704 15632
rect 11756 15580 11762 15632
rect 16224 15629 16252 15660
rect 16592 15660 17224 15688
rect 16209 15623 16267 15629
rect 16209 15589 16221 15623
rect 16255 15589 16267 15623
rect 16209 15583 16267 15589
rect 16390 15580 16396 15632
rect 16448 15620 16454 15632
rect 16592 15629 16620 15660
rect 17218 15648 17224 15660
rect 17276 15648 17282 15700
rect 17770 15648 17776 15700
rect 17828 15688 17834 15700
rect 18969 15691 19027 15697
rect 18969 15688 18981 15691
rect 17828 15660 18981 15688
rect 17828 15648 17834 15660
rect 18969 15657 18981 15660
rect 19015 15657 19027 15691
rect 18969 15651 19027 15657
rect 19352 15660 21404 15688
rect 16577 15623 16635 15629
rect 16577 15620 16589 15623
rect 16448 15592 16589 15620
rect 16448 15580 16454 15592
rect 16577 15589 16589 15592
rect 16623 15589 16635 15623
rect 16577 15583 16635 15589
rect 11609 15555 11667 15561
rect 11609 15552 11621 15555
rect 11440 15524 11621 15552
rect 11609 15521 11621 15524
rect 11655 15521 11667 15555
rect 11716 15552 11744 15580
rect 11936 15555 11994 15561
rect 11936 15552 11948 15555
rect 11716 15524 11948 15552
rect 11609 15515 11667 15521
rect 11936 15521 11948 15524
rect 11982 15521 11994 15555
rect 13817 15555 13875 15561
rect 11936 15515 11994 15521
rect 12268 15524 13768 15552
rect 10336 15456 10916 15484
rect 12115 15487 12173 15493
rect 10336 15348 10364 15456
rect 12115 15453 12127 15487
rect 12161 15484 12173 15487
rect 12268 15484 12296 15524
rect 12161 15456 12296 15484
rect 12345 15487 12403 15493
rect 12161 15453 12173 15456
rect 12115 15447 12173 15453
rect 12345 15453 12357 15487
rect 12391 15484 12403 15487
rect 12526 15484 12532 15496
rect 12391 15456 12532 15484
rect 12391 15453 12403 15456
rect 12345 15447 12403 15453
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 10594 15376 10600 15428
rect 10652 15416 10658 15428
rect 11514 15416 11520 15428
rect 10652 15388 11520 15416
rect 10652 15376 10658 15388
rect 11514 15376 11520 15388
rect 11572 15376 11578 15428
rect 8312 15320 10364 15348
rect 8205 15311 8263 15317
rect 10410 15308 10416 15360
rect 10468 15308 10474 15360
rect 11054 15308 11060 15360
rect 11112 15348 11118 15360
rect 13449 15351 13507 15357
rect 13449 15348 13461 15351
rect 11112 15320 13461 15348
rect 11112 15308 11118 15320
rect 13449 15317 13461 15320
rect 13495 15317 13507 15351
rect 13740 15348 13768 15524
rect 13817 15521 13829 15555
rect 13863 15552 13875 15555
rect 14182 15552 14188 15564
rect 13863 15524 14188 15552
rect 13863 15521 13875 15524
rect 13817 15515 13875 15521
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 14550 15512 14556 15564
rect 14608 15512 14614 15564
rect 15930 15512 15936 15564
rect 15988 15512 15994 15564
rect 17037 15555 17095 15561
rect 17037 15521 17049 15555
rect 17083 15521 17095 15555
rect 17037 15515 17095 15521
rect 17129 15556 17187 15561
rect 17236 15556 17264 15648
rect 17129 15555 17264 15556
rect 17129 15521 17141 15555
rect 17175 15528 17264 15555
rect 17175 15521 17187 15528
rect 17129 15515 17187 15521
rect 14323 15487 14381 15493
rect 14323 15453 14335 15487
rect 14369 15484 14381 15487
rect 17052 15484 17080 15515
rect 18138 15512 18144 15564
rect 18196 15552 18202 15564
rect 19352 15552 19380 15660
rect 21376 15564 21404 15660
rect 21818 15648 21824 15700
rect 21876 15688 21882 15700
rect 23109 15691 23167 15697
rect 23109 15688 23121 15691
rect 21876 15660 23121 15688
rect 21876 15648 21882 15660
rect 23109 15657 23121 15660
rect 23155 15657 23167 15691
rect 23109 15651 23167 15657
rect 23943 15691 24001 15697
rect 23943 15657 23955 15691
rect 23989 15688 24001 15691
rect 24210 15688 24216 15700
rect 23989 15660 24216 15688
rect 23989 15657 24001 15660
rect 23943 15651 24001 15657
rect 24210 15648 24216 15660
rect 24268 15648 24274 15700
rect 27430 15648 27436 15700
rect 27488 15688 27494 15700
rect 28261 15691 28319 15697
rect 28261 15688 28273 15691
rect 27488 15660 28273 15688
rect 27488 15648 27494 15660
rect 28261 15657 28273 15660
rect 28307 15657 28319 15691
rect 28261 15651 28319 15657
rect 29270 15648 29276 15700
rect 29328 15688 29334 15700
rect 30377 15691 30435 15697
rect 30377 15688 30389 15691
rect 29328 15660 30389 15688
rect 29328 15648 29334 15660
rect 30377 15657 30389 15660
rect 30423 15657 30435 15691
rect 30377 15651 30435 15657
rect 25869 15623 25927 15629
rect 25869 15589 25881 15623
rect 25915 15620 25927 15623
rect 25958 15620 25964 15632
rect 25915 15592 25964 15620
rect 25915 15589 25927 15592
rect 25869 15583 25927 15589
rect 25958 15580 25964 15592
rect 26016 15580 26022 15632
rect 26510 15580 26516 15632
rect 26568 15580 26574 15632
rect 18196 15524 19380 15552
rect 18196 15512 18202 15524
rect 19426 15512 19432 15564
rect 19484 15512 19490 15564
rect 21266 15512 21272 15564
rect 21324 15512 21330 15564
rect 21358 15512 21364 15564
rect 21416 15512 21422 15564
rect 22005 15555 22063 15561
rect 22005 15552 22017 15555
rect 21468 15524 22017 15552
rect 17310 15484 17316 15496
rect 14369 15456 16988 15484
rect 17052 15456 17316 15484
rect 14369 15453 14381 15456
rect 14323 15447 14381 15453
rect 16850 15376 16856 15428
rect 16908 15376 16914 15428
rect 16022 15348 16028 15360
rect 13740 15320 16028 15348
rect 13449 15311 13507 15317
rect 16022 15308 16028 15320
rect 16080 15308 16086 15360
rect 16960 15348 16988 15456
rect 17310 15444 17316 15456
rect 17368 15444 17374 15496
rect 17494 15493 17500 15496
rect 17456 15487 17500 15493
rect 17456 15453 17468 15487
rect 17456 15447 17500 15453
rect 17494 15444 17500 15447
rect 17552 15444 17558 15496
rect 17678 15493 17684 15496
rect 17635 15487 17684 15493
rect 17635 15453 17647 15487
rect 17681 15453 17684 15487
rect 17635 15447 17684 15453
rect 17678 15444 17684 15447
rect 17736 15444 17742 15496
rect 17862 15444 17868 15496
rect 17920 15444 17926 15496
rect 19058 15444 19064 15496
rect 19116 15484 19122 15496
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 19116 15456 19717 15484
rect 19116 15444 19122 15456
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 20162 15444 20168 15496
rect 20220 15484 20226 15496
rect 21468 15484 21496 15524
rect 22005 15521 22017 15524
rect 22051 15521 22063 15555
rect 26528 15552 26556 15580
rect 26748 15555 26806 15561
rect 26748 15552 26760 15555
rect 22005 15515 22063 15521
rect 23032 15524 25360 15552
rect 26528 15524 26760 15552
rect 21634 15493 21640 15496
rect 20220 15456 21496 15484
rect 21596 15487 21640 15493
rect 20220 15444 20226 15456
rect 21596 15453 21608 15487
rect 21596 15447 21640 15453
rect 21634 15444 21640 15447
rect 21692 15444 21698 15496
rect 21775 15487 21833 15493
rect 21775 15453 21787 15487
rect 21821 15484 21833 15487
rect 23032 15484 23060 15524
rect 25332 15496 25360 15524
rect 26748 15521 26760 15524
rect 26794 15521 26806 15555
rect 27430 15552 27436 15564
rect 26748 15515 26806 15521
rect 27086 15524 27436 15552
rect 21821 15456 23060 15484
rect 23477 15487 23535 15493
rect 21821 15453 21833 15456
rect 21775 15447 21833 15453
rect 23477 15453 23489 15487
rect 23523 15484 23535 15487
rect 23750 15484 23756 15496
rect 23523 15456 23756 15484
rect 23523 15453 23535 15456
rect 23477 15447 23535 15453
rect 23750 15444 23756 15456
rect 23808 15444 23814 15496
rect 23940 15489 23998 15495
rect 23940 15455 23952 15489
rect 23986 15484 23998 15489
rect 24026 15484 24032 15496
rect 23986 15456 24032 15484
rect 23986 15455 23998 15456
rect 23940 15449 23998 15455
rect 24026 15444 24032 15456
rect 24084 15444 24090 15496
rect 24213 15487 24271 15493
rect 24213 15453 24225 15487
rect 24259 15484 24271 15487
rect 24302 15484 24308 15496
rect 24259 15456 24308 15484
rect 24259 15453 24271 15456
rect 24213 15447 24271 15453
rect 24302 15444 24308 15456
rect 24360 15444 24366 15496
rect 25314 15444 25320 15496
rect 25372 15444 25378 15496
rect 25958 15444 25964 15496
rect 26016 15484 26022 15496
rect 26142 15484 26148 15496
rect 26016 15456 26148 15484
rect 26016 15444 26022 15456
rect 26142 15444 26148 15456
rect 26200 15484 26206 15496
rect 26421 15487 26479 15493
rect 26421 15484 26433 15487
rect 26200 15456 26433 15484
rect 26200 15444 26206 15456
rect 26421 15453 26433 15456
rect 26467 15453 26479 15487
rect 26421 15447 26479 15453
rect 26927 15487 26985 15493
rect 26927 15453 26939 15487
rect 26973 15484 26985 15487
rect 27086 15484 27114 15524
rect 27430 15512 27436 15524
rect 27488 15512 27494 15564
rect 27982 15512 27988 15564
rect 28040 15552 28046 15564
rect 28905 15555 28963 15561
rect 28905 15552 28917 15555
rect 28040 15524 28917 15552
rect 28040 15512 28046 15524
rect 28905 15521 28917 15524
rect 28951 15521 28963 15555
rect 28905 15515 28963 15521
rect 29638 15512 29644 15564
rect 29696 15552 29702 15564
rect 30561 15555 30619 15561
rect 30561 15552 30573 15555
rect 29696 15524 30573 15552
rect 29696 15512 29702 15524
rect 30561 15521 30573 15524
rect 30607 15521 30619 15555
rect 30561 15515 30619 15521
rect 26973 15456 27114 15484
rect 27157 15487 27215 15493
rect 26973 15453 26985 15456
rect 26927 15447 26985 15453
rect 27157 15453 27169 15487
rect 27203 15484 27215 15487
rect 28534 15484 28540 15496
rect 27203 15456 28540 15484
rect 27203 15453 27215 15456
rect 27157 15447 27215 15453
rect 18874 15376 18880 15428
rect 18932 15376 18938 15428
rect 25498 15416 25504 15428
rect 24872 15388 25504 15416
rect 18892 15348 18920 15376
rect 16960 15320 18920 15348
rect 18966 15308 18972 15360
rect 19024 15348 19030 15360
rect 20714 15348 20720 15360
rect 19024 15320 20720 15348
rect 19024 15308 19030 15320
rect 20714 15308 20720 15320
rect 20772 15308 20778 15360
rect 20993 15351 21051 15357
rect 20993 15317 21005 15351
rect 21039 15348 21051 15351
rect 22186 15348 22192 15360
rect 21039 15320 22192 15348
rect 21039 15317 21051 15320
rect 20993 15311 21051 15317
rect 22186 15308 22192 15320
rect 22244 15308 22250 15360
rect 22370 15308 22376 15360
rect 22428 15348 22434 15360
rect 23842 15348 23848 15360
rect 22428 15320 23848 15348
rect 22428 15308 22434 15320
rect 23842 15308 23848 15320
rect 23900 15308 23906 15360
rect 24026 15308 24032 15360
rect 24084 15348 24090 15360
rect 24872 15348 24900 15388
rect 25498 15376 25504 15388
rect 25556 15376 25562 15428
rect 24084 15320 24900 15348
rect 24084 15308 24090 15320
rect 25314 15308 25320 15360
rect 25372 15308 25378 15360
rect 26142 15308 26148 15360
rect 26200 15308 26206 15360
rect 26436 15348 26464 15447
rect 28534 15444 28540 15456
rect 28592 15444 28598 15496
rect 28629 15487 28687 15493
rect 28629 15453 28641 15487
rect 28675 15453 28687 15487
rect 28629 15447 28687 15453
rect 27982 15376 27988 15428
rect 28040 15416 28046 15428
rect 28644 15416 28672 15447
rect 28040 15388 28672 15416
rect 28040 15376 28046 15388
rect 26694 15348 26700 15360
rect 26436 15320 26700 15348
rect 26694 15308 26700 15320
rect 26752 15308 26758 15360
rect 29270 15308 29276 15360
rect 29328 15348 29334 15360
rect 30009 15351 30067 15357
rect 30009 15348 30021 15351
rect 29328 15320 30021 15348
rect 29328 15308 29334 15320
rect 30009 15317 30021 15320
rect 30055 15317 30067 15351
rect 30009 15311 30067 15317
rect 552 15258 30912 15280
rect 552 15206 4193 15258
rect 4245 15206 4257 15258
rect 4309 15206 4321 15258
rect 4373 15206 4385 15258
rect 4437 15206 4449 15258
rect 4501 15206 11783 15258
rect 11835 15206 11847 15258
rect 11899 15206 11911 15258
rect 11963 15206 11975 15258
rect 12027 15206 12039 15258
rect 12091 15206 19373 15258
rect 19425 15206 19437 15258
rect 19489 15206 19501 15258
rect 19553 15206 19565 15258
rect 19617 15206 19629 15258
rect 19681 15206 26963 15258
rect 27015 15206 27027 15258
rect 27079 15206 27091 15258
rect 27143 15206 27155 15258
rect 27207 15206 27219 15258
rect 27271 15206 30912 15258
rect 552 15184 30912 15206
rect 2774 15104 2780 15156
rect 2832 15104 2838 15156
rect 4982 15144 4988 15156
rect 3160 15116 4988 15144
rect 937 15011 995 15017
rect 937 14977 949 15011
rect 983 15008 995 15011
rect 1118 15008 1124 15020
rect 983 14980 1124 15008
rect 983 14977 995 14980
rect 937 14971 995 14977
rect 1118 14968 1124 14980
rect 1176 14968 1182 15020
rect 1443 15011 1501 15017
rect 1443 14977 1455 15011
rect 1489 15008 1501 15011
rect 2958 15008 2964 15020
rect 1489 14980 2964 15008
rect 1489 14977 1501 14980
rect 1443 14971 1501 14977
rect 2958 14968 2964 14980
rect 3016 14968 3022 15020
rect 1673 14943 1731 14949
rect 1673 14909 1685 14943
rect 1719 14940 1731 14943
rect 3160 14940 3188 15116
rect 4982 15104 4988 15116
rect 5040 15104 5046 15156
rect 5813 15147 5871 15153
rect 5813 15113 5825 15147
rect 5859 15144 5871 15147
rect 6362 15144 6368 15156
rect 5859 15116 6368 15144
rect 5859 15113 5871 15116
rect 5813 15107 5871 15113
rect 6362 15104 6368 15116
rect 6420 15104 6426 15156
rect 6454 15104 6460 15156
rect 6512 15144 6518 15156
rect 6512 15116 7972 15144
rect 6512 15104 6518 15116
rect 4295 15011 4353 15017
rect 4295 14977 4307 15011
rect 4341 15008 4353 15011
rect 6270 15008 6276 15020
rect 4341 14980 6276 15008
rect 4341 14977 4353 14980
rect 4295 14971 4353 14977
rect 6270 14968 6276 14980
rect 6328 14968 6334 15020
rect 6546 14968 6552 15020
rect 6604 15017 6610 15020
rect 6604 15011 6653 15017
rect 6604 14977 6607 15011
rect 6641 14977 6653 15011
rect 7006 15008 7012 15020
rect 6604 14971 6653 14977
rect 6748 14980 7012 15008
rect 6604 14968 6610 14971
rect 1719 14912 3188 14940
rect 1719 14909 1731 14912
rect 1673 14903 1731 14909
rect 3234 14900 3240 14952
rect 3292 14900 3298 14952
rect 3786 14900 3792 14952
rect 3844 14900 3850 14952
rect 3878 14900 3884 14952
rect 3936 14900 3942 14952
rect 4522 14900 4528 14952
rect 4580 14900 4586 14952
rect 6086 14900 6092 14952
rect 6144 14900 6150 14952
rect 6748 14940 6776 14980
rect 7006 14968 7012 14980
rect 7064 14968 7070 15020
rect 7944 15008 7972 15116
rect 9490 15104 9496 15156
rect 9548 15144 9554 15156
rect 10318 15144 10324 15156
rect 9548 15116 10324 15144
rect 9548 15104 9554 15116
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 10965 15147 11023 15153
rect 10965 15113 10977 15147
rect 11011 15144 11023 15147
rect 12894 15144 12900 15156
rect 11011 15116 12900 15144
rect 11011 15113 11023 15116
rect 10965 15107 11023 15113
rect 12894 15104 12900 15116
rect 12952 15104 12958 15156
rect 13909 15147 13967 15153
rect 13909 15113 13921 15147
rect 13955 15144 13967 15147
rect 14182 15144 14188 15156
rect 13955 15116 14188 15144
rect 13955 15113 13967 15116
rect 13909 15107 13967 15113
rect 14182 15104 14188 15116
rect 14240 15104 14246 15156
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 15344 15116 15608 15144
rect 15344 15104 15350 15116
rect 10336 15076 10364 15104
rect 10336 15048 11192 15076
rect 8938 15017 8944 15020
rect 8900 15011 8944 15017
rect 8900 15008 8912 15011
rect 7944 14980 8912 15008
rect 8900 14977 8912 14980
rect 8900 14971 8944 14977
rect 8938 14968 8944 14971
rect 8996 14968 9002 15020
rect 9079 15011 9137 15017
rect 9079 14977 9091 15011
rect 9125 15008 9137 15011
rect 10686 15008 10692 15020
rect 9125 14980 10692 15008
rect 9125 14977 9137 14980
rect 9079 14971 9137 14977
rect 10686 14968 10692 14980
rect 10744 14968 10750 15020
rect 6196 14912 6776 14940
rect 6825 14943 6883 14949
rect 3513 14875 3571 14881
rect 3513 14841 3525 14875
rect 3559 14872 3571 14875
rect 3896 14872 3924 14900
rect 3559 14844 3924 14872
rect 3559 14841 3571 14844
rect 3513 14835 3571 14841
rect 1394 14764 1400 14816
rect 1452 14813 1458 14816
rect 1452 14804 1461 14813
rect 3528 14804 3556 14835
rect 1452 14776 3556 14804
rect 3896 14804 3924 14844
rect 5902 14832 5908 14884
rect 5960 14872 5966 14884
rect 6196 14872 6224 14912
rect 6825 14909 6837 14943
rect 6871 14940 6883 14943
rect 6914 14940 6920 14952
rect 6871 14912 6920 14940
rect 6871 14909 6883 14912
rect 6825 14903 6883 14909
rect 6914 14900 6920 14912
rect 6972 14900 6978 14952
rect 7282 14900 7288 14952
rect 7340 14940 7346 14952
rect 7340 14912 8294 14940
rect 7340 14900 7346 14912
rect 5960 14844 6224 14872
rect 5960 14832 5966 14844
rect 4255 14807 4313 14813
rect 4255 14804 4267 14807
rect 3896 14776 4267 14804
rect 1452 14767 1461 14776
rect 4255 14773 4267 14776
rect 4301 14773 4313 14807
rect 4255 14767 4313 14773
rect 1452 14764 1458 14767
rect 6454 14764 6460 14816
rect 6512 14804 6518 14816
rect 6555 14807 6613 14813
rect 6555 14804 6567 14807
rect 6512 14776 6567 14804
rect 6512 14764 6518 14776
rect 6555 14773 6567 14776
rect 6601 14773 6613 14807
rect 6555 14767 6613 14773
rect 6730 14764 6736 14816
rect 6788 14804 6794 14816
rect 7929 14807 7987 14813
rect 7929 14804 7941 14807
rect 6788 14776 7941 14804
rect 6788 14764 6794 14776
rect 7929 14773 7941 14776
rect 7975 14773 7987 14807
rect 8266 14804 8294 14912
rect 8570 14900 8576 14952
rect 8628 14900 8634 14952
rect 9309 14943 9367 14949
rect 9309 14909 9321 14943
rect 9355 14940 9367 14943
rect 9674 14940 9680 14952
rect 9355 14912 9680 14940
rect 9355 14909 9367 14912
rect 9309 14903 9367 14909
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 11164 14949 11192 15048
rect 11238 15036 11244 15088
rect 11296 15036 11302 15088
rect 13078 15036 13084 15088
rect 13136 15036 13142 15088
rect 15580 15076 15608 15116
rect 16022 15104 16028 15156
rect 16080 15104 16086 15156
rect 18233 15147 18291 15153
rect 18233 15144 18245 15147
rect 16132 15116 18245 15144
rect 16132 15076 16160 15116
rect 18233 15113 18245 15116
rect 18279 15113 18291 15147
rect 18233 15107 18291 15113
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 21637 15147 21695 15153
rect 21637 15144 21649 15147
rect 20772 15116 21649 15144
rect 20772 15104 20778 15116
rect 21637 15113 21649 15116
rect 21683 15113 21695 15147
rect 21637 15107 21695 15113
rect 21744 15116 23336 15144
rect 19150 15076 19156 15088
rect 15580 15048 16160 15076
rect 18716 15048 19156 15076
rect 11256 15008 11284 15036
rect 11606 15008 11612 15020
rect 11256 14980 11612 15008
rect 11606 14968 11612 14980
rect 11664 14968 11670 15020
rect 11747 15011 11805 15017
rect 11747 14977 11759 15011
rect 11793 15008 11805 15011
rect 14691 15011 14749 15017
rect 11793 14980 14320 15008
rect 11793 14977 11805 14980
rect 11747 14971 11805 14977
rect 11149 14943 11207 14949
rect 11149 14909 11161 14943
rect 11195 14909 11207 14943
rect 11149 14903 11207 14909
rect 11241 14943 11299 14949
rect 11241 14909 11253 14943
rect 11287 14940 11299 14943
rect 11330 14940 11336 14952
rect 11287 14912 11336 14940
rect 11287 14909 11299 14912
rect 11241 14903 11299 14909
rect 10336 14844 10916 14872
rect 10336 14804 10364 14844
rect 10888 14816 10916 14844
rect 8266 14776 10364 14804
rect 7929 14767 7987 14773
rect 10410 14764 10416 14816
rect 10468 14764 10474 14816
rect 10870 14764 10876 14816
rect 10928 14764 10934 14816
rect 11164 14804 11192 14903
rect 11330 14900 11336 14912
rect 11388 14940 11394 14952
rect 11882 14940 11888 14952
rect 11388 14912 11888 14940
rect 11388 14900 11394 14912
rect 11882 14900 11888 14912
rect 11940 14900 11946 14952
rect 11974 14900 11980 14952
rect 12032 14900 12038 14952
rect 14182 14900 14188 14952
rect 14240 14900 14246 14952
rect 13633 14875 13691 14881
rect 13633 14872 13645 14875
rect 13004 14844 13645 14872
rect 11606 14804 11612 14816
rect 11164 14776 11612 14804
rect 11606 14764 11612 14776
rect 11664 14764 11670 14816
rect 11698 14764 11704 14816
rect 11756 14813 11762 14816
rect 11756 14804 11765 14813
rect 11756 14776 11801 14804
rect 11756 14767 11765 14776
rect 11756 14764 11762 14767
rect 11882 14764 11888 14816
rect 11940 14804 11946 14816
rect 13004 14804 13032 14844
rect 13633 14841 13645 14844
rect 13679 14841 13691 14875
rect 13633 14835 13691 14841
rect 14292 14816 14320 14980
rect 14691 14977 14703 15011
rect 14737 15008 14749 15011
rect 14737 14980 15608 15008
rect 14737 14977 14749 14980
rect 14691 14971 14749 14977
rect 14921 14943 14979 14949
rect 14921 14909 14933 14943
rect 14967 14940 14979 14943
rect 15194 14940 15200 14952
rect 14967 14912 15200 14940
rect 14967 14909 14979 14912
rect 14921 14903 14979 14909
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 11940 14776 13032 14804
rect 11940 14764 11946 14776
rect 14274 14764 14280 14816
rect 14332 14764 14338 14816
rect 14458 14764 14464 14816
rect 14516 14804 14522 14816
rect 14651 14807 14709 14813
rect 14651 14804 14663 14807
rect 14516 14776 14663 14804
rect 14516 14764 14522 14776
rect 14651 14773 14663 14776
rect 14697 14773 14709 14807
rect 15580 14804 15608 14980
rect 16390 14968 16396 15020
rect 16448 14968 16454 15020
rect 16899 15011 16957 15017
rect 16899 14977 16911 15011
rect 16945 15008 16957 15011
rect 18716 15008 18744 15048
rect 19150 15036 19156 15048
rect 19208 15036 19214 15088
rect 21358 15036 21364 15088
rect 21416 15076 21422 15088
rect 21744 15076 21772 15116
rect 21416 15048 21772 15076
rect 21416 15036 21422 15048
rect 16945 14980 18744 15008
rect 16945 14977 16957 14980
rect 16899 14971 16957 14977
rect 18782 14968 18788 15020
rect 18840 15008 18846 15020
rect 22281 15011 22339 15017
rect 18840 14980 19380 15008
rect 18840 14968 18846 14980
rect 17129 14943 17187 14949
rect 17129 14909 17141 14943
rect 17175 14940 17187 14943
rect 17954 14940 17960 14952
rect 17175 14912 17960 14940
rect 17175 14909 17187 14912
rect 17129 14903 17187 14909
rect 17954 14900 17960 14912
rect 18012 14900 18018 14952
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14940 18751 14943
rect 19242 14940 19248 14952
rect 18739 14912 19248 14940
rect 18739 14909 18751 14912
rect 18693 14903 18751 14909
rect 19242 14900 19248 14912
rect 19300 14900 19306 14952
rect 19352 14949 19380 14980
rect 20272 14993 21772 15008
rect 20272 14962 20305 14993
rect 20293 14959 20305 14962
rect 20339 14980 21772 14993
rect 20339 14959 20351 14980
rect 20293 14953 20351 14959
rect 19337 14943 19395 14949
rect 19337 14909 19349 14943
rect 19383 14909 19395 14943
rect 19337 14903 19395 14909
rect 19705 14943 19763 14949
rect 19705 14909 19717 14943
rect 19751 14940 19763 14943
rect 19794 14940 19800 14952
rect 19751 14912 19800 14940
rect 19751 14909 19763 14912
rect 19705 14903 19763 14909
rect 19794 14900 19800 14912
rect 19852 14900 19858 14952
rect 20533 14943 20591 14949
rect 20533 14909 20545 14943
rect 20579 14940 20591 14943
rect 20622 14940 20628 14952
rect 20579 14912 20628 14940
rect 20579 14909 20591 14912
rect 20533 14903 20591 14909
rect 20622 14900 20628 14912
rect 20680 14900 20686 14952
rect 18969 14875 19027 14881
rect 18969 14841 18981 14875
rect 19015 14841 19027 14875
rect 18969 14835 19027 14841
rect 16390 14804 16396 14816
rect 15580 14776 16396 14804
rect 14651 14767 14709 14773
rect 16390 14764 16396 14776
rect 16448 14764 16454 14816
rect 16758 14764 16764 14816
rect 16816 14804 16822 14816
rect 16859 14807 16917 14813
rect 16859 14804 16871 14807
rect 16816 14776 16871 14804
rect 16816 14764 16822 14776
rect 16859 14773 16871 14776
rect 16905 14804 16917 14807
rect 17494 14804 17500 14816
rect 16905 14776 17500 14804
rect 16905 14773 16917 14776
rect 16859 14767 16917 14773
rect 17494 14764 17500 14776
rect 17552 14804 17558 14816
rect 18984 14804 19012 14835
rect 17552 14776 19012 14804
rect 17552 14764 17558 14776
rect 20254 14764 20260 14816
rect 20312 14813 20318 14816
rect 20312 14804 20321 14813
rect 21174 14804 21180 14816
rect 20312 14776 21180 14804
rect 20312 14767 20321 14776
rect 20312 14764 20318 14767
rect 21174 14764 21180 14776
rect 21232 14764 21238 14816
rect 21744 14804 21772 14980
rect 22281 14977 22293 15011
rect 22327 15008 22339 15011
rect 22922 15008 22928 15020
rect 22327 14980 22928 15008
rect 22327 14977 22339 14980
rect 22281 14971 22339 14977
rect 22922 14968 22928 14980
rect 22980 14968 22986 15020
rect 23308 15008 23336 15116
rect 23474 15104 23480 15156
rect 23532 15144 23538 15156
rect 27890 15144 27896 15156
rect 23532 15116 25360 15144
rect 23532 15104 23538 15116
rect 25332 15088 25360 15116
rect 26068 15116 27896 15144
rect 23569 15079 23627 15085
rect 23569 15045 23581 15079
rect 23615 15076 23627 15079
rect 23658 15076 23664 15088
rect 23615 15048 23664 15076
rect 23615 15045 23627 15048
rect 23569 15039 23627 15045
rect 23658 15036 23664 15048
rect 23716 15036 23722 15088
rect 25314 15036 25320 15088
rect 25372 15036 25378 15088
rect 23308 14980 23704 15008
rect 22005 14943 22063 14949
rect 22005 14909 22017 14943
rect 22051 14940 22063 14943
rect 23566 14940 23572 14952
rect 22051 14912 23572 14940
rect 22051 14909 22063 14912
rect 22005 14903 22063 14909
rect 23566 14900 23572 14912
rect 23624 14900 23630 14952
rect 23676 14940 23704 14980
rect 23750 14968 23756 15020
rect 23808 15008 23814 15020
rect 24210 15017 24216 15020
rect 23845 15011 23903 15017
rect 23845 15008 23857 15011
rect 23808 14980 23857 15008
rect 23808 14968 23814 14980
rect 23845 14977 23857 14980
rect 23891 14977 23903 15011
rect 23845 14971 23903 14977
rect 24172 15011 24216 15017
rect 24172 14977 24184 15011
rect 24172 14971 24216 14977
rect 24210 14968 24216 14971
rect 24268 14968 24274 15020
rect 24351 15011 24409 15017
rect 24351 14977 24363 15011
rect 24397 15008 24409 15011
rect 26068 15008 26096 15116
rect 27890 15104 27896 15116
rect 27948 15104 27954 15156
rect 28166 15104 28172 15156
rect 28224 15144 28230 15156
rect 28445 15147 28503 15153
rect 28445 15144 28457 15147
rect 28224 15116 28457 15144
rect 28224 15104 28230 15116
rect 28445 15113 28457 15116
rect 28491 15113 28503 15147
rect 28445 15107 28503 15113
rect 28534 15104 28540 15156
rect 28592 15144 28598 15156
rect 30101 15147 30159 15153
rect 30101 15144 30113 15147
rect 28592 15116 30113 15144
rect 28592 15104 28598 15116
rect 30101 15113 30113 15116
rect 30147 15113 30159 15147
rect 30101 15107 30159 15113
rect 30374 15104 30380 15156
rect 30432 15104 30438 15156
rect 27522 15036 27528 15088
rect 27580 15076 27586 15088
rect 28077 15079 28135 15085
rect 28077 15076 28089 15079
rect 27580 15048 28089 15076
rect 27580 15036 27586 15048
rect 28077 15045 28089 15048
rect 28123 15045 28135 15079
rect 28077 15039 28135 15045
rect 24397 14980 26096 15008
rect 26160 14999 26559 15008
rect 26160 14993 26574 14999
rect 26160 14980 26528 14993
rect 24397 14977 24409 14980
rect 24351 14971 24409 14977
rect 24581 14943 24639 14949
rect 23676 14936 24532 14940
rect 24581 14936 24593 14943
rect 23676 14912 24593 14936
rect 24504 14909 24593 14912
rect 24627 14909 24639 14943
rect 24504 14908 24639 14909
rect 24581 14903 24639 14908
rect 25958 14900 25964 14952
rect 26016 14940 26022 14952
rect 26053 14943 26111 14949
rect 26053 14940 26065 14943
rect 26016 14912 26065 14940
rect 26016 14900 26022 14912
rect 26053 14909 26065 14912
rect 26099 14909 26111 14943
rect 26053 14903 26111 14909
rect 26160 14816 26188 14980
rect 26516 14959 26528 14980
rect 26562 14959 26574 14993
rect 26602 14968 26608 15020
rect 26660 15008 26666 15020
rect 28184 15008 28212 15104
rect 28902 15036 28908 15088
rect 28960 15076 28966 15088
rect 28960 15048 30604 15076
rect 28960 15036 28966 15048
rect 26660 14980 28212 15008
rect 26660 14968 26666 14980
rect 29638 14968 29644 15020
rect 29696 14968 29702 15020
rect 26516 14953 26574 14959
rect 26789 14943 26847 14949
rect 26789 14909 26801 14943
rect 26835 14940 26847 14943
rect 29362 14940 29368 14952
rect 26835 14912 29368 14940
rect 26835 14909 26847 14912
rect 26789 14903 26847 14909
rect 29362 14900 29368 14912
rect 29420 14900 29426 14952
rect 29457 14943 29515 14949
rect 29457 14909 29469 14943
rect 29503 14940 29515 14943
rect 29656 14940 29684 14968
rect 29503 14912 29684 14940
rect 29503 14909 29515 14912
rect 29457 14903 29515 14909
rect 29730 14900 29736 14952
rect 29788 14900 29794 14952
rect 30006 14900 30012 14952
rect 30064 14940 30070 14952
rect 30576 14949 30604 15048
rect 30285 14943 30343 14949
rect 30285 14940 30297 14943
rect 30064 14912 30297 14940
rect 30064 14900 30070 14912
rect 30285 14909 30297 14912
rect 30331 14909 30343 14943
rect 30285 14903 30343 14909
rect 30561 14943 30619 14949
rect 30561 14909 30573 14943
rect 30607 14909 30619 14943
rect 30561 14903 30619 14909
rect 31386 14900 31392 14952
rect 31444 14900 31450 14952
rect 28353 14875 28411 14881
rect 28353 14841 28365 14875
rect 28399 14841 28411 14875
rect 28353 14835 28411 14841
rect 25685 14807 25743 14813
rect 25685 14804 25697 14807
rect 21744 14776 25697 14804
rect 25685 14773 25697 14776
rect 25731 14773 25743 14807
rect 25685 14767 25743 14773
rect 26142 14764 26148 14816
rect 26200 14764 26206 14816
rect 26510 14764 26516 14816
rect 26568 14813 26574 14816
rect 26568 14804 26577 14813
rect 26568 14776 26613 14804
rect 26568 14767 26577 14776
rect 26568 14764 26574 14767
rect 26694 14764 26700 14816
rect 26752 14804 26758 14816
rect 28368 14804 28396 14835
rect 29086 14832 29092 14884
rect 29144 14832 29150 14884
rect 29641 14875 29699 14881
rect 29641 14841 29653 14875
rect 29687 14872 29699 14875
rect 29748 14872 29776 14900
rect 29687 14844 29776 14872
rect 29687 14841 29699 14844
rect 29641 14835 29699 14841
rect 26752 14776 28396 14804
rect 29917 14807 29975 14813
rect 26752 14764 26758 14776
rect 29917 14773 29929 14807
rect 29963 14804 29975 14807
rect 30374 14804 30380 14816
rect 29963 14776 30380 14804
rect 29963 14773 29975 14776
rect 29917 14767 29975 14773
rect 30374 14764 30380 14776
rect 30432 14804 30438 14816
rect 31404 14804 31432 14900
rect 30432 14776 31432 14804
rect 30432 14764 30438 14776
rect 552 14714 31072 14736
rect 552 14662 7988 14714
rect 8040 14662 8052 14714
rect 8104 14662 8116 14714
rect 8168 14662 8180 14714
rect 8232 14662 8244 14714
rect 8296 14662 15578 14714
rect 15630 14662 15642 14714
rect 15694 14662 15706 14714
rect 15758 14662 15770 14714
rect 15822 14662 15834 14714
rect 15886 14662 23168 14714
rect 23220 14662 23232 14714
rect 23284 14662 23296 14714
rect 23348 14662 23360 14714
rect 23412 14662 23424 14714
rect 23476 14662 30758 14714
rect 30810 14662 30822 14714
rect 30874 14662 30886 14714
rect 30938 14662 30950 14714
rect 31002 14662 31014 14714
rect 31066 14662 31072 14714
rect 552 14640 31072 14662
rect 1118 14560 1124 14612
rect 1176 14560 1182 14612
rect 3050 14560 3056 14612
rect 3108 14560 3114 14612
rect 3878 14560 3884 14612
rect 3936 14600 3942 14612
rect 3979 14603 4037 14609
rect 3979 14600 3991 14603
rect 3936 14572 3991 14600
rect 3936 14560 3942 14572
rect 3979 14569 3991 14572
rect 4025 14569 4037 14603
rect 3979 14563 4037 14569
rect 4706 14560 4712 14612
rect 4764 14600 4770 14612
rect 4764 14572 5488 14600
rect 4764 14560 4770 14572
rect 1136 14532 1164 14560
rect 3602 14532 3608 14544
rect 1136 14504 1256 14532
rect 1228 14473 1256 14504
rect 2746 14504 3608 14532
rect 1121 14467 1179 14473
rect 1121 14433 1133 14467
rect 1167 14433 1179 14467
rect 1121 14427 1179 14433
rect 1213 14467 1271 14473
rect 1213 14433 1225 14467
rect 1259 14433 1271 14467
rect 2746 14464 2774 14504
rect 3602 14492 3608 14504
rect 3660 14492 3666 14544
rect 5460 14532 5488 14572
rect 5534 14560 5540 14612
rect 5592 14560 5598 14612
rect 5902 14560 5908 14612
rect 5960 14600 5966 14612
rect 6089 14603 6147 14609
rect 6089 14600 6101 14603
rect 5960 14572 6101 14600
rect 5960 14560 5966 14572
rect 6089 14569 6101 14572
rect 6135 14569 6147 14603
rect 6914 14600 6920 14612
rect 6089 14563 6147 14569
rect 6610 14572 6920 14600
rect 6610 14532 6638 14572
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 7374 14560 7380 14612
rect 7432 14600 7438 14612
rect 7432 14572 9260 14600
rect 7432 14560 7438 14572
rect 5460 14504 6316 14532
rect 6288 14476 6316 14504
rect 6472 14504 6638 14532
rect 1213 14427 1271 14433
rect 1872 14436 2774 14464
rect 3513 14467 3571 14473
rect 1136 14328 1164 14427
rect 1709 14417 1767 14423
rect 1709 14414 1721 14417
rect 1394 14356 1400 14408
rect 1452 14396 1458 14408
rect 1540 14399 1598 14405
rect 1540 14396 1552 14399
rect 1452 14368 1552 14396
rect 1452 14356 1458 14368
rect 1540 14365 1552 14368
rect 1586 14365 1598 14399
rect 1688 14383 1721 14414
rect 1755 14396 1767 14417
rect 1872 14396 1900 14436
rect 3513 14433 3525 14467
rect 3559 14464 3571 14467
rect 3786 14464 3792 14476
rect 3559 14436 3792 14464
rect 3559 14433 3571 14436
rect 3513 14427 3571 14433
rect 3786 14424 3792 14436
rect 3844 14424 3850 14476
rect 5902 14464 5908 14476
rect 3896 14436 5908 14464
rect 1755 14383 1900 14396
rect 1688 14368 1900 14383
rect 1540 14359 1598 14365
rect 1946 14356 1952 14408
rect 2004 14356 2010 14408
rect 3896 14396 3924 14436
rect 5902 14424 5908 14436
rect 5960 14464 5966 14476
rect 5997 14467 6055 14473
rect 5997 14464 6009 14467
rect 5960 14436 6009 14464
rect 5960 14424 5966 14436
rect 5997 14433 6009 14436
rect 6043 14433 6055 14467
rect 5997 14427 6055 14433
rect 6270 14424 6276 14476
rect 6328 14424 6334 14476
rect 2608 14368 3924 14396
rect 4019 14399 4077 14405
rect 1136 14300 1256 14328
rect 934 14220 940 14272
rect 992 14220 998 14272
rect 1228 14260 1256 14300
rect 2608 14260 2636 14368
rect 4019 14365 4031 14399
rect 4065 14396 4077 14399
rect 4154 14396 4160 14408
rect 4065 14368 4160 14396
rect 4065 14365 4077 14368
rect 4019 14359 4077 14365
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14396 4307 14399
rect 4295 14368 6316 14396
rect 4295 14365 4307 14368
rect 4249 14359 4307 14365
rect 1228 14232 2636 14260
rect 3234 14220 3240 14272
rect 3292 14260 3298 14272
rect 5626 14260 5632 14272
rect 3292 14232 5632 14260
rect 3292 14220 3298 14232
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 5810 14220 5816 14272
rect 5868 14220 5874 14272
rect 6288 14260 6316 14368
rect 6365 14331 6423 14337
rect 6365 14297 6377 14331
rect 6411 14328 6423 14331
rect 6472 14328 6500 14504
rect 8938 14492 8944 14544
rect 8996 14532 9002 14544
rect 9125 14535 9183 14541
rect 9125 14532 9137 14535
rect 8996 14504 9137 14532
rect 8996 14492 9002 14504
rect 9125 14501 9137 14504
rect 9171 14501 9183 14535
rect 9232 14532 9260 14572
rect 9306 14560 9312 14612
rect 9364 14600 9370 14612
rect 9401 14603 9459 14609
rect 9401 14600 9413 14603
rect 9364 14572 9413 14600
rect 9364 14560 9370 14572
rect 9401 14569 9413 14572
rect 9447 14569 9459 14603
rect 9401 14563 9459 14569
rect 9674 14560 9680 14612
rect 9732 14560 9738 14612
rect 9950 14560 9956 14612
rect 10008 14560 10014 14612
rect 11057 14603 11115 14609
rect 11057 14569 11069 14603
rect 11103 14600 11115 14603
rect 11238 14600 11244 14612
rect 11103 14572 11244 14600
rect 11103 14569 11115 14572
rect 11057 14563 11115 14569
rect 11238 14560 11244 14572
rect 11296 14560 11302 14612
rect 11333 14603 11391 14609
rect 11333 14569 11345 14603
rect 11379 14600 11391 14603
rect 11974 14600 11980 14612
rect 11379 14572 11980 14600
rect 11379 14569 11391 14572
rect 11333 14563 11391 14569
rect 11974 14560 11980 14572
rect 12032 14560 12038 14612
rect 13446 14560 13452 14612
rect 13504 14560 13510 14612
rect 14283 14603 14341 14609
rect 14283 14569 14295 14603
rect 14329 14600 14341 14603
rect 14458 14600 14464 14612
rect 14329 14572 14464 14600
rect 14329 14569 14341 14572
rect 14283 14563 14341 14569
rect 14458 14560 14464 14572
rect 14516 14560 14522 14612
rect 15657 14603 15715 14609
rect 15657 14569 15669 14603
rect 15703 14569 15715 14603
rect 15657 14563 15715 14569
rect 10505 14535 10563 14541
rect 10505 14532 10517 14535
rect 9232 14504 10517 14532
rect 9125 14495 9183 14501
rect 10505 14501 10517 14504
rect 10551 14501 10563 14535
rect 11422 14532 11428 14544
rect 10505 14495 10563 14501
rect 11256 14504 11428 14532
rect 6546 14424 6552 14476
rect 6604 14424 6610 14476
rect 8754 14424 8760 14476
rect 8812 14464 8818 14476
rect 8849 14467 8907 14473
rect 8849 14464 8861 14467
rect 8812 14436 8861 14464
rect 8812 14424 8818 14436
rect 8849 14433 8861 14436
rect 8895 14433 8907 14467
rect 8849 14427 8907 14433
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 9490 14464 9496 14476
rect 9088 14436 9496 14464
rect 9088 14424 9094 14436
rect 9490 14424 9496 14436
rect 9548 14464 9554 14476
rect 9585 14467 9643 14473
rect 9585 14464 9597 14467
rect 9548 14436 9597 14464
rect 9548 14424 9554 14436
rect 9585 14433 9597 14436
rect 9631 14433 9643 14467
rect 9585 14427 9643 14433
rect 9674 14424 9680 14476
rect 9732 14464 9738 14476
rect 9861 14467 9919 14473
rect 9861 14464 9873 14467
rect 9732 14436 9873 14464
rect 9732 14424 9738 14436
rect 9861 14433 9873 14436
rect 9907 14464 9919 14467
rect 10042 14464 10048 14476
rect 9907 14436 10048 14464
rect 9907 14433 9919 14436
rect 9861 14427 9919 14433
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 10137 14467 10195 14473
rect 10137 14433 10149 14467
rect 10183 14433 10195 14467
rect 10137 14427 10195 14433
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14365 6699 14399
rect 6641 14359 6699 14365
rect 6411 14300 6500 14328
rect 6411 14297 6423 14300
rect 6365 14291 6423 14297
rect 6546 14288 6552 14340
rect 6604 14328 6610 14340
rect 6656 14328 6684 14359
rect 6822 14356 6828 14408
rect 6880 14396 6886 14408
rect 6968 14399 7026 14405
rect 6968 14396 6980 14399
rect 6880 14368 6980 14396
rect 6880 14356 6886 14368
rect 6968 14365 6980 14368
rect 7014 14365 7026 14399
rect 6968 14359 7026 14365
rect 7098 14356 7104 14408
rect 7156 14356 7162 14408
rect 7374 14356 7380 14408
rect 7432 14356 7438 14408
rect 10152 14396 10180 14427
rect 10318 14424 10324 14476
rect 10376 14464 10382 14476
rect 11256 14473 11284 14504
rect 11422 14492 11428 14504
rect 11480 14492 11486 14544
rect 11698 14492 11704 14544
rect 11756 14492 11762 14544
rect 10413 14467 10471 14473
rect 10413 14464 10425 14467
rect 10376 14436 10425 14464
rect 10376 14424 10382 14436
rect 10413 14433 10425 14436
rect 10459 14433 10471 14467
rect 10413 14427 10471 14433
rect 11241 14467 11299 14473
rect 11241 14433 11253 14467
rect 11287 14433 11299 14467
rect 11241 14427 11299 14433
rect 10152 14368 10364 14396
rect 10229 14331 10287 14337
rect 10229 14328 10241 14331
rect 6604 14300 6684 14328
rect 8266 14300 10241 14328
rect 6604 14288 6610 14300
rect 8266 14260 8294 14300
rect 10229 14297 10241 14300
rect 10275 14297 10287 14331
rect 10229 14291 10287 14297
rect 6288 14232 8294 14260
rect 8665 14263 8723 14269
rect 8665 14229 8677 14263
rect 8711 14260 8723 14263
rect 9858 14260 9864 14272
rect 8711 14232 9864 14260
rect 8711 14229 8723 14232
rect 8665 14223 8723 14229
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 10336 14260 10364 14368
rect 10428 14328 10456 14427
rect 11146 14356 11152 14408
rect 11204 14396 11210 14408
rect 11256 14396 11284 14427
rect 11330 14424 11336 14476
rect 11388 14464 11394 14476
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 11388 14436 11529 14464
rect 11388 14424 11394 14436
rect 11517 14433 11529 14436
rect 11563 14433 11575 14467
rect 11716 14464 11744 14492
rect 11936 14467 11994 14473
rect 11936 14464 11948 14467
rect 11716 14436 11948 14464
rect 11517 14427 11575 14433
rect 11936 14433 11948 14436
rect 11982 14433 11994 14467
rect 15672 14464 15700 14563
rect 16482 14560 16488 14612
rect 16540 14600 16546 14612
rect 19705 14603 19763 14609
rect 16540 14572 17080 14600
rect 16540 14560 16546 14572
rect 16942 14532 16948 14544
rect 16224 14504 16948 14532
rect 11936 14427 11994 14433
rect 12268 14436 15700 14464
rect 11204 14368 11284 14396
rect 11609 14399 11667 14405
rect 11204 14356 11210 14368
rect 11609 14365 11621 14399
rect 11655 14396 11667 14399
rect 11790 14396 11796 14408
rect 11655 14368 11796 14396
rect 11655 14365 11667 14368
rect 11609 14359 11667 14365
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 12115 14399 12173 14405
rect 12115 14365 12127 14399
rect 12161 14396 12173 14399
rect 12268 14396 12296 14436
rect 15930 14424 15936 14476
rect 15988 14464 15994 14476
rect 16224 14473 16252 14504
rect 16942 14492 16948 14504
rect 17000 14492 17006 14544
rect 16209 14467 16267 14473
rect 16209 14464 16221 14467
rect 15988 14436 16221 14464
rect 15988 14424 15994 14436
rect 16209 14433 16221 14436
rect 16255 14433 16267 14467
rect 16209 14427 16267 14433
rect 16298 14424 16304 14476
rect 16356 14464 16362 14476
rect 17052 14473 17080 14572
rect 19705 14569 19717 14603
rect 19751 14600 19763 14603
rect 19886 14600 19892 14612
rect 19751 14572 19892 14600
rect 19751 14569 19763 14572
rect 19705 14563 19763 14569
rect 19886 14560 19892 14572
rect 19944 14560 19950 14612
rect 19981 14603 20039 14609
rect 19981 14569 19993 14603
rect 20027 14600 20039 14603
rect 20162 14600 20168 14612
rect 20027 14572 20168 14600
rect 20027 14569 20039 14572
rect 19981 14563 20039 14569
rect 20162 14560 20168 14572
rect 20220 14560 20226 14612
rect 20257 14603 20315 14609
rect 20257 14569 20269 14603
rect 20303 14569 20315 14603
rect 20257 14563 20315 14569
rect 20533 14603 20591 14609
rect 20533 14569 20545 14603
rect 20579 14600 20591 14603
rect 20579 14572 21128 14600
rect 20579 14569 20591 14572
rect 20533 14563 20591 14569
rect 19610 14492 19616 14544
rect 19668 14532 19674 14544
rect 20272 14532 20300 14563
rect 20622 14532 20628 14544
rect 19668 14504 19932 14532
rect 20272 14504 20628 14532
rect 19668 14492 19674 14504
rect 19904 14476 19932 14504
rect 20622 14492 20628 14504
rect 20680 14492 20686 14544
rect 21100 14532 21128 14572
rect 21174 14560 21180 14612
rect 21232 14600 21238 14612
rect 21634 14600 21640 14612
rect 21232 14572 21640 14600
rect 21232 14560 21238 14572
rect 21634 14560 21640 14572
rect 21692 14600 21698 14612
rect 21735 14603 21793 14609
rect 21735 14600 21747 14603
rect 21692 14572 21747 14600
rect 21692 14560 21698 14572
rect 21735 14569 21747 14572
rect 21781 14569 21793 14603
rect 21735 14563 21793 14569
rect 23106 14560 23112 14612
rect 23164 14560 23170 14612
rect 23569 14603 23627 14609
rect 23569 14569 23581 14603
rect 23615 14569 23627 14603
rect 23569 14563 23627 14569
rect 23584 14532 23612 14563
rect 24578 14560 24584 14612
rect 24636 14609 24642 14612
rect 24636 14600 24645 14609
rect 24636 14572 24681 14600
rect 24636 14563 24645 14572
rect 24636 14560 24642 14563
rect 25590 14560 25596 14612
rect 25648 14560 25654 14612
rect 26142 14560 26148 14612
rect 26200 14560 26206 14612
rect 27798 14600 27804 14612
rect 26528 14572 27804 14600
rect 25608 14532 25636 14560
rect 26528 14532 26556 14572
rect 27798 14560 27804 14572
rect 27856 14560 27862 14612
rect 29270 14560 29276 14612
rect 29328 14600 29334 14612
rect 30377 14603 30435 14609
rect 30377 14600 30389 14603
rect 29328 14572 30389 14600
rect 29328 14560 29334 14572
rect 30377 14569 30389 14572
rect 30423 14569 30435 14603
rect 30377 14563 30435 14569
rect 30558 14560 30564 14612
rect 30616 14560 30622 14612
rect 21100 14504 21312 14532
rect 23584 14504 24256 14532
rect 25608 14504 26556 14532
rect 16853 14467 16911 14473
rect 16853 14464 16865 14467
rect 16356 14436 16865 14464
rect 16356 14424 16362 14436
rect 16853 14433 16865 14436
rect 16899 14433 16911 14467
rect 16853 14427 16911 14433
rect 17037 14467 17095 14473
rect 17037 14433 17049 14467
rect 17083 14433 17095 14467
rect 17037 14427 17095 14433
rect 19429 14467 19487 14473
rect 19429 14433 19441 14467
rect 19475 14433 19487 14467
rect 19429 14427 19487 14433
rect 17533 14417 17591 14423
rect 17533 14414 17545 14417
rect 17512 14408 17545 14414
rect 12161 14368 12296 14396
rect 12161 14365 12173 14368
rect 12115 14359 12173 14365
rect 12342 14356 12348 14408
rect 12400 14356 12406 14408
rect 13817 14399 13875 14405
rect 13817 14365 13829 14399
rect 13863 14396 13875 14399
rect 14182 14396 14188 14408
rect 13863 14368 14188 14396
rect 13863 14365 13875 14368
rect 13817 14359 13875 14365
rect 14182 14356 14188 14368
rect 14240 14356 14246 14408
rect 14323 14399 14381 14405
rect 14323 14365 14335 14399
rect 14369 14396 14381 14399
rect 14458 14396 14464 14408
rect 14369 14368 14464 14396
rect 14369 14365 14381 14368
rect 14323 14359 14381 14365
rect 14458 14356 14464 14368
rect 14516 14356 14522 14408
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14396 14611 14399
rect 14599 14368 16712 14396
rect 14599 14365 14611 14368
rect 14553 14359 14611 14365
rect 16684 14337 16712 14368
rect 16758 14356 16764 14408
rect 16816 14396 16822 14408
rect 17364 14399 17422 14405
rect 17364 14396 17376 14399
rect 16816 14368 17376 14396
rect 16816 14356 16822 14368
rect 17364 14365 17376 14368
rect 17410 14365 17422 14399
rect 17364 14359 17422 14365
rect 17494 14356 17500 14408
rect 17579 14383 17591 14417
rect 17552 14377 17591 14383
rect 17773 14399 17831 14405
rect 17552 14356 17558 14377
rect 17773 14365 17785 14399
rect 17819 14396 17831 14399
rect 19444 14396 19472 14427
rect 19886 14424 19892 14476
rect 19944 14424 19950 14476
rect 20162 14424 20168 14476
rect 20220 14424 20226 14476
rect 20441 14467 20499 14473
rect 20441 14433 20453 14467
rect 20487 14464 20499 14467
rect 20530 14464 20536 14476
rect 20487 14436 20536 14464
rect 20487 14433 20499 14436
rect 20441 14427 20499 14433
rect 20530 14424 20536 14436
rect 20588 14424 20594 14476
rect 20717 14467 20775 14473
rect 20717 14433 20729 14467
rect 20763 14464 20775 14467
rect 20993 14467 21051 14473
rect 20763 14436 20852 14464
rect 20763 14433 20775 14436
rect 20717 14427 20775 14433
rect 20824 14408 20852 14436
rect 20993 14433 21005 14467
rect 21039 14433 21051 14467
rect 21284 14464 21312 14504
rect 22005 14467 22063 14473
rect 22005 14464 22017 14467
rect 21284 14436 22017 14464
rect 20993 14427 21051 14433
rect 22005 14433 22017 14436
rect 22051 14433 22063 14467
rect 22005 14427 22063 14433
rect 20806 14396 20812 14408
rect 17819 14368 19288 14396
rect 19444 14368 20812 14396
rect 17819 14365 17831 14368
rect 17773 14359 17831 14365
rect 19260 14337 19288 14368
rect 20806 14356 20812 14368
rect 20864 14356 20870 14408
rect 21008 14340 21036 14427
rect 23566 14424 23572 14476
rect 23624 14424 23630 14476
rect 23750 14424 23756 14476
rect 23808 14464 23814 14476
rect 23934 14464 23940 14476
rect 23808 14436 23940 14464
rect 23808 14424 23814 14436
rect 23934 14424 23940 14436
rect 23992 14424 23998 14476
rect 24026 14424 24032 14476
rect 24084 14424 24090 14476
rect 24228 14464 24256 14504
rect 24857 14467 24915 14473
rect 24857 14464 24869 14467
rect 24228 14436 24869 14464
rect 24857 14433 24869 14436
rect 24903 14433 24915 14467
rect 24857 14427 24915 14433
rect 25958 14424 25964 14476
rect 26016 14464 26022 14476
rect 26421 14467 26479 14473
rect 26421 14464 26433 14467
rect 26016 14436 26433 14464
rect 26016 14424 26022 14436
rect 26421 14433 26433 14436
rect 26467 14464 26479 14467
rect 26510 14464 26516 14476
rect 26467 14436 26516 14464
rect 26467 14433 26479 14436
rect 26421 14427 26479 14433
rect 26510 14424 26516 14436
rect 26568 14424 26574 14476
rect 26697 14467 26755 14473
rect 26697 14433 26709 14467
rect 26743 14464 26755 14467
rect 27338 14464 27344 14476
rect 26743 14436 27344 14464
rect 26743 14433 26755 14436
rect 26697 14427 26755 14433
rect 27338 14424 27344 14436
rect 27396 14424 27402 14476
rect 27706 14424 27712 14476
rect 27764 14464 27770 14476
rect 30576 14473 30604 14560
rect 28496 14467 28554 14473
rect 28496 14464 28508 14467
rect 27764 14436 28508 14464
rect 27764 14424 27770 14436
rect 28496 14433 28508 14436
rect 28542 14433 28554 14467
rect 30561 14467 30619 14473
rect 28496 14427 28554 14433
rect 28828 14436 30512 14464
rect 21266 14356 21272 14408
rect 21324 14356 21330 14408
rect 21775 14399 21833 14405
rect 21775 14365 21787 14399
rect 21821 14396 21833 14399
rect 23584 14396 23612 14424
rect 21821 14368 23612 14396
rect 21821 14365 21833 14368
rect 21775 14359 21833 14365
rect 23842 14356 23848 14408
rect 23900 14396 23906 14408
rect 24121 14399 24179 14405
rect 24121 14396 24133 14399
rect 23900 14368 24133 14396
rect 23900 14356 23906 14368
rect 24121 14365 24133 14368
rect 24167 14365 24179 14399
rect 24121 14359 24179 14365
rect 24627 14399 24685 14405
rect 24627 14365 24639 14399
rect 24673 14396 24685 14399
rect 25682 14396 25688 14408
rect 24673 14368 25688 14396
rect 24673 14365 24685 14368
rect 24627 14359 24685 14365
rect 25682 14356 25688 14368
rect 25740 14356 25746 14408
rect 26878 14356 26884 14408
rect 26936 14396 26942 14408
rect 28169 14399 28227 14405
rect 28169 14396 28181 14399
rect 26936 14368 28181 14396
rect 26936 14356 26942 14368
rect 28169 14365 28181 14368
rect 28215 14365 28227 14399
rect 28169 14359 28227 14365
rect 28675 14399 28733 14405
rect 28675 14365 28687 14399
rect 28721 14396 28733 14399
rect 28828 14396 28856 14436
rect 28721 14368 28856 14396
rect 28905 14399 28963 14405
rect 28721 14365 28733 14368
rect 28675 14359 28733 14365
rect 28905 14365 28917 14399
rect 28951 14396 28963 14399
rect 29270 14396 29276 14408
rect 28951 14368 29276 14396
rect 28951 14365 28963 14368
rect 28905 14359 28963 14365
rect 29270 14356 29276 14368
rect 29328 14356 29334 14408
rect 30484 14396 30512 14436
rect 30561 14433 30573 14467
rect 30607 14433 30619 14467
rect 30561 14427 30619 14433
rect 30650 14396 30656 14408
rect 30484 14368 30656 14396
rect 30650 14356 30656 14368
rect 30708 14356 30714 14408
rect 16669 14331 16727 14337
rect 10428 14300 11284 14328
rect 11256 14272 11284 14300
rect 15212 14300 16436 14328
rect 10870 14260 10876 14272
rect 10336 14232 10876 14260
rect 10870 14220 10876 14232
rect 10928 14220 10934 14272
rect 11238 14220 11244 14272
rect 11296 14220 11302 14272
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 14182 14260 14188 14272
rect 12860 14232 14188 14260
rect 12860 14220 12866 14232
rect 14182 14220 14188 14232
rect 14240 14220 14246 14272
rect 14458 14220 14464 14272
rect 14516 14260 14522 14272
rect 15212 14260 15240 14300
rect 14516 14232 15240 14260
rect 14516 14220 14522 14232
rect 16298 14220 16304 14272
rect 16356 14220 16362 14272
rect 16408 14260 16436 14300
rect 16669 14297 16681 14331
rect 16715 14297 16727 14331
rect 16669 14291 16727 14297
rect 19245 14331 19303 14337
rect 19245 14297 19257 14331
rect 19291 14297 19303 14331
rect 19245 14291 19303 14297
rect 20990 14288 20996 14340
rect 21048 14288 21054 14340
rect 18877 14263 18935 14269
rect 18877 14260 18889 14263
rect 16408 14232 18889 14260
rect 18877 14229 18889 14232
rect 18923 14229 18935 14263
rect 18877 14223 18935 14229
rect 20714 14220 20720 14272
rect 20772 14260 20778 14272
rect 20809 14263 20867 14269
rect 20809 14260 20821 14263
rect 20772 14232 20821 14260
rect 20772 14220 20778 14232
rect 20809 14229 20821 14232
rect 20855 14229 20867 14263
rect 20809 14223 20867 14229
rect 20898 14220 20904 14272
rect 20956 14260 20962 14272
rect 21284 14260 21312 14356
rect 23860 14328 23888 14356
rect 23584 14300 23888 14328
rect 27356 14300 28120 14328
rect 20956 14232 21312 14260
rect 20956 14220 20962 14232
rect 21450 14220 21456 14272
rect 21508 14260 21514 14272
rect 23584 14260 23612 14300
rect 21508 14232 23612 14260
rect 23845 14263 23903 14269
rect 21508 14220 21514 14232
rect 23845 14229 23857 14263
rect 23891 14260 23903 14263
rect 24670 14260 24676 14272
rect 23891 14232 24676 14260
rect 23891 14229 23903 14232
rect 23845 14223 23903 14229
rect 24670 14220 24676 14232
rect 24728 14220 24734 14272
rect 24854 14220 24860 14272
rect 24912 14260 24918 14272
rect 27356 14260 27384 14300
rect 24912 14232 27384 14260
rect 24912 14220 24918 14232
rect 27982 14220 27988 14272
rect 28040 14220 28046 14272
rect 28092 14260 28120 14300
rect 29914 14288 29920 14340
rect 29972 14328 29978 14340
rect 30009 14331 30067 14337
rect 30009 14328 30021 14331
rect 29972 14300 30021 14328
rect 29972 14288 29978 14300
rect 30009 14297 30021 14300
rect 30055 14297 30067 14331
rect 30009 14291 30067 14297
rect 29086 14260 29092 14272
rect 28092 14232 29092 14260
rect 29086 14220 29092 14232
rect 29144 14260 29150 14272
rect 29638 14260 29644 14272
rect 29144 14232 29644 14260
rect 29144 14220 29150 14232
rect 29638 14220 29644 14232
rect 29696 14260 29702 14272
rect 31202 14260 31208 14272
rect 29696 14232 31208 14260
rect 29696 14220 29702 14232
rect 31202 14220 31208 14232
rect 31260 14220 31266 14272
rect 552 14170 30912 14192
rect 552 14118 4193 14170
rect 4245 14118 4257 14170
rect 4309 14118 4321 14170
rect 4373 14118 4385 14170
rect 4437 14118 4449 14170
rect 4501 14118 11783 14170
rect 11835 14118 11847 14170
rect 11899 14118 11911 14170
rect 11963 14118 11975 14170
rect 12027 14118 12039 14170
rect 12091 14118 19373 14170
rect 19425 14118 19437 14170
rect 19489 14118 19501 14170
rect 19553 14118 19565 14170
rect 19617 14118 19629 14170
rect 19681 14118 26963 14170
rect 27015 14118 27027 14170
rect 27079 14118 27091 14170
rect 27143 14118 27155 14170
rect 27207 14118 27219 14170
rect 27271 14118 30912 14170
rect 552 14096 30912 14118
rect 1302 14056 1308 14068
rect 952 14028 1308 14056
rect 750 13880 756 13932
rect 808 13920 814 13932
rect 952 13929 980 14028
rect 1302 14016 1308 14028
rect 1360 14016 1366 14068
rect 4062 14056 4068 14068
rect 3344 14028 4068 14056
rect 3344 13997 3372 14028
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 5810 14016 5816 14068
rect 5868 14056 5874 14068
rect 6730 14056 6736 14068
rect 5868 14028 6736 14056
rect 5868 14016 5874 14028
rect 6730 14016 6736 14028
rect 6788 14016 6794 14068
rect 7650 14016 7656 14068
rect 7708 14056 7714 14068
rect 8389 14059 8447 14065
rect 8389 14056 8401 14059
rect 7708 14028 8401 14056
rect 7708 14016 7714 14028
rect 8389 14025 8401 14028
rect 8435 14025 8447 14059
rect 8665 14059 8723 14065
rect 8665 14056 8677 14059
rect 8389 14019 8447 14025
rect 8496 14028 8677 14056
rect 3329 13991 3387 13997
rect 3329 13957 3341 13991
rect 3375 13957 3387 13991
rect 3329 13951 3387 13957
rect 7834 13948 7840 14000
rect 7892 13988 7898 14000
rect 7929 13991 7987 13997
rect 7929 13988 7941 13991
rect 7892 13960 7941 13988
rect 7892 13948 7898 13960
rect 7929 13957 7941 13960
rect 7975 13957 7987 13991
rect 8496 13988 8524 14028
rect 8665 14025 8677 14028
rect 8711 14025 8723 14059
rect 8665 14019 8723 14025
rect 9033 14059 9091 14065
rect 9033 14025 9045 14059
rect 9079 14056 9091 14059
rect 9214 14056 9220 14068
rect 9079 14028 9220 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 9309 14059 9367 14065
rect 9309 14025 9321 14059
rect 9355 14056 9367 14059
rect 9398 14056 9404 14068
rect 9355 14028 9404 14056
rect 9355 14025 9367 14028
rect 9309 14019 9367 14025
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 9508 14028 12480 14056
rect 8754 13988 8760 14000
rect 7929 13951 7987 13957
rect 8036 13960 8524 13988
rect 8588 13960 8760 13988
rect 937 13923 995 13929
rect 937 13920 949 13923
rect 808 13892 949 13920
rect 808 13880 814 13892
rect 937 13889 949 13892
rect 983 13889 995 13923
rect 937 13883 995 13889
rect 1443 13923 1501 13929
rect 1443 13889 1455 13923
rect 1489 13920 1501 13923
rect 3142 13920 3148 13932
rect 1489 13892 3148 13920
rect 1489 13889 1501 13892
rect 1443 13883 1501 13889
rect 3142 13880 3148 13892
rect 3200 13880 3206 13932
rect 3697 13923 3755 13929
rect 3697 13920 3709 13923
rect 3436 13892 3709 13920
rect 3436 13864 3464 13892
rect 3697 13889 3709 13892
rect 3743 13889 3755 13923
rect 3697 13883 3755 13889
rect 3878 13880 3884 13932
rect 3936 13920 3942 13932
rect 4203 13923 4261 13929
rect 4203 13920 4215 13923
rect 3936 13892 4215 13920
rect 3936 13880 3942 13892
rect 4203 13889 4215 13892
rect 4249 13889 4261 13923
rect 4203 13883 4261 13889
rect 6086 13880 6092 13932
rect 6144 13880 6150 13932
rect 6638 13929 6644 13932
rect 6595 13923 6644 13929
rect 6595 13889 6607 13923
rect 6641 13889 6644 13923
rect 6595 13883 6644 13889
rect 6638 13880 6644 13883
rect 6696 13880 6702 13932
rect 6730 13880 6736 13932
rect 6788 13920 6794 13932
rect 6788 13892 6868 13920
rect 6788 13880 6794 13892
rect 1670 13812 1676 13864
rect 1728 13812 1734 13864
rect 3418 13812 3424 13864
rect 3476 13812 3482 13864
rect 3510 13812 3516 13864
rect 3568 13812 3574 13864
rect 4433 13855 4491 13861
rect 4433 13821 4445 13855
rect 4479 13852 4491 13855
rect 5166 13852 5172 13864
rect 4479 13824 5172 13852
rect 4479 13821 4491 13824
rect 4433 13815 4491 13821
rect 5166 13812 5172 13824
rect 5224 13812 5230 13864
rect 6454 13861 6460 13864
rect 6416 13855 6460 13861
rect 6416 13821 6428 13855
rect 6416 13815 6460 13821
rect 6454 13812 6460 13815
rect 6512 13812 6518 13864
rect 6840 13861 6868 13892
rect 7006 13880 7012 13932
rect 7064 13880 7070 13932
rect 8036 13920 8064 13960
rect 7760 13892 8064 13920
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13821 6883 13855
rect 7024 13852 7052 13880
rect 7760 13852 7788 13892
rect 8588 13861 8616 13960
rect 8754 13948 8760 13960
rect 8812 13988 8818 14000
rect 9508 13988 9536 14028
rect 12158 13988 12164 14000
rect 8812 13960 9536 13988
rect 10980 13960 12164 13988
rect 8812 13948 8818 13960
rect 8662 13880 8668 13932
rect 8720 13920 8726 13932
rect 8720 13892 9536 13920
rect 8720 13880 8726 13892
rect 7024 13824 7788 13852
rect 8573 13855 8631 13861
rect 6825 13815 6883 13821
rect 8573 13821 8585 13855
rect 8619 13821 8631 13855
rect 8680 13852 8708 13880
rect 9508 13861 9536 13892
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 10048 13923 10106 13929
rect 10048 13920 10060 13923
rect 9916 13892 10060 13920
rect 9916 13880 9922 13892
rect 10048 13889 10060 13892
rect 10094 13889 10106 13923
rect 10048 13883 10106 13889
rect 10152 13892 10732 13920
rect 10152 13864 10180 13892
rect 8849 13855 8907 13861
rect 8849 13852 8861 13855
rect 8680 13824 8861 13852
rect 8573 13815 8631 13821
rect 8849 13821 8861 13824
rect 8895 13821 8907 13855
rect 8849 13815 8907 13821
rect 9217 13855 9275 13861
rect 9217 13821 9229 13855
rect 9263 13821 9275 13855
rect 9217 13815 9275 13821
rect 9493 13855 9551 13861
rect 9493 13821 9505 13855
rect 9539 13821 9551 13855
rect 9493 13815 9551 13821
rect 9611 13855 9669 13861
rect 9611 13821 9623 13855
rect 9657 13852 9669 13855
rect 9657 13821 9674 13852
rect 9611 13815 9674 13821
rect 5813 13787 5871 13793
rect 5813 13753 5825 13787
rect 5859 13784 5871 13787
rect 6086 13784 6092 13796
rect 5859 13756 6092 13784
rect 5859 13753 5871 13756
rect 5813 13747 5871 13753
rect 6086 13744 6092 13756
rect 6144 13744 6150 13796
rect 1403 13719 1461 13725
rect 1403 13685 1415 13719
rect 1449 13716 1461 13719
rect 1578 13716 1584 13728
rect 1449 13688 1584 13716
rect 1449 13685 1461 13688
rect 1403 13679 1461 13685
rect 1578 13676 1584 13688
rect 1636 13716 1642 13728
rect 2314 13716 2320 13728
rect 1636 13688 2320 13716
rect 1636 13676 1642 13688
rect 2314 13676 2320 13688
rect 2372 13676 2378 13728
rect 2774 13676 2780 13728
rect 2832 13676 2838 13728
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 4163 13719 4221 13725
rect 4163 13716 4175 13719
rect 4028 13688 4175 13716
rect 4028 13676 4034 13688
rect 4163 13685 4175 13688
rect 4209 13685 4221 13719
rect 4163 13679 4221 13685
rect 5534 13676 5540 13728
rect 5592 13716 5598 13728
rect 8588 13716 8616 13815
rect 5592 13688 8616 13716
rect 9232 13716 9260 13815
rect 9646 13784 9674 13815
rect 10134 13812 10140 13864
rect 10192 13812 10198 13864
rect 10318 13812 10324 13864
rect 10376 13812 10382 13864
rect 10704 13852 10732 13892
rect 10778 13880 10784 13932
rect 10836 13920 10842 13932
rect 10980 13920 11008 13960
rect 12158 13948 12164 13960
rect 12216 13948 12222 14000
rect 12342 13948 12348 14000
rect 12400 13948 12406 14000
rect 12452 13988 12480 14028
rect 12526 14016 12532 14068
rect 12584 14056 12590 14068
rect 12621 14059 12679 14065
rect 12621 14056 12633 14059
rect 12584 14028 12633 14056
rect 12584 14016 12590 14028
rect 12621 14025 12633 14028
rect 12667 14025 12679 14059
rect 12621 14019 12679 14025
rect 13725 14059 13783 14065
rect 13725 14025 13737 14059
rect 13771 14056 13783 14059
rect 13771 14028 15700 14056
rect 13771 14025 13783 14028
rect 13725 14019 13783 14025
rect 13078 13988 13084 14000
rect 12452 13960 13084 13988
rect 10836 13892 11008 13920
rect 11701 13923 11759 13929
rect 10836 13880 10842 13892
rect 11701 13889 11713 13923
rect 11747 13920 11759 13923
rect 12434 13920 12440 13932
rect 11747 13892 12440 13920
rect 11747 13889 11759 13892
rect 11701 13883 11759 13889
rect 12434 13880 12440 13892
rect 12492 13880 12498 13932
rect 11422 13852 11428 13864
rect 10704 13824 11428 13852
rect 11422 13812 11428 13824
rect 11480 13852 11486 13864
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 11480 13824 11805 13852
rect 11480 13812 11486 13824
rect 11793 13821 11805 13824
rect 11839 13821 11851 13855
rect 11793 13815 11851 13821
rect 11882 13812 11888 13864
rect 11940 13852 11946 13864
rect 12069 13855 12127 13861
rect 12069 13852 12081 13855
rect 11940 13824 12081 13852
rect 11940 13812 11946 13824
rect 12069 13821 12081 13824
rect 12115 13821 12127 13855
rect 12069 13815 12127 13821
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13852 12587 13855
rect 12636 13852 12664 13960
rect 13078 13948 13084 13960
rect 13136 13948 13142 14000
rect 13354 13948 13360 14000
rect 13412 13948 13418 14000
rect 13446 13948 13452 14000
rect 13504 13988 13510 14000
rect 13740 13988 13768 14019
rect 15672 14000 15700 14028
rect 16390 14016 16396 14068
rect 16448 14056 16454 14068
rect 16448 14028 17816 14056
rect 16448 14016 16454 14028
rect 13504 13960 13768 13988
rect 13504 13948 13510 13960
rect 15654 13948 15660 14000
rect 15712 13948 15718 14000
rect 17788 13988 17816 14028
rect 17954 14016 17960 14068
rect 18012 14056 18018 14068
rect 18693 14059 18751 14065
rect 18693 14056 18705 14059
rect 18012 14028 18705 14056
rect 18012 14016 18018 14028
rect 18693 14025 18705 14028
rect 18739 14025 18751 14059
rect 21637 14059 21695 14065
rect 21637 14056 21649 14059
rect 18693 14019 18751 14025
rect 19260 14028 21649 14056
rect 18233 13991 18291 13997
rect 18233 13988 18245 13991
rect 17788 13960 18245 13988
rect 18233 13957 18245 13960
rect 18279 13957 18291 13991
rect 18233 13951 18291 13957
rect 14090 13880 14096 13932
rect 14148 13920 14154 13932
rect 14550 13929 14556 13932
rect 14185 13923 14243 13929
rect 14185 13920 14197 13923
rect 14148 13892 14197 13920
rect 14148 13880 14154 13892
rect 14185 13889 14197 13892
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14512 13923 14556 13929
rect 14512 13889 14524 13923
rect 14512 13883 14556 13889
rect 14550 13880 14556 13883
rect 14608 13880 14614 13932
rect 14691 13923 14749 13929
rect 14691 13889 14703 13923
rect 14737 13920 14749 13923
rect 14826 13920 14832 13932
rect 14737 13892 14832 13920
rect 14737 13889 14749 13892
rect 14691 13883 14749 13889
rect 14826 13880 14832 13892
rect 14884 13880 14890 13932
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13920 14979 13923
rect 16022 13920 16028 13932
rect 14967 13892 16028 13920
rect 14967 13889 14979 13892
rect 14921 13883 14979 13889
rect 16022 13880 16028 13892
rect 16080 13880 16086 13932
rect 16758 13929 16764 13932
rect 16720 13923 16764 13929
rect 16720 13889 16732 13923
rect 16720 13883 16764 13889
rect 16758 13880 16764 13883
rect 16816 13880 16822 13932
rect 16899 13923 16957 13929
rect 16899 13889 16911 13923
rect 16945 13920 16957 13923
rect 19260 13920 19288 14028
rect 21637 14025 21649 14028
rect 21683 14025 21695 14059
rect 21637 14019 21695 14025
rect 21726 14016 21732 14068
rect 21784 14056 21790 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 21784 14028 23397 14056
rect 21784 14016 21790 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 27522 14056 27528 14068
rect 23385 14019 23443 14025
rect 24044 14028 25452 14056
rect 19518 13948 19524 14000
rect 19576 13948 19582 14000
rect 23014 13948 23020 14000
rect 23072 13988 23078 14000
rect 24044 13988 24072 14028
rect 23072 13960 24072 13988
rect 23072 13948 23078 13960
rect 20162 13920 20168 13932
rect 16945 13892 19288 13920
rect 19720 13892 20168 13920
rect 16945 13889 16957 13892
rect 16899 13883 16957 13889
rect 12575 13824 12664 13852
rect 12805 13855 12863 13861
rect 12575 13821 12587 13824
rect 12529 13815 12587 13821
rect 12805 13821 12817 13855
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 9646 13756 9720 13784
rect 9398 13716 9404 13728
rect 9232 13688 9404 13716
rect 5592 13676 5598 13688
rect 9398 13676 9404 13688
rect 9456 13676 9462 13728
rect 9582 13676 9588 13728
rect 9640 13716 9646 13728
rect 9692 13716 9720 13756
rect 11514 13744 11520 13796
rect 11572 13784 11578 13796
rect 11698 13784 11704 13796
rect 11572 13756 11704 13784
rect 11572 13744 11578 13756
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 12820 13784 12848 13815
rect 12894 13812 12900 13864
rect 12952 13812 12958 13864
rect 13170 13812 13176 13864
rect 13228 13852 13234 13864
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 13228 13824 13553 13852
rect 13228 13812 13234 13824
rect 13541 13821 13553 13824
rect 13587 13821 13599 13855
rect 13541 13815 13599 13821
rect 14274 13812 14280 13864
rect 14332 13852 14338 13864
rect 16301 13855 16359 13861
rect 16301 13852 16313 13855
rect 14332 13824 16313 13852
rect 14332 13812 14338 13824
rect 16301 13821 16313 13824
rect 16347 13821 16359 13855
rect 16301 13815 16359 13821
rect 16393 13855 16451 13861
rect 16393 13821 16405 13855
rect 16439 13852 16451 13855
rect 16482 13852 16488 13864
rect 16439 13824 16488 13852
rect 16439 13821 16451 13824
rect 16393 13815 16451 13821
rect 16482 13812 16488 13824
rect 16540 13812 16546 13864
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17494 13852 17500 13864
rect 17175 13824 17500 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17494 13812 17500 13824
rect 17552 13812 17558 13864
rect 18874 13812 18880 13864
rect 18932 13812 18938 13864
rect 19150 13812 19156 13864
rect 19208 13812 19214 13864
rect 19720 13861 19748 13892
rect 20162 13880 20168 13892
rect 20220 13880 20226 13932
rect 20303 13923 20361 13929
rect 20303 13889 20315 13923
rect 20349 13920 20361 13923
rect 20438 13920 20444 13932
rect 20349 13892 20444 13920
rect 20349 13889 20361 13892
rect 20303 13883 20361 13889
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 20533 13923 20591 13929
rect 20533 13889 20545 13923
rect 20579 13920 20591 13923
rect 20714 13920 20720 13932
rect 20579 13892 20720 13920
rect 20579 13889 20591 13892
rect 20533 13883 20591 13889
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 20990 13880 20996 13932
rect 21048 13920 21054 13932
rect 21818 13920 21824 13932
rect 21048 13892 21824 13920
rect 21048 13880 21054 13892
rect 21818 13880 21824 13892
rect 21876 13920 21882 13932
rect 21876 13892 22140 13920
rect 21876 13880 21882 13892
rect 19705 13855 19763 13861
rect 19705 13821 19717 13855
rect 19751 13821 19763 13855
rect 19705 13815 19763 13821
rect 19794 13812 19800 13864
rect 19852 13852 19858 13864
rect 20898 13852 20904 13864
rect 19852 13824 20904 13852
rect 19852 13812 19858 13824
rect 20898 13812 20904 13824
rect 20956 13812 20962 13864
rect 22002 13861 22008 13864
rect 21994 13855 22008 13861
rect 21994 13852 22006 13855
rect 21963 13824 22006 13852
rect 21994 13821 22006 13824
rect 21994 13815 22008 13821
rect 22002 13812 22008 13815
rect 22060 13812 22066 13864
rect 22112 13852 22140 13892
rect 22186 13880 22192 13932
rect 22244 13920 22250 13932
rect 22281 13923 22339 13929
rect 22281 13920 22293 13923
rect 22244 13892 22293 13920
rect 22244 13880 22250 13892
rect 22281 13889 22293 13892
rect 22327 13889 22339 13923
rect 22281 13883 22339 13889
rect 23842 13880 23848 13932
rect 23900 13920 23906 13932
rect 23900 13892 24072 13920
rect 23900 13880 23906 13892
rect 23934 13852 23940 13864
rect 22112 13824 23940 13852
rect 23934 13812 23940 13824
rect 23992 13812 23998 13864
rect 24044 13861 24072 13892
rect 24210 13880 24216 13932
rect 24268 13920 24274 13932
rect 24492 13923 24550 13929
rect 24492 13920 24504 13923
rect 24268 13892 24504 13920
rect 24268 13880 24274 13892
rect 24492 13889 24504 13892
rect 24538 13889 24550 13923
rect 24492 13883 24550 13889
rect 24578 13880 24584 13932
rect 24636 13880 24642 13932
rect 24670 13880 24676 13932
rect 24728 13920 24734 13932
rect 24765 13923 24823 13929
rect 24765 13920 24777 13923
rect 24728 13892 24777 13920
rect 24728 13880 24734 13892
rect 24765 13889 24777 13892
rect 24811 13889 24823 13923
rect 25424 13920 25452 14028
rect 26344 14028 27528 14056
rect 25498 13948 25504 14000
rect 25556 13988 25562 14000
rect 26237 13991 26295 13997
rect 26237 13988 26249 13991
rect 25556 13960 26249 13988
rect 25556 13948 25562 13960
rect 26237 13957 26249 13960
rect 26283 13957 26295 13991
rect 26237 13951 26295 13957
rect 26344 13920 26372 14028
rect 27522 14016 27528 14028
rect 27580 14016 27586 14068
rect 27614 14016 27620 14068
rect 27672 14056 27678 14068
rect 28537 14059 28595 14065
rect 28537 14056 28549 14059
rect 27672 14028 28549 14056
rect 27672 14016 27678 14028
rect 28537 14025 28549 14028
rect 28583 14025 28595 14059
rect 28537 14019 28595 14025
rect 28994 14016 29000 14068
rect 29052 14056 29058 14068
rect 29273 14059 29331 14065
rect 29273 14056 29285 14059
rect 29052 14028 29285 14056
rect 29052 14016 29058 14028
rect 29273 14025 29285 14028
rect 29319 14025 29331 14059
rect 29273 14019 29331 14025
rect 29546 14016 29552 14068
rect 29604 14016 29610 14068
rect 29825 14059 29883 14065
rect 29825 14056 29837 14059
rect 29656 14028 29837 14056
rect 25424 13892 26372 13920
rect 26697 13923 26755 13929
rect 24765 13883 24823 13889
rect 26697 13889 26709 13923
rect 26743 13920 26755 13923
rect 26878 13920 26884 13932
rect 26743 13892 26884 13920
rect 26743 13889 26755 13892
rect 26697 13883 26755 13889
rect 26878 13880 26884 13892
rect 26936 13880 26942 13932
rect 27062 13880 27068 13932
rect 27120 13880 27126 13932
rect 27338 13920 27344 13932
rect 27172 13905 27344 13920
rect 24029 13855 24087 13861
rect 24029 13821 24041 13855
rect 24075 13852 24087 13855
rect 24118 13852 24124 13864
rect 24075 13824 24124 13852
rect 24075 13821 24087 13824
rect 24029 13815 24087 13821
rect 24118 13812 24124 13824
rect 24176 13812 24182 13864
rect 24356 13855 24414 13861
rect 24356 13821 24368 13855
rect 24402 13852 24414 13855
rect 24596 13852 24624 13880
rect 26418 13861 26424 13864
rect 26413 13852 26424 13861
rect 24402 13824 24624 13852
rect 26379 13824 26424 13852
rect 24402 13821 24414 13824
rect 24356 13815 24414 13821
rect 26413 13815 26424 13824
rect 26418 13812 26424 13815
rect 26476 13812 26482 13864
rect 27080 13852 27108 13880
rect 27172 13874 27205 13905
rect 27193 13871 27205 13874
rect 27239 13892 27344 13905
rect 27239 13871 27251 13892
rect 27338 13880 27344 13892
rect 27396 13880 27402 13932
rect 27614 13880 27620 13932
rect 27672 13920 27678 13932
rect 29656 13920 29684 14028
rect 29825 14025 29837 14028
rect 29871 14025 29883 14059
rect 29825 14019 29883 14025
rect 30098 14016 30104 14068
rect 30156 14016 30162 14068
rect 30282 14016 30288 14068
rect 30340 14016 30346 14068
rect 29914 13988 29920 14000
rect 27672 13892 29684 13920
rect 29748 13960 29920 13988
rect 27672 13880 27678 13892
rect 27193 13865 27251 13871
rect 26528 13824 27108 13852
rect 12986 13784 12992 13796
rect 12544 13756 12992 13784
rect 9640 13688 9720 13716
rect 9640 13676 9646 13688
rect 10042 13676 10048 13728
rect 10100 13725 10106 13728
rect 10100 13679 10109 13725
rect 10100 13676 10106 13679
rect 10686 13676 10692 13728
rect 10744 13716 10750 13728
rect 12544 13716 12572 13756
rect 12986 13744 12992 13756
rect 13044 13744 13050 13796
rect 19242 13784 19248 13796
rect 17788 13756 19248 13784
rect 10744 13688 12572 13716
rect 10744 13676 10750 13688
rect 12618 13676 12624 13728
rect 12676 13716 12682 13728
rect 13170 13716 13176 13728
rect 12676 13688 13176 13716
rect 12676 13676 12682 13688
rect 13170 13676 13176 13688
rect 13228 13676 13234 13728
rect 13814 13676 13820 13728
rect 13872 13676 13878 13728
rect 14182 13676 14188 13728
rect 14240 13716 14246 13728
rect 15010 13716 15016 13728
rect 14240 13688 15016 13716
rect 14240 13676 14246 13688
rect 15010 13676 15016 13688
rect 15068 13716 15074 13728
rect 17788 13716 17816 13756
rect 19242 13744 19248 13756
rect 19300 13744 19306 13796
rect 26145 13787 26203 13793
rect 26145 13753 26157 13787
rect 26191 13784 26203 13787
rect 26528 13784 26556 13824
rect 27430 13812 27436 13864
rect 27488 13812 27494 13864
rect 27798 13812 27804 13864
rect 27856 13852 27862 13864
rect 27856 13824 29040 13852
rect 27856 13812 27862 13824
rect 26191 13756 26556 13784
rect 29012 13784 29040 13824
rect 29086 13812 29092 13864
rect 29144 13852 29150 13864
rect 29748 13861 29776 13960
rect 29914 13948 29920 13960
rect 29972 13988 29978 14000
rect 30300 13988 30328 14016
rect 29972 13960 30328 13988
rect 29972 13948 29978 13960
rect 29181 13855 29239 13861
rect 29181 13852 29193 13855
rect 29144 13824 29193 13852
rect 29144 13812 29150 13824
rect 29181 13821 29193 13824
rect 29227 13821 29239 13855
rect 29181 13815 29239 13821
rect 29457 13855 29515 13861
rect 29457 13821 29469 13855
rect 29503 13821 29515 13855
rect 29457 13815 29515 13821
rect 29733 13855 29791 13861
rect 29733 13821 29745 13855
rect 29779 13821 29791 13855
rect 29733 13815 29791 13821
rect 29472 13784 29500 13815
rect 29822 13812 29828 13864
rect 29880 13852 29886 13864
rect 30009 13855 30067 13861
rect 30009 13852 30021 13855
rect 29880 13824 30021 13852
rect 29880 13812 29886 13824
rect 30009 13821 30021 13824
rect 30055 13821 30067 13855
rect 30009 13815 30067 13821
rect 30285 13855 30343 13861
rect 30285 13821 30297 13855
rect 30331 13852 30343 13855
rect 30374 13852 30380 13864
rect 30331 13824 30380 13852
rect 30331 13821 30343 13824
rect 30285 13815 30343 13821
rect 30374 13812 30380 13824
rect 30432 13852 30438 13864
rect 30561 13855 30619 13861
rect 30561 13852 30573 13855
rect 30432 13824 30573 13852
rect 30432 13812 30438 13824
rect 30561 13821 30573 13824
rect 30607 13821 30619 13855
rect 30561 13815 30619 13821
rect 30098 13784 30104 13796
rect 29012 13756 29132 13784
rect 29472 13756 30104 13784
rect 26191 13753 26203 13756
rect 26145 13747 26203 13753
rect 15068 13688 17816 13716
rect 15068 13676 15074 13688
rect 18138 13676 18144 13728
rect 18196 13716 18202 13728
rect 19702 13716 19708 13728
rect 18196 13688 19708 13716
rect 18196 13676 18202 13688
rect 19702 13676 19708 13688
rect 19760 13676 19766 13728
rect 20254 13676 20260 13728
rect 20312 13725 20318 13728
rect 20312 13679 20321 13725
rect 20312 13676 20318 13679
rect 21174 13676 21180 13728
rect 21232 13716 21238 13728
rect 26234 13716 26240 13728
rect 21232 13688 26240 13716
rect 21232 13676 21238 13688
rect 26234 13676 26240 13688
rect 26292 13676 26298 13728
rect 26786 13676 26792 13728
rect 26844 13716 26850 13728
rect 27163 13719 27221 13725
rect 27163 13716 27175 13719
rect 26844 13688 27175 13716
rect 26844 13676 26850 13688
rect 27163 13685 27175 13688
rect 27209 13716 27221 13719
rect 27706 13716 27712 13728
rect 27209 13688 27712 13716
rect 27209 13685 27221 13688
rect 27163 13679 27221 13685
rect 27706 13676 27712 13688
rect 27764 13676 27770 13728
rect 28994 13676 29000 13728
rect 29052 13676 29058 13728
rect 29104 13716 29132 13756
rect 30098 13744 30104 13756
rect 30156 13784 30162 13796
rect 30156 13756 30604 13784
rect 30156 13744 30162 13756
rect 30576 13728 30604 13756
rect 30377 13719 30435 13725
rect 30377 13716 30389 13719
rect 29104 13688 30389 13716
rect 30377 13685 30389 13688
rect 30423 13685 30435 13719
rect 30377 13679 30435 13685
rect 30558 13676 30564 13728
rect 30616 13676 30622 13728
rect 552 13626 31072 13648
rect 552 13574 7988 13626
rect 8040 13574 8052 13626
rect 8104 13574 8116 13626
rect 8168 13574 8180 13626
rect 8232 13574 8244 13626
rect 8296 13574 15578 13626
rect 15630 13574 15642 13626
rect 15694 13574 15706 13626
rect 15758 13574 15770 13626
rect 15822 13574 15834 13626
rect 15886 13574 23168 13626
rect 23220 13574 23232 13626
rect 23284 13574 23296 13626
rect 23348 13574 23360 13626
rect 23412 13574 23424 13626
rect 23476 13574 30758 13626
rect 30810 13574 30822 13626
rect 30874 13574 30886 13626
rect 30938 13574 30950 13626
rect 31002 13574 31014 13626
rect 31066 13574 31072 13626
rect 552 13552 31072 13574
rect 3970 13472 3976 13524
rect 4028 13521 4034 13524
rect 4028 13512 4037 13521
rect 4028 13484 4073 13512
rect 4028 13475 4037 13484
rect 4028 13472 4034 13475
rect 5166 13472 5172 13524
rect 5224 13512 5230 13524
rect 5813 13515 5871 13521
rect 5813 13512 5825 13515
rect 5224 13484 5825 13512
rect 5224 13472 5230 13484
rect 5813 13481 5825 13484
rect 5859 13481 5871 13515
rect 5813 13475 5871 13481
rect 6181 13515 6239 13521
rect 6181 13481 6193 13515
rect 6227 13512 6239 13515
rect 7282 13512 7288 13524
rect 6227 13484 7288 13512
rect 6227 13481 6239 13484
rect 6181 13475 6239 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 8386 13472 8392 13524
rect 8444 13512 8450 13524
rect 8570 13512 8576 13524
rect 8444 13484 8576 13512
rect 8444 13472 8450 13484
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 8938 13472 8944 13524
rect 8996 13472 9002 13524
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 9401 13515 9459 13521
rect 9401 13512 9413 13515
rect 9180 13484 9413 13512
rect 9180 13472 9186 13484
rect 9401 13481 9413 13484
rect 9447 13481 9459 13515
rect 9401 13475 9459 13481
rect 9766 13472 9772 13524
rect 9824 13512 9830 13524
rect 9953 13515 10011 13521
rect 9953 13512 9965 13515
rect 9824 13484 9965 13512
rect 9824 13472 9830 13484
rect 9953 13481 9965 13484
rect 9999 13481 10011 13515
rect 9953 13475 10011 13481
rect 10318 13472 10324 13524
rect 10376 13512 10382 13524
rect 10965 13515 11023 13521
rect 10965 13512 10977 13515
rect 10376 13484 10977 13512
rect 10376 13472 10382 13484
rect 10965 13481 10977 13484
rect 11011 13481 11023 13515
rect 10965 13475 11023 13481
rect 11422 13472 11428 13524
rect 11480 13512 11486 13524
rect 12802 13512 12808 13524
rect 11480 13484 12808 13512
rect 11480 13472 11486 13484
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 12995 13515 13053 13521
rect 12995 13481 13007 13515
rect 13041 13512 13053 13515
rect 13630 13512 13636 13524
rect 13041 13484 13636 13512
rect 13041 13481 13053 13484
rect 12995 13475 13053 13481
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 15473 13515 15531 13521
rect 15473 13512 15485 13515
rect 15252 13484 15485 13512
rect 15252 13472 15258 13484
rect 15473 13481 15485 13484
rect 15519 13481 15531 13515
rect 15473 13475 15531 13481
rect 15749 13515 15807 13521
rect 15749 13481 15761 13515
rect 15795 13481 15807 13515
rect 15749 13475 15807 13481
rect 952 13416 1446 13444
rect 952 13388 980 13416
rect 934 13336 940 13388
rect 992 13336 998 13388
rect 1213 13379 1271 13385
rect 1213 13345 1225 13379
rect 1259 13345 1271 13379
rect 1418 13376 1446 13416
rect 6270 13404 6276 13456
rect 6328 13404 6334 13456
rect 6730 13444 6736 13456
rect 6656 13416 6736 13444
rect 2041 13379 2099 13385
rect 2041 13376 2053 13379
rect 1418 13348 2053 13376
rect 1213 13339 1271 13345
rect 2041 13345 2053 13348
rect 2087 13345 2099 13379
rect 2041 13339 2099 13345
rect 3421 13379 3479 13385
rect 3421 13345 3433 13379
rect 3467 13376 3479 13379
rect 5997 13379 6055 13385
rect 3467 13348 4019 13376
rect 3467 13345 3479 13348
rect 3421 13339 3479 13345
rect 842 13268 848 13320
rect 900 13308 906 13320
rect 1228 13308 1256 13339
rect 900 13280 1256 13308
rect 900 13268 906 13280
rect 1302 13268 1308 13320
rect 1360 13268 1366 13320
rect 1670 13317 1676 13320
rect 1632 13311 1676 13317
rect 1632 13277 1644 13311
rect 1632 13271 1676 13277
rect 1670 13268 1676 13271
rect 1728 13268 1734 13320
rect 1811 13313 1869 13319
rect 1811 13279 1823 13313
rect 1857 13308 1869 13313
rect 2222 13308 2228 13320
rect 1857 13280 2228 13308
rect 1857 13279 1869 13280
rect 1811 13273 1869 13279
rect 2222 13268 2228 13280
rect 2280 13268 2286 13320
rect 3991 13319 4019 13348
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 6288 13376 6316 13404
rect 6656 13385 6684 13416
rect 6730 13404 6736 13416
rect 6788 13404 6794 13456
rect 6822 13404 6828 13456
rect 6880 13404 6886 13456
rect 8849 13447 8907 13453
rect 8849 13413 8861 13447
rect 8895 13444 8907 13447
rect 9858 13444 9864 13456
rect 8895 13416 9864 13444
rect 8895 13413 8907 13416
rect 8849 13407 8907 13413
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 11514 13444 11520 13456
rect 10244 13416 11520 13444
rect 6365 13379 6423 13385
rect 6365 13376 6377 13379
rect 6043 13348 6377 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 6365 13345 6377 13348
rect 6411 13345 6423 13379
rect 6365 13339 6423 13345
rect 6641 13379 6699 13385
rect 6641 13345 6653 13379
rect 6687 13345 6699 13379
rect 6641 13339 6699 13345
rect 3513 13311 3571 13317
rect 3513 13308 3525 13311
rect 3436 13280 3525 13308
rect 3436 13184 3464 13280
rect 3513 13277 3525 13280
rect 3559 13277 3571 13311
rect 3513 13271 3571 13277
rect 3976 13313 4034 13319
rect 3976 13279 3988 13313
rect 4022 13279 4034 13313
rect 3976 13273 4034 13279
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13308 4307 13311
rect 5810 13308 5816 13320
rect 4295 13280 5816 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 6178 13268 6184 13320
rect 6236 13308 6242 13320
rect 6546 13308 6552 13320
rect 6236 13280 6552 13308
rect 6236 13268 6242 13280
rect 6546 13268 6552 13280
rect 6604 13308 6610 13320
rect 6733 13311 6791 13317
rect 6733 13308 6745 13311
rect 6604 13280 6745 13308
rect 6604 13268 6610 13280
rect 6733 13277 6745 13280
rect 6779 13277 6791 13311
rect 6840 13308 6868 13404
rect 9125 13379 9183 13385
rect 9125 13345 9137 13379
rect 9171 13345 9183 13379
rect 9125 13339 9183 13345
rect 6914 13308 6920 13320
rect 6840 13280 6920 13308
rect 6733 13271 6791 13277
rect 6914 13268 6920 13280
rect 6972 13308 6978 13320
rect 7060 13311 7118 13317
rect 7060 13308 7072 13311
rect 6972 13280 7072 13308
rect 6972 13268 6978 13280
rect 7060 13277 7072 13280
rect 7106 13277 7118 13311
rect 7060 13271 7118 13277
rect 7190 13268 7196 13320
rect 7248 13268 7254 13320
rect 7466 13268 7472 13320
rect 7524 13268 7530 13320
rect 4982 13200 4988 13252
rect 5040 13240 5046 13252
rect 9140 13240 9168 13339
rect 9214 13336 9220 13388
rect 9272 13336 9278 13388
rect 9306 13336 9312 13388
rect 9364 13336 9370 13388
rect 9398 13336 9404 13388
rect 9456 13376 9462 13388
rect 9769 13379 9827 13385
rect 9769 13376 9781 13379
rect 9456 13348 9781 13376
rect 9456 13336 9462 13348
rect 9769 13345 9781 13348
rect 9815 13376 9827 13379
rect 10244 13376 10272 13416
rect 11514 13404 11520 13416
rect 11572 13404 11578 13456
rect 11606 13404 11612 13456
rect 11664 13444 11670 13456
rect 11664 13416 11836 13444
rect 11664 13404 11670 13416
rect 9815 13348 10272 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 10318 13336 10324 13388
rect 10376 13336 10382 13388
rect 10502 13336 10508 13388
rect 10560 13376 10566 13388
rect 10597 13379 10655 13385
rect 10597 13376 10609 13379
rect 10560 13348 10609 13376
rect 10560 13336 10566 13348
rect 10597 13345 10609 13348
rect 10643 13376 10655 13379
rect 10686 13376 10692 13388
rect 10643 13348 10692 13376
rect 10643 13345 10655 13348
rect 10597 13339 10655 13345
rect 10686 13336 10692 13348
rect 10744 13336 10750 13388
rect 10962 13336 10968 13388
rect 11020 13376 11026 13388
rect 11808 13385 11836 13416
rect 15378 13404 15384 13456
rect 15436 13444 15442 13456
rect 15764 13444 15792 13475
rect 16022 13472 16028 13524
rect 16080 13472 16086 13524
rect 16574 13472 16580 13524
rect 16632 13472 16638 13524
rect 16761 13515 16819 13521
rect 16761 13481 16773 13515
rect 16807 13481 16819 13515
rect 16761 13475 16819 13481
rect 15436 13416 15792 13444
rect 16040 13444 16068 13472
rect 16776 13444 16804 13475
rect 17494 13472 17500 13524
rect 17552 13512 17558 13524
rect 17865 13515 17923 13521
rect 17865 13512 17877 13515
rect 17552 13484 17877 13512
rect 17552 13472 17558 13484
rect 17865 13481 17877 13484
rect 17911 13481 17923 13515
rect 17865 13475 17923 13481
rect 20622 13472 20628 13524
rect 20680 13472 20686 13524
rect 20806 13472 20812 13524
rect 20864 13472 20870 13524
rect 20901 13515 20959 13521
rect 20901 13481 20913 13515
rect 20947 13512 20959 13515
rect 21082 13512 21088 13524
rect 20947 13484 21088 13512
rect 20947 13481 20959 13484
rect 20901 13475 20959 13481
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 21637 13515 21695 13521
rect 21637 13481 21649 13515
rect 21683 13512 21695 13515
rect 22379 13515 22437 13521
rect 21683 13484 21864 13512
rect 21683 13481 21695 13484
rect 21637 13475 21695 13481
rect 20824 13444 20852 13472
rect 21836 13444 21864 13484
rect 22379 13481 22391 13515
rect 22425 13512 22437 13515
rect 23842 13512 23848 13524
rect 22425 13484 23848 13512
rect 22425 13481 22437 13484
rect 22379 13475 22437 13481
rect 23842 13472 23848 13484
rect 23900 13472 23906 13524
rect 24578 13472 24584 13524
rect 24636 13521 24642 13524
rect 24636 13512 24645 13521
rect 26418 13512 26424 13524
rect 24636 13484 26424 13512
rect 24636 13475 24645 13484
rect 24636 13472 24642 13475
rect 26418 13472 26424 13484
rect 26476 13512 26482 13524
rect 26887 13515 26945 13521
rect 26887 13512 26899 13515
rect 26476 13484 26899 13512
rect 26476 13472 26482 13484
rect 26887 13481 26899 13484
rect 26933 13512 26945 13515
rect 27798 13512 27804 13524
rect 26933 13484 27804 13512
rect 26933 13481 26945 13484
rect 26887 13475 26945 13481
rect 27798 13472 27804 13484
rect 27856 13472 27862 13524
rect 28994 13512 29000 13524
rect 27908 13484 29000 13512
rect 24029 13447 24087 13453
rect 16040 13416 16804 13444
rect 16960 13416 18460 13444
rect 20824 13416 21588 13444
rect 21836 13416 22048 13444
rect 15436 13404 15442 13416
rect 11149 13379 11207 13385
rect 11149 13376 11161 13379
rect 11020 13348 11161 13376
rect 11020 13336 11026 13348
rect 11149 13345 11161 13348
rect 11195 13345 11207 13379
rect 11149 13339 11207 13345
rect 11241 13379 11299 13385
rect 11241 13345 11253 13379
rect 11287 13345 11299 13379
rect 11241 13339 11299 13345
rect 11793 13379 11851 13385
rect 11793 13345 11805 13379
rect 11839 13345 11851 13379
rect 11793 13339 11851 13345
rect 9324 13308 9352 13336
rect 9493 13311 9551 13317
rect 9493 13308 9505 13311
rect 9324 13280 9505 13308
rect 9493 13277 9505 13280
rect 9539 13277 9551 13311
rect 11256 13308 11284 13339
rect 12066 13336 12072 13388
rect 12124 13336 12130 13388
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 14921 13379 14979 13385
rect 12216 13348 12664 13376
rect 12216 13336 12222 13348
rect 11422 13308 11428 13320
rect 9493 13271 9551 13277
rect 9646 13280 11428 13308
rect 9646 13240 9674 13280
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13308 11575 13311
rect 11882 13308 11888 13320
rect 11563 13280 11888 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 12526 13268 12532 13320
rect 12584 13268 12590 13320
rect 12636 13308 12664 13348
rect 14921 13345 14933 13379
rect 14967 13376 14979 13379
rect 15010 13376 15016 13388
rect 14967 13348 15016 13376
rect 14967 13345 14979 13348
rect 14921 13339 14979 13345
rect 15010 13336 15016 13348
rect 15068 13336 15074 13388
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 15933 13379 15991 13385
rect 15933 13345 15945 13379
rect 15979 13376 15991 13379
rect 16758 13376 16764 13388
rect 15979 13348 16764 13376
rect 15979 13345 15991 13348
rect 15933 13339 15991 13345
rect 12992 13311 13050 13317
rect 12992 13308 13004 13311
rect 12636 13280 13004 13308
rect 12992 13277 13004 13280
rect 13038 13277 13050 13311
rect 12992 13271 13050 13277
rect 13262 13268 13268 13320
rect 13320 13268 13326 13320
rect 14550 13268 14556 13320
rect 14608 13308 14614 13320
rect 15105 13311 15163 13317
rect 15105 13308 15117 13311
rect 14608 13280 15117 13308
rect 14608 13268 14614 13280
rect 15105 13277 15117 13280
rect 15151 13277 15163 13311
rect 15672 13308 15700 13339
rect 16758 13336 16764 13348
rect 16816 13336 16822 13388
rect 16960 13385 16988 13416
rect 16945 13379 17003 13385
rect 16945 13345 16957 13379
rect 16991 13345 17003 13379
rect 16945 13339 17003 13345
rect 17034 13336 17040 13388
rect 17092 13376 17098 13388
rect 17221 13379 17279 13385
rect 17221 13376 17233 13379
rect 17092 13348 17233 13376
rect 17092 13336 17098 13348
rect 17221 13345 17233 13348
rect 17267 13345 17279 13379
rect 17221 13339 17279 13345
rect 17678 13336 17684 13388
rect 17736 13376 17742 13388
rect 17773 13379 17831 13385
rect 17773 13376 17785 13379
rect 17736 13348 17785 13376
rect 17736 13336 17742 13348
rect 17773 13345 17785 13348
rect 17819 13345 17831 13379
rect 17773 13339 17831 13345
rect 18049 13379 18107 13385
rect 18049 13345 18061 13379
rect 18095 13376 18107 13379
rect 18138 13376 18144 13388
rect 18095 13348 18144 13376
rect 18095 13345 18107 13348
rect 18049 13339 18107 13345
rect 16574 13308 16580 13320
rect 15672 13280 16580 13308
rect 15105 13271 15163 13277
rect 16574 13268 16580 13280
rect 16632 13268 16638 13320
rect 18064 13308 18092 13339
rect 18138 13336 18144 13348
rect 18196 13336 18202 13388
rect 18432 13376 18460 13416
rect 20530 13376 20536 13388
rect 18432 13348 20536 13376
rect 20530 13336 20536 13348
rect 20588 13336 20594 13388
rect 20801 13379 20859 13385
rect 20801 13376 20813 13379
rect 20732 13348 20813 13376
rect 20732 13320 20760 13348
rect 20801 13345 20813 13348
rect 20847 13345 20859 13379
rect 20801 13339 20859 13345
rect 20898 13336 20904 13388
rect 20956 13376 20962 13388
rect 21560 13385 21588 13416
rect 21085 13379 21143 13385
rect 21085 13376 21097 13379
rect 20956 13348 21097 13376
rect 20956 13336 20962 13348
rect 21085 13345 21097 13348
rect 21131 13345 21143 13379
rect 21085 13339 21143 13345
rect 21545 13379 21603 13385
rect 21545 13345 21557 13379
rect 21591 13376 21603 13379
rect 21591 13348 21772 13376
rect 21591 13345 21603 13348
rect 21545 13339 21603 13345
rect 17512 13280 18092 13308
rect 5040 13212 6776 13240
rect 9140 13212 9674 13240
rect 5040 13200 5046 13212
rect 1029 13175 1087 13181
rect 1029 13141 1041 13175
rect 1075 13172 1087 13175
rect 1578 13172 1584 13184
rect 1075 13144 1584 13172
rect 1075 13141 1087 13144
rect 1029 13135 1087 13141
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 2222 13132 2228 13184
rect 2280 13172 2286 13184
rect 2498 13172 2504 13184
rect 2280 13144 2504 13172
rect 2280 13132 2286 13144
rect 2498 13132 2504 13144
rect 2556 13132 2562 13184
rect 3418 13132 3424 13184
rect 3476 13132 3482 13184
rect 3786 13132 3792 13184
rect 3844 13172 3850 13184
rect 5442 13172 5448 13184
rect 3844 13144 5448 13172
rect 3844 13132 3850 13144
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 5537 13175 5595 13181
rect 5537 13141 5549 13175
rect 5583 13172 5595 13175
rect 6362 13172 6368 13184
rect 5583 13144 6368 13172
rect 5583 13141 5595 13144
rect 5537 13135 5595 13141
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 6457 13175 6515 13181
rect 6457 13141 6469 13175
rect 6503 13172 6515 13175
rect 6638 13172 6644 13184
rect 6503 13144 6644 13172
rect 6503 13141 6515 13144
rect 6457 13135 6515 13141
rect 6638 13132 6644 13144
rect 6696 13132 6702 13184
rect 6748 13172 6776 13212
rect 9398 13172 9404 13184
rect 6748 13144 9404 13172
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 9490 13132 9496 13184
rect 9548 13172 9554 13184
rect 9646 13172 9674 13212
rect 10318 13200 10324 13252
rect 10376 13200 10382 13252
rect 10410 13200 10416 13252
rect 10468 13200 10474 13252
rect 10594 13200 10600 13252
rect 10652 13200 10658 13252
rect 11238 13200 11244 13252
rect 11296 13240 11302 13252
rect 11296 13212 12112 13240
rect 11296 13200 11302 13212
rect 9548 13144 9674 13172
rect 9548 13132 9554 13144
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 10042 13172 10048 13184
rect 9824 13144 10048 13172
rect 9824 13132 9830 13144
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 10134 13132 10140 13184
rect 10192 13132 10198 13184
rect 10336 13172 10364 13200
rect 10502 13172 10508 13184
rect 10336 13144 10508 13172
rect 10502 13132 10508 13144
rect 10560 13132 10566 13184
rect 10612 13172 10640 13200
rect 11425 13175 11483 13181
rect 11425 13172 11437 13175
rect 10612 13144 11437 13172
rect 11425 13141 11437 13144
rect 11471 13141 11483 13175
rect 11425 13135 11483 13141
rect 11974 13132 11980 13184
rect 12032 13132 12038 13184
rect 12084 13172 12112 13212
rect 14292 13212 15516 13240
rect 12802 13172 12808 13184
rect 12084 13144 12808 13172
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 13170 13132 13176 13184
rect 13228 13172 13234 13184
rect 14292 13172 14320 13212
rect 13228 13144 14320 13172
rect 13228 13132 13234 13144
rect 14366 13132 14372 13184
rect 14424 13132 14430 13184
rect 15488 13172 15516 13212
rect 17512 13172 17540 13280
rect 18322 13268 18328 13320
rect 18380 13268 18386 13320
rect 18690 13317 18696 13320
rect 18652 13311 18696 13317
rect 18652 13277 18664 13311
rect 18652 13271 18696 13277
rect 18690 13268 18696 13271
rect 18748 13268 18754 13320
rect 18782 13268 18788 13320
rect 18840 13268 18846 13320
rect 19061 13311 19119 13317
rect 19061 13277 19073 13311
rect 19107 13308 19119 13311
rect 19978 13308 19984 13320
rect 19107 13280 19984 13308
rect 19107 13277 19119 13280
rect 19061 13271 19119 13277
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 20990 13308 20996 13320
rect 20772 13280 20996 13308
rect 20772 13268 20778 13280
rect 20990 13268 20996 13280
rect 21048 13268 21054 13320
rect 17589 13243 17647 13249
rect 17589 13209 17601 13243
rect 17635 13240 17647 13243
rect 17862 13240 17868 13252
rect 17635 13212 17868 13240
rect 17635 13209 17647 13212
rect 17589 13203 17647 13209
rect 17862 13200 17868 13212
rect 17920 13200 17926 13252
rect 21100 13240 21128 13339
rect 21744 13252 21772 13348
rect 21818 13336 21824 13388
rect 21876 13336 21882 13388
rect 22020 13376 22048 13416
rect 24029 13413 24041 13447
rect 24075 13444 24087 13447
rect 24210 13444 24216 13456
rect 24075 13416 24216 13444
rect 24075 13413 24087 13416
rect 24029 13407 24087 13413
rect 24210 13404 24216 13416
rect 24268 13404 24274 13456
rect 26237 13447 26295 13453
rect 26237 13413 26249 13447
rect 26283 13444 26295 13447
rect 26326 13444 26332 13456
rect 26283 13416 26332 13444
rect 26283 13413 26295 13416
rect 26237 13407 26295 13413
rect 26326 13404 26332 13416
rect 26384 13404 26390 13456
rect 22649 13379 22707 13385
rect 22649 13376 22661 13379
rect 22020 13348 22661 13376
rect 22649 13345 22661 13348
rect 22695 13345 22707 13379
rect 22649 13339 22707 13345
rect 24118 13336 24124 13388
rect 24176 13336 24182 13388
rect 24857 13379 24915 13385
rect 24857 13345 24869 13379
rect 24903 13376 24915 13379
rect 25498 13376 25504 13388
rect 24903 13348 25504 13376
rect 24903 13345 24915 13348
rect 24857 13339 24915 13345
rect 25498 13336 25504 13348
rect 25556 13336 25562 13388
rect 26050 13336 26056 13388
rect 26108 13376 26114 13388
rect 27157 13379 27215 13385
rect 26108 13348 26740 13376
rect 26108 13336 26114 13348
rect 21913 13311 21971 13317
rect 21913 13277 21925 13311
rect 21959 13308 21971 13311
rect 22278 13308 22284 13320
rect 21959 13280 22284 13308
rect 21959 13277 21971 13280
rect 21913 13271 21971 13277
rect 22278 13268 22284 13280
rect 22336 13268 22342 13320
rect 22419 13311 22477 13317
rect 22419 13277 22431 13311
rect 22465 13308 22477 13311
rect 22554 13308 22560 13320
rect 22465 13280 22560 13308
rect 22465 13277 22477 13280
rect 22419 13271 22477 13277
rect 22554 13268 22560 13280
rect 22612 13268 22618 13320
rect 21542 13240 21548 13252
rect 20272 13212 20760 13240
rect 21100 13212 21548 13240
rect 15488 13144 17540 13172
rect 17678 13132 17684 13184
rect 17736 13172 17742 13184
rect 20272 13172 20300 13212
rect 17736 13144 20300 13172
rect 17736 13132 17742 13144
rect 20346 13132 20352 13184
rect 20404 13132 20410 13184
rect 20732 13172 20760 13212
rect 21542 13200 21548 13212
rect 21600 13200 21606 13252
rect 21726 13200 21732 13252
rect 21784 13200 21790 13252
rect 21266 13172 21272 13184
rect 20732 13144 21272 13172
rect 21266 13132 21272 13144
rect 21324 13132 21330 13184
rect 21361 13175 21419 13181
rect 21361 13141 21373 13175
rect 21407 13172 21419 13175
rect 21910 13172 21916 13184
rect 21407 13144 21916 13172
rect 21407 13141 21419 13144
rect 21361 13135 21419 13141
rect 21910 13132 21916 13144
rect 21968 13132 21974 13184
rect 22278 13132 22284 13184
rect 22336 13172 22342 13184
rect 23658 13172 23664 13184
rect 22336 13144 23664 13172
rect 22336 13132 22342 13144
rect 23658 13132 23664 13144
rect 23716 13132 23722 13184
rect 24136 13172 24164 13336
rect 24627 13311 24685 13317
rect 24627 13277 24639 13311
rect 24673 13308 24685 13311
rect 25314 13308 25320 13320
rect 24673 13280 25320 13308
rect 24673 13277 24685 13280
rect 24627 13271 24685 13277
rect 25314 13268 25320 13280
rect 25372 13268 25378 13320
rect 26421 13311 26479 13317
rect 26421 13308 26433 13311
rect 25516 13280 26433 13308
rect 25516 13172 25544 13280
rect 26421 13277 26433 13280
rect 26467 13308 26479 13311
rect 26602 13308 26608 13320
rect 26467 13280 26608 13308
rect 26467 13277 26479 13280
rect 26421 13271 26479 13277
rect 26602 13268 26608 13280
rect 26660 13268 26666 13320
rect 26712 13308 26740 13348
rect 27157 13345 27169 13379
rect 27203 13376 27215 13379
rect 27908 13376 27936 13484
rect 28994 13472 29000 13484
rect 29052 13472 29058 13524
rect 29362 13472 29368 13524
rect 29420 13512 29426 13524
rect 30377 13515 30435 13521
rect 30377 13512 30389 13515
rect 29420 13484 30389 13512
rect 29420 13472 29426 13484
rect 30377 13481 30389 13484
rect 30423 13481 30435 13515
rect 30377 13475 30435 13481
rect 27203 13348 27936 13376
rect 27203 13345 27215 13348
rect 27157 13339 27215 13345
rect 27982 13336 27988 13388
rect 28040 13376 28046 13388
rect 28905 13379 28963 13385
rect 28905 13376 28917 13379
rect 28040 13348 28917 13376
rect 28040 13336 28046 13348
rect 28905 13345 28917 13348
rect 28951 13345 28963 13379
rect 28905 13339 28963 13345
rect 29362 13336 29368 13388
rect 29420 13376 29426 13388
rect 29546 13376 29552 13388
rect 29420 13348 29552 13376
rect 29420 13336 29426 13348
rect 29546 13336 29552 13348
rect 29604 13336 29610 13388
rect 30561 13379 30619 13385
rect 30561 13345 30573 13379
rect 30607 13345 30619 13379
rect 30561 13339 30619 13345
rect 26884 13329 26942 13335
rect 26884 13308 26896 13329
rect 26712 13295 26896 13308
rect 26930 13295 26942 13329
rect 26712 13289 26942 13295
rect 28629 13311 28687 13317
rect 26712 13280 26924 13289
rect 28629 13277 28641 13311
rect 28675 13277 28687 13311
rect 28629 13271 28687 13277
rect 28258 13200 28264 13252
rect 28316 13200 28322 13252
rect 24136 13144 25544 13172
rect 25958 13132 25964 13184
rect 26016 13172 26022 13184
rect 28644 13172 28672 13271
rect 29086 13268 29092 13320
rect 29144 13308 29150 13320
rect 30576 13308 30604 13339
rect 29144 13280 30604 13308
rect 29144 13268 29150 13280
rect 26016 13144 28672 13172
rect 26016 13132 26022 13144
rect 28902 13132 28908 13184
rect 28960 13172 28966 13184
rect 30009 13175 30067 13181
rect 30009 13172 30021 13175
rect 28960 13144 30021 13172
rect 28960 13132 28966 13144
rect 30009 13141 30021 13144
rect 30055 13141 30067 13175
rect 30009 13135 30067 13141
rect 552 13082 30912 13104
rect 552 13030 4193 13082
rect 4245 13030 4257 13082
rect 4309 13030 4321 13082
rect 4373 13030 4385 13082
rect 4437 13030 4449 13082
rect 4501 13030 11783 13082
rect 11835 13030 11847 13082
rect 11899 13030 11911 13082
rect 11963 13030 11975 13082
rect 12027 13030 12039 13082
rect 12091 13030 19373 13082
rect 19425 13030 19437 13082
rect 19489 13030 19501 13082
rect 19553 13030 19565 13082
rect 19617 13030 19629 13082
rect 19681 13030 26963 13082
rect 27015 13030 27027 13082
rect 27079 13030 27091 13082
rect 27143 13030 27155 13082
rect 27207 13030 27219 13082
rect 27271 13030 30912 13082
rect 552 13008 30912 13030
rect 842 12928 848 12980
rect 900 12968 906 12980
rect 2961 12971 3019 12977
rect 900 12940 2774 12968
rect 900 12928 906 12940
rect 2746 12900 2774 12940
rect 2961 12937 2973 12971
rect 3007 12968 3019 12971
rect 4246 12968 4252 12980
rect 3007 12940 4252 12968
rect 3007 12937 3019 12940
rect 2961 12931 3019 12937
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 7190 12968 7196 12980
rect 5951 12940 7196 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 7466 12928 7472 12980
rect 7524 12968 7530 12980
rect 8757 12971 8815 12977
rect 8757 12968 8769 12971
rect 7524 12940 8769 12968
rect 7524 12928 7530 12940
rect 8757 12937 8769 12940
rect 8803 12937 8815 12971
rect 8757 12931 8815 12937
rect 8846 12928 8852 12980
rect 8904 12968 8910 12980
rect 9217 12971 9275 12977
rect 9217 12968 9229 12971
rect 8904 12940 9229 12968
rect 8904 12928 8910 12940
rect 9217 12937 9229 12940
rect 9263 12937 9275 12971
rect 12897 12971 12955 12977
rect 9217 12931 9275 12937
rect 9514 12940 12848 12968
rect 3605 12903 3663 12909
rect 2746 12872 3556 12900
rect 3050 12832 3056 12844
rect 1418 12817 3056 12832
rect 1418 12786 1445 12817
rect 1433 12783 1445 12786
rect 1479 12804 3056 12817
rect 1479 12783 1491 12804
rect 3050 12792 3056 12804
rect 3108 12832 3114 12844
rect 3421 12835 3479 12841
rect 3421 12832 3433 12835
rect 3108 12804 3433 12832
rect 3108 12792 3114 12804
rect 3421 12801 3433 12804
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 1433 12777 1491 12783
rect 937 12767 995 12773
rect 937 12733 949 12767
rect 983 12764 995 12767
rect 1302 12764 1308 12776
rect 983 12736 1308 12764
rect 983 12733 995 12736
rect 937 12727 995 12733
rect 1302 12724 1308 12736
rect 1360 12724 1366 12776
rect 1578 12724 1584 12776
rect 1636 12764 1642 12776
rect 1673 12767 1731 12773
rect 1673 12764 1685 12767
rect 1636 12736 1685 12764
rect 1636 12724 1642 12736
rect 1673 12733 1685 12736
rect 1719 12733 1731 12767
rect 3528 12764 3556 12872
rect 3605 12869 3617 12903
rect 3651 12869 3663 12903
rect 8573 12903 8631 12909
rect 8573 12900 8585 12903
rect 3605 12863 3663 12869
rect 7484 12872 8585 12900
rect 3620 12832 3648 12863
rect 3620 12804 4200 12832
rect 3786 12764 3792 12776
rect 3528 12736 3792 12764
rect 1673 12727 1731 12733
rect 3786 12724 3792 12736
rect 3844 12724 3850 12776
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12733 3939 12767
rect 4172 12764 4200 12804
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4344 12835 4402 12841
rect 4344 12832 4356 12835
rect 4304 12804 4356 12832
rect 4304 12792 4310 12804
rect 4344 12801 4356 12804
rect 4390 12801 4402 12835
rect 4344 12795 4402 12801
rect 5626 12792 5632 12844
rect 5684 12832 5690 12844
rect 6552 12835 6610 12841
rect 6552 12832 6564 12835
rect 5684 12804 6564 12832
rect 5684 12792 5690 12804
rect 6552 12801 6564 12804
rect 6598 12801 6610 12835
rect 6552 12795 6610 12801
rect 6730 12792 6736 12844
rect 6788 12832 6794 12844
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6788 12804 6837 12832
rect 6788 12792 6794 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 4617 12767 4675 12773
rect 4617 12764 4629 12767
rect 4172 12736 4629 12764
rect 3881 12727 3939 12733
rect 4617 12733 4629 12736
rect 4663 12733 4675 12767
rect 4617 12727 4675 12733
rect 6089 12767 6147 12773
rect 6089 12733 6101 12767
rect 6135 12764 6147 12767
rect 6178 12764 6184 12776
rect 6135 12736 6184 12764
rect 6135 12733 6147 12736
rect 6089 12727 6147 12733
rect 3418 12656 3424 12708
rect 3476 12696 3482 12708
rect 3896 12696 3924 12727
rect 6178 12724 6184 12736
rect 6236 12764 6242 12776
rect 6638 12764 6644 12776
rect 6236 12736 6644 12764
rect 6236 12724 6242 12736
rect 6638 12724 6644 12736
rect 6696 12724 6702 12776
rect 3476 12668 3924 12696
rect 3476 12656 3482 12668
rect 1403 12631 1461 12637
rect 1403 12597 1415 12631
rect 1449 12628 1461 12631
rect 1670 12628 1676 12640
rect 1449 12600 1676 12628
rect 1449 12597 1461 12600
rect 1403 12591 1461 12597
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 3970 12588 3976 12640
rect 4028 12628 4034 12640
rect 4347 12631 4405 12637
rect 4347 12628 4359 12631
rect 4028 12600 4359 12628
rect 4028 12588 4034 12600
rect 4347 12597 4359 12600
rect 4393 12597 4405 12631
rect 4347 12591 4405 12597
rect 6454 12588 6460 12640
rect 6512 12628 6518 12640
rect 6555 12631 6613 12637
rect 6555 12628 6567 12631
rect 6512 12600 6567 12628
rect 6512 12588 6518 12600
rect 6555 12597 6567 12600
rect 6601 12597 6613 12631
rect 6555 12591 6613 12597
rect 6730 12588 6736 12640
rect 6788 12628 6794 12640
rect 7484 12628 7512 12872
rect 8573 12869 8585 12872
rect 8619 12869 8631 12903
rect 9030 12900 9036 12912
rect 8573 12863 8631 12869
rect 8680 12872 9036 12900
rect 8389 12767 8447 12773
rect 8389 12733 8401 12767
rect 8435 12764 8447 12767
rect 8680 12764 8708 12872
rect 9030 12860 9036 12872
rect 9088 12860 9094 12912
rect 9306 12860 9312 12912
rect 9364 12860 9370 12912
rect 8754 12792 8760 12844
rect 8812 12792 8818 12844
rect 8435 12736 8708 12764
rect 8772 12764 8800 12792
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 8772 12736 8953 12764
rect 8435 12733 8447 12736
rect 8389 12727 8447 12733
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 9033 12767 9091 12773
rect 9033 12733 9045 12767
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 7834 12656 7840 12708
rect 7892 12696 7898 12708
rect 9048 12696 9076 12727
rect 9398 12724 9404 12776
rect 9456 12724 9462 12776
rect 9514 12773 9542 12940
rect 11238 12860 11244 12912
rect 11296 12900 11302 12912
rect 11977 12903 12035 12909
rect 11977 12900 11989 12903
rect 11296 12872 11989 12900
rect 11296 12860 11302 12872
rect 11977 12869 11989 12872
rect 12023 12869 12035 12903
rect 11977 12863 12035 12869
rect 9582 12792 9588 12844
rect 9640 12792 9646 12844
rect 9766 12792 9772 12844
rect 9824 12832 9830 12844
rect 9912 12835 9970 12841
rect 10134 12839 10140 12844
rect 9912 12832 9924 12835
rect 9824 12804 9924 12832
rect 9824 12792 9830 12804
rect 9912 12801 9924 12804
rect 9958 12801 9970 12835
rect 9912 12795 9970 12801
rect 10091 12833 10140 12839
rect 10091 12799 10103 12833
rect 10137 12799 10140 12833
rect 10091 12793 10140 12799
rect 10134 12792 10140 12793
rect 10192 12792 10198 12844
rect 10321 12835 10379 12841
rect 10321 12801 10333 12835
rect 10367 12832 10379 12835
rect 10410 12832 10416 12844
rect 10367 12804 10416 12832
rect 10367 12801 10379 12804
rect 10321 12795 10379 12801
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 10686 12792 10692 12844
rect 10744 12832 10750 12844
rect 11701 12835 11759 12841
rect 10744 12804 11376 12832
rect 10744 12792 10750 12804
rect 9493 12767 9551 12773
rect 9493 12733 9505 12767
rect 9539 12733 9551 12767
rect 11238 12764 11244 12776
rect 9493 12727 9551 12733
rect 9600 12736 11244 12764
rect 9214 12696 9220 12708
rect 7892 12668 8987 12696
rect 9048 12668 9220 12696
rect 7892 12656 7898 12668
rect 6788 12600 7512 12628
rect 8113 12631 8171 12637
rect 6788 12588 6794 12600
rect 8113 12597 8125 12631
rect 8159 12628 8171 12631
rect 8662 12628 8668 12640
rect 8159 12600 8668 12628
rect 8159 12597 8171 12600
rect 8113 12591 8171 12597
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 8959 12628 8987 12668
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 9416 12696 9444 12724
rect 9600 12696 9628 12736
rect 11238 12724 11244 12736
rect 11296 12724 11302 12776
rect 9416 12668 9628 12696
rect 11348 12696 11376 12804
rect 11701 12801 11713 12835
rect 11747 12832 11759 12835
rect 12618 12832 12624 12844
rect 11747 12804 12624 12832
rect 11747 12801 11759 12804
rect 11701 12795 11759 12801
rect 12618 12792 12624 12804
rect 12676 12792 12682 12844
rect 12820 12832 12848 12940
rect 12897 12937 12909 12971
rect 12943 12968 12955 12971
rect 13262 12968 13268 12980
rect 12943 12940 13268 12968
rect 12943 12937 12955 12940
rect 12897 12931 12955 12937
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 15102 12928 15108 12980
rect 15160 12968 15166 12980
rect 16482 12968 16488 12980
rect 15160 12940 16488 12968
rect 15160 12928 15166 12940
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 17586 12928 17592 12980
rect 17644 12928 17650 12980
rect 19794 12968 19800 12980
rect 18248 12940 19800 12968
rect 12986 12860 12992 12912
rect 13044 12900 13050 12912
rect 18248 12909 18276 12940
rect 19794 12928 19800 12940
rect 19852 12928 19858 12980
rect 22925 12971 22983 12977
rect 22925 12937 22937 12971
rect 22971 12968 22983 12971
rect 22971 12940 23888 12968
rect 22971 12937 22983 12940
rect 22925 12931 22983 12937
rect 18233 12903 18291 12909
rect 13044 12872 13400 12900
rect 13044 12860 13050 12872
rect 13372 12832 13400 12872
rect 18233 12869 18245 12903
rect 18279 12869 18291 12903
rect 18233 12863 18291 12869
rect 23109 12903 23167 12909
rect 23109 12869 23121 12903
rect 23155 12900 23167 12903
rect 23382 12900 23388 12912
rect 23155 12872 23388 12900
rect 23155 12869 23167 12872
rect 23109 12863 23167 12869
rect 23382 12860 23388 12872
rect 23440 12860 23446 12912
rect 23750 12900 23756 12912
rect 23584 12872 23756 12900
rect 13722 12832 13728 12844
rect 12820 12804 13124 12832
rect 11422 12724 11428 12776
rect 11480 12764 11486 12776
rect 11793 12767 11851 12773
rect 11793 12764 11805 12767
rect 11480 12736 11805 12764
rect 11480 12724 11486 12736
rect 11793 12733 11805 12736
rect 11839 12733 11851 12767
rect 11793 12727 11851 12733
rect 12250 12724 12256 12776
rect 12308 12724 12314 12776
rect 12802 12724 12808 12776
rect 12860 12724 12866 12776
rect 12986 12724 12992 12776
rect 13044 12764 13050 12776
rect 13096 12773 13124 12804
rect 13372 12804 13728 12832
rect 13372 12773 13400 12804
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 13814 12792 13820 12844
rect 13872 12832 13878 12844
rect 14004 12835 14062 12841
rect 14004 12832 14016 12835
rect 13872 12804 14016 12832
rect 13872 12792 13878 12804
rect 14004 12801 14016 12804
rect 14050 12801 14062 12835
rect 14004 12795 14062 12801
rect 16206 12792 16212 12844
rect 16264 12839 16270 12844
rect 16264 12833 16286 12839
rect 16274 12799 16286 12833
rect 16264 12793 16286 12799
rect 16264 12792 16270 12793
rect 18322 12792 18328 12844
rect 18380 12832 18386 12844
rect 18693 12835 18751 12841
rect 18693 12832 18705 12835
rect 18380 12804 18705 12832
rect 18380 12792 18386 12804
rect 18693 12801 18705 12804
rect 18739 12801 18751 12835
rect 18693 12795 18751 12801
rect 19058 12792 19064 12844
rect 19116 12832 19122 12844
rect 19156 12835 19214 12841
rect 19156 12832 19168 12835
rect 19116 12804 19168 12832
rect 19116 12792 19122 12804
rect 19156 12801 19168 12804
rect 19202 12801 19214 12835
rect 19156 12795 19214 12801
rect 19306 12804 19564 12832
rect 13081 12767 13139 12773
rect 13081 12764 13093 12767
rect 13044 12736 13093 12764
rect 13044 12724 13050 12736
rect 13081 12733 13093 12736
rect 13127 12733 13139 12767
rect 13081 12727 13139 12733
rect 13357 12767 13415 12773
rect 13357 12733 13369 12767
rect 13403 12733 13415 12767
rect 13357 12727 13415 12733
rect 13538 12724 13544 12776
rect 13596 12724 13602 12776
rect 14277 12767 14335 12773
rect 14277 12764 14289 12767
rect 13648 12736 14289 12764
rect 12345 12699 12403 12705
rect 12345 12696 12357 12699
rect 11348 12668 12357 12696
rect 12345 12665 12357 12668
rect 12391 12665 12403 12699
rect 13648 12696 13676 12736
rect 14277 12733 14289 12736
rect 14323 12733 14335 12767
rect 14277 12727 14335 12733
rect 14550 12724 14556 12776
rect 14608 12764 14614 12776
rect 15749 12767 15807 12773
rect 15749 12764 15761 12767
rect 14608 12736 15761 12764
rect 14608 12724 14614 12736
rect 15749 12733 15761 12736
rect 15795 12733 15807 12767
rect 16076 12767 16134 12773
rect 16076 12764 16088 12767
rect 15749 12727 15807 12733
rect 15856 12736 16088 12764
rect 12345 12659 12403 12665
rect 12636 12668 13676 12696
rect 10686 12628 10692 12640
rect 8959 12600 10692 12628
rect 10686 12588 10692 12600
rect 10744 12588 10750 12640
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 12636 12637 12664 12668
rect 15470 12656 15476 12708
rect 15528 12696 15534 12708
rect 15856 12696 15884 12736
rect 16076 12733 16088 12736
rect 16122 12733 16134 12767
rect 16076 12727 16134 12733
rect 16482 12724 16488 12776
rect 16540 12724 16546 12776
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 18417 12767 18475 12773
rect 16632 12736 18276 12764
rect 16632 12724 16638 12736
rect 15528 12668 15884 12696
rect 18248 12696 18276 12736
rect 18417 12733 18429 12767
rect 18463 12764 18475 12767
rect 19306 12764 19334 12804
rect 18463 12736 19334 12764
rect 18463 12733 18475 12736
rect 18417 12727 18475 12733
rect 18432 12696 18460 12727
rect 19426 12724 19432 12776
rect 19484 12724 19490 12776
rect 19536 12764 19564 12804
rect 20346 12792 20352 12844
rect 20404 12832 20410 12844
rect 21364 12835 21422 12841
rect 21364 12832 21376 12835
rect 20404 12804 21376 12832
rect 20404 12792 20410 12804
rect 21364 12801 21376 12804
rect 21410 12801 21422 12835
rect 21364 12795 21422 12801
rect 21542 12792 21548 12844
rect 21600 12832 21606 12844
rect 21600 12804 23336 12832
rect 21600 12792 21606 12804
rect 23308 12776 23336 12804
rect 20714 12764 20720 12776
rect 19536 12736 20720 12764
rect 20714 12724 20720 12736
rect 20772 12724 20778 12776
rect 20898 12724 20904 12776
rect 20956 12724 20962 12776
rect 21637 12767 21695 12773
rect 21637 12764 21649 12767
rect 21008 12736 21649 12764
rect 18248 12668 18460 12696
rect 15528 12656 15534 12668
rect 18690 12656 18696 12708
rect 18748 12656 18754 12708
rect 20622 12656 20628 12708
rect 20680 12696 20686 12708
rect 21008 12696 21036 12736
rect 21637 12733 21649 12736
rect 21683 12733 21695 12767
rect 21637 12727 21695 12733
rect 23290 12724 23296 12776
rect 23348 12724 23354 12776
rect 23584 12773 23612 12872
rect 23750 12860 23756 12872
rect 23808 12860 23814 12912
rect 23658 12792 23664 12844
rect 23716 12792 23722 12844
rect 23860 12832 23888 12940
rect 25682 12928 25688 12980
rect 25740 12928 25746 12980
rect 26878 12968 26884 12980
rect 26620 12940 26884 12968
rect 24026 12832 24032 12844
rect 23860 12804 24032 12832
rect 24026 12792 24032 12804
rect 24084 12792 24090 12844
rect 24210 12792 24216 12844
rect 24268 12832 24274 12844
rect 24308 12835 24366 12841
rect 24308 12832 24320 12835
rect 24268 12804 24320 12832
rect 24268 12792 24274 12804
rect 24308 12801 24320 12804
rect 24354 12801 24366 12835
rect 24308 12795 24366 12801
rect 26329 12835 26387 12841
rect 26329 12801 26341 12835
rect 26375 12832 26387 12835
rect 26418 12832 26424 12844
rect 26375 12804 26424 12832
rect 26375 12801 26387 12804
rect 26329 12795 26387 12801
rect 26418 12792 26424 12804
rect 26476 12792 26482 12844
rect 23569 12767 23627 12773
rect 23569 12733 23581 12767
rect 23615 12733 23627 12767
rect 23676 12764 23704 12792
rect 26620 12776 26648 12940
rect 26878 12928 26884 12940
rect 26936 12968 26942 12980
rect 27706 12968 27712 12980
rect 26936 12940 27712 12968
rect 26936 12928 26942 12940
rect 27706 12928 27712 12940
rect 27764 12928 27770 12980
rect 28442 12928 28448 12980
rect 28500 12928 28506 12980
rect 28810 12928 28816 12980
rect 28868 12968 28874 12980
rect 30285 12971 30343 12977
rect 30285 12968 30297 12971
rect 28868 12940 30297 12968
rect 28868 12928 28874 12940
rect 30285 12937 30297 12940
rect 30331 12937 30343 12971
rect 30285 12931 30343 12937
rect 30469 12971 30527 12977
rect 30469 12937 30481 12971
rect 30515 12968 30527 12971
rect 31294 12968 31300 12980
rect 30515 12940 31300 12968
rect 30515 12937 30527 12940
rect 30469 12931 30527 12937
rect 31294 12928 31300 12940
rect 31352 12928 31358 12980
rect 29549 12903 29607 12909
rect 29549 12869 29561 12903
rect 29595 12869 29607 12903
rect 30098 12900 30104 12912
rect 29549 12863 29607 12869
rect 29748 12872 30104 12900
rect 26786 12792 26792 12844
rect 26844 12832 26850 12844
rect 26932 12835 26990 12841
rect 26932 12832 26944 12835
rect 26844 12804 26944 12832
rect 26844 12792 26850 12804
rect 26932 12801 26944 12804
rect 26978 12801 26990 12835
rect 26932 12795 26990 12801
rect 27111 12835 27169 12841
rect 27111 12801 27123 12835
rect 27157 12832 27169 12835
rect 27341 12835 27399 12841
rect 27157 12804 27292 12832
rect 27157 12801 27169 12804
rect 27111 12795 27169 12801
rect 23845 12767 23903 12773
rect 23845 12764 23857 12767
rect 23676 12736 23857 12764
rect 23569 12727 23627 12733
rect 23845 12733 23857 12736
rect 23891 12733 23903 12767
rect 24581 12767 24639 12773
rect 24581 12764 24593 12767
rect 23845 12727 23903 12733
rect 23958 12736 24593 12764
rect 23958 12696 23986 12736
rect 24581 12733 24593 12736
rect 24627 12733 24639 12767
rect 24581 12727 24639 12733
rect 25406 12724 25412 12776
rect 25464 12764 25470 12776
rect 26053 12767 26111 12773
rect 26053 12764 26065 12767
rect 25464 12736 26065 12764
rect 25464 12724 25470 12736
rect 26053 12733 26065 12736
rect 26099 12764 26111 12767
rect 26142 12764 26148 12776
rect 26099 12736 26148 12764
rect 26099 12733 26111 12736
rect 26053 12727 26111 12733
rect 26142 12724 26148 12736
rect 26200 12724 26206 12776
rect 26602 12724 26608 12776
rect 26660 12724 26666 12776
rect 27264 12764 27292 12804
rect 27341 12801 27353 12835
rect 27387 12832 27399 12835
rect 29564 12832 29592 12863
rect 27387 12804 29592 12832
rect 27387 12801 27399 12804
rect 27341 12795 27399 12801
rect 27264 12736 28028 12764
rect 20680 12668 21036 12696
rect 23408 12668 23986 12696
rect 20680 12656 20686 12668
rect 12069 12631 12127 12637
rect 12069 12628 12081 12631
rect 11296 12600 12081 12628
rect 11296 12588 11302 12600
rect 12069 12597 12081 12600
rect 12115 12597 12127 12631
rect 12069 12591 12127 12597
rect 12621 12631 12679 12637
rect 12621 12597 12633 12631
rect 12667 12597 12679 12631
rect 12621 12591 12679 12597
rect 13170 12588 13176 12640
rect 13228 12588 13234 12640
rect 13630 12588 13636 12640
rect 13688 12628 13694 12640
rect 14007 12631 14065 12637
rect 14007 12628 14019 12631
rect 13688 12600 14019 12628
rect 13688 12588 13694 12600
rect 14007 12597 14019 12600
rect 14053 12597 14065 12631
rect 14007 12591 14065 12597
rect 14182 12588 14188 12640
rect 14240 12628 14246 12640
rect 15381 12631 15439 12637
rect 15381 12628 15393 12631
rect 14240 12600 15393 12628
rect 14240 12588 14246 12600
rect 15381 12597 15393 12600
rect 15427 12597 15439 12631
rect 18708 12628 18736 12656
rect 19150 12628 19156 12640
rect 19208 12637 19214 12640
rect 18708 12600 19156 12628
rect 15381 12591 15439 12597
rect 19150 12588 19156 12600
rect 19208 12591 19217 12637
rect 19208 12588 19214 12591
rect 20714 12588 20720 12640
rect 20772 12588 20778 12640
rect 21367 12631 21425 12637
rect 21367 12597 21379 12631
rect 21413 12628 21425 12631
rect 21634 12628 21640 12640
rect 21413 12600 21640 12628
rect 21413 12597 21425 12600
rect 21367 12591 21425 12597
rect 21634 12588 21640 12600
rect 21692 12588 21698 12640
rect 23408 12637 23436 12668
rect 28000 12640 28028 12736
rect 28994 12724 29000 12776
rect 29052 12764 29058 12776
rect 29748 12773 29776 12872
rect 30098 12860 30104 12872
rect 30156 12860 30162 12912
rect 29733 12767 29791 12773
rect 29733 12764 29745 12767
rect 29052 12736 29745 12764
rect 29052 12724 29058 12736
rect 29733 12733 29745 12736
rect 29779 12733 29791 12767
rect 29733 12727 29791 12733
rect 29822 12724 29828 12776
rect 29880 12724 29886 12776
rect 29914 12724 29920 12776
rect 29972 12764 29978 12776
rect 30101 12767 30159 12773
rect 30101 12764 30113 12767
rect 29972 12736 30113 12764
rect 29972 12724 29978 12736
rect 30101 12733 30113 12736
rect 30147 12733 30159 12767
rect 30101 12727 30159 12733
rect 30377 12767 30435 12773
rect 30377 12733 30389 12767
rect 30423 12733 30435 12767
rect 30377 12727 30435 12733
rect 28166 12656 28172 12708
rect 28224 12696 28230 12708
rect 29089 12699 29147 12705
rect 29089 12696 29101 12699
rect 28224 12668 29101 12696
rect 28224 12656 28230 12668
rect 29089 12665 29101 12668
rect 29135 12665 29147 12699
rect 29089 12659 29147 12665
rect 29546 12656 29552 12708
rect 29604 12696 29610 12708
rect 30392 12696 30420 12727
rect 29604 12668 30420 12696
rect 29604 12656 29610 12668
rect 23385 12631 23443 12637
rect 23385 12597 23397 12631
rect 23431 12597 23443 12631
rect 23385 12591 23443 12597
rect 24118 12588 24124 12640
rect 24176 12628 24182 12640
rect 24311 12631 24369 12637
rect 24311 12628 24323 12631
rect 24176 12600 24323 12628
rect 24176 12588 24182 12600
rect 24311 12597 24323 12600
rect 24357 12597 24369 12631
rect 24311 12591 24369 12597
rect 26326 12588 26332 12640
rect 26384 12628 26390 12640
rect 26694 12628 26700 12640
rect 26384 12600 26700 12628
rect 26384 12588 26390 12600
rect 26694 12588 26700 12600
rect 26752 12588 26758 12640
rect 27982 12588 27988 12640
rect 28040 12588 28046 12640
rect 28074 12588 28080 12640
rect 28132 12628 28138 12640
rect 29181 12631 29239 12637
rect 29181 12628 29193 12631
rect 28132 12600 29193 12628
rect 28132 12588 28138 12600
rect 29181 12597 29193 12600
rect 29227 12597 29239 12631
rect 29181 12591 29239 12597
rect 30006 12588 30012 12640
rect 30064 12588 30070 12640
rect 552 12538 31072 12560
rect 552 12486 7988 12538
rect 8040 12486 8052 12538
rect 8104 12486 8116 12538
rect 8168 12486 8180 12538
rect 8232 12486 8244 12538
rect 8296 12486 15578 12538
rect 15630 12486 15642 12538
rect 15694 12486 15706 12538
rect 15758 12486 15770 12538
rect 15822 12486 15834 12538
rect 15886 12486 23168 12538
rect 23220 12486 23232 12538
rect 23284 12486 23296 12538
rect 23348 12486 23360 12538
rect 23412 12486 23424 12538
rect 23476 12486 30758 12538
rect 30810 12486 30822 12538
rect 30874 12486 30886 12538
rect 30938 12486 30950 12538
rect 31002 12486 31014 12538
rect 31066 12486 31072 12538
rect 552 12464 31072 12486
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 1771 12427 1829 12433
rect 1771 12424 1783 12427
rect 1728 12396 1783 12424
rect 1728 12384 1734 12396
rect 1771 12393 1783 12396
rect 1817 12393 1829 12427
rect 1771 12387 1829 12393
rect 2682 12384 2688 12436
rect 2740 12424 2746 12436
rect 5537 12427 5595 12433
rect 2740 12396 5488 12424
rect 2740 12384 2746 12396
rect 3510 12356 3516 12368
rect 3344 12328 3516 12356
rect 1213 12291 1271 12297
rect 1213 12257 1225 12291
rect 1259 12288 1271 12291
rect 3344 12288 3372 12328
rect 3510 12316 3516 12328
rect 3568 12316 3574 12368
rect 5460 12356 5488 12396
rect 5537 12393 5549 12427
rect 5583 12424 5595 12427
rect 5626 12424 5632 12436
rect 5583 12396 5632 12424
rect 5583 12393 5595 12396
rect 5537 12387 5595 12393
rect 5626 12384 5632 12396
rect 5684 12384 5690 12436
rect 5810 12384 5816 12436
rect 5868 12384 5874 12436
rect 7926 12424 7932 12436
rect 6104 12396 7932 12424
rect 6104 12356 6132 12396
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 8481 12427 8539 12433
rect 8481 12393 8493 12427
rect 8527 12424 8539 12427
rect 10226 12424 10232 12436
rect 8527 12396 10232 12424
rect 8527 12393 8539 12396
rect 8481 12387 8539 12393
rect 10226 12384 10232 12396
rect 10284 12384 10290 12436
rect 10965 12427 11023 12433
rect 10965 12393 10977 12427
rect 11011 12393 11023 12427
rect 10965 12387 11023 12393
rect 11241 12427 11299 12433
rect 11241 12393 11253 12427
rect 11287 12393 11299 12427
rect 11241 12387 11299 12393
rect 6546 12356 6552 12368
rect 5460 12328 6132 12356
rect 6472 12328 6552 12356
rect 1259 12260 3372 12288
rect 3421 12291 3479 12297
rect 1259 12257 1271 12260
rect 1213 12251 1271 12257
rect 3421 12257 3433 12291
rect 3467 12288 3479 12291
rect 3840 12292 3898 12297
rect 3840 12291 3975 12292
rect 3467 12260 3743 12288
rect 3467 12257 3479 12260
rect 3421 12251 3479 12257
rect 1302 12180 1308 12232
rect 1360 12180 1366 12232
rect 1811 12225 1869 12231
rect 1811 12191 1823 12225
rect 1857 12220 1869 12225
rect 1946 12220 1952 12232
rect 1857 12192 1952 12220
rect 1857 12191 1869 12192
rect 1811 12185 1869 12191
rect 1946 12180 1952 12192
rect 2004 12180 2010 12232
rect 2038 12180 2044 12232
rect 2096 12180 2102 12232
rect 3513 12223 3571 12229
rect 3513 12220 3525 12223
rect 3436 12192 3525 12220
rect 3436 12164 3464 12192
rect 3513 12189 3525 12192
rect 3559 12189 3571 12223
rect 3715 12220 3743 12260
rect 3840 12257 3852 12291
rect 3886 12288 3975 12291
rect 3886 12264 4108 12288
rect 3886 12257 3898 12264
rect 3947 12260 4108 12264
rect 3840 12251 3898 12257
rect 4080 12232 4108 12260
rect 4154 12248 4160 12300
rect 4212 12288 4218 12300
rect 4249 12291 4307 12297
rect 4249 12288 4261 12291
rect 4212 12260 4261 12288
rect 4212 12248 4218 12260
rect 4249 12257 4261 12260
rect 4295 12257 4307 12291
rect 4249 12251 4307 12257
rect 5902 12248 5908 12300
rect 5960 12288 5966 12300
rect 6472 12297 6500 12328
rect 6546 12316 6552 12328
rect 6604 12316 6610 12368
rect 8662 12316 8668 12368
rect 8720 12316 8726 12368
rect 10686 12316 10692 12368
rect 10744 12356 10750 12368
rect 10980 12356 11008 12387
rect 11256 12356 11284 12387
rect 11698 12384 11704 12436
rect 11756 12424 11762 12436
rect 12069 12427 12127 12433
rect 12069 12424 12081 12427
rect 11756 12396 12081 12424
rect 11756 12384 11762 12396
rect 12069 12393 12081 12396
rect 12115 12393 12127 12427
rect 12069 12387 12127 12393
rect 12618 12384 12624 12436
rect 12676 12384 12682 12436
rect 13998 12384 14004 12436
rect 14056 12424 14062 12436
rect 15010 12424 15016 12436
rect 14056 12396 15016 12424
rect 14056 12384 14062 12396
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 16669 12427 16727 12433
rect 16669 12393 16681 12427
rect 16715 12424 16727 12427
rect 18969 12427 19027 12433
rect 16715 12396 17080 12424
rect 16715 12393 16727 12396
rect 16669 12387 16727 12393
rect 10744 12328 11008 12356
rect 11072 12328 11284 12356
rect 10744 12316 10750 12328
rect 6822 12297 6828 12300
rect 5997 12291 6055 12297
rect 5997 12288 6009 12291
rect 5960 12260 6009 12288
rect 5960 12248 5966 12260
rect 5997 12257 6009 12260
rect 6043 12288 6055 12291
rect 6365 12291 6423 12297
rect 6365 12288 6377 12291
rect 6043 12260 6377 12288
rect 6043 12257 6055 12260
rect 5997 12251 6055 12257
rect 6365 12257 6377 12260
rect 6411 12257 6423 12291
rect 6365 12251 6423 12257
rect 6457 12291 6515 12297
rect 6457 12257 6469 12291
rect 6503 12257 6515 12291
rect 6784 12291 6828 12297
rect 6784 12288 6796 12291
rect 6457 12251 6515 12257
rect 6567 12260 6796 12288
rect 3976 12225 4034 12231
rect 3976 12220 3988 12225
rect 3715 12192 3988 12220
rect 3513 12183 3571 12189
rect 3976 12191 3988 12192
rect 4022 12191 4034 12225
rect 3976 12185 4034 12191
rect 4062 12180 4068 12232
rect 4120 12180 4126 12232
rect 6567 12220 6595 12260
rect 6784 12257 6796 12260
rect 6784 12251 6828 12257
rect 6822 12248 6828 12251
rect 6880 12248 6886 12300
rect 8680 12288 8708 12316
rect 9030 12297 9036 12300
rect 8992 12291 9036 12297
rect 6932 12260 7103 12288
rect 8680 12260 8800 12288
rect 6932 12229 6960 12260
rect 7075 12232 7103 12260
rect 6472 12192 6595 12220
rect 6920 12223 6978 12229
rect 6472 12164 6500 12192
rect 6920 12189 6932 12223
rect 6966 12189 6978 12223
rect 7075 12192 7104 12232
rect 6920 12183 6978 12189
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 7190 12180 7196 12232
rect 7248 12180 7254 12232
rect 8662 12180 8668 12232
rect 8720 12180 8726 12232
rect 8772 12220 8800 12260
rect 8992 12257 9004 12291
rect 8992 12251 9036 12257
rect 9030 12248 9036 12251
rect 9088 12248 9094 12300
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 9401 12291 9459 12297
rect 9401 12288 9413 12291
rect 9364 12260 9413 12288
rect 9364 12248 9370 12260
rect 9401 12257 9413 12260
rect 9447 12257 9459 12291
rect 9401 12251 9459 12257
rect 9128 12223 9186 12229
rect 9128 12220 9140 12223
rect 8772 12192 9140 12220
rect 9128 12189 9140 12192
rect 9174 12189 9186 12223
rect 9128 12183 9186 12189
rect 10410 12180 10416 12232
rect 10468 12220 10474 12232
rect 11072 12220 11100 12328
rect 11330 12316 11336 12368
rect 11388 12356 11394 12368
rect 11388 12328 11744 12356
rect 11388 12316 11394 12328
rect 11146 12248 11152 12300
rect 11204 12248 11210 12300
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12288 11483 12291
rect 11514 12288 11520 12300
rect 11471 12260 11520 12288
rect 11471 12257 11483 12260
rect 11425 12251 11483 12257
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 11716 12297 11744 12328
rect 11790 12316 11796 12368
rect 11848 12356 11854 12368
rect 11848 12328 12020 12356
rect 11848 12316 11854 12328
rect 11992 12297 12020 12328
rect 12434 12316 12440 12368
rect 12492 12316 12498 12368
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12257 11759 12291
rect 11701 12251 11759 12257
rect 11977 12291 12035 12297
rect 11977 12257 11989 12291
rect 12023 12288 12035 12291
rect 12066 12288 12072 12300
rect 12023 12260 12072 12288
rect 12023 12257 12035 12260
rect 11977 12251 12035 12257
rect 12066 12248 12072 12260
rect 12124 12248 12130 12300
rect 12250 12248 12256 12300
rect 12308 12288 12314 12300
rect 12452 12288 12480 12316
rect 12308 12260 12480 12288
rect 12529 12291 12587 12297
rect 12308 12248 12314 12260
rect 12529 12257 12541 12291
rect 12575 12257 12587 12291
rect 12636 12288 12664 12384
rect 16758 12316 16764 12368
rect 16816 12316 16822 12368
rect 12636 12260 13127 12288
rect 12529 12251 12587 12257
rect 10468 12192 11100 12220
rect 11164 12220 11192 12248
rect 12544 12220 12572 12251
rect 11164 12192 12572 12220
rect 12621 12223 12679 12229
rect 10468 12180 10474 12192
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 3418 12112 3424 12164
rect 3476 12112 3482 12164
rect 6454 12112 6460 12164
rect 6512 12112 6518 12164
rect 10689 12155 10747 12161
rect 10689 12121 10701 12155
rect 10735 12152 10747 12155
rect 10778 12152 10784 12164
rect 10735 12124 10784 12152
rect 10735 12121 10747 12124
rect 10689 12115 10747 12121
rect 10778 12112 10784 12124
rect 10836 12112 10842 12164
rect 10962 12112 10968 12164
rect 11020 12152 11026 12164
rect 11020 12124 11744 12152
rect 11020 12112 11026 12124
rect 11716 12096 11744 12124
rect 11974 12112 11980 12164
rect 12032 12112 12038 12164
rect 1029 12087 1087 12093
rect 1029 12053 1041 12087
rect 1075 12084 1087 12087
rect 2038 12084 2044 12096
rect 1075 12056 2044 12084
rect 1075 12053 1087 12056
rect 1029 12047 1087 12053
rect 2038 12044 2044 12056
rect 2096 12044 2102 12096
rect 6181 12087 6239 12093
rect 6181 12053 6193 12087
rect 6227 12084 6239 12087
rect 7190 12084 7196 12096
rect 6227 12056 7196 12084
rect 6227 12053 6239 12056
rect 6181 12047 6239 12053
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 7558 12044 7564 12096
rect 7616 12084 7622 12096
rect 11517 12087 11575 12093
rect 11517 12084 11529 12087
rect 7616 12056 11529 12084
rect 7616 12044 7622 12056
rect 11517 12053 11529 12056
rect 11563 12053 11575 12087
rect 11517 12047 11575 12053
rect 11698 12044 11704 12096
rect 11756 12044 11762 12096
rect 11793 12087 11851 12093
rect 11793 12053 11805 12087
rect 11839 12084 11851 12087
rect 11992 12084 12020 12112
rect 11839 12056 12020 12084
rect 11839 12053 11851 12056
rect 11793 12047 11851 12053
rect 12342 12044 12348 12096
rect 12400 12044 12406 12096
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 12636 12084 12664 12183
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 13099 12231 13127 12260
rect 13262 12248 13268 12300
rect 13320 12288 13326 12300
rect 13357 12291 13415 12297
rect 13357 12288 13369 12291
rect 13320 12260 13369 12288
rect 13320 12248 13326 12260
rect 13357 12257 13369 12260
rect 13403 12257 13415 12291
rect 13357 12251 13415 12257
rect 13630 12248 13636 12300
rect 13688 12248 13694 12300
rect 13998 12248 14004 12300
rect 14056 12288 14062 12300
rect 14829 12291 14887 12297
rect 14829 12288 14841 12291
rect 14056 12260 14841 12288
rect 14056 12248 14062 12260
rect 14829 12257 14841 12260
rect 14875 12257 14887 12291
rect 16776 12288 16804 12316
rect 16853 12291 16911 12297
rect 16853 12288 16865 12291
rect 16776 12260 16865 12288
rect 14829 12251 14887 12257
rect 16853 12257 16865 12260
rect 16899 12257 16911 12291
rect 17052 12288 17080 12396
rect 18969 12393 18981 12427
rect 19015 12424 19027 12427
rect 19058 12424 19064 12436
rect 19015 12396 19064 12424
rect 19015 12393 19027 12396
rect 18969 12387 19027 12393
rect 19058 12384 19064 12396
rect 19116 12384 19122 12436
rect 19150 12384 19156 12436
rect 19208 12384 19214 12436
rect 19426 12384 19432 12436
rect 19484 12424 19490 12436
rect 19705 12427 19763 12433
rect 19705 12424 19717 12427
rect 19484 12396 19717 12424
rect 19484 12384 19490 12396
rect 19705 12393 19717 12396
rect 19751 12393 19763 12427
rect 19705 12387 19763 12393
rect 19978 12384 19984 12436
rect 20036 12384 20042 12436
rect 20530 12384 20536 12436
rect 20588 12384 20594 12436
rect 20622 12384 20628 12436
rect 20680 12384 20686 12436
rect 21266 12424 21272 12436
rect 20824 12396 21272 12424
rect 19168 12356 19196 12384
rect 20548 12356 20576 12384
rect 19168 12328 19288 12356
rect 17681 12291 17739 12297
rect 17681 12288 17693 12291
rect 17052 12260 17693 12288
rect 16853 12251 16911 12257
rect 17681 12257 17693 12260
rect 17727 12257 17739 12291
rect 17681 12251 17739 12257
rect 12948 12223 13006 12229
rect 12948 12220 12960 12223
rect 12860 12192 12960 12220
rect 12860 12180 12866 12192
rect 12948 12189 12960 12192
rect 12994 12189 13006 12223
rect 13099 12225 13158 12231
rect 13099 12194 13112 12225
rect 12948 12183 13006 12189
rect 13100 12191 13112 12194
rect 13146 12191 13158 12225
rect 13648 12220 13676 12248
rect 15013 12223 15071 12229
rect 15013 12220 15025 12223
rect 13648 12192 15025 12220
rect 13100 12185 13158 12191
rect 15013 12189 15025 12192
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 15657 12223 15715 12229
rect 15657 12189 15669 12223
rect 15703 12220 15715 12223
rect 16298 12220 16304 12232
rect 15703 12192 16304 12220
rect 15703 12189 15715 12192
rect 15657 12183 15715 12189
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 13538 12084 13544 12096
rect 12584 12056 13544 12084
rect 12584 12044 12590 12056
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 14458 12044 14464 12096
rect 14516 12044 14522 12096
rect 16868 12084 16896 12251
rect 19150 12248 19156 12300
rect 19208 12248 19214 12300
rect 16942 12180 16948 12232
rect 17000 12180 17006 12232
rect 17310 12229 17316 12232
rect 17272 12223 17316 12229
rect 17272 12189 17284 12223
rect 17272 12183 17316 12189
rect 17310 12180 17316 12183
rect 17368 12180 17374 12232
rect 17451 12223 17509 12229
rect 17451 12189 17463 12223
rect 17497 12220 17509 12223
rect 18046 12220 18052 12232
rect 17497 12192 18052 12220
rect 17497 12189 17509 12192
rect 17451 12183 17509 12189
rect 18046 12180 18052 12192
rect 18104 12180 18110 12232
rect 19260 12220 19288 12328
rect 19720 12328 20116 12356
rect 19720 12300 19748 12328
rect 19702 12248 19708 12300
rect 19760 12248 19766 12300
rect 19886 12248 19892 12300
rect 19944 12248 19950 12300
rect 19337 12223 19395 12229
rect 19337 12220 19349 12223
rect 19260 12192 19349 12220
rect 19150 12112 19156 12164
rect 19208 12152 19214 12164
rect 19260 12152 19288 12192
rect 19337 12189 19349 12192
rect 19383 12189 19395 12223
rect 19337 12183 19395 12189
rect 19208 12124 19288 12152
rect 19208 12112 19214 12124
rect 19904 12084 19932 12248
rect 20088 12220 20116 12328
rect 20180 12328 20576 12356
rect 20180 12297 20208 12328
rect 20824 12297 20852 12396
rect 21266 12384 21272 12396
rect 21324 12384 21330 12436
rect 22646 12384 22652 12436
rect 22704 12424 22710 12436
rect 23109 12427 23167 12433
rect 23109 12424 23121 12427
rect 22704 12396 23121 12424
rect 22704 12384 22710 12396
rect 23109 12393 23121 12396
rect 23155 12393 23167 12427
rect 24026 12424 24032 12436
rect 23109 12387 23167 12393
rect 23584 12396 24032 12424
rect 23584 12368 23612 12396
rect 24026 12384 24032 12396
rect 24084 12384 24090 12436
rect 24118 12384 24124 12436
rect 24176 12424 24182 12436
rect 24176 12396 24900 12424
rect 24176 12384 24182 12396
rect 21174 12356 21180 12368
rect 21100 12328 21180 12356
rect 21100 12297 21128 12328
rect 21174 12316 21180 12328
rect 21232 12316 21238 12368
rect 23566 12316 23572 12368
rect 23624 12316 23630 12368
rect 24872 12356 24900 12396
rect 25314 12384 25320 12436
rect 25372 12384 25378 12436
rect 26142 12384 26148 12436
rect 26200 12424 26206 12436
rect 26200 12396 27108 12424
rect 26200 12384 26206 12396
rect 25961 12359 26019 12365
rect 25961 12356 25973 12359
rect 24872 12328 25973 12356
rect 25961 12325 25973 12328
rect 26007 12356 26019 12359
rect 26786 12356 26792 12368
rect 26007 12328 26792 12356
rect 26007 12325 26019 12328
rect 25961 12319 26019 12325
rect 26786 12316 26792 12328
rect 26844 12316 26850 12368
rect 26878 12316 26884 12368
rect 26936 12316 26942 12368
rect 20165 12291 20223 12297
rect 20165 12257 20177 12291
rect 20211 12257 20223 12291
rect 20165 12251 20223 12257
rect 20533 12291 20591 12297
rect 20533 12257 20545 12291
rect 20579 12257 20591 12291
rect 20533 12251 20591 12257
rect 20809 12291 20867 12297
rect 20809 12257 20821 12291
rect 20855 12257 20867 12291
rect 20809 12251 20867 12257
rect 21085 12291 21143 12297
rect 21085 12257 21097 12291
rect 21131 12257 21143 12291
rect 21085 12251 21143 12257
rect 20548 12220 20576 12251
rect 21266 12248 21272 12300
rect 21324 12248 21330 12300
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 21376 12260 22017 12288
rect 21376 12220 21404 12260
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 24118 12248 24124 12300
rect 24176 12288 24182 12300
rect 24213 12291 24271 12297
rect 24213 12288 24225 12291
rect 24176 12260 24225 12288
rect 24176 12248 24182 12260
rect 24213 12257 24225 12260
rect 24259 12257 24271 12291
rect 24213 12251 24271 12257
rect 24302 12248 24308 12300
rect 24360 12288 24366 12300
rect 25685 12291 25743 12297
rect 24360 12260 25636 12288
rect 24360 12248 24366 12260
rect 21634 12229 21640 12232
rect 20088 12192 20576 12220
rect 21284 12192 21404 12220
rect 21596 12223 21640 12229
rect 20349 12155 20407 12161
rect 20349 12121 20361 12155
rect 20395 12152 20407 12155
rect 21284 12152 21312 12192
rect 21596 12189 21608 12223
rect 21596 12183 21640 12189
rect 21634 12180 21640 12183
rect 21692 12180 21698 12232
rect 21818 12229 21824 12232
rect 21775 12223 21824 12229
rect 21775 12189 21787 12223
rect 21821 12189 21824 12223
rect 21775 12183 21824 12189
rect 21818 12180 21824 12183
rect 21876 12180 21882 12232
rect 23477 12223 23535 12229
rect 23477 12189 23489 12223
rect 23523 12220 23535 12223
rect 23658 12220 23664 12232
rect 23523 12192 23664 12220
rect 23523 12189 23535 12192
rect 23477 12183 23535 12189
rect 23658 12180 23664 12192
rect 23716 12180 23722 12232
rect 23842 12229 23848 12232
rect 23804 12223 23848 12229
rect 23804 12189 23816 12223
rect 23804 12183 23848 12189
rect 23842 12180 23848 12183
rect 23900 12180 23906 12232
rect 23934 12180 23940 12232
rect 23992 12220 23998 12232
rect 25608 12220 25636 12260
rect 25685 12257 25697 12291
rect 25731 12288 25743 12291
rect 25774 12288 25780 12300
rect 25731 12260 25780 12288
rect 25731 12257 25743 12260
rect 25685 12251 25743 12257
rect 25774 12248 25780 12260
rect 25832 12288 25838 12300
rect 26142 12288 26148 12300
rect 25832 12260 26148 12288
rect 25832 12248 25838 12260
rect 26142 12248 26148 12260
rect 26200 12248 26206 12300
rect 26513 12291 26571 12297
rect 26513 12257 26525 12291
rect 26559 12288 26571 12291
rect 26602 12288 26608 12300
rect 26559 12260 26608 12288
rect 26559 12257 26571 12260
rect 26513 12251 26571 12257
rect 26528 12220 26556 12251
rect 26602 12248 26608 12260
rect 26660 12248 26666 12300
rect 26694 12248 26700 12300
rect 26752 12248 26758 12300
rect 27080 12297 27108 12396
rect 27154 12384 27160 12436
rect 27212 12424 27218 12436
rect 28543 12427 28601 12433
rect 28543 12424 28555 12427
rect 27212 12396 28555 12424
rect 27212 12384 27218 12396
rect 28543 12393 28555 12396
rect 28589 12393 28601 12427
rect 28543 12387 28601 12393
rect 29178 12384 29184 12436
rect 29236 12424 29242 12436
rect 29917 12427 29975 12433
rect 29917 12424 29929 12427
rect 29236 12396 29929 12424
rect 29236 12384 29242 12396
rect 29917 12393 29929 12396
rect 29963 12393 29975 12427
rect 29917 12387 29975 12393
rect 27065 12291 27123 12297
rect 27065 12257 27077 12291
rect 27111 12257 27123 12291
rect 27065 12251 27123 12257
rect 27525 12291 27583 12297
rect 27525 12257 27537 12291
rect 27571 12257 27583 12291
rect 27525 12251 27583 12257
rect 23992 12192 24037 12220
rect 25608 12192 26556 12220
rect 26712 12220 26740 12248
rect 27540 12220 27568 12251
rect 27706 12248 27712 12300
rect 27764 12288 27770 12300
rect 28074 12288 28080 12300
rect 27764 12260 28080 12288
rect 27764 12248 27770 12260
rect 28074 12248 28080 12260
rect 28132 12248 28138 12300
rect 28511 12260 28994 12288
rect 28511 12220 28539 12260
rect 28966 12232 28994 12260
rect 30374 12248 30380 12300
rect 30432 12248 30438 12300
rect 26712 12192 28539 12220
rect 28583 12223 28641 12229
rect 23992 12180 23998 12192
rect 28583 12189 28595 12223
rect 28629 12220 28641 12223
rect 28718 12220 28724 12232
rect 28629 12192 28724 12220
rect 28629 12189 28641 12192
rect 28583 12183 28641 12189
rect 28718 12180 28724 12192
rect 28776 12180 28782 12232
rect 28810 12180 28816 12232
rect 28868 12180 28874 12232
rect 28966 12192 29000 12232
rect 28994 12180 29000 12192
rect 29052 12180 29058 12232
rect 27709 12155 27767 12161
rect 27709 12152 27721 12155
rect 20395 12124 21312 12152
rect 24872 12124 27721 12152
rect 20395 12121 20407 12124
rect 20349 12115 20407 12121
rect 16868 12056 19932 12084
rect 20901 12087 20959 12093
rect 20901 12053 20913 12087
rect 20947 12084 20959 12087
rect 21542 12084 21548 12096
rect 20947 12056 21548 12084
rect 20947 12053 20959 12056
rect 20901 12047 20959 12053
rect 21542 12044 21548 12056
rect 21600 12044 21606 12096
rect 21726 12044 21732 12096
rect 21784 12084 21790 12096
rect 23014 12084 23020 12096
rect 21784 12056 23020 12084
rect 21784 12044 21790 12056
rect 23014 12044 23020 12056
rect 23072 12044 23078 12096
rect 23382 12044 23388 12096
rect 23440 12084 23446 12096
rect 24872 12084 24900 12124
rect 27709 12121 27721 12124
rect 27755 12121 27767 12155
rect 27709 12115 27767 12121
rect 23440 12056 24900 12084
rect 23440 12044 23446 12056
rect 25866 12044 25872 12096
rect 25924 12084 25930 12096
rect 27157 12087 27215 12093
rect 27157 12084 27169 12087
rect 25924 12056 27169 12084
rect 25924 12044 25930 12056
rect 27157 12053 27169 12056
rect 27203 12053 27215 12087
rect 27157 12047 27215 12053
rect 28350 12044 28356 12096
rect 28408 12084 28414 12096
rect 30561 12087 30619 12093
rect 30561 12084 30573 12087
rect 28408 12056 30573 12084
rect 28408 12044 28414 12056
rect 30561 12053 30573 12056
rect 30607 12053 30619 12087
rect 30561 12047 30619 12053
rect 552 11994 30912 12016
rect 552 11942 4193 11994
rect 4245 11942 4257 11994
rect 4309 11942 4321 11994
rect 4373 11942 4385 11994
rect 4437 11942 4449 11994
rect 4501 11942 11783 11994
rect 11835 11942 11847 11994
rect 11899 11942 11911 11994
rect 11963 11942 11975 11994
rect 12027 11942 12039 11994
rect 12091 11942 19373 11994
rect 19425 11942 19437 11994
rect 19489 11942 19501 11994
rect 19553 11942 19565 11994
rect 19617 11942 19629 11994
rect 19681 11942 26963 11994
rect 27015 11942 27027 11994
rect 27079 11942 27091 11994
rect 27143 11942 27155 11994
rect 27207 11942 27219 11994
rect 27271 11942 30912 11994
rect 552 11920 30912 11942
rect 1118 11880 1124 11892
rect 952 11852 1124 11880
rect 952 11753 980 11852
rect 1118 11840 1124 11852
rect 1176 11880 1182 11892
rect 1302 11880 1308 11892
rect 1176 11852 1308 11880
rect 1176 11840 1182 11852
rect 1302 11840 1308 11852
rect 1360 11840 1366 11892
rect 2961 11883 3019 11889
rect 2961 11849 2973 11883
rect 3007 11880 3019 11883
rect 3878 11880 3884 11892
rect 3007 11852 3884 11880
rect 3007 11849 3019 11852
rect 2961 11843 3019 11849
rect 3878 11840 3884 11852
rect 3936 11840 3942 11892
rect 5353 11883 5411 11889
rect 5353 11849 5365 11883
rect 5399 11880 5411 11883
rect 7006 11880 7012 11892
rect 5399 11852 7012 11880
rect 5399 11849 5411 11852
rect 5353 11843 5411 11849
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 7466 11840 7472 11892
rect 7524 11880 7530 11892
rect 7745 11883 7803 11889
rect 7745 11880 7757 11883
rect 7524 11852 7757 11880
rect 7524 11840 7530 11852
rect 7745 11849 7757 11852
rect 7791 11849 7803 11883
rect 7745 11843 7803 11849
rect 7926 11840 7932 11892
rect 7984 11880 7990 11892
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 7984 11852 8861 11880
rect 7984 11840 7990 11852
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 8849 11843 8907 11849
rect 9030 11840 9036 11892
rect 9088 11880 9094 11892
rect 9674 11880 9680 11892
rect 9088 11852 9680 11880
rect 9088 11840 9094 11852
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 11974 11840 11980 11892
rect 12032 11880 12038 11892
rect 12161 11883 12219 11889
rect 12161 11880 12173 11883
rect 12032 11852 12173 11880
rect 12032 11840 12038 11852
rect 12161 11849 12173 11852
rect 12207 11849 12219 11883
rect 12161 11843 12219 11849
rect 12986 11840 12992 11892
rect 13044 11880 13050 11892
rect 13265 11883 13323 11889
rect 13265 11880 13277 11883
rect 13044 11852 13277 11880
rect 13044 11840 13050 11852
rect 13265 11849 13277 11852
rect 13311 11880 13323 11883
rect 13354 11880 13360 11892
rect 13311 11852 13360 11880
rect 13311 11849 13323 11852
rect 13265 11843 13323 11849
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 14918 11840 14924 11892
rect 14976 11880 14982 11892
rect 18874 11880 18880 11892
rect 14976 11852 18880 11880
rect 14976 11840 14982 11852
rect 18874 11840 18880 11852
rect 18932 11840 18938 11892
rect 19058 11840 19064 11892
rect 19116 11880 19122 11892
rect 22925 11883 22983 11889
rect 19116 11852 22879 11880
rect 19116 11840 19122 11852
rect 7650 11772 7656 11824
rect 7708 11812 7714 11824
rect 8573 11815 8631 11821
rect 8573 11812 8585 11815
rect 7708 11784 8585 11812
rect 7708 11772 7714 11784
rect 8573 11781 8585 11784
rect 8619 11781 8631 11815
rect 8573 11775 8631 11781
rect 11517 11815 11575 11821
rect 11517 11781 11529 11815
rect 11563 11812 11575 11815
rect 22851 11812 22879 11852
rect 22925 11849 22937 11883
rect 22971 11880 22983 11883
rect 24210 11880 24216 11892
rect 22971 11852 24216 11880
rect 22971 11849 22983 11852
rect 22925 11843 22983 11849
rect 24210 11840 24216 11852
rect 24268 11840 24274 11892
rect 25961 11883 26019 11889
rect 25961 11849 25973 11883
rect 26007 11880 26019 11883
rect 26050 11880 26056 11892
rect 26007 11852 26056 11880
rect 26007 11849 26019 11852
rect 25961 11843 26019 11849
rect 26050 11840 26056 11852
rect 26108 11840 26114 11892
rect 26786 11880 26792 11892
rect 26160 11852 26792 11880
rect 11563 11784 13216 11812
rect 22851 11784 23336 11812
rect 11563 11781 11575 11784
rect 11517 11775 11575 11781
rect 1302 11753 1308 11756
rect 937 11747 995 11753
rect 937 11713 949 11747
rect 983 11713 995 11747
rect 937 11707 995 11713
rect 1264 11747 1308 11753
rect 1264 11713 1276 11747
rect 1264 11707 1308 11713
rect 1302 11704 1308 11707
rect 1360 11704 1366 11756
rect 1443 11747 1501 11753
rect 1443 11713 1455 11747
rect 1489 11744 1501 11747
rect 2498 11744 2504 11756
rect 1489 11716 2504 11744
rect 1489 11713 1501 11716
rect 1443 11707 1501 11713
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 3792 11747 3850 11753
rect 3792 11744 3804 11747
rect 3620 11716 3804 11744
rect 3620 11688 3648 11716
rect 3792 11713 3804 11716
rect 3838 11713 3850 11747
rect 3792 11707 3850 11713
rect 4356 11716 5764 11744
rect 4356 11688 4384 11716
rect 1673 11679 1731 11685
rect 1673 11676 1685 11679
rect 1044 11648 1685 11676
rect 1044 11540 1072 11648
rect 1673 11645 1685 11648
rect 1719 11645 1731 11679
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 1673 11639 1731 11645
rect 2746 11648 3341 11676
rect 1210 11540 1216 11552
rect 1044 11512 1216 11540
rect 1210 11500 1216 11512
rect 1268 11500 1274 11552
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 2746 11540 2774 11648
rect 3329 11645 3341 11648
rect 3375 11676 3387 11679
rect 3418 11676 3424 11688
rect 3375 11648 3424 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 3602 11636 3608 11688
rect 3660 11636 3666 11688
rect 4062 11636 4068 11688
rect 4120 11636 4126 11688
rect 4338 11636 4344 11688
rect 4396 11636 4402 11688
rect 5537 11679 5595 11685
rect 5537 11645 5549 11679
rect 5583 11676 5595 11679
rect 5626 11676 5632 11688
rect 5583 11648 5632 11676
rect 5583 11645 5595 11648
rect 5537 11639 5595 11645
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 5736 11676 5764 11716
rect 5810 11704 5816 11756
rect 5868 11744 5874 11756
rect 6000 11747 6058 11753
rect 6000 11744 6012 11747
rect 5868 11716 6012 11744
rect 5868 11704 5874 11716
rect 6000 11713 6012 11716
rect 6046 11713 6058 11747
rect 6000 11707 6058 11713
rect 6104 11716 6408 11744
rect 6104 11676 6132 11716
rect 5736 11648 6132 11676
rect 6178 11636 6184 11688
rect 6236 11676 6242 11688
rect 6273 11679 6331 11685
rect 6273 11676 6285 11679
rect 6236 11648 6285 11676
rect 6236 11636 6242 11648
rect 6273 11645 6285 11648
rect 6319 11645 6331 11679
rect 6380 11676 6408 11716
rect 7834 11704 7840 11756
rect 7892 11744 7898 11756
rect 8938 11744 8944 11756
rect 7892 11716 8248 11744
rect 7892 11704 7898 11716
rect 8220 11685 8248 11716
rect 8404 11716 8944 11744
rect 8404 11685 8432 11716
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 9677 11747 9735 11753
rect 9677 11744 9689 11747
rect 9640 11716 9689 11744
rect 9640 11704 9646 11716
rect 9677 11713 9689 11716
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 9858 11704 9864 11756
rect 9916 11744 9922 11756
rect 10140 11747 10198 11753
rect 10140 11744 10152 11747
rect 9916 11716 10152 11744
rect 9916 11704 9922 11716
rect 10140 11713 10152 11716
rect 10186 11713 10198 11747
rect 10140 11707 10198 11713
rect 10318 11704 10324 11756
rect 10376 11744 10382 11756
rect 10413 11747 10471 11753
rect 10413 11744 10425 11747
rect 10376 11716 10425 11744
rect 10376 11704 10382 11716
rect 10413 11713 10425 11716
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 10870 11704 10876 11756
rect 10928 11744 10934 11756
rect 12434 11744 12440 11756
rect 10928 11716 12440 11744
rect 10928 11704 10934 11716
rect 12434 11704 12440 11716
rect 12492 11704 12498 11756
rect 13078 11744 13084 11756
rect 12544 11716 13084 11744
rect 7929 11679 7987 11685
rect 7929 11676 7941 11679
rect 6380 11648 7941 11676
rect 6273 11639 6331 11645
rect 7929 11645 7941 11648
rect 7975 11645 7987 11679
rect 7929 11639 7987 11645
rect 8205 11679 8263 11685
rect 8205 11645 8217 11679
rect 8251 11645 8263 11679
rect 8205 11639 8263 11645
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11645 8447 11679
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 8389 11639 8447 11645
rect 8496 11648 8677 11676
rect 8496 11620 8524 11648
rect 8665 11645 8677 11648
rect 8711 11676 8723 11679
rect 9122 11676 9128 11688
rect 8711 11648 9128 11676
rect 8711 11645 8723 11648
rect 8665 11639 8723 11645
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11676 9275 11679
rect 9306 11676 9312 11688
rect 9263 11648 9312 11676
rect 9263 11645 9275 11648
rect 9217 11639 9275 11645
rect 9306 11636 9312 11648
rect 9364 11636 9370 11688
rect 11422 11676 11428 11688
rect 9646 11648 11428 11676
rect 7190 11568 7196 11620
rect 7248 11608 7254 11620
rect 7248 11580 8432 11608
rect 7248 11568 7254 11580
rect 1636 11512 2774 11540
rect 3795 11543 3853 11549
rect 1636 11500 1642 11512
rect 3795 11509 3807 11543
rect 3841 11540 3853 11543
rect 3970 11540 3976 11552
rect 3841 11512 3976 11540
rect 3841 11509 3853 11512
rect 3795 11503 3853 11509
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 6003 11543 6061 11549
rect 6003 11509 6015 11543
rect 6049 11540 6061 11543
rect 6546 11540 6552 11552
rect 6049 11512 6552 11540
rect 6049 11509 6061 11512
rect 6003 11503 6061 11509
rect 6546 11500 6552 11512
rect 6604 11500 6610 11552
rect 6914 11500 6920 11552
rect 6972 11540 6978 11552
rect 7377 11543 7435 11549
rect 7377 11540 7389 11543
rect 6972 11512 7389 11540
rect 6972 11500 6978 11512
rect 7377 11509 7389 11512
rect 7423 11509 7435 11543
rect 7377 11503 7435 11509
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 8021 11543 8079 11549
rect 8021 11540 8033 11543
rect 7892 11512 8033 11540
rect 7892 11500 7898 11512
rect 8021 11509 8033 11512
rect 8067 11509 8079 11543
rect 8404 11540 8432 11580
rect 8478 11568 8484 11620
rect 8536 11568 8542 11620
rect 9646 11608 9674 11648
rect 11422 11636 11428 11648
rect 11480 11636 11486 11688
rect 11514 11636 11520 11688
rect 11572 11676 11578 11688
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11572 11648 12081 11676
rect 11572 11636 11578 11648
rect 12069 11645 12081 11648
rect 12115 11676 12127 11679
rect 12250 11676 12256 11688
rect 12115 11648 12256 11676
rect 12115 11645 12127 11648
rect 12069 11639 12127 11645
rect 12250 11636 12256 11648
rect 12308 11636 12314 11688
rect 12544 11685 12572 11716
rect 13078 11704 13084 11716
rect 13136 11704 13142 11756
rect 13188 11744 13216 11784
rect 14004 11747 14062 11753
rect 14004 11744 14016 11747
rect 13188 11716 14016 11744
rect 14004 11713 14016 11716
rect 14050 11713 14062 11747
rect 14004 11707 14062 11713
rect 14090 11704 14096 11756
rect 14148 11744 14154 11756
rect 14148 11716 16804 11744
rect 14148 11704 14154 11716
rect 12345 11679 12403 11685
rect 12345 11645 12357 11679
rect 12391 11676 12403 11679
rect 12529 11679 12587 11685
rect 12529 11676 12541 11679
rect 12391 11648 12541 11676
rect 12391 11645 12403 11648
rect 12345 11639 12403 11645
rect 12529 11645 12541 11648
rect 12575 11645 12587 11679
rect 12989 11679 13047 11685
rect 12989 11676 13001 11679
rect 12529 11639 12587 11645
rect 12728 11648 13001 11676
rect 8680 11580 9674 11608
rect 8680 11540 8708 11580
rect 9766 11568 9772 11620
rect 9824 11568 9830 11620
rect 12728 11608 12756 11648
rect 12989 11645 13001 11648
rect 13035 11645 13047 11679
rect 12989 11639 13047 11645
rect 13096 11648 13492 11676
rect 13096 11608 13124 11648
rect 11348 11580 12756 11608
rect 12820 11580 13124 11608
rect 8404 11512 8708 11540
rect 8021 11503 8079 11509
rect 8754 11500 8760 11552
rect 8812 11540 8818 11552
rect 9122 11540 9128 11552
rect 8812 11512 9128 11540
rect 8812 11500 8818 11512
rect 9122 11500 9128 11512
rect 9180 11540 9186 11552
rect 9309 11543 9367 11549
rect 9309 11540 9321 11543
rect 9180 11512 9321 11540
rect 9180 11500 9186 11512
rect 9309 11509 9321 11512
rect 9355 11540 9367 11543
rect 9582 11540 9588 11552
rect 9355 11512 9588 11540
rect 9355 11509 9367 11512
rect 9309 11503 9367 11509
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 9784 11540 9812 11568
rect 10042 11540 10048 11552
rect 9784 11512 10048 11540
rect 10042 11500 10048 11512
rect 10100 11540 10106 11552
rect 10143 11543 10201 11549
rect 10143 11540 10155 11543
rect 10100 11512 10155 11540
rect 10100 11500 10106 11512
rect 10143 11509 10155 11512
rect 10189 11509 10201 11543
rect 10143 11503 10201 11509
rect 10502 11500 10508 11552
rect 10560 11540 10566 11552
rect 11348 11540 11376 11580
rect 10560 11512 11376 11540
rect 10560 11500 10566 11512
rect 11422 11500 11428 11552
rect 11480 11540 11486 11552
rect 11885 11543 11943 11549
rect 11885 11540 11897 11543
rect 11480 11512 11897 11540
rect 11480 11500 11486 11512
rect 11885 11509 11897 11512
rect 11931 11509 11943 11543
rect 11885 11503 11943 11509
rect 12618 11500 12624 11552
rect 12676 11500 12682 11552
rect 12820 11549 12848 11580
rect 13170 11568 13176 11620
rect 13228 11568 13234 11620
rect 13464 11608 13492 11648
rect 13538 11636 13544 11688
rect 13596 11636 13602 11688
rect 14277 11679 14335 11685
rect 14277 11676 14289 11679
rect 13648 11648 14289 11676
rect 13648 11608 13676 11648
rect 14277 11645 14289 11648
rect 14323 11645 14335 11679
rect 14277 11639 14335 11645
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11676 16451 11679
rect 16482 11676 16488 11688
rect 16439 11648 16488 11676
rect 16439 11645 16451 11648
rect 16393 11639 16451 11645
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 16776 11676 16804 11716
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 19058 11744 19064 11756
rect 16908 11716 16953 11744
rect 17052 11716 19064 11744
rect 16908 11704 16914 11716
rect 17052 11676 17080 11716
rect 19058 11704 19064 11716
rect 19116 11704 19122 11756
rect 19156 11745 19214 11751
rect 19156 11711 19168 11745
rect 19202 11711 19214 11745
rect 19156 11705 19214 11711
rect 19429 11747 19487 11753
rect 19429 11713 19441 11747
rect 19475 11744 19487 11747
rect 19794 11744 19800 11756
rect 19475 11716 19800 11744
rect 19475 11713 19487 11716
rect 19429 11707 19487 11713
rect 16776 11648 17080 11676
rect 17129 11679 17187 11685
rect 17129 11645 17141 11679
rect 17175 11676 17187 11679
rect 17586 11676 17592 11688
rect 17175 11648 17592 11676
rect 17175 11645 17187 11648
rect 17129 11639 17187 11645
rect 17586 11636 17592 11648
rect 17644 11636 17650 11688
rect 18322 11636 18328 11688
rect 18380 11676 18386 11688
rect 18693 11679 18751 11685
rect 18693 11676 18705 11679
rect 18380 11648 18705 11676
rect 18380 11636 18386 11648
rect 18693 11645 18705 11648
rect 18739 11645 18751 11679
rect 18693 11639 18751 11645
rect 18966 11636 18972 11688
rect 19024 11676 19030 11688
rect 19171 11676 19199 11705
rect 19794 11704 19800 11716
rect 19852 11704 19858 11756
rect 20714 11704 20720 11756
rect 20772 11744 20778 11756
rect 21364 11747 21422 11753
rect 21364 11744 21376 11747
rect 20772 11716 21376 11744
rect 20772 11704 20778 11716
rect 21364 11713 21376 11716
rect 21410 11713 21422 11747
rect 21364 11707 21422 11713
rect 21542 11704 21548 11756
rect 21600 11744 21606 11756
rect 21637 11747 21695 11753
rect 21637 11744 21649 11747
rect 21600 11716 21649 11744
rect 21600 11704 21606 11716
rect 21637 11713 21649 11716
rect 21683 11713 21695 11747
rect 21637 11707 21695 11713
rect 21818 11704 21824 11756
rect 21876 11704 21882 11756
rect 19024 11648 19199 11676
rect 19024 11636 19030 11648
rect 20898 11636 20904 11688
rect 20956 11636 20962 11688
rect 21836 11676 21864 11704
rect 23308 11688 23336 11784
rect 23382 11772 23388 11824
rect 23440 11772 23446 11824
rect 23477 11815 23535 11821
rect 23477 11781 23489 11815
rect 23523 11781 23535 11815
rect 23477 11775 23535 11781
rect 21008 11648 21864 11676
rect 13464 11580 13676 11608
rect 15010 11568 15016 11620
rect 15068 11608 15074 11620
rect 20809 11611 20867 11617
rect 15068 11580 16068 11608
rect 15068 11568 15074 11580
rect 12805 11543 12863 11549
rect 12805 11509 12817 11543
rect 12851 11509 12863 11543
rect 12805 11503 12863 11509
rect 12894 11500 12900 11552
rect 12952 11540 12958 11552
rect 13630 11540 13636 11552
rect 12952 11512 13636 11540
rect 12952 11500 12958 11512
rect 13630 11500 13636 11512
rect 13688 11540 13694 11552
rect 14007 11543 14065 11549
rect 14007 11540 14019 11543
rect 13688 11512 14019 11540
rect 13688 11500 13694 11512
rect 14007 11509 14019 11512
rect 14053 11509 14065 11543
rect 14007 11503 14065 11509
rect 14918 11500 14924 11552
rect 14976 11540 14982 11552
rect 16040 11549 16068 11580
rect 20809 11577 20821 11611
rect 20855 11608 20867 11611
rect 21008 11608 21036 11648
rect 23290 11636 23296 11688
rect 23348 11636 23354 11688
rect 23400 11685 23428 11772
rect 23492 11744 23520 11775
rect 23658 11772 23664 11824
rect 23716 11812 23722 11824
rect 23934 11812 23940 11824
rect 23716 11784 23940 11812
rect 23716 11772 23722 11784
rect 23934 11772 23940 11784
rect 23992 11772 23998 11824
rect 24486 11751 24492 11756
rect 24443 11745 24492 11751
rect 23492 11716 24399 11744
rect 23385 11679 23443 11685
rect 23385 11645 23397 11679
rect 23431 11645 23443 11679
rect 23385 11639 23443 11645
rect 23661 11679 23719 11685
rect 23661 11645 23673 11679
rect 23707 11676 23719 11679
rect 23707 11648 23796 11676
rect 23707 11645 23719 11648
rect 23661 11639 23719 11645
rect 23768 11620 23796 11648
rect 23934 11636 23940 11688
rect 23992 11636 23998 11688
rect 24264 11679 24322 11685
rect 24264 11676 24276 11679
rect 24044 11648 24276 11676
rect 23750 11608 23756 11620
rect 20855 11580 21036 11608
rect 22296 11580 23756 11608
rect 20855 11577 20867 11580
rect 20809 11571 20867 11577
rect 22296 11552 22324 11580
rect 23750 11568 23756 11580
rect 23808 11568 23814 11620
rect 23842 11568 23848 11620
rect 23900 11608 23906 11620
rect 24044 11608 24072 11648
rect 24264 11645 24276 11648
rect 24310 11645 24322 11679
rect 24371 11676 24399 11716
rect 24443 11711 24455 11745
rect 24489 11711 24492 11745
rect 24443 11705 24492 11711
rect 24486 11704 24492 11705
rect 24544 11704 24550 11756
rect 24673 11679 24731 11685
rect 24673 11676 24685 11679
rect 24371 11648 24685 11676
rect 24264 11639 24322 11645
rect 24673 11645 24685 11648
rect 24719 11645 24731 11679
rect 24673 11639 24731 11645
rect 25314 11636 25320 11688
rect 25372 11676 25378 11688
rect 26160 11685 26188 11852
rect 26786 11840 26792 11852
rect 26844 11840 26850 11892
rect 27522 11840 27528 11892
rect 27580 11840 27586 11892
rect 27982 11840 27988 11892
rect 28040 11840 28046 11892
rect 28629 11883 28687 11889
rect 28629 11849 28641 11883
rect 28675 11880 28687 11883
rect 28810 11880 28816 11892
rect 28675 11852 28816 11880
rect 28675 11849 28687 11852
rect 28629 11843 28687 11849
rect 28810 11840 28816 11852
rect 28868 11840 28874 11892
rect 29270 11840 29276 11892
rect 29328 11880 29334 11892
rect 29549 11883 29607 11889
rect 29549 11880 29561 11883
rect 29328 11852 29561 11880
rect 29328 11840 29334 11852
rect 29549 11849 29561 11852
rect 29595 11849 29607 11883
rect 29549 11843 29607 11849
rect 27540 11812 27568 11840
rect 28353 11815 28411 11821
rect 28353 11812 28365 11815
rect 27540 11784 28365 11812
rect 28353 11781 28365 11784
rect 28399 11781 28411 11815
rect 29730 11812 29736 11824
rect 28353 11775 28411 11781
rect 29288 11784 29736 11812
rect 29288 11756 29316 11784
rect 29730 11772 29736 11784
rect 29788 11772 29794 11824
rect 26694 11751 26700 11756
rect 26651 11745 26700 11751
rect 26651 11711 26663 11745
rect 26697 11711 26700 11745
rect 26651 11705 26700 11711
rect 26694 11704 26700 11705
rect 26752 11704 26758 11756
rect 29270 11744 29276 11756
rect 27172 11716 29276 11744
rect 27172 11688 27200 11716
rect 26145 11679 26203 11685
rect 26145 11676 26157 11679
rect 25372 11648 26157 11676
rect 25372 11636 25378 11648
rect 26145 11645 26157 11648
rect 26191 11645 26203 11679
rect 26881 11679 26939 11685
rect 26881 11676 26893 11679
rect 26145 11639 26203 11645
rect 26252 11648 26893 11676
rect 23900 11580 24072 11608
rect 23900 11568 23906 11580
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 14976 11512 15393 11540
rect 14976 11500 14982 11512
rect 15381 11509 15393 11512
rect 15427 11509 15439 11543
rect 15381 11503 15439 11509
rect 16025 11543 16083 11549
rect 16025 11509 16037 11543
rect 16071 11540 16083 11543
rect 16666 11540 16672 11552
rect 16071 11512 16672 11540
rect 16071 11509 16083 11512
rect 16025 11503 16083 11509
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 16859 11543 16917 11549
rect 16859 11509 16871 11543
rect 16905 11540 16917 11543
rect 17034 11540 17040 11552
rect 16905 11512 17040 11540
rect 16905 11509 16917 11512
rect 16859 11503 16917 11509
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 18414 11500 18420 11552
rect 18472 11500 18478 11552
rect 19150 11540 19156 11552
rect 19208 11549 19214 11552
rect 19117 11512 19156 11540
rect 19150 11500 19156 11512
rect 19208 11540 19217 11549
rect 21174 11540 21180 11552
rect 19208 11512 21180 11540
rect 19208 11503 19217 11512
rect 19208 11500 19214 11503
rect 21174 11500 21180 11512
rect 21232 11500 21238 11552
rect 21367 11543 21425 11549
rect 21367 11509 21379 11543
rect 21413 11540 21425 11543
rect 21634 11540 21640 11552
rect 21413 11512 21640 11540
rect 21413 11509 21425 11512
rect 21367 11503 21425 11509
rect 21634 11500 21640 11512
rect 21692 11540 21698 11552
rect 22094 11540 22100 11552
rect 21692 11512 22100 11540
rect 21692 11500 21698 11512
rect 22094 11500 22100 11512
rect 22152 11500 22158 11552
rect 22278 11500 22284 11552
rect 22336 11500 22342 11552
rect 23201 11543 23259 11549
rect 23201 11509 23213 11543
rect 23247 11540 23259 11543
rect 26252 11540 26280 11648
rect 26881 11645 26893 11648
rect 26927 11645 26939 11679
rect 26881 11639 26939 11645
rect 27154 11636 27160 11688
rect 27212 11636 27218 11688
rect 28828 11685 28856 11716
rect 29270 11704 29276 11716
rect 29328 11704 29334 11756
rect 28537 11679 28595 11685
rect 28537 11645 28549 11679
rect 28583 11645 28595 11679
rect 28537 11639 28595 11645
rect 28813 11679 28871 11685
rect 28813 11645 28825 11679
rect 28859 11676 28871 11679
rect 29733 11679 29791 11685
rect 28859 11648 28893 11676
rect 28859 11645 28871 11648
rect 28813 11639 28871 11645
rect 29733 11645 29745 11679
rect 29779 11676 29791 11679
rect 29779 11648 30144 11676
rect 29779 11645 29791 11648
rect 29733 11639 29791 11645
rect 23247 11512 26280 11540
rect 23247 11509 23259 11512
rect 23201 11503 23259 11509
rect 26602 11500 26608 11552
rect 26660 11549 26666 11552
rect 26660 11540 26669 11549
rect 28552 11540 28580 11639
rect 29089 11611 29147 11617
rect 29089 11577 29101 11611
rect 29135 11608 29147 11611
rect 29638 11608 29644 11620
rect 29135 11580 29644 11608
rect 29135 11577 29147 11580
rect 29089 11571 29147 11577
rect 29638 11568 29644 11580
rect 29696 11608 29702 11620
rect 29914 11608 29920 11620
rect 29696 11580 29920 11608
rect 29696 11568 29702 11580
rect 29914 11568 29920 11580
rect 29972 11568 29978 11620
rect 30116 11552 30144 11648
rect 29178 11540 29184 11552
rect 26660 11512 26705 11540
rect 28552 11512 29184 11540
rect 26660 11503 26669 11512
rect 26660 11500 26666 11503
rect 29178 11500 29184 11512
rect 29236 11500 29242 11552
rect 30098 11500 30104 11552
rect 30156 11500 30162 11552
rect 552 11450 31072 11472
rect 552 11398 7988 11450
rect 8040 11398 8052 11450
rect 8104 11398 8116 11450
rect 8168 11398 8180 11450
rect 8232 11398 8244 11450
rect 8296 11398 15578 11450
rect 15630 11398 15642 11450
rect 15694 11398 15706 11450
rect 15758 11398 15770 11450
rect 15822 11398 15834 11450
rect 15886 11398 23168 11450
rect 23220 11398 23232 11450
rect 23284 11398 23296 11450
rect 23348 11398 23360 11450
rect 23412 11398 23424 11450
rect 23476 11398 30758 11450
rect 30810 11398 30822 11450
rect 30874 11398 30886 11450
rect 30938 11398 30950 11450
rect 31002 11398 31014 11450
rect 31066 11398 31072 11450
rect 552 11376 31072 11398
rect 1118 11296 1124 11348
rect 1176 11296 1182 11348
rect 3513 11339 3571 11345
rect 3513 11305 3525 11339
rect 3559 11336 3571 11339
rect 3602 11336 3608 11348
rect 3559 11308 3608 11336
rect 3559 11305 3571 11308
rect 3513 11299 3571 11305
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4249 11339 4307 11345
rect 4249 11336 4261 11339
rect 4120 11308 4261 11336
rect 4120 11296 4126 11308
rect 4249 11305 4261 11308
rect 4295 11305 4307 11339
rect 4249 11299 4307 11305
rect 4522 11296 4528 11348
rect 4580 11336 4586 11348
rect 5077 11339 5135 11345
rect 5077 11336 5089 11339
rect 4580 11308 5089 11336
rect 4580 11296 4586 11308
rect 5077 11305 5089 11308
rect 5123 11305 5135 11339
rect 5077 11299 5135 11305
rect 5350 11296 5356 11348
rect 5408 11296 5414 11348
rect 5994 11296 6000 11348
rect 6052 11296 6058 11348
rect 6270 11296 6276 11348
rect 6328 11296 6334 11348
rect 8754 11336 8760 11348
rect 6472 11308 8760 11336
rect 1029 11271 1087 11277
rect 1029 11237 1041 11271
rect 1075 11268 1087 11271
rect 1578 11268 1584 11280
rect 1075 11240 1584 11268
rect 1075 11237 1087 11240
rect 1029 11231 1087 11237
rect 1578 11228 1584 11240
rect 1636 11228 1642 11280
rect 4338 11268 4344 11280
rect 3344 11240 4344 11268
rect 2225 11203 2283 11209
rect 2225 11200 2237 11203
rect 1044 11172 2237 11200
rect 1044 11144 1072 11172
rect 2225 11169 2237 11172
rect 2271 11169 2283 11203
rect 2225 11163 2283 11169
rect 1026 11092 1032 11144
rect 1084 11092 1090 11144
rect 1118 11092 1124 11144
rect 1176 11132 1182 11144
rect 1489 11135 1547 11141
rect 1489 11132 1501 11135
rect 1176 11104 1501 11132
rect 1176 11092 1182 11104
rect 1489 11101 1501 11104
rect 1535 11101 1547 11135
rect 1489 11095 1547 11101
rect 1670 11092 1676 11144
rect 1728 11132 1734 11144
rect 1816 11135 1874 11141
rect 1816 11132 1828 11135
rect 1728 11104 1828 11132
rect 1728 11092 1734 11104
rect 1816 11101 1828 11104
rect 1862 11101 1874 11135
rect 1816 11095 1874 11101
rect 1995 11137 2053 11143
rect 1995 11103 2007 11137
rect 2041 11132 2053 11137
rect 2958 11132 2964 11144
rect 2041 11104 2964 11132
rect 2041 11103 2053 11104
rect 1995 11097 2053 11103
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 658 11024 664 11076
rect 716 11024 722 11076
rect 676 10996 704 11024
rect 3344 10996 3372 11240
rect 4338 11228 4344 11240
rect 4396 11268 4402 11280
rect 6288 11268 6316 11296
rect 4396 11228 4430 11268
rect 3697 11203 3755 11209
rect 3697 11169 3709 11203
rect 3743 11200 3755 11203
rect 3786 11200 3792 11212
rect 3743 11172 3792 11200
rect 3743 11169 3755 11172
rect 3697 11163 3755 11169
rect 3786 11160 3792 11172
rect 3844 11160 3850 11212
rect 3970 11160 3976 11212
rect 4028 11160 4034 11212
rect 4402 11209 4430 11228
rect 5276 11240 6316 11268
rect 5276 11209 5304 11240
rect 4402 11203 4467 11209
rect 4402 11172 4421 11203
rect 4409 11169 4421 11172
rect 4455 11169 4467 11203
rect 4409 11163 4467 11169
rect 4617 11203 4675 11209
rect 4617 11169 4629 11203
rect 4663 11200 4675 11203
rect 5261 11203 5319 11209
rect 4663 11172 5212 11200
rect 4663 11169 4675 11172
rect 4617 11163 4675 11169
rect 3418 11092 3424 11144
rect 3476 11132 3482 11144
rect 4893 11135 4951 11141
rect 4893 11132 4905 11135
rect 3476 11104 4905 11132
rect 3476 11092 3482 11104
rect 4893 11101 4905 11104
rect 4939 11101 4951 11135
rect 5184 11132 5212 11172
rect 5261 11169 5273 11203
rect 5307 11169 5319 11203
rect 5261 11163 5319 11169
rect 5534 11160 5540 11212
rect 5592 11160 5598 11212
rect 6472 11209 6500 11308
rect 8754 11296 8760 11308
rect 8812 11336 8818 11348
rect 9214 11336 9220 11348
rect 8812 11308 9220 11336
rect 8812 11296 8818 11308
rect 9214 11296 9220 11308
rect 9272 11296 9278 11348
rect 9398 11296 9404 11348
rect 9456 11296 9462 11348
rect 9490 11296 9496 11348
rect 9548 11296 9554 11348
rect 9677 11339 9735 11345
rect 9677 11305 9689 11339
rect 9723 11336 9735 11339
rect 9950 11336 9956 11348
rect 9723 11308 9956 11336
rect 9723 11305 9735 11308
rect 9677 11299 9735 11305
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 10318 11296 10324 11348
rect 10376 11336 10382 11348
rect 10965 11339 11023 11345
rect 10965 11336 10977 11339
rect 10376 11308 10977 11336
rect 10376 11296 10382 11308
rect 10965 11305 10977 11308
rect 11011 11305 11023 11339
rect 10965 11299 11023 11305
rect 11330 11296 11336 11348
rect 11388 11296 11394 11348
rect 12158 11296 12164 11348
rect 12216 11336 12222 11348
rect 13170 11336 13176 11348
rect 12216 11308 13176 11336
rect 12216 11296 12222 11308
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 15470 11296 15476 11348
rect 15528 11336 15534 11348
rect 16298 11336 16304 11348
rect 15528 11308 16304 11336
rect 15528 11296 15534 11308
rect 16298 11296 16304 11308
rect 16356 11296 16362 11348
rect 16669 11339 16727 11345
rect 16669 11305 16681 11339
rect 16715 11336 16727 11339
rect 16715 11308 17080 11336
rect 16715 11305 16727 11308
rect 16669 11299 16727 11305
rect 6546 11228 6552 11280
rect 6604 11268 6610 11280
rect 6604 11240 6776 11268
rect 6604 11228 6610 11240
rect 6457 11203 6515 11209
rect 6457 11169 6469 11203
rect 6503 11169 6515 11203
rect 6457 11163 6515 11169
rect 6638 11160 6644 11212
rect 6696 11160 6702 11212
rect 6748 11200 6776 11240
rect 8570 11228 8576 11280
rect 8628 11228 8634 11280
rect 9508 11268 9536 11296
rect 10778 11268 10784 11280
rect 8864 11240 9536 11268
rect 6968 11203 7026 11209
rect 6968 11200 6980 11203
rect 6748 11172 6980 11200
rect 6968 11169 6980 11172
rect 7014 11169 7026 11203
rect 6968 11163 7026 11169
rect 7282 11160 7288 11212
rect 7340 11200 7346 11212
rect 7377 11203 7435 11209
rect 7377 11200 7389 11203
rect 7340 11172 7389 11200
rect 7340 11160 7346 11172
rect 7377 11169 7389 11172
rect 7423 11169 7435 11203
rect 7377 11163 7435 11169
rect 5626 11132 5632 11144
rect 5184 11104 5632 11132
rect 4893 11095 4951 11101
rect 5626 11092 5632 11104
rect 5684 11092 5690 11144
rect 5718 11092 5724 11144
rect 5776 11092 5782 11144
rect 6086 11092 6092 11144
rect 6144 11132 6150 11144
rect 7104 11135 7162 11141
rect 7104 11132 7116 11135
rect 6144 11104 7116 11132
rect 6144 11092 6150 11104
rect 7104 11101 7116 11104
rect 7150 11101 7162 11135
rect 8588 11132 8616 11228
rect 8864 11209 8892 11240
rect 8849 11203 8907 11209
rect 8849 11169 8861 11203
rect 8895 11169 8907 11203
rect 8849 11163 8907 11169
rect 8938 11160 8944 11212
rect 8996 11200 9002 11212
rect 9508 11209 9536 11240
rect 10244 11240 10784 11268
rect 10244 11212 10272 11240
rect 10778 11228 10784 11240
rect 10836 11268 10842 11280
rect 11348 11268 11376 11296
rect 10836 11240 11192 11268
rect 10836 11228 10842 11240
rect 9217 11203 9275 11209
rect 9217 11200 9229 11203
rect 8996 11172 9229 11200
rect 8996 11160 9002 11172
rect 9217 11169 9229 11172
rect 9263 11169 9275 11203
rect 9217 11163 9275 11169
rect 9493 11203 9551 11209
rect 9493 11169 9505 11203
rect 9539 11169 9551 11203
rect 9493 11163 9551 11169
rect 9769 11203 9827 11209
rect 9769 11169 9781 11203
rect 9815 11200 9827 11203
rect 10226 11200 10232 11212
rect 9815 11172 10232 11200
rect 9815 11169 9827 11172
rect 9769 11163 9827 11169
rect 10226 11160 10232 11172
rect 10284 11160 10290 11212
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 10502 11200 10508 11212
rect 10367 11172 10508 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 10502 11160 10508 11172
rect 10560 11160 10566 11212
rect 11164 11209 11192 11240
rect 11348 11240 11836 11268
rect 10597 11203 10655 11209
rect 10597 11169 10609 11203
rect 10643 11169 10655 11203
rect 10597 11163 10655 11169
rect 11149 11203 11207 11209
rect 11149 11169 11161 11203
rect 11195 11169 11207 11203
rect 11348 11200 11376 11240
rect 11425 11203 11483 11209
rect 11425 11200 11437 11203
rect 11348 11172 11437 11200
rect 11149 11163 11207 11169
rect 11425 11169 11437 11172
rect 11471 11169 11483 11203
rect 11425 11163 11483 11169
rect 8757 11135 8815 11141
rect 8588 11104 8708 11132
rect 7104 11095 7162 11101
rect 5736 11064 5764 11092
rect 6273 11067 6331 11073
rect 6273 11064 6285 11067
rect 5736 11036 6285 11064
rect 6273 11033 6285 11036
rect 6319 11033 6331 11067
rect 6273 11027 6331 11033
rect 8570 11024 8576 11076
rect 8628 11024 8634 11076
rect 8680 11064 8708 11104
rect 8757 11101 8769 11135
rect 8803 11132 8815 11135
rect 9858 11132 9864 11144
rect 8803 11104 9864 11132
rect 8803 11101 8815 11104
rect 8757 11095 8815 11101
rect 9858 11092 9864 11104
rect 9916 11092 9922 11144
rect 10612 11132 10640 11163
rect 11698 11160 11704 11212
rect 11756 11160 11762 11212
rect 11808 11209 11836 11240
rect 12250 11228 12256 11280
rect 12308 11228 12314 11280
rect 14826 11228 14832 11280
rect 14884 11228 14890 11280
rect 11793 11203 11851 11209
rect 11793 11169 11805 11203
rect 11839 11169 11851 11203
rect 11793 11163 11851 11169
rect 12802 11160 12808 11212
rect 12860 11209 12866 11212
rect 12860 11203 12914 11209
rect 12860 11169 12868 11203
rect 12902 11169 12914 11203
rect 12860 11163 12914 11169
rect 12860 11160 12866 11163
rect 13906 11160 13912 11212
rect 13964 11200 13970 11212
rect 15473 11203 15531 11209
rect 15473 11200 15485 11203
rect 13964 11172 15485 11200
rect 13964 11160 13970 11172
rect 15473 11169 15485 11172
rect 15519 11169 15531 11203
rect 15473 11163 15531 11169
rect 16574 11160 16580 11212
rect 16632 11160 16638 11212
rect 16853 11203 16911 11209
rect 16853 11169 16865 11203
rect 16899 11169 16911 11203
rect 16853 11163 16911 11169
rect 12434 11132 12440 11144
rect 9968 11104 10548 11132
rect 10612 11104 12440 11132
rect 9968 11064 9996 11104
rect 8680 11036 9996 11064
rect 10410 11024 10416 11076
rect 10468 11024 10474 11076
rect 10520 11064 10548 11104
rect 12434 11092 12440 11104
rect 12492 11092 12498 11144
rect 12526 11092 12532 11144
rect 12584 11092 12590 11144
rect 12986 11092 12992 11144
rect 13044 11092 13050 11144
rect 13262 11092 13268 11144
rect 13320 11092 13326 11144
rect 13446 11092 13452 11144
rect 13504 11132 13510 11144
rect 14642 11132 14648 11144
rect 13504 11104 14648 11132
rect 13504 11092 13510 11104
rect 14642 11092 14648 11104
rect 14700 11092 14706 11144
rect 15105 11135 15163 11141
rect 15105 11101 15117 11135
rect 15151 11132 15163 11135
rect 16868 11132 16896 11163
rect 16942 11160 16948 11212
rect 17000 11160 17006 11212
rect 17052 11200 17080 11308
rect 17218 11296 17224 11348
rect 17276 11336 17282 11348
rect 17276 11308 18368 11336
rect 17276 11296 17282 11308
rect 18340 11268 18368 11308
rect 18782 11296 18788 11348
rect 18840 11296 18846 11348
rect 19242 11296 19248 11348
rect 19300 11336 19306 11348
rect 21082 11336 21088 11348
rect 19300 11308 21088 11336
rect 19300 11296 19306 11308
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 21266 11296 21272 11348
rect 21324 11336 21330 11348
rect 21324 11308 22416 11336
rect 21324 11296 21330 11308
rect 21358 11268 21364 11280
rect 18340 11240 21364 11268
rect 21358 11228 21364 11240
rect 21416 11228 21422 11280
rect 22278 11268 22284 11280
rect 21468 11240 22284 11268
rect 17681 11203 17739 11209
rect 17681 11200 17693 11203
rect 17052 11172 17693 11200
rect 17681 11169 17693 11172
rect 17727 11169 17739 11203
rect 17681 11163 17739 11169
rect 18322 11160 18328 11212
rect 18380 11200 18386 11212
rect 19242 11200 19248 11212
rect 18380 11172 19248 11200
rect 18380 11160 18386 11172
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 19978 11160 19984 11212
rect 20036 11160 20042 11212
rect 20622 11160 20628 11212
rect 20680 11200 20686 11212
rect 21468 11209 21496 11240
rect 22278 11228 22284 11240
rect 22336 11228 22342 11280
rect 22388 11209 22416 11308
rect 22830 11296 22836 11348
rect 22888 11345 22894 11348
rect 22888 11336 22897 11345
rect 22888 11308 22933 11336
rect 22888 11299 22897 11308
rect 22888 11296 22894 11299
rect 24394 11296 24400 11348
rect 24452 11296 24458 11348
rect 24486 11296 24492 11348
rect 24544 11336 24550 11348
rect 29362 11336 29368 11348
rect 24544 11308 29368 11336
rect 24544 11296 24550 11308
rect 29362 11296 29368 11308
rect 29420 11296 29426 11348
rect 25314 11228 25320 11280
rect 25372 11228 25378 11280
rect 26234 11228 26240 11280
rect 26292 11268 26298 11280
rect 26292 11240 26562 11268
rect 26292 11228 26298 11240
rect 21453 11203 21511 11209
rect 21453 11200 21465 11203
rect 20680 11172 21465 11200
rect 20680 11160 20686 11172
rect 21453 11169 21465 11172
rect 21499 11169 21511 11203
rect 21453 11163 21511 11169
rect 22373 11203 22431 11209
rect 22373 11169 22385 11203
rect 22419 11200 22431 11203
rect 22462 11200 22468 11212
rect 22419 11172 22468 11200
rect 22419 11169 22431 11172
rect 22373 11163 22431 11169
rect 22462 11160 22468 11172
rect 22520 11160 22526 11212
rect 22922 11160 22928 11212
rect 22980 11200 22986 11212
rect 23109 11203 23167 11209
rect 23109 11200 23121 11203
rect 22980 11172 23121 11200
rect 22980 11160 22986 11172
rect 23109 11169 23121 11172
rect 23155 11169 23167 11203
rect 23109 11163 23167 11169
rect 23198 11160 23204 11212
rect 23256 11200 23262 11212
rect 24673 11203 24731 11209
rect 24673 11200 24685 11203
rect 23256 11172 24685 11200
rect 23256 11160 23262 11172
rect 24673 11169 24685 11172
rect 24719 11200 24731 11203
rect 24854 11200 24860 11212
rect 24719 11172 24860 11200
rect 24719 11169 24731 11172
rect 24673 11163 24731 11169
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 25225 11203 25283 11209
rect 25225 11169 25237 11203
rect 25271 11200 25283 11203
rect 25332 11200 25360 11228
rect 25271 11172 25360 11200
rect 25777 11203 25835 11209
rect 25271 11169 25283 11172
rect 25225 11163 25283 11169
rect 25777 11169 25789 11203
rect 25823 11200 25835 11203
rect 25866 11200 25872 11212
rect 25823 11172 25872 11200
rect 25823 11169 25835 11172
rect 25777 11163 25835 11169
rect 17126 11132 17132 11144
rect 15151 11104 15516 11132
rect 16868 11104 17132 11132
rect 15151 11101 15163 11104
rect 15105 11095 15163 11101
rect 10520 11036 11008 11064
rect 676 10968 3372 10996
rect 8588 10996 8616 11024
rect 9033 10999 9091 11005
rect 9033 10996 9045 10999
rect 8588 10968 9045 10996
rect 9033 10965 9045 10968
rect 9079 10965 9091 10999
rect 9033 10959 9091 10965
rect 9950 10956 9956 11008
rect 10008 10956 10014 11008
rect 10134 10956 10140 11008
rect 10192 10956 10198 11008
rect 10980 10996 11008 11036
rect 11054 11024 11060 11076
rect 11112 11064 11118 11076
rect 11241 11067 11299 11073
rect 11241 11064 11253 11067
rect 11112 11036 11253 11064
rect 11112 11024 11118 11036
rect 11241 11033 11253 11036
rect 11287 11033 11299 11067
rect 11517 11067 11575 11073
rect 11517 11064 11529 11067
rect 11241 11027 11299 11033
rect 11348 11036 11529 11064
rect 11348 10996 11376 11036
rect 11517 11033 11529 11036
rect 11563 11033 11575 11067
rect 11517 11027 11575 11033
rect 11977 11067 12035 11073
rect 11977 11033 11989 11067
rect 12023 11064 12035 11067
rect 12544 11064 12572 11092
rect 15488 11076 15516 11104
rect 17126 11092 17132 11104
rect 17184 11092 17190 11144
rect 17310 11141 17316 11144
rect 17272 11135 17316 11141
rect 17272 11101 17284 11135
rect 17272 11095 17316 11101
rect 17310 11092 17316 11095
rect 17368 11092 17374 11144
rect 17451 11135 17509 11141
rect 17451 11101 17463 11135
rect 17497 11132 17509 11135
rect 20530 11132 20536 11144
rect 17497 11104 20536 11132
rect 17497 11101 17509 11104
rect 17451 11095 17509 11101
rect 20530 11092 20536 11104
rect 20588 11092 20594 11144
rect 22836 11137 22894 11143
rect 22836 11103 22848 11137
rect 22882 11132 22894 11137
rect 23290 11132 23296 11144
rect 22882 11104 23296 11132
rect 22882 11103 22894 11104
rect 22836 11097 22894 11103
rect 23290 11092 23296 11104
rect 23348 11092 23354 11144
rect 23750 11092 23756 11144
rect 23808 11132 23814 11144
rect 24946 11132 24952 11144
rect 23808 11104 24952 11132
rect 23808 11092 23814 11104
rect 24946 11092 24952 11104
rect 25004 11092 25010 11144
rect 25498 11092 25504 11144
rect 25556 11132 25562 11144
rect 25792 11132 25820 11163
rect 25866 11160 25872 11172
rect 25924 11160 25930 11212
rect 26142 11160 26148 11212
rect 26200 11200 26206 11212
rect 26421 11203 26479 11209
rect 26421 11200 26433 11203
rect 26200 11172 26433 11200
rect 26200 11160 26206 11172
rect 26421 11169 26433 11172
rect 26467 11169 26479 11203
rect 26534 11200 26562 11240
rect 26534 11172 26791 11200
rect 26421 11163 26479 11169
rect 25556 11104 25820 11132
rect 26053 11135 26111 11141
rect 25556 11092 25562 11104
rect 26053 11101 26065 11135
rect 26099 11132 26111 11135
rect 26602 11132 26608 11144
rect 26099 11104 26608 11132
rect 26099 11101 26111 11104
rect 26053 11095 26111 11101
rect 12023 11036 12204 11064
rect 12023 11033 12035 11036
rect 11977 11027 12035 11033
rect 12176 11008 12204 11036
rect 12406 11036 12572 11064
rect 10980 10968 11376 10996
rect 12158 10956 12164 11008
rect 12216 10956 12222 11008
rect 12250 10956 12256 11008
rect 12308 10996 12314 11008
rect 12406 10996 12434 11036
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 15289 11067 15347 11073
rect 15289 11064 15301 11067
rect 14884 11036 15301 11064
rect 14884 11024 14890 11036
rect 15289 11033 15301 11036
rect 15335 11033 15347 11067
rect 15289 11027 15347 11033
rect 15470 11024 15476 11076
rect 15528 11024 15534 11076
rect 15746 11024 15752 11076
rect 15804 11024 15810 11076
rect 16393 11067 16451 11073
rect 16393 11033 16405 11067
rect 16439 11064 16451 11067
rect 16850 11064 16856 11076
rect 16439 11036 16856 11064
rect 16439 11033 16451 11036
rect 16393 11027 16451 11033
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 18414 11024 18420 11076
rect 18472 11064 18478 11076
rect 22370 11064 22376 11076
rect 18472 11036 22376 11064
rect 18472 11024 18478 11036
rect 22370 11024 22376 11036
rect 22428 11024 22434 11076
rect 26068 11064 26096 11095
rect 26602 11092 26608 11104
rect 26660 11092 26666 11144
rect 26763 11141 26791 11172
rect 26947 11172 27568 11200
rect 26947 11159 26975 11172
rect 26917 11153 26975 11159
rect 26748 11135 26806 11141
rect 26748 11101 26760 11135
rect 26794 11101 26806 11135
rect 26917 11119 26929 11153
rect 26963 11119 26975 11153
rect 27540 11144 27568 11172
rect 27890 11160 27896 11212
rect 27948 11200 27954 11212
rect 28442 11200 28448 11212
rect 27948 11172 28448 11200
rect 27948 11160 27954 11172
rect 28442 11160 28448 11172
rect 28500 11200 28506 11212
rect 28629 11203 28687 11209
rect 28629 11200 28641 11203
rect 28500 11172 28641 11200
rect 28500 11160 28506 11172
rect 28629 11169 28641 11172
rect 28675 11169 28687 11203
rect 28629 11163 28687 11169
rect 28902 11160 28908 11212
rect 28960 11160 28966 11212
rect 26917 11113 26975 11119
rect 27157 11135 27215 11141
rect 26748 11095 26806 11101
rect 27157 11101 27169 11135
rect 27203 11132 27215 11135
rect 27338 11132 27344 11144
rect 27203 11104 27344 11132
rect 27203 11101 27215 11104
rect 27157 11095 27215 11101
rect 27338 11092 27344 11104
rect 27396 11092 27402 11144
rect 27522 11092 27528 11144
rect 27580 11092 27586 11144
rect 23768 11036 26096 11064
rect 12308 10968 12434 10996
rect 12308 10956 12314 10968
rect 14366 10956 14372 11008
rect 14424 10956 14430 11008
rect 16942 10956 16948 11008
rect 17000 10996 17006 11008
rect 19521 10999 19579 11005
rect 19521 10996 19533 10999
rect 17000 10968 19533 10996
rect 17000 10956 17006 10968
rect 19521 10965 19533 10968
rect 19567 10996 19579 10999
rect 19978 10996 19984 11008
rect 19567 10968 19984 10996
rect 19567 10965 19579 10968
rect 19521 10959 19579 10965
rect 19978 10956 19984 10968
rect 20036 10956 20042 11008
rect 21269 10999 21327 11005
rect 21269 10965 21281 10999
rect 21315 10996 21327 10999
rect 22002 10996 22008 11008
rect 21315 10968 22008 10996
rect 21315 10965 21327 10968
rect 21269 10959 21327 10965
rect 22002 10956 22008 10968
rect 22060 10956 22066 11008
rect 22094 10956 22100 11008
rect 22152 10996 22158 11008
rect 22738 10996 22744 11008
rect 22152 10968 22744 10996
rect 22152 10956 22158 10968
rect 22738 10956 22744 10968
rect 22796 10996 22802 11008
rect 23768 10996 23796 11036
rect 28074 11024 28080 11076
rect 28132 11064 28138 11076
rect 28261 11067 28319 11073
rect 28261 11064 28273 11067
rect 28132 11036 28273 11064
rect 28132 11024 28138 11036
rect 28261 11033 28273 11036
rect 28307 11033 28319 11067
rect 28261 11027 28319 11033
rect 30006 11024 30012 11076
rect 30064 11024 30070 11076
rect 22796 10968 23796 10996
rect 24857 10999 24915 11005
rect 22796 10956 22802 10968
rect 24857 10965 24869 10999
rect 24903 10996 24915 10999
rect 24946 10996 24952 11008
rect 24903 10968 24952 10996
rect 24903 10965 24915 10968
rect 24857 10959 24915 10965
rect 24946 10956 24952 10968
rect 25004 10956 25010 11008
rect 25314 10956 25320 11008
rect 25372 10956 25378 11008
rect 552 10906 30912 10928
rect 552 10854 4193 10906
rect 4245 10854 4257 10906
rect 4309 10854 4321 10906
rect 4373 10854 4385 10906
rect 4437 10854 4449 10906
rect 4501 10854 11783 10906
rect 11835 10854 11847 10906
rect 11899 10854 11911 10906
rect 11963 10854 11975 10906
rect 12027 10854 12039 10906
rect 12091 10854 19373 10906
rect 19425 10854 19437 10906
rect 19489 10854 19501 10906
rect 19553 10854 19565 10906
rect 19617 10854 19629 10906
rect 19681 10854 26963 10906
rect 27015 10854 27027 10906
rect 27079 10854 27091 10906
rect 27143 10854 27155 10906
rect 27207 10854 27219 10906
rect 27271 10854 30912 10906
rect 552 10832 30912 10854
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10792 5319 10795
rect 5810 10792 5816 10804
rect 5307 10764 5816 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 6086 10752 6092 10804
rect 6144 10792 6150 10804
rect 6638 10792 6644 10804
rect 6144 10764 6644 10792
rect 6144 10752 6150 10764
rect 6638 10752 6644 10764
rect 6696 10792 6702 10804
rect 7929 10795 7987 10801
rect 7929 10792 7941 10795
rect 6696 10764 7941 10792
rect 6696 10752 6702 10764
rect 7929 10761 7941 10764
rect 7975 10761 7987 10795
rect 11609 10795 11667 10801
rect 7929 10755 7987 10761
rect 8404 10764 11560 10792
rect 937 10659 995 10665
rect 937 10625 949 10659
rect 983 10656 995 10659
rect 1118 10656 1124 10668
rect 983 10628 1124 10656
rect 983 10625 995 10628
rect 937 10619 995 10625
rect 1118 10616 1124 10628
rect 1176 10616 1182 10668
rect 1443 10659 1501 10665
rect 1443 10625 1455 10659
rect 1489 10656 1501 10659
rect 2130 10656 2136 10668
rect 1489 10628 2136 10656
rect 1489 10625 1501 10628
rect 1443 10619 1501 10625
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3700 10659 3758 10665
rect 3700 10656 3712 10659
rect 3099 10628 3712 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3700 10625 3712 10628
rect 3746 10625 3758 10659
rect 3700 10619 3758 10625
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 6000 10659 6058 10665
rect 6000 10656 6012 10659
rect 5500 10628 6012 10656
rect 5500 10616 5506 10628
rect 6000 10625 6012 10628
rect 6046 10625 6058 10659
rect 6000 10619 6058 10625
rect 6196 10628 6592 10656
rect 1578 10548 1584 10600
rect 1636 10588 1642 10600
rect 1673 10591 1731 10597
rect 1673 10588 1685 10591
rect 1636 10560 1685 10588
rect 1636 10548 1642 10560
rect 1673 10557 1685 10560
rect 1719 10557 1731 10591
rect 1673 10551 1731 10557
rect 3237 10591 3295 10597
rect 3237 10557 3249 10591
rect 3283 10588 3295 10591
rect 3326 10588 3332 10600
rect 3283 10560 3332 10588
rect 3283 10557 3295 10560
rect 3237 10551 3295 10557
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 3973 10591 4031 10597
rect 3973 10557 3985 10591
rect 4019 10588 4031 10591
rect 4890 10588 4896 10600
rect 4019 10560 4896 10588
rect 4019 10557 4031 10560
rect 3973 10551 4031 10557
rect 4890 10548 4896 10560
rect 4948 10548 4954 10600
rect 5537 10591 5595 10597
rect 5537 10557 5549 10591
rect 5583 10588 5595 10591
rect 5626 10588 5632 10600
rect 5583 10560 5632 10588
rect 5583 10557 5595 10560
rect 5537 10551 5595 10557
rect 1394 10412 1400 10464
rect 1452 10461 1458 10464
rect 1452 10452 1461 10461
rect 1670 10452 1676 10464
rect 1452 10424 1676 10452
rect 1452 10415 1461 10424
rect 1452 10412 1458 10415
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 3703 10455 3761 10461
rect 3703 10421 3715 10455
rect 3749 10452 3761 10455
rect 3970 10452 3976 10464
rect 3749 10424 3976 10452
rect 3749 10421 3761 10424
rect 3703 10415 3761 10421
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 5552 10452 5580 10551
rect 5626 10548 5632 10560
rect 5684 10548 5690 10600
rect 5902 10597 5908 10600
rect 5864 10591 5908 10597
rect 5864 10557 5876 10591
rect 5960 10588 5966 10600
rect 6196 10588 6224 10628
rect 6564 10600 6592 10628
rect 5960 10560 6224 10588
rect 5864 10551 5908 10557
rect 5902 10548 5908 10551
rect 5960 10548 5966 10560
rect 6270 10548 6276 10600
rect 6328 10548 6334 10600
rect 6546 10548 6552 10600
rect 6604 10548 6610 10600
rect 8404 10597 8432 10764
rect 8938 10684 8944 10736
rect 8996 10684 9002 10736
rect 11532 10724 11560 10764
rect 11609 10761 11621 10795
rect 11655 10792 11667 10795
rect 12986 10792 12992 10804
rect 11655 10764 12992 10792
rect 11655 10761 11667 10764
rect 11609 10755 11667 10761
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 13541 10795 13599 10801
rect 13541 10761 13553 10795
rect 13587 10792 13599 10795
rect 14550 10792 14556 10804
rect 13587 10764 14556 10792
rect 13587 10761 13599 10764
rect 13541 10755 13599 10761
rect 14550 10752 14556 10764
rect 14608 10752 14614 10804
rect 14642 10752 14648 10804
rect 14700 10792 14706 10804
rect 14700 10764 16252 10792
rect 14700 10752 14706 10764
rect 12894 10724 12900 10736
rect 11532 10696 12900 10724
rect 12894 10684 12900 10696
rect 12952 10724 12958 10736
rect 13354 10724 13360 10736
rect 12952 10696 13360 10724
rect 12952 10684 12958 10696
rect 13354 10684 13360 10696
rect 13412 10684 13418 10736
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 8956 10656 8984 10684
rect 8711 10628 8984 10656
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 9030 10616 9036 10668
rect 9088 10656 9094 10668
rect 9306 10656 9312 10668
rect 9088 10628 9312 10656
rect 9088 10616 9094 10628
rect 9306 10616 9312 10628
rect 9364 10656 9370 10668
rect 9364 10628 9720 10656
rect 9364 10616 9370 10628
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10557 8447 10591
rect 8389 10551 8447 10557
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 8941 10591 8999 10597
rect 8941 10588 8953 10591
rect 8812 10560 8953 10588
rect 8812 10548 8818 10560
rect 8941 10557 8953 10560
rect 8987 10557 8999 10591
rect 8941 10551 8999 10557
rect 9122 10548 9128 10600
rect 9180 10548 9186 10600
rect 9398 10548 9404 10600
rect 9456 10588 9462 10600
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 9456 10560 9505 10588
rect 9456 10548 9462 10560
rect 9493 10557 9505 10560
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10557 9643 10591
rect 9692 10588 9720 10628
rect 9858 10616 9864 10668
rect 9916 10656 9922 10668
rect 10048 10659 10106 10665
rect 10048 10656 10060 10659
rect 9916 10628 10060 10656
rect 9916 10616 9922 10628
rect 10048 10625 10060 10628
rect 10094 10625 10106 10659
rect 10048 10619 10106 10625
rect 10321 10659 10379 10665
rect 10321 10625 10333 10659
rect 10367 10656 10379 10659
rect 10686 10656 10692 10668
rect 10367 10628 10692 10656
rect 10367 10625 10379 10628
rect 10321 10619 10379 10625
rect 10686 10616 10692 10628
rect 10744 10616 10750 10668
rect 13814 10656 13820 10668
rect 11900 10628 13820 10656
rect 11900 10597 11928 10628
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 14280 10657 14338 10663
rect 14280 10623 14292 10657
rect 14326 10656 14338 10657
rect 14366 10656 14372 10668
rect 14326 10628 14372 10656
rect 14326 10623 14338 10628
rect 14280 10617 14338 10623
rect 14366 10616 14372 10628
rect 14424 10616 14430 10668
rect 11885 10591 11943 10597
rect 9692 10560 11008 10588
rect 9585 10551 9643 10557
rect 7650 10480 7656 10532
rect 7708 10480 7714 10532
rect 7742 10480 7748 10532
rect 7800 10520 7806 10532
rect 7837 10523 7895 10529
rect 7837 10520 7849 10523
rect 7800 10492 7849 10520
rect 7800 10480 7806 10492
rect 7837 10489 7849 10492
rect 7883 10520 7895 10523
rect 9140 10520 9168 10548
rect 9600 10520 9628 10551
rect 7883 10492 9628 10520
rect 10980 10520 11008 10560
rect 11885 10557 11897 10591
rect 11931 10557 11943 10591
rect 11885 10551 11943 10557
rect 11974 10548 11980 10600
rect 12032 10588 12038 10600
rect 12032 10560 12848 10588
rect 12032 10548 12038 10560
rect 12250 10520 12256 10532
rect 10980 10492 12256 10520
rect 7883 10489 7895 10492
rect 7837 10483 7895 10489
rect 12250 10480 12256 10492
rect 12308 10480 12314 10532
rect 12437 10523 12495 10529
rect 12437 10489 12449 10523
rect 12483 10489 12495 10523
rect 12820 10520 12848 10560
rect 12894 10548 12900 10600
rect 12952 10548 12958 10600
rect 13722 10548 13728 10600
rect 13780 10548 13786 10600
rect 14090 10588 14096 10600
rect 13832 10560 14096 10588
rect 13173 10523 13231 10529
rect 13173 10520 13185 10523
rect 12820 10492 13185 10520
rect 12437 10483 12495 10489
rect 13173 10489 13185 10492
rect 13219 10520 13231 10523
rect 13832 10520 13860 10560
rect 14090 10548 14096 10560
rect 14148 10597 14154 10600
rect 14148 10591 14202 10597
rect 14148 10557 14156 10591
rect 14190 10557 14202 10591
rect 14148 10551 14202 10557
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10588 14611 10591
rect 16114 10588 16120 10600
rect 14599 10560 16120 10588
rect 14599 10557 14611 10560
rect 14553 10551 14611 10557
rect 14148 10548 14154 10551
rect 16114 10548 16120 10560
rect 16172 10548 16178 10600
rect 16224 10597 16252 10764
rect 22738 10752 22744 10804
rect 22796 10752 22802 10804
rect 23477 10795 23535 10801
rect 23477 10761 23489 10795
rect 23523 10792 23535 10795
rect 24486 10792 24492 10804
rect 23523 10764 24492 10792
rect 23523 10761 23535 10764
rect 23477 10755 23535 10761
rect 24486 10752 24492 10764
rect 24544 10752 24550 10804
rect 25958 10752 25964 10804
rect 26016 10792 26022 10804
rect 26016 10764 29224 10792
rect 26016 10752 26022 10764
rect 19613 10727 19671 10733
rect 19613 10693 19625 10727
rect 19659 10724 19671 10727
rect 19794 10724 19800 10736
rect 19659 10696 19800 10724
rect 19659 10693 19671 10696
rect 19613 10687 19671 10693
rect 19794 10684 19800 10696
rect 19852 10684 19858 10736
rect 23566 10684 23572 10736
rect 23624 10684 23630 10736
rect 28997 10727 29055 10733
rect 28997 10693 29009 10727
rect 29043 10693 29055 10727
rect 28997 10687 29055 10693
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 16856 10659 16914 10665
rect 16856 10656 16868 10659
rect 16632 10628 16868 10656
rect 16632 10616 16638 10628
rect 16856 10625 16868 10628
rect 16902 10625 16914 10659
rect 16856 10619 16914 10625
rect 17494 10616 17500 10668
rect 17552 10656 17558 10668
rect 20487 10659 20545 10665
rect 17552 10628 20351 10656
rect 17552 10616 17558 10628
rect 20323 10600 20351 10628
rect 20487 10625 20499 10659
rect 20533 10656 20545 10659
rect 22738 10656 22744 10668
rect 20533 10628 22744 10656
rect 20533 10625 20545 10628
rect 20487 10619 20545 10625
rect 22738 10616 22744 10628
rect 22796 10616 22802 10668
rect 23584 10656 23612 10684
rect 22851 10628 23612 10656
rect 16209 10591 16267 10597
rect 16209 10557 16221 10591
rect 16255 10557 16267 10591
rect 16209 10551 16267 10557
rect 16393 10591 16451 10597
rect 16393 10557 16405 10591
rect 16439 10588 16451 10591
rect 16482 10588 16488 10600
rect 16439 10560 16488 10588
rect 16439 10557 16451 10560
rect 16393 10551 16451 10557
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 17129 10591 17187 10597
rect 17129 10557 17141 10591
rect 17175 10588 17187 10591
rect 17770 10588 17776 10600
rect 17175 10560 17776 10588
rect 17175 10557 17187 10560
rect 17129 10551 17187 10557
rect 17770 10548 17776 10560
rect 17828 10548 17834 10600
rect 18877 10591 18935 10597
rect 18877 10557 18889 10591
rect 18923 10588 18935 10591
rect 18923 10560 19104 10588
rect 18923 10557 18935 10560
rect 18877 10551 18935 10557
rect 13219 10492 13860 10520
rect 15933 10523 15991 10529
rect 13219 10489 13231 10492
rect 13173 10483 13231 10489
rect 15933 10489 15945 10523
rect 15979 10520 15991 10523
rect 15979 10492 16528 10520
rect 15979 10489 15991 10492
rect 15933 10483 15991 10489
rect 6086 10452 6092 10464
rect 5552 10424 6092 10452
rect 6086 10412 6092 10424
rect 6144 10412 6150 10464
rect 6546 10412 6552 10464
rect 6604 10452 6610 10464
rect 7558 10452 7564 10464
rect 6604 10424 7564 10452
rect 6604 10412 6610 10424
rect 7558 10412 7564 10424
rect 7616 10452 7622 10464
rect 9125 10455 9183 10461
rect 9125 10452 9137 10455
rect 7616 10424 9137 10452
rect 7616 10412 7622 10424
rect 9125 10421 9137 10424
rect 9171 10421 9183 10455
rect 9125 10415 9183 10421
rect 9309 10455 9367 10461
rect 9309 10421 9321 10455
rect 9355 10452 9367 10455
rect 9950 10452 9956 10464
rect 9355 10424 9956 10452
rect 9355 10421 9367 10424
rect 9309 10415 9367 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10042 10412 10048 10464
rect 10100 10461 10106 10464
rect 10100 10452 10109 10461
rect 10100 10424 10145 10452
rect 10100 10415 10109 10424
rect 10100 10412 10106 10415
rect 11606 10412 11612 10464
rect 11664 10452 11670 10464
rect 12452 10452 12480 10483
rect 11664 10424 12480 10452
rect 12713 10455 12771 10461
rect 11664 10412 11670 10424
rect 12713 10421 12725 10455
rect 12759 10452 12771 10455
rect 13906 10452 13912 10464
rect 12759 10424 13912 10452
rect 12759 10421 12771 10424
rect 12713 10415 12771 10421
rect 13906 10412 13912 10424
rect 13964 10412 13970 10464
rect 16022 10412 16028 10464
rect 16080 10412 16086 10464
rect 16500 10452 16528 10492
rect 18506 10480 18512 10532
rect 18564 10480 18570 10532
rect 19076 10464 19104 10560
rect 19978 10548 19984 10600
rect 20036 10548 20042 10600
rect 20323 10597 20352 10600
rect 20308 10591 20352 10597
rect 20308 10557 20320 10591
rect 20308 10551 20352 10557
rect 20346 10548 20352 10551
rect 20404 10548 20410 10600
rect 20714 10548 20720 10600
rect 20772 10548 20778 10600
rect 21358 10548 21364 10600
rect 21416 10588 21422 10600
rect 22465 10591 22523 10597
rect 22465 10588 22477 10591
rect 21416 10560 22477 10588
rect 21416 10548 21422 10560
rect 22465 10557 22477 10560
rect 22511 10588 22523 10591
rect 22646 10588 22652 10600
rect 22511 10560 22652 10588
rect 22511 10557 22523 10560
rect 22465 10551 22523 10557
rect 22646 10548 22652 10560
rect 22704 10588 22710 10600
rect 22851 10588 22879 10628
rect 22704 10560 22879 10588
rect 22925 10591 22983 10597
rect 22704 10548 22710 10560
rect 22925 10557 22937 10591
rect 22971 10588 22983 10591
rect 23198 10588 23204 10600
rect 22971 10560 23204 10588
rect 22971 10557 22983 10560
rect 22925 10551 22983 10557
rect 23198 10548 23204 10560
rect 23256 10548 23262 10600
rect 23584 10588 23612 10628
rect 24302 10616 24308 10668
rect 24360 10656 24366 10668
rect 26472 10659 26530 10665
rect 26472 10656 26484 10659
rect 24360 10628 24405 10656
rect 25056 10628 26484 10656
rect 24360 10616 24366 10628
rect 25056 10600 25084 10628
rect 26252 10600 26280 10628
rect 26472 10625 26484 10628
rect 26518 10625 26530 10659
rect 26472 10619 26530 10625
rect 26651 10659 26709 10665
rect 26651 10625 26663 10659
rect 26697 10656 26709 10659
rect 26881 10659 26939 10665
rect 26697 10628 26832 10656
rect 26697 10625 26709 10628
rect 26651 10619 26709 10625
rect 23661 10591 23719 10597
rect 23661 10588 23673 10591
rect 23584 10560 23673 10588
rect 23661 10557 23673 10560
rect 23707 10557 23719 10591
rect 23661 10551 23719 10557
rect 23842 10548 23848 10600
rect 23900 10548 23906 10600
rect 24210 10597 24216 10600
rect 24172 10591 24216 10597
rect 24172 10557 24184 10591
rect 24172 10551 24216 10557
rect 24210 10548 24216 10551
rect 24268 10548 24274 10600
rect 24578 10548 24584 10600
rect 24636 10548 24642 10600
rect 25038 10548 25044 10600
rect 25096 10548 25102 10600
rect 25314 10548 25320 10600
rect 25372 10588 25378 10600
rect 26142 10588 26148 10600
rect 25372 10560 26148 10588
rect 25372 10548 25378 10560
rect 26142 10548 26148 10560
rect 26200 10548 26206 10600
rect 26234 10548 26240 10600
rect 26292 10548 26298 10600
rect 26804 10588 26832 10628
rect 26881 10625 26893 10659
rect 26927 10656 26939 10659
rect 29012 10656 29040 10687
rect 26927 10628 29040 10656
rect 26927 10625 26939 10628
rect 26881 10619 26939 10625
rect 29196 10597 29224 10764
rect 29270 10616 29276 10668
rect 29328 10616 29334 10668
rect 29181 10591 29239 10597
rect 26804 10560 27752 10588
rect 16666 10452 16672 10464
rect 16500 10424 16672 10452
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 16859 10455 16917 10461
rect 16859 10421 16871 10455
rect 16905 10452 16917 10455
rect 17034 10452 17040 10464
rect 16905 10424 17040 10452
rect 16905 10421 16917 10424
rect 16859 10415 16917 10421
rect 17034 10412 17040 10424
rect 17092 10412 17098 10464
rect 18322 10412 18328 10464
rect 18380 10452 18386 10464
rect 18693 10455 18751 10461
rect 18693 10452 18705 10455
rect 18380 10424 18705 10452
rect 18380 10412 18386 10424
rect 18693 10421 18705 10424
rect 18739 10421 18751 10455
rect 18693 10415 18751 10421
rect 19058 10412 19064 10464
rect 19116 10412 19122 10464
rect 19150 10412 19156 10464
rect 19208 10412 19214 10464
rect 19996 10452 20024 10548
rect 27724 10464 27752 10560
rect 29181 10557 29193 10591
rect 29227 10557 29239 10591
rect 29288 10588 29316 10616
rect 29457 10591 29515 10597
rect 29457 10588 29469 10591
rect 29288 10560 29469 10588
rect 29181 10551 29239 10557
rect 29457 10557 29469 10560
rect 29503 10557 29515 10591
rect 29457 10551 29515 10557
rect 29733 10591 29791 10597
rect 29733 10557 29745 10591
rect 29779 10557 29791 10591
rect 29733 10551 29791 10557
rect 30009 10591 30067 10597
rect 30009 10557 30021 10591
rect 30055 10588 30067 10591
rect 30055 10560 30144 10588
rect 30055 10557 30067 10560
rect 30009 10551 30067 10557
rect 28445 10523 28503 10529
rect 28445 10489 28457 10523
rect 28491 10520 28503 10523
rect 28491 10492 28672 10520
rect 28491 10489 28503 10492
rect 28445 10483 28503 10489
rect 20438 10452 20444 10464
rect 19996 10424 20444 10452
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 21726 10412 21732 10464
rect 21784 10452 21790 10464
rect 21821 10455 21879 10461
rect 21821 10452 21833 10455
rect 21784 10424 21833 10452
rect 21784 10412 21790 10424
rect 21821 10421 21833 10424
rect 21867 10421 21879 10455
rect 21821 10415 21879 10421
rect 22281 10455 22339 10461
rect 22281 10421 22293 10455
rect 22327 10452 22339 10455
rect 24578 10452 24584 10464
rect 22327 10424 24584 10452
rect 22327 10421 22339 10424
rect 22281 10415 22339 10421
rect 24578 10412 24584 10424
rect 24636 10412 24642 10464
rect 25682 10412 25688 10464
rect 25740 10412 25746 10464
rect 27706 10412 27712 10464
rect 27764 10412 27770 10464
rect 28166 10412 28172 10464
rect 28224 10412 28230 10464
rect 28534 10412 28540 10464
rect 28592 10412 28598 10464
rect 28644 10452 28672 10492
rect 28718 10480 28724 10532
rect 28776 10520 28782 10532
rect 29748 10520 29776 10551
rect 29914 10520 29920 10532
rect 28776 10492 29592 10520
rect 29748 10492 29920 10520
rect 28776 10480 28782 10492
rect 28902 10452 28908 10464
rect 28644 10424 28908 10452
rect 28902 10412 28908 10424
rect 28960 10412 28966 10464
rect 29270 10412 29276 10464
rect 29328 10412 29334 10464
rect 29564 10461 29592 10492
rect 29914 10480 29920 10492
rect 29972 10480 29978 10532
rect 30116 10464 30144 10560
rect 29549 10455 29607 10461
rect 29549 10421 29561 10455
rect 29595 10421 29607 10455
rect 29549 10415 29607 10421
rect 29638 10412 29644 10464
rect 29696 10452 29702 10464
rect 29825 10455 29883 10461
rect 29825 10452 29837 10455
rect 29696 10424 29837 10452
rect 29696 10412 29702 10424
rect 29825 10421 29837 10424
rect 29871 10421 29883 10455
rect 29825 10415 29883 10421
rect 30098 10412 30104 10464
rect 30156 10412 30162 10464
rect 552 10362 31072 10384
rect 552 10310 7988 10362
rect 8040 10310 8052 10362
rect 8104 10310 8116 10362
rect 8168 10310 8180 10362
rect 8232 10310 8244 10362
rect 8296 10310 15578 10362
rect 15630 10310 15642 10362
rect 15694 10310 15706 10362
rect 15758 10310 15770 10362
rect 15822 10310 15834 10362
rect 15886 10310 23168 10362
rect 23220 10310 23232 10362
rect 23284 10310 23296 10362
rect 23348 10310 23360 10362
rect 23412 10310 23424 10362
rect 23476 10310 30758 10362
rect 30810 10310 30822 10362
rect 30874 10310 30886 10362
rect 30938 10310 30950 10362
rect 31002 10310 31014 10362
rect 31066 10310 31072 10362
rect 552 10288 31072 10310
rect 658 10208 664 10260
rect 716 10208 722 10260
rect 1394 10208 1400 10260
rect 1452 10248 1458 10260
rect 1587 10251 1645 10257
rect 1587 10248 1599 10251
rect 1452 10220 1599 10248
rect 1452 10208 1458 10220
rect 1587 10217 1599 10220
rect 1633 10217 1645 10251
rect 1587 10211 1645 10217
rect 2958 10208 2964 10260
rect 3016 10248 3022 10260
rect 3694 10248 3700 10260
rect 3016 10220 3700 10248
rect 3016 10208 3022 10220
rect 3694 10208 3700 10220
rect 3752 10208 3758 10260
rect 3795 10251 3853 10257
rect 3795 10217 3807 10251
rect 3841 10248 3853 10251
rect 3970 10248 3976 10260
rect 3841 10220 3976 10248
rect 3841 10217 3853 10220
rect 3795 10211 3853 10217
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 6454 10208 6460 10260
rect 6512 10208 6518 10260
rect 6923 10251 6981 10257
rect 6923 10217 6935 10251
rect 6969 10248 6981 10251
rect 7466 10248 7472 10260
rect 6969 10220 7472 10248
rect 6969 10217 6981 10220
rect 6923 10211 6981 10217
rect 7466 10208 7472 10220
rect 7524 10248 7530 10260
rect 8938 10248 8944 10260
rect 7524 10220 8944 10248
rect 7524 10208 7530 10220
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9131 10251 9189 10257
rect 9131 10217 9143 10251
rect 9177 10248 9189 10251
rect 9306 10248 9312 10260
rect 9177 10220 9312 10248
rect 9177 10217 9189 10220
rect 9131 10211 9189 10217
rect 9306 10208 9312 10220
rect 9364 10248 9370 10260
rect 9490 10248 9496 10260
rect 9364 10220 9496 10248
rect 9364 10208 9370 10220
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 11606 10208 11612 10260
rect 11664 10257 11670 10260
rect 11664 10248 11673 10257
rect 11974 10248 11980 10260
rect 11664 10220 11980 10248
rect 11664 10211 11673 10220
rect 11664 10208 11670 10211
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 14090 10208 14096 10260
rect 14148 10248 14154 10260
rect 14283 10251 14341 10257
rect 14283 10248 14295 10251
rect 14148 10220 14295 10248
rect 14148 10208 14154 10220
rect 14283 10217 14295 10220
rect 14329 10217 14341 10251
rect 17227 10251 17285 10257
rect 17227 10248 17239 10251
rect 14283 10211 14341 10217
rect 16500 10220 17239 10248
rect 676 10112 704 10208
rect 5442 10140 5448 10192
rect 5500 10140 5506 10192
rect 6086 10180 6092 10192
rect 5920 10152 6092 10180
rect 1029 10115 1087 10121
rect 1029 10112 1041 10115
rect 676 10084 1041 10112
rect 1029 10081 1041 10084
rect 1075 10081 1087 10115
rect 1029 10075 1087 10081
rect 1118 10072 1124 10124
rect 1176 10072 1182 10124
rect 3237 10115 3295 10121
rect 1786 10084 3188 10112
rect 1617 10065 1675 10071
rect 1617 10062 1629 10065
rect 1596 10031 1629 10062
rect 1663 10044 1675 10065
rect 1786 10044 1814 10084
rect 1663 10031 1814 10044
rect 1596 10016 1814 10031
rect 1854 10004 1860 10056
rect 1912 10004 1918 10056
rect 845 9911 903 9917
rect 845 9877 857 9911
rect 891 9908 903 9911
rect 3050 9908 3056 9920
rect 891 9880 3056 9908
rect 891 9877 903 9880
rect 845 9871 903 9877
rect 3050 9868 3056 9880
rect 3108 9868 3114 9920
rect 3160 9908 3188 10084
rect 3237 10081 3249 10115
rect 3283 10112 3295 10115
rect 3283 10084 3832 10112
rect 3283 10081 3295 10084
rect 3237 10075 3295 10081
rect 3326 10004 3332 10056
rect 3384 10004 3390 10056
rect 3804 10053 3832 10084
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 5920 10121 5948 10152
rect 6086 10140 6092 10152
rect 6144 10140 6150 10192
rect 6181 10183 6239 10189
rect 6181 10149 6193 10183
rect 6227 10180 6239 10183
rect 6472 10180 6500 10208
rect 16500 10189 16528 10220
rect 17227 10217 17239 10220
rect 17273 10248 17285 10251
rect 17494 10248 17500 10260
rect 17273 10220 17500 10248
rect 17273 10217 17285 10220
rect 17227 10211 17285 10217
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 20349 10251 20407 10257
rect 20349 10217 20361 10251
rect 20395 10248 20407 10251
rect 20714 10248 20720 10260
rect 20395 10220 20720 10248
rect 20395 10217 20407 10220
rect 20349 10211 20407 10217
rect 20714 10208 20720 10220
rect 20772 10208 20778 10260
rect 21174 10208 21180 10260
rect 21232 10248 21238 10260
rect 21735 10251 21793 10257
rect 21735 10248 21747 10251
rect 21232 10220 21747 10248
rect 21232 10208 21238 10220
rect 21735 10217 21747 10220
rect 21781 10248 21793 10251
rect 21781 10220 22968 10248
rect 21781 10217 21793 10220
rect 21735 10211 21793 10217
rect 6227 10152 6500 10180
rect 16485 10183 16543 10189
rect 6227 10149 6239 10152
rect 6181 10143 6239 10149
rect 16485 10149 16497 10183
rect 16531 10149 16543 10183
rect 16485 10143 16543 10149
rect 18877 10183 18935 10189
rect 18877 10149 18889 10183
rect 18923 10180 18935 10183
rect 18966 10180 18972 10192
rect 18923 10152 18972 10180
rect 18923 10149 18935 10152
rect 18877 10143 18935 10149
rect 18966 10140 18972 10152
rect 19024 10140 19030 10192
rect 21358 10180 21364 10192
rect 19812 10152 21364 10180
rect 5905 10115 5963 10121
rect 5905 10112 5917 10115
rect 3936 10084 5917 10112
rect 3936 10072 3942 10084
rect 5905 10081 5917 10084
rect 5951 10081 5963 10115
rect 5905 10075 5963 10081
rect 8573 10115 8631 10121
rect 8573 10081 8585 10115
rect 8619 10112 8631 10115
rect 9401 10115 9459 10121
rect 8619 10084 9171 10112
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 3792 10047 3850 10053
rect 3792 10013 3804 10047
rect 3838 10013 3850 10047
rect 3792 10007 3850 10013
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10044 4123 10047
rect 5718 10044 5724 10056
rect 4111 10016 5724 10044
rect 4111 10013 4123 10016
rect 4065 10007 4123 10013
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 6454 10004 6460 10056
rect 6512 10004 6518 10056
rect 6920 10049 6978 10055
rect 6920 10015 6932 10049
rect 6966 10044 6978 10049
rect 7006 10044 7012 10056
rect 6966 10016 7012 10044
rect 6966 10015 6978 10016
rect 6920 10009 6978 10015
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10044 7251 10047
rect 7558 10044 7564 10056
rect 7239 10016 7564 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 7558 10004 7564 10016
rect 7616 10004 7622 10056
rect 8665 10047 8723 10053
rect 8665 10013 8677 10047
rect 8711 10044 8723 10047
rect 9030 10044 9036 10056
rect 8711 10016 9036 10044
rect 8711 10013 8723 10016
rect 8665 10007 8723 10013
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 9143 10055 9171 10084
rect 9401 10081 9413 10115
rect 9447 10112 9459 10115
rect 10134 10112 10140 10124
rect 9447 10084 10140 10112
rect 9447 10081 9459 10084
rect 9401 10075 9459 10081
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 10962 10072 10968 10124
rect 11020 10112 11026 10124
rect 11020 10084 11284 10112
rect 11020 10072 11026 10084
rect 9128 10049 9186 10055
rect 9128 10015 9140 10049
rect 9174 10015 9186 10049
rect 9128 10009 9186 10015
rect 11146 10004 11152 10056
rect 11204 10004 11210 10056
rect 11256 10044 11284 10084
rect 12250 10072 12256 10124
rect 12308 10112 12314 10124
rect 13541 10115 13599 10121
rect 13541 10112 13553 10115
rect 12308 10084 13553 10112
rect 12308 10072 12314 10084
rect 13541 10081 13553 10084
rect 13587 10081 13599 10115
rect 13541 10075 13599 10081
rect 13814 10072 13820 10124
rect 13872 10072 13878 10124
rect 14458 10072 14464 10124
rect 14516 10072 14522 10124
rect 14550 10072 14556 10124
rect 14608 10072 14614 10124
rect 16209 10115 16267 10121
rect 16209 10081 16221 10115
rect 16255 10081 16267 10115
rect 16209 10075 16267 10081
rect 11612 10065 11670 10071
rect 11612 10044 11624 10065
rect 11256 10031 11624 10044
rect 11658 10031 11670 10065
rect 11256 10025 11670 10031
rect 11885 10047 11943 10053
rect 11256 10016 11652 10025
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 12526 10044 12532 10056
rect 11931 10016 12532 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 12526 10004 12532 10016
rect 12584 10004 12590 10056
rect 14323 10047 14381 10053
rect 14323 10013 14335 10047
rect 14369 10044 14381 10047
rect 14476 10044 14504 10072
rect 14369 10016 14504 10044
rect 14369 10013 14381 10016
rect 14323 10007 14381 10013
rect 16224 9976 16252 10075
rect 16850 10072 16856 10124
rect 16908 10112 16914 10124
rect 17497 10115 17555 10121
rect 17497 10112 17509 10115
rect 16908 10084 17509 10112
rect 16908 10072 16914 10084
rect 17497 10081 17509 10084
rect 17543 10081 17555 10115
rect 17497 10075 17555 10081
rect 18598 10072 18604 10124
rect 18656 10112 18662 10124
rect 19150 10112 19156 10124
rect 18656 10084 19156 10112
rect 18656 10072 18662 10084
rect 19150 10072 19156 10084
rect 19208 10112 19214 10124
rect 19812 10121 19840 10152
rect 21358 10140 21364 10152
rect 21416 10140 21422 10192
rect 19337 10115 19395 10121
rect 19337 10112 19349 10115
rect 19208 10084 19349 10112
rect 19208 10072 19214 10084
rect 19337 10081 19349 10084
rect 19383 10081 19395 10115
rect 19337 10075 19395 10081
rect 19797 10115 19855 10121
rect 19797 10081 19809 10115
rect 19843 10081 19855 10115
rect 19797 10075 19855 10081
rect 20073 10115 20131 10121
rect 20073 10081 20085 10115
rect 20119 10112 20131 10115
rect 20533 10115 20591 10121
rect 20533 10112 20545 10115
rect 20119 10084 20545 10112
rect 20119 10081 20131 10084
rect 20073 10075 20131 10081
rect 20533 10081 20545 10084
rect 20579 10112 20591 10115
rect 20622 10112 20628 10124
rect 20579 10084 20628 10112
rect 20579 10081 20591 10084
rect 20533 10075 20591 10081
rect 20622 10072 20628 10084
rect 20680 10072 20686 10124
rect 20717 10115 20775 10121
rect 20717 10081 20729 10115
rect 20763 10081 20775 10115
rect 20717 10075 20775 10081
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10044 16819 10047
rect 16942 10044 16948 10056
rect 16807 10016 16948 10044
rect 16807 10013 16819 10016
rect 16761 10007 16819 10013
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17267 10047 17325 10053
rect 17267 10013 17279 10047
rect 17313 10044 17325 10047
rect 18782 10044 18788 10056
rect 17313 10016 18788 10044
rect 17313 10013 17325 10016
rect 17267 10007 17325 10013
rect 18782 10004 18788 10016
rect 18840 10004 18846 10056
rect 20438 10004 20444 10056
rect 20496 10044 20502 10056
rect 20732 10044 20760 10075
rect 21082 10072 21088 10124
rect 21140 10112 21146 10124
rect 21269 10115 21327 10121
rect 21269 10112 21281 10115
rect 21140 10084 21281 10112
rect 21140 10072 21146 10084
rect 21269 10081 21281 10084
rect 21315 10112 21327 10115
rect 21315 10084 21864 10112
rect 21315 10081 21327 10084
rect 21269 10075 21327 10081
rect 21726 10044 21732 10056
rect 20496 10016 20760 10044
rect 21690 10016 21732 10044
rect 20496 10004 20502 10016
rect 21726 10004 21732 10016
rect 21784 10004 21790 10056
rect 21836 10044 21864 10084
rect 22002 10072 22008 10124
rect 22060 10072 22066 10124
rect 22940 10112 22968 10220
rect 23014 10208 23020 10260
rect 23072 10248 23078 10260
rect 23109 10251 23167 10257
rect 23109 10248 23121 10251
rect 23072 10220 23121 10248
rect 23072 10208 23078 10220
rect 23109 10217 23121 10220
rect 23155 10217 23167 10251
rect 25038 10248 25044 10260
rect 23109 10211 23167 10217
rect 23676 10220 25044 10248
rect 23676 10112 23704 10220
rect 25038 10208 25044 10220
rect 25096 10208 25102 10260
rect 25682 10208 25688 10260
rect 25740 10208 25746 10260
rect 25866 10208 25872 10260
rect 25924 10248 25930 10260
rect 30009 10251 30067 10257
rect 30009 10248 30021 10251
rect 25924 10220 30021 10248
rect 25924 10208 25930 10220
rect 30009 10217 30021 10220
rect 30055 10217 30067 10251
rect 30009 10211 30067 10217
rect 23896 10115 23954 10121
rect 23896 10112 23908 10115
rect 22940 10084 23908 10112
rect 23896 10081 23908 10084
rect 23942 10081 23954 10115
rect 25700 10112 25728 10208
rect 28258 10140 28264 10192
rect 28316 10180 28322 10192
rect 28316 10152 28764 10180
rect 28316 10140 28322 10152
rect 23896 10075 23954 10081
rect 24228 10084 25728 10112
rect 25961 10115 26019 10121
rect 23569 10047 23627 10053
rect 23569 10044 23581 10047
rect 21836 10016 23581 10044
rect 23569 10013 23581 10016
rect 23615 10013 23627 10047
rect 23569 10007 23627 10013
rect 24075 10047 24133 10053
rect 24075 10013 24087 10047
rect 24121 10044 24133 10047
rect 24228 10044 24256 10084
rect 25961 10081 25973 10115
rect 26007 10081 26019 10115
rect 25961 10075 26019 10081
rect 24121 10016 24256 10044
rect 24305 10047 24363 10053
rect 24121 10013 24133 10016
rect 24075 10007 24133 10013
rect 24305 10013 24317 10047
rect 24351 10044 24363 10047
rect 24486 10044 24492 10056
rect 24351 10016 24492 10044
rect 24351 10013 24363 10016
rect 24305 10007 24363 10013
rect 19613 9979 19671 9985
rect 10060 9948 11192 9976
rect 16224 9948 16804 9976
rect 10060 9908 10088 9948
rect 3160 9880 10088 9908
rect 10689 9911 10747 9917
rect 10689 9877 10701 9911
rect 10735 9908 10747 9911
rect 11054 9908 11060 9920
rect 10735 9880 11060 9908
rect 10735 9877 10747 9880
rect 10689 9871 10747 9877
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11164 9908 11192 9948
rect 16776 9920 16804 9948
rect 19613 9945 19625 9979
rect 19659 9976 19671 9979
rect 19659 9948 21312 9976
rect 19659 9945 19671 9948
rect 19613 9939 19671 9945
rect 12250 9908 12256 9920
rect 11164 9880 12256 9908
rect 12250 9868 12256 9880
rect 12308 9868 12314 9920
rect 12342 9868 12348 9920
rect 12400 9908 12406 9920
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12400 9880 13001 9908
rect 12400 9868 12406 9880
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 12989 9871 13047 9877
rect 15010 9868 15016 9920
rect 15068 9908 15074 9920
rect 15657 9911 15715 9917
rect 15657 9908 15669 9911
rect 15068 9880 15669 9908
rect 15068 9868 15074 9880
rect 15657 9877 15669 9880
rect 15703 9877 15715 9911
rect 15657 9871 15715 9877
rect 16758 9868 16764 9920
rect 16816 9868 16822 9920
rect 18138 9868 18144 9920
rect 18196 9908 18202 9920
rect 19153 9911 19211 9917
rect 19153 9908 19165 9911
rect 18196 9880 19165 9908
rect 18196 9868 18202 9880
rect 19153 9877 19165 9880
rect 19199 9877 19211 9911
rect 19153 9871 19211 9877
rect 19889 9911 19947 9917
rect 19889 9877 19901 9911
rect 19935 9908 19947 9911
rect 20714 9908 20720 9920
rect 19935 9880 20720 9908
rect 19935 9877 19947 9880
rect 19889 9871 19947 9877
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 20806 9868 20812 9920
rect 20864 9868 20870 9920
rect 21284 9908 21312 9948
rect 21910 9908 21916 9920
rect 21284 9880 21916 9908
rect 21910 9868 21916 9880
rect 21968 9868 21974 9920
rect 23584 9908 23612 10007
rect 24486 10004 24492 10016
rect 24544 10004 24550 10056
rect 25130 10004 25136 10056
rect 25188 10044 25194 10056
rect 25976 10044 26004 10075
rect 26142 10072 26148 10124
rect 26200 10112 26206 10124
rect 26421 10115 26479 10121
rect 26421 10112 26433 10115
rect 26200 10084 26433 10112
rect 26200 10072 26206 10084
rect 26421 10081 26433 10084
rect 26467 10081 26479 10115
rect 26421 10075 26479 10081
rect 27157 10115 27215 10121
rect 27157 10081 27169 10115
rect 27203 10112 27215 10115
rect 28350 10112 28356 10124
rect 27203 10084 28356 10112
rect 27203 10081 27215 10084
rect 27157 10075 27215 10081
rect 28350 10072 28356 10084
rect 28408 10072 28414 10124
rect 28442 10072 28448 10124
rect 28500 10112 28506 10124
rect 28629 10115 28687 10121
rect 28629 10112 28641 10115
rect 28500 10084 28641 10112
rect 28500 10072 28506 10084
rect 28629 10081 28641 10084
rect 28675 10081 28687 10115
rect 28736 10112 28764 10152
rect 28905 10115 28963 10121
rect 28905 10112 28917 10115
rect 28736 10084 28917 10112
rect 28629 10075 28687 10081
rect 28905 10081 28917 10084
rect 28951 10081 28963 10115
rect 28905 10075 28963 10081
rect 26050 10044 26056 10056
rect 25188 10016 26056 10044
rect 25188 10004 25194 10016
rect 26050 10004 26056 10016
rect 26108 10004 26114 10056
rect 26234 10004 26240 10056
rect 26292 10044 26298 10056
rect 26748 10047 26806 10053
rect 26748 10044 26760 10047
rect 26292 10016 26760 10044
rect 26292 10004 26298 10016
rect 26748 10013 26760 10016
rect 26794 10013 26806 10047
rect 26748 10007 26806 10013
rect 26878 10004 26884 10056
rect 26936 10004 26942 10056
rect 25314 9976 25320 9988
rect 24970 9948 25320 9976
rect 24970 9908 24998 9948
rect 25314 9936 25320 9948
rect 25372 9936 25378 9988
rect 25593 9979 25651 9985
rect 25593 9945 25605 9979
rect 25639 9976 25651 9979
rect 25639 9948 26464 9976
rect 25639 9945 25651 9948
rect 25593 9939 25651 9945
rect 23584 9880 24998 9908
rect 25038 9868 25044 9920
rect 25096 9908 25102 9920
rect 25958 9908 25964 9920
rect 25096 9880 25964 9908
rect 25096 9868 25102 9880
rect 25958 9868 25964 9880
rect 26016 9908 26022 9920
rect 26145 9911 26203 9917
rect 26145 9908 26157 9911
rect 26016 9880 26157 9908
rect 26016 9868 26022 9880
rect 26145 9877 26157 9880
rect 26191 9877 26203 9911
rect 26436 9908 26464 9948
rect 26694 9908 26700 9920
rect 26436 9880 26700 9908
rect 26145 9871 26203 9877
rect 26694 9868 26700 9880
rect 26752 9868 26758 9920
rect 28258 9868 28264 9920
rect 28316 9868 28322 9920
rect 28902 9868 28908 9920
rect 28960 9908 28966 9920
rect 30098 9908 30104 9920
rect 28960 9880 30104 9908
rect 28960 9868 28966 9880
rect 30098 9868 30104 9880
rect 30156 9868 30162 9920
rect 552 9818 30912 9840
rect 552 9766 4193 9818
rect 4245 9766 4257 9818
rect 4309 9766 4321 9818
rect 4373 9766 4385 9818
rect 4437 9766 4449 9818
rect 4501 9766 11783 9818
rect 11835 9766 11847 9818
rect 11899 9766 11911 9818
rect 11963 9766 11975 9818
rect 12027 9766 12039 9818
rect 12091 9766 19373 9818
rect 19425 9766 19437 9818
rect 19489 9766 19501 9818
rect 19553 9766 19565 9818
rect 19617 9766 19629 9818
rect 19681 9766 26963 9818
rect 27015 9766 27027 9818
rect 27079 9766 27091 9818
rect 27143 9766 27155 9818
rect 27207 9766 27219 9818
rect 27271 9766 30912 9818
rect 552 9744 30912 9766
rect 842 9664 848 9716
rect 900 9704 906 9716
rect 1854 9704 1860 9716
rect 900 9676 1860 9704
rect 900 9664 906 9676
rect 1854 9664 1860 9676
rect 1912 9664 1918 9716
rect 2682 9664 2688 9716
rect 2740 9704 2746 9716
rect 2740 9664 2774 9704
rect 3050 9664 3056 9716
rect 3108 9704 3114 9716
rect 5258 9704 5264 9716
rect 3108 9676 5264 9704
rect 3108 9664 3114 9676
rect 5258 9664 5264 9676
rect 5316 9664 5322 9716
rect 5813 9707 5871 9713
rect 5813 9673 5825 9707
rect 5859 9704 5871 9707
rect 6270 9704 6276 9716
rect 5859 9676 6276 9704
rect 5859 9673 5871 9676
rect 5813 9667 5871 9673
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 6638 9664 6644 9716
rect 6696 9704 6702 9716
rect 9122 9704 9128 9716
rect 6696 9676 7512 9704
rect 6696 9664 6702 9676
rect 2746 9648 2774 9664
rect 2746 9608 2780 9648
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 3234 9636 3240 9648
rect 2884 9608 3240 9636
rect 937 9571 995 9577
rect 937 9537 949 9571
rect 983 9568 995 9571
rect 1118 9568 1124 9580
rect 983 9540 1124 9568
rect 983 9537 995 9540
rect 937 9531 995 9537
rect 1118 9528 1124 9540
rect 1176 9528 1182 9580
rect 1443 9571 1501 9577
rect 1443 9537 1455 9571
rect 1489 9568 1501 9571
rect 2884 9568 2912 9608
rect 3234 9596 3240 9608
rect 3292 9636 3298 9648
rect 3421 9639 3479 9645
rect 3421 9636 3433 9639
rect 3292 9608 3433 9636
rect 3292 9596 3298 9608
rect 3421 9605 3433 9608
rect 3467 9605 3479 9639
rect 7484 9636 7512 9676
rect 8312 9676 9128 9704
rect 8312 9636 8340 9676
rect 9122 9664 9128 9676
rect 9180 9704 9186 9716
rect 9180 9676 10916 9704
rect 9180 9664 9186 9676
rect 7484 9608 8340 9636
rect 3421 9599 3479 9605
rect 8386 9596 8392 9648
rect 8444 9636 8450 9648
rect 8573 9639 8631 9645
rect 8573 9636 8585 9639
rect 8444 9608 8585 9636
rect 8444 9596 8450 9608
rect 8573 9605 8585 9608
rect 8619 9605 8631 9639
rect 10888 9636 10916 9676
rect 10962 9664 10968 9716
rect 11020 9664 11026 9716
rect 13906 9704 13912 9716
rect 11072 9676 13912 9704
rect 11072 9636 11100 9676
rect 13906 9664 13912 9676
rect 13964 9664 13970 9716
rect 16114 9664 16120 9716
rect 16172 9664 16178 9716
rect 16758 9664 16764 9716
rect 16816 9704 16822 9716
rect 17034 9704 17040 9716
rect 16816 9676 17040 9704
rect 16816 9664 16822 9676
rect 17034 9664 17040 9676
rect 17092 9664 17098 9716
rect 19886 9704 19892 9716
rect 17926 9676 19892 9704
rect 10888 9608 11100 9636
rect 8573 9599 8631 9605
rect 1489 9540 2912 9568
rect 3053 9571 3111 9577
rect 1489 9537 1501 9540
rect 1443 9531 1501 9537
rect 3053 9537 3065 9571
rect 3099 9568 3111 9571
rect 4068 9571 4126 9577
rect 4068 9568 4080 9571
rect 3099 9540 4080 9568
rect 3099 9537 3111 9540
rect 3053 9531 3111 9537
rect 4068 9537 4080 9540
rect 4114 9537 4126 9571
rect 4068 9531 4126 9537
rect 6089 9571 6147 9577
rect 6089 9537 6101 9571
rect 6135 9568 6147 9571
rect 6362 9568 6368 9580
rect 6135 9540 6368 9568
rect 6135 9537 6147 9540
rect 6089 9531 6147 9537
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 6595 9571 6653 9577
rect 6595 9537 6607 9571
rect 6641 9568 6653 9571
rect 6914 9568 6920 9580
rect 6641 9540 6920 9568
rect 6641 9537 6653 9540
rect 6595 9531 6653 9537
rect 6914 9528 6920 9540
rect 6972 9528 6978 9580
rect 8588 9568 8616 9599
rect 9306 9577 9312 9580
rect 9268 9571 9312 9577
rect 8588 9540 9168 9568
rect 1670 9460 1676 9512
rect 1728 9460 1734 9512
rect 3326 9460 3332 9512
rect 3384 9500 3390 9512
rect 3970 9509 3976 9512
rect 3605 9503 3663 9509
rect 3605 9500 3617 9503
rect 3384 9472 3617 9500
rect 3384 9460 3390 9472
rect 3605 9469 3617 9472
rect 3651 9469 3663 9503
rect 3605 9463 3663 9469
rect 3932 9503 3976 9509
rect 3932 9469 3944 9503
rect 3932 9463 3976 9469
rect 3970 9460 3976 9463
rect 4028 9460 4034 9512
rect 4338 9460 4344 9512
rect 4396 9460 4402 9512
rect 5997 9503 6055 9509
rect 5997 9500 6009 9503
rect 5276 9472 6009 9500
rect 5276 9376 5304 9472
rect 5997 9469 6009 9472
rect 6043 9500 6055 9503
rect 6454 9500 6460 9512
rect 6043 9472 6460 9500
rect 6043 9469 6055 9472
rect 5997 9463 6055 9469
rect 6454 9460 6460 9472
rect 6512 9460 6518 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 7098 9500 7104 9512
rect 6871 9472 7104 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 8389 9503 8447 9509
rect 8389 9469 8401 9503
rect 8435 9500 8447 9503
rect 8478 9500 8484 9512
rect 8435 9472 8484 9500
rect 8435 9469 8447 9472
rect 8389 9463 8447 9469
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9500 8999 9503
rect 9030 9500 9036 9512
rect 8987 9472 9036 9500
rect 8987 9469 8999 9472
rect 8941 9463 8999 9469
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9140 9500 9168 9540
rect 9268 9537 9280 9571
rect 9268 9531 9312 9537
rect 9306 9528 9312 9531
rect 9364 9528 9370 9580
rect 9404 9569 9462 9575
rect 9404 9535 9416 9569
rect 9450 9568 9462 9569
rect 9490 9568 9496 9580
rect 9450 9540 9496 9568
rect 9450 9535 9462 9540
rect 9404 9529 9462 9535
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 9677 9571 9735 9577
rect 9677 9537 9689 9571
rect 9723 9568 9735 9571
rect 10410 9568 10416 9580
rect 9723 9540 10416 9568
rect 9723 9537 9735 9540
rect 9677 9531 9735 9537
rect 10410 9528 10416 9540
rect 10468 9528 10474 9580
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 14090 9577 14096 9580
rect 11612 9571 11670 9577
rect 11612 9568 11624 9571
rect 11112 9540 11624 9568
rect 11112 9528 11118 9540
rect 11612 9537 11624 9540
rect 11658 9537 11670 9571
rect 14052 9571 14096 9577
rect 11612 9531 11670 9537
rect 11716 9540 13676 9568
rect 9140 9472 10456 9500
rect 5442 9392 5448 9444
rect 5500 9432 5506 9444
rect 5721 9435 5779 9441
rect 5721 9432 5733 9435
rect 5500 9404 5733 9432
rect 5500 9392 5506 9404
rect 5721 9401 5733 9404
rect 5767 9401 5779 9435
rect 5721 9395 5779 9401
rect 8205 9435 8263 9441
rect 8205 9401 8217 9435
rect 8251 9432 8263 9435
rect 8754 9432 8760 9444
rect 8251 9404 8760 9432
rect 8251 9401 8263 9404
rect 8205 9395 8263 9401
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 1394 9324 1400 9376
rect 1452 9373 1458 9376
rect 1452 9364 1461 9373
rect 1452 9336 1497 9364
rect 1452 9327 1461 9336
rect 1452 9324 1458 9327
rect 2038 9324 2044 9376
rect 2096 9364 2102 9376
rect 2958 9364 2964 9376
rect 2096 9336 2964 9364
rect 2096 9324 2102 9336
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 4246 9324 4252 9376
rect 4304 9364 4310 9376
rect 5258 9364 5264 9376
rect 4304 9336 5264 9364
rect 4304 9324 4310 9336
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 6555 9367 6613 9373
rect 6555 9333 6567 9367
rect 6601 9364 6613 9367
rect 7466 9364 7472 9376
rect 6601 9336 7472 9364
rect 6601 9333 6613 9336
rect 6555 9327 6613 9333
rect 7466 9324 7472 9336
rect 7524 9324 7530 9376
rect 9048 9364 9076 9460
rect 9582 9364 9588 9376
rect 9048 9336 9588 9364
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 10428 9364 10456 9472
rect 11146 9460 11152 9512
rect 11204 9460 11210 9512
rect 11716 9500 11744 9540
rect 11256 9472 11744 9500
rect 10502 9392 10508 9444
rect 10560 9432 10566 9444
rect 11256 9432 11284 9472
rect 11882 9460 11888 9512
rect 11940 9460 11946 9512
rect 10560 9404 11284 9432
rect 10560 9392 10566 9404
rect 11238 9364 11244 9376
rect 10428 9336 11244 9364
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 11606 9324 11612 9376
rect 11664 9373 11670 9376
rect 11664 9364 11673 9373
rect 11664 9336 11709 9364
rect 11664 9327 11673 9336
rect 11664 9324 11670 9327
rect 12618 9324 12624 9376
rect 12676 9364 12682 9376
rect 12989 9367 13047 9373
rect 12989 9364 13001 9367
rect 12676 9336 13001 9364
rect 12676 9324 12682 9336
rect 12989 9333 13001 9336
rect 13035 9333 13047 9367
rect 13648 9364 13676 9540
rect 14052 9537 14064 9571
rect 14052 9531 14096 9537
rect 14090 9528 14096 9531
rect 14148 9528 14154 9580
rect 14231 9571 14289 9577
rect 14231 9537 14243 9571
rect 14277 9568 14289 9571
rect 14918 9568 14924 9580
rect 14277 9540 14924 9568
rect 14277 9537 14289 9540
rect 14231 9531 14289 9537
rect 14918 9528 14924 9540
rect 14976 9528 14982 9580
rect 16899 9571 16957 9577
rect 16899 9537 16911 9571
rect 16945 9568 16957 9571
rect 17926 9568 17954 9676
rect 19886 9664 19892 9676
rect 19944 9664 19950 9716
rect 20438 9664 20444 9716
rect 20496 9704 20502 9716
rect 20496 9676 22692 9704
rect 20496 9664 20502 9676
rect 18046 9596 18052 9648
rect 18104 9636 18110 9648
rect 18233 9639 18291 9645
rect 18233 9636 18245 9639
rect 18104 9608 18245 9636
rect 18104 9596 18110 9608
rect 18233 9605 18245 9608
rect 18279 9605 18291 9639
rect 18233 9599 18291 9605
rect 20530 9596 20536 9648
rect 20588 9596 20594 9648
rect 22664 9636 22692 9676
rect 22738 9664 22744 9716
rect 22796 9664 22802 9716
rect 23842 9704 23848 9716
rect 22848 9676 23848 9704
rect 22848 9636 22876 9676
rect 23842 9664 23848 9676
rect 23900 9664 23906 9716
rect 26421 9707 26479 9713
rect 26421 9673 26433 9707
rect 26467 9704 26479 9707
rect 26878 9704 26884 9716
rect 26467 9676 26884 9704
rect 26467 9673 26479 9676
rect 26421 9667 26479 9673
rect 26878 9664 26884 9676
rect 26936 9664 26942 9716
rect 27706 9664 27712 9716
rect 27764 9704 27770 9716
rect 28445 9707 28503 9713
rect 28445 9704 28457 9707
rect 27764 9676 28457 9704
rect 27764 9664 27770 9676
rect 28445 9673 28457 9676
rect 28491 9673 28503 9707
rect 28997 9707 29055 9713
rect 28997 9704 29009 9707
rect 28445 9667 28503 9673
rect 28552 9676 29009 9704
rect 22664 9608 22876 9636
rect 23860 9636 23888 9664
rect 23860 9608 24256 9636
rect 16945 9540 17954 9568
rect 16945 9537 16957 9540
rect 16899 9531 16957 9537
rect 19150 9528 19156 9580
rect 19208 9528 19214 9580
rect 20714 9528 20720 9580
rect 20772 9568 20778 9580
rect 20772 9540 21036 9568
rect 20772 9528 20778 9540
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9500 13783 9503
rect 13814 9500 13820 9512
rect 13771 9472 13820 9500
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 14458 9460 14464 9512
rect 14516 9460 14522 9512
rect 15470 9460 15476 9512
rect 15528 9500 15534 9512
rect 16301 9503 16359 9509
rect 16301 9500 16313 9503
rect 15528 9472 16313 9500
rect 15528 9460 15534 9472
rect 16301 9469 16313 9472
rect 16347 9469 16359 9503
rect 16301 9463 16359 9469
rect 16390 9460 16396 9512
rect 16448 9460 16454 9512
rect 17129 9503 17187 9509
rect 17129 9469 17141 9503
rect 17175 9500 17187 9503
rect 18322 9500 18328 9512
rect 17175 9472 18328 9500
rect 17175 9469 17187 9472
rect 17129 9463 17187 9469
rect 18322 9460 18328 9472
rect 18380 9460 18386 9512
rect 18693 9503 18751 9509
rect 18693 9469 18705 9503
rect 18739 9469 18751 9503
rect 18693 9463 18751 9469
rect 19429 9503 19487 9509
rect 19429 9469 19441 9503
rect 19475 9500 19487 9503
rect 19794 9500 19800 9512
rect 19475 9472 19800 9500
rect 19475 9469 19487 9472
rect 19429 9463 19487 9469
rect 18046 9392 18052 9444
rect 18104 9432 18110 9444
rect 18708 9432 18736 9463
rect 19794 9460 19800 9472
rect 19852 9460 19858 9512
rect 20806 9460 20812 9512
rect 20864 9500 20870 9512
rect 20901 9503 20959 9509
rect 20901 9500 20913 9503
rect 20864 9472 20913 9500
rect 20864 9460 20870 9472
rect 20901 9469 20913 9472
rect 20947 9469 20959 9503
rect 21008 9500 21036 9540
rect 21082 9528 21088 9580
rect 21140 9568 21146 9580
rect 21364 9571 21422 9577
rect 21364 9568 21376 9571
rect 21140 9540 21376 9568
rect 21140 9528 21146 9540
rect 21364 9537 21376 9540
rect 21410 9537 21422 9571
rect 21364 9531 21422 9537
rect 21450 9528 21456 9580
rect 21508 9568 21514 9580
rect 22554 9568 22560 9580
rect 21508 9540 22560 9568
rect 21508 9528 21514 9540
rect 22554 9528 22560 9540
rect 22612 9568 22618 9580
rect 22612 9540 24072 9568
rect 22612 9528 22618 9540
rect 21637 9503 21695 9509
rect 21637 9500 21649 9503
rect 21008 9472 21649 9500
rect 20901 9463 20959 9469
rect 21637 9469 21649 9472
rect 21683 9469 21695 9503
rect 21637 9463 21695 9469
rect 22002 9460 22008 9512
rect 22060 9500 22066 9512
rect 24044 9509 24072 9540
rect 24228 9550 24256 9608
rect 28350 9596 28356 9648
rect 28408 9636 28414 9648
rect 28552 9636 28580 9676
rect 28997 9673 29009 9676
rect 29043 9673 29055 9707
rect 28997 9667 29055 9673
rect 28408 9608 28580 9636
rect 28408 9596 28414 9608
rect 24397 9571 24455 9577
rect 24397 9550 24409 9571
rect 24228 9537 24409 9550
rect 24443 9568 24455 9571
rect 24762 9568 24768 9580
rect 24443 9540 24768 9568
rect 24443 9537 24455 9540
rect 24228 9531 24455 9537
rect 24228 9522 24440 9531
rect 24762 9528 24768 9540
rect 24820 9528 24826 9580
rect 24854 9528 24860 9580
rect 24912 9568 24918 9580
rect 27068 9571 27126 9577
rect 27068 9568 27080 9571
rect 24912 9540 24957 9568
rect 25884 9540 27080 9568
rect 24912 9528 24918 9540
rect 23477 9503 23535 9509
rect 23477 9500 23489 9503
rect 22060 9472 23489 9500
rect 22060 9460 22066 9472
rect 23477 9469 23489 9472
rect 23523 9469 23535 9503
rect 23477 9463 23535 9469
rect 24029 9503 24087 9509
rect 24029 9469 24041 9503
rect 24075 9500 24087 9503
rect 24118 9500 24124 9512
rect 24075 9472 24124 9500
rect 24075 9469 24087 9472
rect 24029 9463 24087 9469
rect 23492 9432 23520 9463
rect 24118 9460 24124 9472
rect 24176 9460 24182 9512
rect 25133 9503 25191 9509
rect 24305 9479 24363 9485
rect 24305 9445 24317 9479
rect 24351 9445 24363 9479
rect 25133 9469 25145 9503
rect 25179 9500 25191 9503
rect 25406 9500 25412 9512
rect 25179 9472 25412 9500
rect 25179 9469 25191 9472
rect 25133 9463 25191 9469
rect 25406 9460 25412 9472
rect 25464 9460 25470 9512
rect 23658 9432 23664 9444
rect 18104 9404 18736 9432
rect 20088 9404 20668 9432
rect 23492 9404 23664 9432
rect 18104 9392 18110 9404
rect 15102 9364 15108 9376
rect 13648 9336 15108 9364
rect 12989 9327 13047 9333
rect 15102 9324 15108 9336
rect 15160 9324 15166 9376
rect 15378 9324 15384 9376
rect 15436 9364 15442 9376
rect 15565 9367 15623 9373
rect 15565 9364 15577 9367
rect 15436 9336 15577 9364
rect 15436 9324 15442 9336
rect 15565 9333 15577 9336
rect 15611 9333 15623 9367
rect 15565 9327 15623 9333
rect 16859 9367 16917 9373
rect 16859 9333 16871 9367
rect 16905 9364 16917 9367
rect 17034 9364 17040 9376
rect 16905 9336 17040 9364
rect 16905 9333 16917 9336
rect 16859 9327 16917 9333
rect 17034 9324 17040 9336
rect 17092 9364 17098 9376
rect 19159 9367 19217 9373
rect 19159 9364 19171 9367
rect 17092 9336 19171 9364
rect 17092 9324 17098 9336
rect 19159 9333 19171 9336
rect 19205 9364 19217 9367
rect 20088 9364 20116 9404
rect 19205 9336 20116 9364
rect 20640 9364 20668 9404
rect 23658 9392 23664 9404
rect 23716 9392 23722 9444
rect 24305 9439 24363 9445
rect 25884 9444 25912 9540
rect 27068 9537 27080 9540
rect 27114 9537 27126 9571
rect 27068 9531 27126 9537
rect 28534 9528 28540 9580
rect 28592 9568 28598 9580
rect 28592 9540 29500 9568
rect 28592 9528 28598 9540
rect 26050 9460 26056 9512
rect 26108 9500 26114 9512
rect 26605 9503 26663 9509
rect 26605 9500 26617 9503
rect 26108 9472 26617 9500
rect 26108 9460 26114 9472
rect 26605 9469 26617 9472
rect 26651 9469 26663 9503
rect 26605 9463 26663 9469
rect 26694 9460 26700 9512
rect 26752 9500 26758 9512
rect 27341 9503 27399 9509
rect 27341 9500 27353 9503
rect 26752 9472 27353 9500
rect 26752 9460 26758 9472
rect 27341 9469 27353 9472
rect 27387 9469 27399 9503
rect 29178 9500 29184 9512
rect 27341 9463 27399 9469
rect 29012 9472 29184 9500
rect 29012 9444 29040 9472
rect 29178 9460 29184 9472
rect 29236 9460 29242 9512
rect 29472 9509 29500 9540
rect 29457 9503 29515 9509
rect 29457 9469 29469 9503
rect 29503 9469 29515 9503
rect 29457 9463 29515 9469
rect 24326 9376 24354 9439
rect 25866 9392 25872 9444
rect 25924 9392 25930 9444
rect 28994 9392 29000 9444
rect 29052 9392 29058 9444
rect 29472 9376 29500 9463
rect 21367 9367 21425 9373
rect 21367 9364 21379 9367
rect 20640 9336 21379 9364
rect 19205 9333 19217 9336
rect 19159 9327 19217 9333
rect 21367 9333 21379 9336
rect 21413 9364 21425 9367
rect 21542 9364 21548 9376
rect 21413 9336 21548 9364
rect 21413 9333 21425 9336
rect 21367 9327 21425 9333
rect 21542 9324 21548 9336
rect 21600 9324 21606 9376
rect 23293 9367 23351 9373
rect 23293 9333 23305 9367
rect 23339 9364 23351 9367
rect 23750 9364 23756 9376
rect 23339 9336 23756 9364
rect 23339 9333 23351 9336
rect 23293 9327 23351 9333
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 23845 9367 23903 9373
rect 23845 9333 23857 9367
rect 23891 9364 23903 9367
rect 23934 9364 23940 9376
rect 23891 9336 23940 9364
rect 23891 9333 23903 9336
rect 23845 9327 23903 9333
rect 23934 9324 23940 9336
rect 23992 9324 23998 9376
rect 24118 9324 24124 9376
rect 24176 9324 24182 9376
rect 24302 9324 24308 9376
rect 24360 9324 24366 9376
rect 24394 9324 24400 9376
rect 24452 9364 24458 9376
rect 24863 9367 24921 9373
rect 24863 9364 24875 9367
rect 24452 9336 24875 9364
rect 24452 9324 24458 9336
rect 24863 9333 24875 9336
rect 24909 9364 24921 9367
rect 26878 9364 26884 9376
rect 24909 9336 26884 9364
rect 24909 9333 24921 9336
rect 24863 9327 24921 9333
rect 26878 9324 26884 9336
rect 26936 9364 26942 9376
rect 27071 9367 27129 9373
rect 27071 9364 27083 9367
rect 26936 9336 27083 9364
rect 26936 9324 26942 9336
rect 27071 9333 27083 9336
rect 27117 9333 27129 9367
rect 27071 9327 27129 9333
rect 27338 9324 27344 9376
rect 27396 9364 27402 9376
rect 29273 9367 29331 9373
rect 29273 9364 29285 9367
rect 27396 9336 29285 9364
rect 27396 9324 27402 9336
rect 29273 9333 29285 9336
rect 29319 9333 29331 9367
rect 29273 9327 29331 9333
rect 29454 9324 29460 9376
rect 29512 9324 29518 9376
rect 552 9274 31072 9296
rect 552 9222 7988 9274
rect 8040 9222 8052 9274
rect 8104 9222 8116 9274
rect 8168 9222 8180 9274
rect 8232 9222 8244 9274
rect 8296 9222 15578 9274
rect 15630 9222 15642 9274
rect 15694 9222 15706 9274
rect 15758 9222 15770 9274
rect 15822 9222 15834 9274
rect 15886 9222 23168 9274
rect 23220 9222 23232 9274
rect 23284 9222 23296 9274
rect 23348 9222 23360 9274
rect 23412 9222 23424 9274
rect 23476 9222 30758 9274
rect 30810 9222 30822 9274
rect 30874 9222 30886 9274
rect 30938 9222 30950 9274
rect 31002 9222 31014 9274
rect 31066 9222 31072 9274
rect 552 9200 31072 9222
rect 842 9120 848 9172
rect 900 9120 906 9172
rect 4246 9160 4252 9172
rect 1044 9132 4252 9160
rect 750 8984 756 9036
rect 808 8984 814 9036
rect 1044 9033 1072 9132
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 4617 9163 4675 9169
rect 4617 9160 4629 9163
rect 4396 9132 4629 9160
rect 4396 9120 4402 9132
rect 4617 9129 4629 9132
rect 4663 9129 4675 9163
rect 4617 9123 4675 9129
rect 4890 9120 4896 9172
rect 4948 9120 4954 9172
rect 5166 9120 5172 9172
rect 5224 9120 5230 9172
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 6178 9160 6184 9172
rect 5491 9132 6184 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 7377 9163 7435 9169
rect 7377 9160 7389 9163
rect 7156 9132 7389 9160
rect 7156 9120 7162 9132
rect 7377 9129 7389 9132
rect 7423 9129 7435 9163
rect 7377 9123 7435 9129
rect 7466 9120 7472 9172
rect 7524 9120 7530 9172
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 8110 9160 8116 9172
rect 7708 9132 8116 9160
rect 7708 9120 7714 9132
rect 8110 9120 8116 9132
rect 8168 9120 8174 9172
rect 9490 9120 9496 9172
rect 9548 9120 9554 9172
rect 9861 9163 9919 9169
rect 9861 9129 9873 9163
rect 9907 9160 9919 9163
rect 10502 9160 10508 9172
rect 9907 9132 10508 9160
rect 9907 9129 9919 9132
rect 9861 9123 9919 9129
rect 10502 9120 10508 9132
rect 10560 9120 10566 9172
rect 10597 9163 10655 9169
rect 10597 9129 10609 9163
rect 10643 9160 10655 9163
rect 11882 9160 11888 9172
rect 10643 9132 11888 9160
rect 10643 9129 10655 9132
rect 10597 9123 10655 9129
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 14090 9120 14096 9172
rect 14148 9160 14154 9172
rect 14283 9163 14341 9169
rect 14283 9160 14295 9163
rect 14148 9132 14295 9160
rect 14148 9120 14154 9132
rect 14283 9129 14295 9132
rect 14329 9129 14341 9163
rect 14283 9123 14341 9129
rect 14458 9120 14464 9172
rect 14516 9160 14522 9172
rect 16117 9163 16175 9169
rect 16117 9160 16129 9163
rect 14516 9132 16129 9160
rect 14516 9120 14522 9132
rect 16117 9129 16129 9132
rect 16163 9129 16175 9163
rect 16117 9123 16175 9129
rect 16390 9120 16396 9172
rect 16448 9120 16454 9172
rect 17034 9120 17040 9172
rect 17092 9160 17098 9172
rect 17871 9163 17929 9169
rect 17871 9160 17883 9163
rect 17092 9132 17883 9160
rect 17092 9120 17098 9132
rect 1394 9052 1400 9104
rect 1452 9092 1458 9104
rect 1949 9095 2007 9101
rect 1949 9092 1961 9095
rect 1452 9064 1961 9092
rect 1452 9052 1458 9064
rect 1949 9061 1961 9064
rect 1995 9061 2007 9095
rect 7484 9092 7512 9120
rect 1949 9055 2007 9061
rect 4816 9064 6040 9092
rect 1029 9027 1087 9033
rect 1029 8993 1041 9027
rect 1075 8993 1087 9027
rect 1029 8987 1087 8993
rect 1121 9027 1179 9033
rect 1121 8993 1133 9027
rect 1167 9024 1179 9027
rect 1673 9027 1731 9033
rect 1673 9024 1685 9027
rect 1167 8996 1685 9024
rect 1167 8993 1179 8996
rect 1121 8987 1179 8993
rect 1673 8993 1685 8996
rect 1719 9024 1731 9027
rect 2038 9024 2044 9036
rect 1719 8996 2044 9024
rect 1719 8993 1731 8996
rect 1673 8987 1731 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 2314 8984 2320 9036
rect 2372 9024 2378 9036
rect 2552 9027 2610 9033
rect 2552 9024 2564 9027
rect 2372 8996 2564 9024
rect 2372 8984 2378 8996
rect 2552 8993 2564 8996
rect 2598 9024 2610 9027
rect 3602 9024 3608 9036
rect 2598 8996 3608 9024
rect 2598 8993 2610 8996
rect 2552 8987 2610 8993
rect 3602 8984 3608 8996
rect 3660 8984 3666 9036
rect 4816 9033 4844 9064
rect 4801 9027 4859 9033
rect 4801 9024 4813 9027
rect 4080 8996 4813 9024
rect 768 8888 796 8984
rect 4080 8968 4108 8996
rect 4801 8993 4813 8996
rect 4847 8993 4859 9027
rect 4801 8987 4859 8993
rect 5077 9027 5135 9033
rect 5077 8993 5089 9027
rect 5123 8993 5135 9027
rect 5077 8987 5135 8993
rect 1394 8916 1400 8968
rect 1452 8916 1458 8968
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 2731 8959 2789 8965
rect 2731 8925 2743 8959
rect 2777 8956 2789 8959
rect 2866 8956 2872 8968
rect 2777 8928 2872 8956
rect 2777 8925 2789 8928
rect 2731 8919 2789 8925
rect 2240 8888 2268 8919
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 2958 8916 2964 8968
rect 3016 8916 3022 8968
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 3108 8928 4022 8956
rect 3108 8916 3114 8928
rect 768 8860 2268 8888
rect 3994 8888 4022 8928
rect 4062 8916 4068 8968
rect 4120 8916 4126 8968
rect 5092 8956 5120 8987
rect 5350 8984 5356 9036
rect 5408 8984 5414 9036
rect 6012 9033 6040 9064
rect 6380 9064 7420 9092
rect 7484 9064 7788 9092
rect 6380 9033 6408 9064
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 8993 5687 9027
rect 5629 8987 5687 8993
rect 5997 9027 6055 9033
rect 5997 8993 6009 9027
rect 6043 8993 6055 9027
rect 5997 8987 6055 8993
rect 6365 9027 6423 9033
rect 6365 8993 6377 9027
rect 6411 8993 6423 9027
rect 6365 8987 6423 8993
rect 5644 8956 5672 8987
rect 5092 8928 5672 8956
rect 6012 8956 6040 8987
rect 6086 8956 6092 8968
rect 6012 8928 6092 8956
rect 5092 8888 5120 8928
rect 3994 8860 5120 8888
rect 5644 8888 5672 8928
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 6380 8888 6408 8987
rect 6638 8984 6644 9036
rect 6696 8984 6702 9036
rect 6914 8984 6920 9036
rect 6972 8984 6978 9036
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 9024 7251 9027
rect 7282 9024 7288 9036
rect 7239 8996 7288 9024
rect 7239 8993 7251 8996
rect 7193 8987 7251 8993
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 7392 9024 7420 9064
rect 7466 9024 7472 9036
rect 7392 8996 7472 9024
rect 7466 8984 7472 8996
rect 7524 9024 7530 9036
rect 7561 9027 7619 9033
rect 7561 9024 7573 9027
rect 7524 8996 7573 9024
rect 7524 8984 7530 8996
rect 7561 8993 7573 8996
rect 7607 8993 7619 9027
rect 7561 8987 7619 8993
rect 7650 8984 7656 9036
rect 7708 8984 7714 9036
rect 7760 9024 7788 9064
rect 9398 9052 9404 9104
rect 9456 9092 9462 9104
rect 11238 9092 11244 9104
rect 9456 9064 11244 9092
rect 9456 9052 9462 9064
rect 7980 9027 8038 9033
rect 7980 9024 7992 9027
rect 7760 8996 7992 9024
rect 7980 8993 7992 8996
rect 8026 8993 8038 9027
rect 7980 8987 8038 8993
rect 8202 8984 8208 9036
rect 8260 9024 8266 9036
rect 8389 9027 8447 9033
rect 8389 9024 8401 9027
rect 8260 8996 8401 9024
rect 8260 8984 8266 8996
rect 8389 8993 8401 8996
rect 8435 8993 8447 9027
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 8389 8987 8447 8993
rect 9784 8996 10057 9024
rect 6454 8916 6460 8968
rect 6512 8956 6518 8968
rect 7668 8956 7696 8984
rect 6512 8928 7696 8956
rect 6512 8916 6518 8928
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 8168 8928 8213 8956
rect 8168 8916 8174 8928
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 9490 8956 9496 8968
rect 8812 8928 9496 8956
rect 8812 8916 8818 8928
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 9784 8900 9812 8996
rect 10045 8993 10057 8996
rect 10091 9024 10103 9027
rect 10226 9024 10232 9036
rect 10091 8996 10232 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 10520 9033 10548 9064
rect 11238 9052 11244 9064
rect 11296 9052 11302 9104
rect 13449 9095 13507 9101
rect 13449 9061 13461 9095
rect 13495 9092 13507 9095
rect 13495 9064 13952 9092
rect 13495 9061 13507 9064
rect 13449 9055 13507 9061
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 10778 8984 10784 9036
rect 10836 8984 10842 9036
rect 11885 9027 11943 9033
rect 11885 9024 11897 9027
rect 11072 8996 11897 9024
rect 5644 8860 6408 8888
rect 6932 8860 7236 8888
rect 2240 8820 2268 8860
rect 6932 8832 6960 8860
rect 2774 8820 2780 8832
rect 2240 8792 2780 8820
rect 2774 8780 2780 8792
rect 2832 8780 2838 8832
rect 3326 8780 3332 8832
rect 3384 8820 3390 8832
rect 4065 8823 4123 8829
rect 4065 8820 4077 8823
rect 3384 8792 4077 8820
rect 3384 8780 3390 8792
rect 4065 8789 4077 8792
rect 4111 8789 4123 8823
rect 4065 8783 4123 8789
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 5626 8820 5632 8832
rect 5408 8792 5632 8820
rect 5408 8780 5414 8792
rect 5626 8780 5632 8792
rect 5684 8780 5690 8832
rect 5810 8780 5816 8832
rect 5868 8780 5874 8832
rect 5994 8780 6000 8832
rect 6052 8820 6058 8832
rect 6181 8823 6239 8829
rect 6181 8820 6193 8823
rect 6052 8792 6193 8820
rect 6052 8780 6058 8792
rect 6181 8789 6193 8792
rect 6227 8789 6239 8823
rect 6181 8783 6239 8789
rect 6454 8780 6460 8832
rect 6512 8780 6518 8832
rect 6733 8823 6791 8829
rect 6733 8789 6745 8823
rect 6779 8820 6791 8823
rect 6822 8820 6828 8832
rect 6779 8792 6828 8820
rect 6779 8789 6791 8792
rect 6733 8783 6791 8789
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 6914 8780 6920 8832
rect 6972 8780 6978 8832
rect 7009 8823 7067 8829
rect 7009 8789 7021 8823
rect 7055 8820 7067 8823
rect 7098 8820 7104 8832
rect 7055 8792 7104 8820
rect 7055 8789 7067 8792
rect 7009 8783 7067 8789
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 7208 8820 7236 8860
rect 9766 8848 9772 8900
rect 9824 8848 9830 8900
rect 10321 8891 10379 8897
rect 10321 8857 10333 8891
rect 10367 8888 10379 8891
rect 11072 8888 11100 8996
rect 11885 8993 11897 8996
rect 11931 8993 11943 9027
rect 11885 8987 11943 8993
rect 13814 8984 13820 9036
rect 13872 8984 13878 9036
rect 13924 9024 13952 9064
rect 15930 9052 15936 9104
rect 15988 9092 15994 9104
rect 16408 9092 16436 9120
rect 17144 9101 17172 9132
rect 17871 9129 17883 9132
rect 17917 9129 17929 9163
rect 17871 9123 17929 9129
rect 18046 9120 18052 9172
rect 18104 9160 18110 9172
rect 18104 9132 19288 9160
rect 18104 9120 18110 9132
rect 17129 9095 17187 9101
rect 15988 9064 16344 9092
rect 16408 9064 17080 9092
rect 15988 9052 15994 9064
rect 14553 9027 14611 9033
rect 13924 8996 14044 9024
rect 14016 8968 14044 8996
rect 14553 8993 14565 9027
rect 14599 9024 14611 9027
rect 16022 9024 16028 9036
rect 14599 8996 16028 9024
rect 14599 8993 14611 8996
rect 14553 8987 14611 8993
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 16316 9033 16344 9064
rect 16301 9027 16359 9033
rect 16301 8993 16313 9027
rect 16347 8993 16359 9027
rect 16301 8987 16359 8993
rect 16577 9027 16635 9033
rect 16577 8993 16589 9027
rect 16623 8993 16635 9027
rect 16577 8987 16635 8993
rect 14313 8977 14371 8983
rect 14313 8974 14325 8977
rect 11146 8916 11152 8968
rect 11204 8916 11210 8968
rect 11514 8965 11520 8968
rect 11476 8959 11520 8965
rect 11476 8925 11488 8959
rect 11476 8919 11520 8925
rect 11514 8916 11520 8919
rect 11572 8916 11578 8968
rect 11612 8961 11670 8967
rect 11612 8927 11624 8961
rect 11658 8956 11670 8961
rect 11698 8956 11704 8968
rect 11658 8928 11704 8956
rect 11658 8927 11670 8928
rect 11612 8921 11670 8927
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 13998 8916 14004 8968
rect 14056 8916 14062 8968
rect 14298 8943 14325 8974
rect 14359 8968 14371 8977
rect 14359 8943 14372 8968
rect 14298 8928 14372 8943
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 15470 8916 15476 8968
rect 15528 8956 15534 8968
rect 16592 8956 16620 8987
rect 16850 8984 16856 9036
rect 16908 8984 16914 9036
rect 17052 9024 17080 9064
rect 17129 9061 17141 9095
rect 17175 9061 17187 9095
rect 19260 9092 19288 9132
rect 21542 9120 21548 9172
rect 21600 9160 21606 9172
rect 21735 9163 21793 9169
rect 21735 9160 21747 9163
rect 21600 9132 21747 9160
rect 21600 9120 21606 9132
rect 21735 9129 21747 9132
rect 21781 9160 21793 9163
rect 21781 9132 22876 9160
rect 21781 9129 21793 9132
rect 21735 9123 21793 9129
rect 19705 9095 19763 9101
rect 19705 9092 19717 9095
rect 19260 9064 19717 9092
rect 17129 9055 17187 9061
rect 19705 9061 19717 9064
rect 19751 9092 19763 9095
rect 20806 9092 20812 9104
rect 19751 9064 20812 9092
rect 19751 9061 19763 9064
rect 19705 9055 19763 9061
rect 20806 9052 20812 9064
rect 20864 9092 20870 9104
rect 20864 9064 21312 9092
rect 20864 9052 20870 9064
rect 17405 9027 17463 9033
rect 17405 9024 17417 9027
rect 17052 8996 17417 9024
rect 17405 8993 17417 8996
rect 17451 9024 17463 9027
rect 18046 9024 18052 9036
rect 17451 8996 18052 9024
rect 17451 8993 17463 8996
rect 17405 8987 17463 8993
rect 18046 8984 18052 8996
rect 18104 8984 18110 9036
rect 18138 8984 18144 9036
rect 18196 8984 18202 9036
rect 21284 9033 21312 9064
rect 21269 9027 21327 9033
rect 21269 8993 21281 9027
rect 21315 8993 21327 9027
rect 22848 9024 22876 9132
rect 22922 9120 22928 9172
rect 22980 9160 22986 9172
rect 23109 9163 23167 9169
rect 23109 9160 23121 9163
rect 22980 9132 23121 9160
rect 22980 9120 22986 9132
rect 23109 9129 23121 9132
rect 23155 9129 23167 9163
rect 23109 9123 23167 9129
rect 23750 9120 23756 9172
rect 23808 9160 23814 9172
rect 24210 9160 24216 9172
rect 23808 9132 24216 9160
rect 23808 9120 23814 9132
rect 24210 9120 24216 9132
rect 24268 9120 24274 9172
rect 24854 9120 24860 9172
rect 24912 9160 24918 9172
rect 25317 9163 25375 9169
rect 25317 9160 25329 9163
rect 24912 9132 25329 9160
rect 24912 9120 24918 9132
rect 25317 9129 25329 9132
rect 25363 9129 25375 9163
rect 25317 9123 25375 9129
rect 25406 9120 25412 9172
rect 25464 9160 25470 9172
rect 25685 9163 25743 9169
rect 25685 9160 25697 9163
rect 25464 9132 25697 9160
rect 25464 9120 25470 9132
rect 25685 9129 25697 9132
rect 25731 9129 25743 9163
rect 25685 9123 25743 9129
rect 25961 9163 26019 9169
rect 25961 9129 25973 9163
rect 26007 9160 26019 9163
rect 26694 9160 26700 9172
rect 26007 9132 26700 9160
rect 26007 9129 26019 9132
rect 25961 9123 26019 9129
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 26878 9120 26884 9172
rect 26936 9169 26942 9172
rect 26936 9160 26945 9169
rect 26936 9132 26981 9160
rect 26936 9123 26945 9132
rect 26936 9120 26942 9123
rect 27522 9120 27528 9172
rect 27580 9160 27586 9172
rect 28261 9163 28319 9169
rect 28261 9160 28273 9163
rect 27580 9132 28273 9160
rect 27580 9120 27586 9132
rect 28261 9129 28273 9132
rect 28307 9129 28319 9163
rect 28261 9123 28319 9129
rect 30193 9163 30251 9169
rect 30193 9129 30205 9163
rect 30239 9160 30251 9163
rect 30466 9160 30472 9172
rect 30239 9132 30472 9160
rect 30239 9129 30251 9132
rect 30193 9123 30251 9129
rect 30466 9120 30472 9132
rect 30524 9120 30530 9172
rect 26050 9052 26056 9104
rect 26108 9092 26114 9104
rect 26108 9064 26464 9092
rect 26108 9052 26114 9064
rect 22848 8996 23612 9024
rect 21269 8987 21327 8993
rect 15528 8928 16620 8956
rect 17911 8959 17969 8965
rect 15528 8916 15534 8928
rect 17911 8925 17923 8959
rect 17957 8956 17969 8959
rect 20162 8956 20168 8968
rect 17957 8928 20168 8956
rect 17957 8925 17969 8928
rect 17911 8919 17969 8925
rect 20162 8916 20168 8928
rect 20220 8916 20226 8968
rect 10367 8860 11100 8888
rect 10367 8857 10379 8860
rect 10321 8851 10379 8857
rect 11054 8820 11060 8832
rect 7208 8792 11060 8820
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 11164 8820 11192 8916
rect 18966 8848 18972 8900
rect 19024 8888 19030 8900
rect 19981 8891 20039 8897
rect 19981 8888 19993 8891
rect 19024 8860 19993 8888
rect 19024 8848 19030 8860
rect 19981 8857 19993 8860
rect 20027 8888 20039 8891
rect 20027 8860 20760 8888
rect 20027 8857 20039 8860
rect 19981 8851 20039 8857
rect 20732 8832 20760 8860
rect 12250 8820 12256 8832
rect 11164 8792 12256 8820
rect 12250 8780 12256 8792
rect 12308 8780 12314 8832
rect 12986 8780 12992 8832
rect 13044 8780 13050 8832
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 13412 8792 13553 8820
rect 13412 8780 13418 8792
rect 13541 8789 13553 8792
rect 13587 8789 13599 8823
rect 13541 8783 13599 8789
rect 14366 8780 14372 8832
rect 14424 8820 14430 8832
rect 15657 8823 15715 8829
rect 15657 8820 15669 8823
rect 14424 8792 15669 8820
rect 14424 8780 14430 8792
rect 15657 8789 15669 8792
rect 15703 8789 15715 8823
rect 15657 8783 15715 8789
rect 16022 8780 16028 8832
rect 16080 8820 16086 8832
rect 16393 8823 16451 8829
rect 16393 8820 16405 8823
rect 16080 8792 16405 8820
rect 16080 8780 16086 8792
rect 16393 8789 16405 8792
rect 16439 8789 16451 8823
rect 16393 8783 16451 8789
rect 18782 8780 18788 8832
rect 18840 8820 18846 8832
rect 19245 8823 19303 8829
rect 19245 8820 19257 8823
rect 18840 8792 19257 8820
rect 18840 8780 18846 8792
rect 19245 8789 19257 8792
rect 19291 8789 19303 8823
rect 19245 8783 19303 8789
rect 20441 8823 20499 8829
rect 20441 8789 20453 8823
rect 20487 8820 20499 8823
rect 20622 8820 20628 8832
rect 20487 8792 20628 8820
rect 20487 8789 20499 8792
rect 20441 8783 20499 8789
rect 20622 8780 20628 8792
rect 20680 8780 20686 8832
rect 20714 8780 20720 8832
rect 20772 8780 20778 8832
rect 21284 8820 21312 8987
rect 21818 8967 21824 8968
rect 21775 8961 21824 8967
rect 21775 8927 21787 8961
rect 21821 8927 21824 8961
rect 21775 8921 21824 8927
rect 21818 8916 21824 8921
rect 21876 8916 21882 8968
rect 21910 8916 21916 8968
rect 21968 8956 21974 8968
rect 22005 8959 22063 8965
rect 22005 8956 22017 8959
rect 21968 8928 22017 8956
rect 21968 8916 21974 8928
rect 22005 8925 22017 8928
rect 22051 8925 22063 8959
rect 23467 8959 23525 8965
rect 23467 8956 23479 8959
rect 22005 8919 22063 8925
rect 23400 8928 23479 8956
rect 23400 8820 23428 8928
rect 23467 8925 23479 8928
rect 23513 8925 23525 8959
rect 23584 8956 23612 8996
rect 24210 8984 24216 9036
rect 24268 8984 24274 9036
rect 25869 9027 25927 9033
rect 25869 8993 25881 9027
rect 25915 8993 25927 9027
rect 25869 8987 25927 8993
rect 23658 8956 23664 8968
rect 23584 8928 23664 8956
rect 23467 8919 23525 8925
rect 23658 8916 23664 8928
rect 23716 8956 23722 8968
rect 24026 8965 24032 8968
rect 23804 8959 23862 8965
rect 23804 8956 23816 8959
rect 23716 8928 23816 8956
rect 23716 8916 23722 8928
rect 23804 8925 23816 8928
rect 23850 8925 23862 8959
rect 23804 8919 23862 8925
rect 23983 8959 24032 8965
rect 23983 8925 23995 8959
rect 24029 8925 24032 8959
rect 23983 8919 24032 8925
rect 24026 8916 24032 8919
rect 24084 8916 24090 8968
rect 23474 8820 23480 8832
rect 21284 8792 23480 8820
rect 23474 8780 23480 8792
rect 23532 8780 23538 8832
rect 23750 8780 23756 8832
rect 23808 8820 23814 8832
rect 25884 8820 25912 8987
rect 25958 8984 25964 9036
rect 26016 9024 26022 9036
rect 26436 9033 26464 9064
rect 26145 9027 26203 9033
rect 26145 9024 26157 9027
rect 26016 8996 26157 9024
rect 26016 8984 26022 8996
rect 26145 8993 26157 8996
rect 26191 8993 26203 9027
rect 26145 8987 26203 8993
rect 26421 9027 26479 9033
rect 26421 8993 26433 9027
rect 26467 8993 26479 9027
rect 26421 8987 26479 8993
rect 26160 8956 26188 8987
rect 26510 8984 26516 9036
rect 26568 9024 26574 9036
rect 27157 9027 27215 9033
rect 27157 9024 27169 9027
rect 26568 8996 27169 9024
rect 26568 8984 26574 8996
rect 27157 8993 27169 8996
rect 27203 8993 27215 9027
rect 27157 8987 27215 8993
rect 28626 8984 28632 9036
rect 28684 8984 28690 9036
rect 28905 9027 28963 9033
rect 28905 8993 28917 9027
rect 28951 9024 28963 9027
rect 30006 9024 30012 9036
rect 28951 8996 30012 9024
rect 28951 8993 28963 8996
rect 28905 8987 28963 8993
rect 30006 8984 30012 8996
rect 30064 8984 30070 9036
rect 26694 8956 26700 8968
rect 26160 8928 26700 8956
rect 26694 8916 26700 8928
rect 26752 8916 26758 8968
rect 26878 8916 26884 8968
rect 26936 8916 26942 8968
rect 27338 8916 27344 8968
rect 27396 8956 27402 8968
rect 28534 8956 28540 8968
rect 27396 8928 28540 8956
rect 27396 8916 27402 8928
rect 28534 8916 28540 8928
rect 28592 8916 28598 8968
rect 28994 8820 29000 8832
rect 23808 8792 29000 8820
rect 23808 8780 23814 8792
rect 28994 8780 29000 8792
rect 29052 8780 29058 8832
rect 552 8730 30912 8752
rect 552 8678 4193 8730
rect 4245 8678 4257 8730
rect 4309 8678 4321 8730
rect 4373 8678 4385 8730
rect 4437 8678 4449 8730
rect 4501 8678 11783 8730
rect 11835 8678 11847 8730
rect 11899 8678 11911 8730
rect 11963 8678 11975 8730
rect 12027 8678 12039 8730
rect 12091 8678 19373 8730
rect 19425 8678 19437 8730
rect 19489 8678 19501 8730
rect 19553 8678 19565 8730
rect 19617 8678 19629 8730
rect 19681 8678 26963 8730
rect 27015 8678 27027 8730
rect 27079 8678 27091 8730
rect 27143 8678 27155 8730
rect 27207 8678 27219 8730
rect 27271 8678 30912 8730
rect 552 8656 30912 8678
rect 1118 8576 1124 8628
rect 1176 8616 1182 8628
rect 1176 8588 2820 8616
rect 1176 8576 1182 8588
rect 2792 8548 2820 8588
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 5077 8619 5135 8625
rect 5077 8616 5089 8619
rect 2924 8588 5089 8616
rect 2924 8576 2930 8588
rect 5077 8585 5089 8588
rect 5123 8585 5135 8619
rect 6638 8616 6644 8628
rect 5077 8579 5135 8585
rect 5552 8588 6644 8616
rect 3050 8548 3056 8560
rect 2792 8520 3056 8548
rect 3050 8508 3056 8520
rect 3108 8508 3114 8560
rect 1443 8483 1501 8489
rect 1443 8449 1455 8483
rect 1489 8480 1501 8483
rect 1489 8452 3372 8480
rect 1489 8449 1501 8452
rect 1443 8443 1501 8449
rect 937 8415 995 8421
rect 937 8381 949 8415
rect 983 8412 995 8415
rect 1210 8412 1216 8424
rect 983 8384 1216 8412
rect 983 8381 995 8384
rect 937 8375 995 8381
rect 1210 8372 1216 8384
rect 1268 8372 1274 8424
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 1762 8412 1768 8424
rect 1719 8384 1768 8412
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 1762 8372 1768 8384
rect 1820 8372 1826 8424
rect 2130 8372 2136 8424
rect 2188 8412 2194 8424
rect 2682 8412 2688 8424
rect 2188 8384 2688 8412
rect 2188 8372 2194 8384
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 3237 8415 3295 8421
rect 3237 8412 3249 8415
rect 2832 8384 3249 8412
rect 2832 8372 2838 8384
rect 3237 8381 3249 8384
rect 3283 8381 3295 8415
rect 3344 8412 3372 8452
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 3700 8483 3758 8489
rect 3700 8480 3712 8483
rect 3476 8452 3712 8480
rect 3476 8440 3482 8452
rect 3700 8449 3712 8452
rect 3746 8449 3758 8483
rect 5552 8480 5580 8588
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 7006 8576 7012 8628
rect 7064 8616 7070 8628
rect 7377 8619 7435 8625
rect 7377 8616 7389 8619
rect 7064 8588 7389 8616
rect 7064 8576 7070 8588
rect 7377 8585 7389 8588
rect 7423 8585 7435 8619
rect 7377 8579 7435 8585
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7616 8588 8033 8616
rect 7616 8576 7622 8588
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 10042 8616 10048 8628
rect 8021 8579 8079 8585
rect 8680 8588 9076 8616
rect 7190 8508 7196 8560
rect 7248 8548 7254 8560
rect 8389 8551 8447 8557
rect 8389 8548 8401 8551
rect 7248 8520 8401 8548
rect 7248 8508 7254 8520
rect 8389 8517 8401 8520
rect 8435 8517 8447 8551
rect 8680 8548 8708 8588
rect 9048 8560 9076 8588
rect 9232 8588 10048 8616
rect 8389 8511 8447 8517
rect 8588 8520 8708 8548
rect 6000 8483 6058 8489
rect 6000 8480 6012 8483
rect 3700 8443 3758 8449
rect 3804 8452 5580 8480
rect 5644 8452 6012 8480
rect 3804 8412 3832 8452
rect 3344 8384 3832 8412
rect 3973 8415 4031 8421
rect 3237 8375 3295 8381
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 5350 8412 5356 8424
rect 4019 8384 5356 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 5442 8372 5448 8424
rect 5500 8372 5506 8424
rect 5534 8372 5540 8424
rect 5592 8372 5598 8424
rect 3050 8304 3056 8356
rect 3108 8304 3114 8356
rect 3326 8344 3332 8356
rect 3160 8316 3332 8344
rect 1394 8236 1400 8288
rect 1452 8285 1458 8288
rect 1452 8276 1461 8285
rect 1452 8248 1497 8276
rect 1452 8239 1461 8248
rect 1452 8236 1458 8239
rect 2314 8236 2320 8288
rect 2372 8276 2378 8288
rect 3160 8276 3188 8316
rect 3326 8304 3332 8316
rect 3384 8304 3390 8356
rect 5460 8344 5488 8372
rect 5644 8344 5672 8452
rect 6000 8449 6012 8452
rect 6046 8449 6058 8483
rect 6000 8443 6058 8449
rect 6086 8440 6092 8492
rect 6144 8480 6150 8492
rect 6144 8452 8248 8480
rect 6144 8440 6150 8452
rect 5902 8421 5908 8424
rect 5864 8415 5908 8421
rect 5864 8381 5876 8415
rect 5864 8375 5908 8381
rect 5902 8372 5908 8375
rect 5960 8372 5966 8424
rect 6178 8372 6184 8424
rect 6236 8412 6242 8424
rect 8220 8421 8248 8452
rect 6273 8415 6331 8421
rect 6273 8412 6285 8415
rect 6236 8384 6285 8412
rect 6236 8372 6242 8384
rect 6273 8381 6285 8384
rect 6319 8381 6331 8415
rect 6273 8375 6331 8381
rect 7929 8415 7987 8421
rect 7929 8381 7941 8415
rect 7975 8412 7987 8415
rect 8205 8415 8263 8421
rect 7975 8384 8156 8412
rect 7975 8381 7987 8384
rect 7929 8375 7987 8381
rect 5460 8316 5672 8344
rect 8128 8344 8156 8384
rect 8205 8381 8217 8415
rect 8251 8412 8263 8415
rect 8386 8412 8392 8424
rect 8251 8384 8392 8412
rect 8251 8381 8263 8384
rect 8205 8375 8263 8381
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 8588 8421 8616 8520
rect 8846 8508 8852 8560
rect 8904 8508 8910 8560
rect 9030 8508 9036 8560
rect 9088 8508 9094 8560
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 8665 8415 8723 8421
rect 8665 8381 8677 8415
rect 8711 8412 8723 8415
rect 9232 8412 9260 8588
rect 10042 8576 10048 8588
rect 10100 8616 10106 8628
rect 10778 8616 10784 8628
rect 10100 8588 10784 8616
rect 10100 8576 10106 8588
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 11698 8576 11704 8628
rect 11756 8576 11762 8628
rect 19242 8576 19248 8628
rect 19300 8616 19306 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 19300 8588 20545 8616
rect 19300 8576 19306 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 20533 8579 20591 8585
rect 23400 8588 25452 8616
rect 9306 8508 9312 8560
rect 9364 8548 9370 8560
rect 9401 8551 9459 8557
rect 9401 8548 9413 8551
rect 9364 8520 9413 8548
rect 9364 8508 9370 8520
rect 9401 8517 9413 8520
rect 9447 8517 9459 8551
rect 9401 8511 9459 8517
rect 9490 8508 9496 8560
rect 9548 8548 9554 8560
rect 21269 8551 21327 8557
rect 9548 8520 9674 8548
rect 9548 8508 9554 8520
rect 9646 8480 9674 8520
rect 12176 8520 13124 8548
rect 12176 8492 12204 8520
rect 10140 8483 10198 8489
rect 10140 8480 10152 8483
rect 9646 8452 10152 8480
rect 10140 8449 10152 8452
rect 10186 8449 10198 8483
rect 10140 8443 10198 8449
rect 12158 8440 12164 8492
rect 12216 8440 12222 8492
rect 12710 8440 12716 8492
rect 12768 8440 12774 8492
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 8711 8384 8892 8412
rect 9232 8384 9321 8412
rect 8711 8381 8723 8384
rect 8665 8375 8723 8381
rect 8864 8344 8892 8384
rect 9309 8381 9321 8384
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 9398 8372 9404 8424
rect 9456 8372 9462 8424
rect 9490 8372 9496 8424
rect 9548 8412 9554 8424
rect 9585 8415 9643 8421
rect 9585 8412 9597 8415
rect 9548 8384 9597 8412
rect 9548 8372 9554 8384
rect 9585 8381 9597 8384
rect 9631 8381 9643 8415
rect 9585 8375 9643 8381
rect 9674 8372 9680 8424
rect 9732 8372 9738 8424
rect 9950 8372 9956 8424
rect 10008 8412 10014 8424
rect 10413 8415 10471 8421
rect 10413 8412 10425 8415
rect 10008 8384 10425 8412
rect 10008 8372 10014 8384
rect 10413 8381 10425 8384
rect 10459 8381 10471 8415
rect 10413 8375 10471 8381
rect 12529 8415 12587 8421
rect 12529 8381 12541 8415
rect 12575 8412 12587 8415
rect 12728 8412 12756 8440
rect 13096 8421 13124 8520
rect 21269 8517 21281 8551
rect 21315 8517 21327 8551
rect 21269 8511 21327 8517
rect 13630 8440 13636 8492
rect 13688 8480 13694 8492
rect 14090 8489 14096 8492
rect 14052 8483 14096 8489
rect 13688 8452 13952 8480
rect 13688 8440 13694 8452
rect 12805 8415 12863 8421
rect 12805 8412 12817 8415
rect 12575 8384 12609 8412
rect 12728 8384 12817 8412
rect 12575 8381 12587 8384
rect 12529 8375 12587 8381
rect 12805 8381 12817 8384
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 13081 8415 13139 8421
rect 13081 8381 13093 8415
rect 13127 8381 13139 8415
rect 13081 8375 13139 8381
rect 8128 8316 8892 8344
rect 9416 8344 9444 8372
rect 12161 8347 12219 8353
rect 9416 8316 9812 8344
rect 8864 8288 8892 8316
rect 2372 8248 3188 8276
rect 2372 8236 2378 8248
rect 3234 8236 3240 8288
rect 3292 8276 3298 8288
rect 3703 8279 3761 8285
rect 3703 8276 3715 8279
rect 3292 8248 3715 8276
rect 3292 8236 3298 8248
rect 3703 8245 3715 8248
rect 3749 8245 3761 8279
rect 3703 8239 3761 8245
rect 5810 8236 5816 8288
rect 5868 8276 5874 8288
rect 6178 8276 6184 8288
rect 5868 8248 6184 8276
rect 5868 8236 5874 8248
rect 6178 8236 6184 8248
rect 6236 8236 6242 8288
rect 7742 8236 7748 8288
rect 7800 8236 7806 8288
rect 8846 8236 8852 8288
rect 8904 8236 8910 8288
rect 9125 8279 9183 8285
rect 9125 8245 9137 8279
rect 9171 8276 9183 8279
rect 9398 8276 9404 8288
rect 9171 8248 9404 8276
rect 9171 8245 9183 8248
rect 9125 8239 9183 8245
rect 9398 8236 9404 8248
rect 9456 8236 9462 8288
rect 9784 8276 9812 8316
rect 12161 8313 12173 8347
rect 12207 8313 12219 8347
rect 12161 8307 12219 8313
rect 10143 8279 10201 8285
rect 10143 8276 10155 8279
rect 9784 8248 10155 8276
rect 10143 8245 10155 8248
rect 10189 8245 10201 8279
rect 10143 8239 10201 8245
rect 11974 8236 11980 8288
rect 12032 8276 12038 8288
rect 12176 8276 12204 8307
rect 12250 8304 12256 8356
rect 12308 8344 12314 8356
rect 12544 8344 12572 8375
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 13357 8415 13415 8421
rect 13357 8412 13369 8415
rect 13320 8384 13369 8412
rect 13320 8372 13326 8384
rect 13357 8381 13369 8384
rect 13403 8381 13415 8415
rect 13357 8375 13415 8381
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8412 13783 8415
rect 13814 8412 13820 8424
rect 13771 8384 13820 8412
rect 13771 8381 13783 8384
rect 13725 8375 13783 8381
rect 13740 8344 13768 8375
rect 13814 8372 13820 8384
rect 13872 8372 13878 8424
rect 13924 8412 13952 8452
rect 14052 8449 14064 8483
rect 14052 8443 14096 8449
rect 14090 8440 14096 8443
rect 14148 8440 14154 8492
rect 14182 8440 14188 8492
rect 14240 8440 14246 8492
rect 14461 8483 14519 8489
rect 14461 8449 14473 8483
rect 14507 8480 14519 8483
rect 14826 8480 14832 8492
rect 14507 8452 14832 8480
rect 14507 8449 14519 8452
rect 14461 8443 14519 8449
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 15841 8483 15899 8489
rect 15841 8449 15853 8483
rect 15887 8480 15899 8483
rect 16396 8483 16454 8489
rect 16396 8480 16408 8483
rect 15887 8452 16408 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 16396 8449 16408 8452
rect 16442 8449 16454 8483
rect 16396 8443 16454 8449
rect 18598 8440 18604 8492
rect 18656 8440 18662 8492
rect 19242 8480 19248 8492
rect 19174 8465 19248 8480
rect 13924 8384 15148 8412
rect 12308 8316 13768 8344
rect 15120 8344 15148 8384
rect 15194 8372 15200 8424
rect 15252 8412 15258 8424
rect 15933 8415 15991 8421
rect 15933 8412 15945 8415
rect 15252 8384 15945 8412
rect 15252 8372 15258 8384
rect 15933 8381 15945 8384
rect 15979 8381 15991 8415
rect 16669 8415 16727 8421
rect 16669 8412 16681 8415
rect 15933 8375 15991 8381
rect 16040 8384 16681 8412
rect 16040 8344 16068 8384
rect 16669 8381 16681 8384
rect 16715 8381 16727 8415
rect 16669 8375 16727 8381
rect 18325 8415 18383 8421
rect 18325 8381 18337 8415
rect 18371 8412 18383 8415
rect 18616 8412 18644 8440
rect 19174 8434 19201 8465
rect 19189 8431 19201 8434
rect 19235 8440 19248 8465
rect 19300 8440 19306 8492
rect 21284 8480 21312 8511
rect 22051 8483 22109 8489
rect 21284 8452 21680 8480
rect 19235 8431 19247 8440
rect 19189 8425 19247 8431
rect 18371 8384 18644 8412
rect 18693 8415 18751 8421
rect 18371 8381 18383 8384
rect 18325 8375 18383 8381
rect 18693 8381 18705 8415
rect 18739 8412 18751 8415
rect 18966 8412 18972 8424
rect 18739 8384 18972 8412
rect 18739 8381 18751 8384
rect 18693 8375 18751 8381
rect 18966 8372 18972 8384
rect 19024 8372 19030 8424
rect 19429 8415 19487 8421
rect 19429 8381 19441 8415
rect 19475 8412 19487 8415
rect 20806 8412 20812 8424
rect 19475 8384 20812 8412
rect 19475 8381 19487 8384
rect 19429 8375 19487 8381
rect 20806 8372 20812 8384
rect 20864 8372 20870 8424
rect 21450 8372 21456 8424
rect 21508 8372 21514 8424
rect 21545 8415 21603 8421
rect 21545 8381 21557 8415
rect 21591 8381 21603 8415
rect 21652 8412 21680 8452
rect 22051 8449 22063 8483
rect 22097 8480 22109 8483
rect 23400 8480 23428 8588
rect 25424 8560 25452 8588
rect 25866 8576 25872 8628
rect 25924 8576 25930 8628
rect 26053 8619 26111 8625
rect 26053 8585 26065 8619
rect 26099 8616 26111 8619
rect 26510 8616 26516 8628
rect 26099 8588 26516 8616
rect 26099 8585 26111 8588
rect 26053 8579 26111 8585
rect 26510 8576 26516 8588
rect 26568 8576 26574 8628
rect 27338 8616 27344 8628
rect 26718 8588 27344 8616
rect 23474 8508 23480 8560
rect 23532 8548 23538 8560
rect 23532 8520 23612 8548
rect 23532 8508 23538 8520
rect 22097 8452 23428 8480
rect 22097 8449 22109 8452
rect 22051 8443 22109 8449
rect 22281 8415 22339 8421
rect 22281 8412 22293 8415
rect 21652 8384 22293 8412
rect 21545 8375 21603 8381
rect 22281 8381 22293 8384
rect 22327 8381 22339 8415
rect 23584 8412 23612 8520
rect 25406 8508 25412 8560
rect 25464 8508 25470 8560
rect 26718 8548 26746 8588
rect 27338 8576 27344 8588
rect 27396 8576 27402 8628
rect 27430 8576 27436 8628
rect 27488 8616 27494 8628
rect 28537 8619 28595 8625
rect 28537 8616 28549 8619
rect 27488 8588 28549 8616
rect 27488 8576 27494 8588
rect 28537 8585 28549 8588
rect 28583 8585 28595 8619
rect 28537 8579 28595 8585
rect 26252 8520 26746 8548
rect 23661 8483 23719 8489
rect 23661 8449 23673 8483
rect 23707 8480 23719 8483
rect 24308 8483 24366 8489
rect 24308 8480 24320 8483
rect 23707 8452 24320 8480
rect 23707 8449 23719 8452
rect 23661 8443 23719 8449
rect 24308 8449 24320 8452
rect 24354 8449 24366 8483
rect 24308 8443 24366 8449
rect 24394 8440 24400 8492
rect 24452 8480 24458 8492
rect 24452 8452 25360 8480
rect 24452 8440 24458 8452
rect 25332 8424 25360 8452
rect 23842 8412 23848 8424
rect 23584 8384 23848 8412
rect 22281 8375 22339 8381
rect 15120 8316 16068 8344
rect 12308 8304 12314 8316
rect 18046 8304 18052 8356
rect 18104 8304 18110 8356
rect 20714 8304 20720 8356
rect 20772 8344 20778 8356
rect 21560 8344 21588 8375
rect 23842 8372 23848 8384
rect 23900 8372 23906 8424
rect 23934 8372 23940 8424
rect 23992 8412 23998 8424
rect 24581 8415 24639 8421
rect 24581 8412 24593 8415
rect 23992 8384 24593 8412
rect 23992 8372 23998 8384
rect 24581 8381 24593 8384
rect 24627 8381 24639 8415
rect 24581 8375 24639 8381
rect 25314 8372 25320 8424
rect 25372 8412 25378 8424
rect 26252 8421 26280 8520
rect 26602 8440 26608 8492
rect 26660 8480 26666 8492
rect 27062 8489 27068 8492
rect 27024 8483 27068 8489
rect 27024 8480 27036 8483
rect 26660 8452 27036 8480
rect 26660 8440 26666 8452
rect 27024 8449 27036 8452
rect 27024 8443 27068 8449
rect 27062 8440 27068 8443
rect 27120 8440 27126 8492
rect 27203 8483 27261 8489
rect 27203 8449 27215 8483
rect 27249 8480 27261 8483
rect 28258 8480 28264 8492
rect 27249 8452 28264 8480
rect 27249 8449 27261 8452
rect 27203 8443 27261 8449
rect 28258 8440 28264 8452
rect 28316 8440 28322 8492
rect 28718 8440 28724 8492
rect 28776 8440 28782 8492
rect 26237 8415 26295 8421
rect 26237 8412 26249 8415
rect 25372 8384 26249 8412
rect 25372 8372 25378 8384
rect 26237 8381 26249 8384
rect 26283 8381 26295 8415
rect 26237 8375 26295 8381
rect 26697 8415 26755 8421
rect 26697 8381 26709 8415
rect 26743 8412 26755 8415
rect 26786 8412 26792 8424
rect 26743 8384 26792 8412
rect 26743 8381 26755 8384
rect 26697 8375 26755 8381
rect 20772 8316 21588 8344
rect 20772 8304 20778 8316
rect 21468 8288 21496 8316
rect 23658 8304 23664 8356
rect 23716 8344 23722 8356
rect 23716 8316 23888 8344
rect 23716 8304 23722 8316
rect 12434 8276 12440 8288
rect 12032 8248 12440 8276
rect 12032 8236 12038 8248
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 12526 8236 12532 8288
rect 12584 8276 12590 8288
rect 12621 8279 12679 8285
rect 12621 8276 12633 8279
rect 12584 8248 12633 8276
rect 12584 8236 12590 8248
rect 12621 8245 12633 8248
rect 12667 8245 12679 8279
rect 12621 8239 12679 8245
rect 12710 8236 12716 8288
rect 12768 8276 12774 8288
rect 12897 8279 12955 8285
rect 12897 8276 12909 8279
rect 12768 8248 12909 8276
rect 12768 8236 12774 8248
rect 12897 8245 12909 8248
rect 12943 8245 12955 8279
rect 12897 8239 12955 8245
rect 13170 8236 13176 8288
rect 13228 8236 13234 8288
rect 16390 8236 16396 8288
rect 16448 8285 16454 8288
rect 16448 8239 16457 8285
rect 16448 8236 16454 8239
rect 18138 8236 18144 8288
rect 18196 8236 18202 8288
rect 18782 8236 18788 8288
rect 18840 8276 18846 8288
rect 19159 8279 19217 8285
rect 19159 8276 19171 8279
rect 18840 8248 19171 8276
rect 18840 8236 18846 8248
rect 19159 8245 19171 8248
rect 19205 8245 19217 8279
rect 19159 8239 19217 8245
rect 20990 8236 20996 8288
rect 21048 8276 21054 8288
rect 21085 8279 21143 8285
rect 21085 8276 21097 8279
rect 21048 8248 21097 8276
rect 21048 8236 21054 8248
rect 21085 8245 21097 8248
rect 21131 8245 21143 8279
rect 21085 8239 21143 8245
rect 21450 8236 21456 8288
rect 21508 8236 21514 8288
rect 21634 8236 21640 8288
rect 21692 8276 21698 8288
rect 22011 8279 22069 8285
rect 22011 8276 22023 8279
rect 21692 8248 22023 8276
rect 21692 8236 21698 8248
rect 22011 8245 22023 8248
rect 22057 8276 22069 8279
rect 23750 8276 23756 8288
rect 22057 8248 23756 8276
rect 22057 8245 22069 8248
rect 22011 8239 22069 8245
rect 23750 8236 23756 8248
rect 23808 8236 23814 8288
rect 23860 8276 23888 8316
rect 24302 8276 24308 8288
rect 24360 8285 24366 8288
rect 23860 8248 24308 8276
rect 24302 8236 24308 8248
rect 24360 8239 24369 8285
rect 26712 8276 26740 8375
rect 26786 8372 26792 8384
rect 26844 8372 26850 8424
rect 27433 8415 27491 8421
rect 27433 8381 27445 8415
rect 27479 8412 27491 8415
rect 28736 8412 28764 8440
rect 27479 8384 28764 8412
rect 27479 8381 27491 8384
rect 27433 8375 27491 8381
rect 29086 8372 29092 8424
rect 29144 8412 29150 8424
rect 29144 8384 29776 8412
rect 29144 8372 29150 8384
rect 29748 8356 29776 8384
rect 29546 8304 29552 8356
rect 29604 8344 29610 8356
rect 29641 8347 29699 8353
rect 29641 8344 29653 8347
rect 29604 8316 29653 8344
rect 29604 8304 29610 8316
rect 29641 8313 29653 8316
rect 29687 8313 29699 8347
rect 29641 8307 29699 8313
rect 29730 8304 29736 8356
rect 29788 8304 29794 8356
rect 27798 8276 27804 8288
rect 26712 8248 27804 8276
rect 24360 8236 24366 8239
rect 27798 8236 27804 8248
rect 27856 8236 27862 8288
rect 29178 8236 29184 8288
rect 29236 8236 29242 8288
rect 29917 8279 29975 8285
rect 29917 8245 29929 8279
rect 29963 8276 29975 8279
rect 30006 8276 30012 8288
rect 29963 8248 30012 8276
rect 29963 8245 29975 8248
rect 29917 8239 29975 8245
rect 30006 8236 30012 8248
rect 30064 8236 30070 8288
rect 552 8186 31072 8208
rect 552 8134 7988 8186
rect 8040 8134 8052 8186
rect 8104 8134 8116 8186
rect 8168 8134 8180 8186
rect 8232 8134 8244 8186
rect 8296 8134 15578 8186
rect 15630 8134 15642 8186
rect 15694 8134 15706 8186
rect 15758 8134 15770 8186
rect 15822 8134 15834 8186
rect 15886 8134 23168 8186
rect 23220 8134 23232 8186
rect 23284 8134 23296 8186
rect 23348 8134 23360 8186
rect 23412 8134 23424 8186
rect 23476 8134 30758 8186
rect 30810 8134 30822 8186
rect 30874 8134 30886 8186
rect 30938 8134 30950 8186
rect 31002 8134 31014 8186
rect 31066 8134 31072 8186
rect 552 8112 31072 8134
rect 845 8075 903 8081
rect 845 8041 857 8075
rect 891 8072 903 8075
rect 1670 8072 1676 8084
rect 891 8044 1676 8072
rect 891 8041 903 8044
rect 845 8035 903 8041
rect 1670 8032 1676 8044
rect 1728 8032 1734 8084
rect 10505 8075 10563 8081
rect 10505 8072 10517 8075
rect 2746 8044 10517 8072
rect 1026 7896 1032 7948
rect 1084 7896 1090 7948
rect 2746 7936 2774 8044
rect 10505 8041 10517 8044
rect 10551 8041 10563 8075
rect 10505 8035 10563 8041
rect 12075 8075 12133 8081
rect 12075 8041 12087 8075
rect 12121 8072 12133 8075
rect 12121 8044 13124 8072
rect 12121 8041 12133 8044
rect 12075 8035 12133 8041
rect 6454 7964 6460 8016
rect 6512 7964 6518 8016
rect 1872 7908 2774 7936
rect 1709 7889 1767 7895
rect 1709 7886 1721 7889
rect 1213 7871 1271 7877
rect 1213 7837 1225 7871
rect 1259 7837 1271 7871
rect 1213 7831 1271 7837
rect 1228 7744 1256 7831
rect 1394 7828 1400 7880
rect 1452 7868 1458 7880
rect 1540 7871 1598 7877
rect 1540 7868 1552 7871
rect 1452 7840 1552 7868
rect 1452 7828 1458 7840
rect 1540 7837 1552 7840
rect 1586 7837 1598 7871
rect 1688 7855 1721 7886
rect 1755 7868 1767 7889
rect 1872 7868 1900 7908
rect 3326 7896 3332 7948
rect 3384 7896 3390 7948
rect 3510 7896 3516 7948
rect 3568 7936 3574 7948
rect 5905 7939 5963 7945
rect 5905 7936 5917 7939
rect 3568 7908 5917 7936
rect 3568 7896 3574 7908
rect 5905 7905 5917 7908
rect 5951 7905 5963 7939
rect 6472 7936 6500 7964
rect 6784 7939 6842 7945
rect 6784 7936 6796 7939
rect 6472 7908 6796 7936
rect 5905 7899 5963 7905
rect 6784 7905 6796 7908
rect 6830 7905 6842 7939
rect 6784 7899 6842 7905
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 7156 7908 7205 7936
rect 7156 7896 7162 7908
rect 7193 7905 7205 7908
rect 7239 7905 7251 7939
rect 7193 7899 7251 7905
rect 7650 7896 7656 7948
rect 7708 7936 7714 7948
rect 8665 7939 8723 7945
rect 7708 7908 8432 7936
rect 7708 7896 7714 7908
rect 1755 7855 1900 7868
rect 1688 7840 1900 7855
rect 1540 7831 1598 7837
rect 1946 7828 1952 7880
rect 2004 7828 2010 7880
rect 3528 7800 3556 7896
rect 3694 7828 3700 7880
rect 3752 7868 3758 7880
rect 3840 7871 3898 7877
rect 3840 7868 3852 7871
rect 3752 7840 3852 7868
rect 3752 7828 3758 7840
rect 3840 7837 3852 7840
rect 3886 7837 3898 7871
rect 3840 7831 3898 7837
rect 4019 7871 4077 7877
rect 4019 7837 4031 7871
rect 4065 7868 4077 7871
rect 4154 7868 4160 7880
rect 4065 7840 4160 7868
rect 4065 7837 4077 7840
rect 4019 7831 4077 7837
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 5810 7868 5816 7880
rect 4295 7840 5816 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 5810 7828 5816 7840
rect 5868 7828 5874 7880
rect 6181 7871 6239 7877
rect 6181 7837 6193 7871
rect 6227 7868 6239 7871
rect 6362 7868 6368 7880
rect 6227 7840 6368 7868
rect 6227 7837 6239 7840
rect 6181 7831 6239 7837
rect 6362 7828 6368 7840
rect 6420 7868 6426 7880
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 6420 7840 6469 7868
rect 6420 7828 6426 7840
rect 6457 7837 6469 7840
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 6963 7871 7021 7877
rect 6963 7837 6975 7871
rect 7009 7868 7021 7871
rect 8202 7868 8208 7880
rect 7009 7840 8208 7868
rect 7009 7837 7021 7840
rect 6963 7831 7021 7837
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 2608 7772 3556 7800
rect 4908 7772 6040 7800
rect 1210 7692 1216 7744
rect 1268 7732 1274 7744
rect 2608 7732 2636 7772
rect 1268 7704 2636 7732
rect 1268 7692 1274 7704
rect 3326 7692 3332 7744
rect 3384 7732 3390 7744
rect 4062 7732 4068 7744
rect 3384 7704 4068 7732
rect 3384 7692 3390 7704
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 4154 7692 4160 7744
rect 4212 7732 4218 7744
rect 4908 7732 4936 7772
rect 4212 7704 4936 7732
rect 5537 7735 5595 7741
rect 4212 7692 4218 7704
rect 5537 7701 5549 7735
rect 5583 7732 5595 7735
rect 5902 7732 5908 7744
rect 5583 7704 5908 7732
rect 5583 7701 5595 7704
rect 5537 7695 5595 7701
rect 5902 7692 5908 7704
rect 5960 7692 5966 7744
rect 6012 7732 6040 7772
rect 6730 7732 6736 7744
rect 6012 7704 6736 7732
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 6914 7692 6920 7744
rect 6972 7732 6978 7744
rect 8297 7735 8355 7741
rect 8297 7732 8309 7735
rect 6972 7704 8309 7732
rect 6972 7692 6978 7704
rect 8297 7701 8309 7704
rect 8343 7701 8355 7735
rect 8404 7732 8432 7908
rect 8665 7905 8677 7939
rect 8711 7936 8723 7939
rect 8754 7936 8760 7948
rect 8711 7908 8760 7936
rect 8711 7905 8723 7908
rect 8665 7899 8723 7905
rect 8754 7896 8760 7908
rect 8812 7936 8818 7948
rect 9508 7936 9542 7940
rect 11057 7939 11115 7945
rect 11057 7936 11069 7939
rect 8812 7908 11069 7936
rect 8812 7896 8818 7908
rect 11057 7905 11069 7908
rect 11103 7905 11115 7939
rect 11057 7899 11115 7905
rect 11422 7896 11428 7948
rect 11480 7936 11486 7948
rect 11609 7939 11667 7945
rect 11609 7936 11621 7939
rect 11480 7908 11621 7936
rect 11480 7896 11486 7908
rect 11609 7905 11621 7908
rect 11655 7936 11667 7939
rect 11974 7936 11980 7948
rect 11655 7908 11980 7936
rect 11655 7905 11667 7908
rect 11609 7899 11667 7905
rect 11974 7896 11980 7908
rect 12032 7896 12038 7948
rect 12345 7939 12403 7945
rect 12345 7905 12357 7939
rect 12391 7936 12403 7939
rect 12710 7936 12716 7948
rect 12391 7908 12716 7936
rect 12391 7905 12403 7908
rect 12345 7899 12403 7905
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 13096 7880 13124 8044
rect 18782 8032 18788 8084
rect 18840 8081 18846 8084
rect 18840 8072 18849 8081
rect 18840 8044 20116 8072
rect 18840 8035 18849 8044
rect 18840 8032 18846 8035
rect 20088 8004 20116 8044
rect 20162 8032 20168 8084
rect 20220 8032 20226 8084
rect 20806 8032 20812 8084
rect 20864 8032 20870 8084
rect 21818 8032 21824 8084
rect 21876 8072 21882 8084
rect 23109 8075 23167 8081
rect 23109 8072 23121 8075
rect 21876 8044 23121 8072
rect 21876 8032 21882 8044
rect 23109 8041 23121 8044
rect 23155 8041 23167 8075
rect 23109 8035 23167 8041
rect 23750 8032 23756 8084
rect 23808 8072 23814 8084
rect 23943 8075 24001 8081
rect 23943 8072 23955 8075
rect 23808 8044 23955 8072
rect 23808 8032 23814 8044
rect 23943 8041 23955 8044
rect 23989 8041 24001 8075
rect 23943 8035 24001 8041
rect 27062 8032 27068 8084
rect 27120 8072 27126 8084
rect 27982 8072 27988 8084
rect 27120 8044 27988 8072
rect 27120 8032 27126 8044
rect 27982 8032 27988 8044
rect 28040 8072 28046 8084
rect 28083 8075 28141 8081
rect 28083 8072 28095 8075
rect 28040 8044 28095 8072
rect 28040 8032 28046 8044
rect 28083 8041 28095 8044
rect 28129 8041 28141 8075
rect 28083 8035 28141 8041
rect 28810 8032 28816 8084
rect 28868 8072 28874 8084
rect 29457 8075 29515 8081
rect 29457 8072 29469 8075
rect 28868 8044 29469 8072
rect 28868 8032 28874 8044
rect 29457 8041 29469 8044
rect 29503 8041 29515 8075
rect 29457 8035 29515 8041
rect 20088 7976 21128 8004
rect 13817 7939 13875 7945
rect 13817 7905 13829 7939
rect 13863 7936 13875 7939
rect 13906 7936 13912 7948
rect 13863 7908 13912 7936
rect 13863 7905 13875 7908
rect 13817 7899 13875 7905
rect 13906 7896 13912 7908
rect 13964 7896 13970 7948
rect 14144 7939 14202 7945
rect 14144 7936 14156 7939
rect 14016 7908 14156 7936
rect 8938 7828 8944 7880
rect 8996 7877 9002 7880
rect 8996 7871 9050 7877
rect 8996 7837 9004 7871
rect 9038 7837 9050 7871
rect 8996 7831 9050 7837
rect 8996 7828 9002 7831
rect 9122 7828 9128 7880
rect 9180 7877 9186 7880
rect 9180 7871 9229 7877
rect 9180 7837 9183 7871
rect 9217 7837 9229 7871
rect 9180 7831 9229 7837
rect 9180 7828 9186 7831
rect 9398 7828 9404 7880
rect 9456 7828 9462 7880
rect 9582 7828 9588 7880
rect 9640 7868 9646 7880
rect 12115 7871 12173 7877
rect 9640 7840 11284 7868
rect 9640 7828 9646 7840
rect 11146 7732 11152 7744
rect 8404 7704 11152 7732
rect 8297 7695 8355 7701
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 11256 7732 11284 7840
rect 12115 7837 12127 7871
rect 12161 7868 12173 7871
rect 12986 7868 12992 7880
rect 12161 7840 12992 7868
rect 12161 7837 12173 7840
rect 12115 7831 12173 7837
rect 12986 7828 12992 7840
rect 13044 7828 13050 7880
rect 13078 7828 13084 7880
rect 13136 7868 13142 7880
rect 14016 7868 14044 7908
rect 14144 7905 14156 7908
rect 14190 7936 14202 7939
rect 14458 7936 14464 7948
rect 14190 7908 14464 7936
rect 14190 7905 14202 7908
rect 14144 7899 14202 7905
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 14553 7939 14611 7945
rect 14553 7905 14565 7939
rect 14599 7936 14611 7939
rect 18138 7936 18144 7948
rect 14599 7908 18144 7936
rect 14599 7905 14611 7908
rect 14553 7899 14611 7905
rect 18138 7896 18144 7908
rect 18196 7896 18202 7948
rect 20622 7936 20628 7948
rect 18984 7908 20628 7936
rect 13136 7840 14044 7868
rect 14323 7871 14381 7877
rect 13136 7828 13142 7840
rect 14323 7837 14335 7871
rect 14369 7868 14381 7871
rect 15010 7868 15016 7880
rect 14369 7840 15016 7868
rect 14369 7837 14381 7840
rect 14323 7831 14381 7837
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 16117 7871 16175 7877
rect 16117 7868 16129 7871
rect 15252 7840 16129 7868
rect 15252 7828 15258 7840
rect 16117 7837 16129 7840
rect 16163 7837 16175 7871
rect 16117 7831 16175 7837
rect 16298 7828 16304 7880
rect 16356 7868 16362 7880
rect 16444 7871 16502 7877
rect 16444 7868 16456 7871
rect 16356 7840 16456 7868
rect 16356 7828 16362 7840
rect 16444 7837 16456 7840
rect 16490 7837 16502 7871
rect 16444 7831 16502 7837
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 16853 7871 16911 7877
rect 16632 7840 16677 7868
rect 16632 7828 16638 7840
rect 16853 7837 16865 7871
rect 16899 7868 16911 7871
rect 17494 7868 17500 7880
rect 16899 7840 17500 7868
rect 16899 7837 16911 7840
rect 16853 7831 16911 7837
rect 17494 7828 17500 7840
rect 17552 7828 17558 7880
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 18831 7871 18889 7877
rect 18831 7837 18843 7871
rect 18877 7868 18889 7871
rect 18984 7868 19012 7908
rect 20622 7896 20628 7908
rect 20680 7896 20686 7948
rect 20717 7939 20775 7945
rect 20717 7905 20729 7939
rect 20763 7905 20775 7939
rect 20993 7939 21051 7945
rect 20993 7936 21005 7939
rect 20717 7899 20775 7905
rect 20916 7908 21005 7936
rect 18877 7840 19012 7868
rect 18877 7837 18889 7840
rect 18831 7831 18889 7837
rect 13372 7772 13584 7800
rect 13372 7732 13400 7772
rect 11256 7704 13400 7732
rect 13446 7692 13452 7744
rect 13504 7692 13510 7744
rect 13556 7732 13584 7772
rect 15657 7735 15715 7741
rect 15657 7732 15669 7735
rect 13556 7704 15669 7732
rect 15657 7701 15669 7704
rect 15703 7701 15715 7735
rect 15657 7695 15715 7701
rect 17954 7692 17960 7744
rect 18012 7692 18018 7744
rect 18340 7732 18368 7831
rect 19058 7828 19064 7880
rect 19116 7828 19122 7880
rect 19150 7828 19156 7880
rect 19208 7868 19214 7880
rect 20732 7868 20760 7899
rect 20916 7880 20944 7908
rect 20993 7905 21005 7908
rect 21039 7905 21051 7939
rect 21100 7936 21128 7976
rect 22738 7964 22744 8016
rect 22796 8004 22802 8016
rect 22796 7976 23612 8004
rect 22796 7964 22802 7976
rect 23584 7948 23612 7976
rect 21634 7945 21640 7948
rect 21596 7939 21640 7945
rect 21596 7936 21608 7939
rect 21100 7908 21608 7936
rect 20993 7899 21051 7905
rect 21596 7905 21608 7908
rect 21596 7899 21640 7905
rect 21634 7896 21640 7899
rect 21692 7896 21698 7948
rect 23477 7939 23535 7945
rect 23477 7936 23489 7939
rect 21780 7908 22692 7936
rect 19208 7840 20760 7868
rect 19208 7828 19214 7840
rect 20732 7800 20760 7840
rect 20898 7828 20904 7880
rect 20956 7828 20962 7880
rect 21269 7871 21327 7877
rect 21269 7837 21281 7871
rect 21315 7868 21327 7871
rect 21450 7868 21456 7880
rect 21315 7840 21456 7868
rect 21315 7837 21327 7840
rect 21269 7831 21327 7837
rect 21450 7828 21456 7840
rect 21508 7828 21514 7880
rect 21780 7879 21808 7908
rect 21765 7873 21823 7879
rect 21765 7839 21777 7873
rect 21811 7839 21823 7873
rect 21765 7833 21823 7839
rect 21910 7828 21916 7880
rect 21968 7868 21974 7880
rect 22005 7871 22063 7877
rect 22005 7868 22017 7871
rect 21968 7840 22017 7868
rect 21968 7828 21974 7840
rect 22005 7837 22017 7840
rect 22051 7837 22063 7871
rect 22005 7831 22063 7837
rect 21174 7800 21180 7812
rect 20732 7772 21180 7800
rect 21174 7760 21180 7772
rect 21232 7760 21238 7812
rect 22664 7800 22692 7908
rect 23124 7908 23489 7936
rect 22738 7828 22744 7880
rect 22796 7868 22802 7880
rect 23124 7868 23152 7908
rect 23477 7905 23489 7908
rect 23523 7905 23535 7939
rect 23477 7899 23535 7905
rect 23566 7896 23572 7948
rect 23624 7936 23630 7948
rect 23624 7908 24348 7936
rect 23624 7896 23630 7908
rect 23750 7868 23756 7880
rect 22796 7840 23152 7868
rect 23492 7840 23756 7868
rect 22796 7828 22802 7840
rect 22830 7800 22836 7812
rect 22664 7772 22836 7800
rect 22830 7760 22836 7772
rect 22888 7760 22894 7812
rect 23492 7800 23520 7840
rect 23750 7828 23756 7840
rect 23808 7828 23814 7880
rect 23934 7828 23940 7880
rect 23992 7828 23998 7880
rect 24210 7828 24216 7880
rect 24268 7828 24274 7880
rect 24320 7868 24348 7908
rect 25682 7896 25688 7948
rect 25740 7896 25746 7948
rect 26605 7939 26663 7945
rect 26605 7936 26617 7939
rect 25792 7908 26617 7936
rect 25792 7868 25820 7908
rect 26605 7905 26617 7908
rect 26651 7905 26663 7939
rect 26605 7899 26663 7905
rect 26694 7896 26700 7948
rect 26752 7936 26758 7948
rect 27249 7939 27307 7945
rect 27249 7936 27261 7939
rect 26752 7908 27261 7936
rect 26752 7896 26758 7908
rect 27249 7905 27261 7908
rect 27295 7905 27307 7939
rect 27249 7899 27307 7905
rect 27525 7939 27583 7945
rect 27525 7905 27537 7939
rect 27571 7936 27583 7939
rect 28353 7939 28411 7945
rect 27571 7908 27936 7936
rect 27571 7905 27583 7908
rect 27525 7899 27583 7905
rect 27908 7880 27936 7908
rect 28353 7905 28365 7939
rect 28399 7936 28411 7939
rect 29270 7936 29276 7948
rect 28399 7908 29276 7936
rect 28399 7905 28411 7908
rect 28353 7899 28411 7905
rect 29270 7896 29276 7908
rect 29328 7896 29334 7948
rect 30006 7896 30012 7948
rect 30064 7896 30070 7948
rect 28113 7889 28171 7895
rect 28113 7886 28125 7889
rect 24320 7840 25820 7868
rect 25866 7828 25872 7880
rect 25924 7828 25930 7880
rect 25958 7828 25964 7880
rect 26016 7868 26022 7880
rect 27617 7871 27675 7877
rect 26016 7840 27568 7868
rect 26016 7828 26022 7840
rect 27065 7803 27123 7809
rect 23308 7772 23520 7800
rect 24872 7772 25544 7800
rect 18966 7732 18972 7744
rect 18340 7704 18972 7732
rect 18966 7692 18972 7704
rect 19024 7692 19030 7744
rect 20530 7692 20536 7744
rect 20588 7692 20594 7744
rect 20622 7692 20628 7744
rect 20680 7732 20686 7744
rect 23308 7732 23336 7772
rect 20680 7704 23336 7732
rect 20680 7692 20686 7704
rect 23382 7692 23388 7744
rect 23440 7732 23446 7744
rect 24872 7732 24900 7772
rect 25516 7744 25544 7772
rect 27065 7769 27077 7803
rect 27111 7800 27123 7803
rect 27430 7800 27436 7812
rect 27111 7772 27436 7800
rect 27111 7769 27123 7772
rect 27065 7763 27123 7769
rect 27430 7760 27436 7772
rect 27488 7760 27494 7812
rect 23440 7704 24900 7732
rect 23440 7692 23446 7704
rect 25314 7692 25320 7744
rect 25372 7692 25378 7744
rect 25498 7692 25504 7744
rect 25556 7692 25562 7744
rect 25590 7692 25596 7744
rect 25648 7732 25654 7744
rect 26421 7735 26479 7741
rect 26421 7732 26433 7735
rect 25648 7704 26433 7732
rect 25648 7692 25654 7704
rect 26421 7701 26433 7704
rect 26467 7701 26479 7735
rect 26421 7695 26479 7701
rect 27338 7692 27344 7744
rect 27396 7692 27402 7744
rect 27540 7732 27568 7840
rect 27617 7837 27629 7871
rect 27663 7868 27675 7871
rect 27798 7868 27804 7880
rect 27663 7840 27804 7868
rect 27663 7837 27675 7840
rect 27617 7831 27675 7837
rect 27798 7828 27804 7840
rect 27856 7828 27862 7880
rect 27890 7828 27896 7880
rect 27948 7828 27954 7880
rect 28098 7855 28125 7886
rect 28159 7880 28171 7889
rect 28159 7855 28172 7880
rect 28098 7840 28172 7855
rect 28166 7828 28172 7840
rect 28224 7828 28230 7880
rect 29362 7732 29368 7744
rect 27540 7704 29368 7732
rect 29362 7692 29368 7704
rect 29420 7692 29426 7744
rect 29822 7692 29828 7744
rect 29880 7692 29886 7744
rect 552 7642 30912 7664
rect 552 7590 4193 7642
rect 4245 7590 4257 7642
rect 4309 7590 4321 7642
rect 4373 7590 4385 7642
rect 4437 7590 4449 7642
rect 4501 7590 11783 7642
rect 11835 7590 11847 7642
rect 11899 7590 11911 7642
rect 11963 7590 11975 7642
rect 12027 7590 12039 7642
rect 12091 7590 19373 7642
rect 19425 7590 19437 7642
rect 19489 7590 19501 7642
rect 19553 7590 19565 7642
rect 19617 7590 19629 7642
rect 19681 7590 26963 7642
rect 27015 7590 27027 7642
rect 27079 7590 27091 7642
rect 27143 7590 27155 7642
rect 27207 7590 27219 7642
rect 27271 7590 30912 7642
rect 552 7568 30912 7590
rect 5353 7531 5411 7537
rect 5353 7528 5365 7531
rect 3068 7500 5365 7528
rect 2406 7420 2412 7472
rect 2464 7460 2470 7472
rect 3068 7460 3096 7500
rect 5353 7497 5365 7500
rect 5399 7497 5411 7531
rect 5353 7491 5411 7497
rect 5718 7488 5724 7540
rect 5776 7488 5782 7540
rect 13446 7528 13452 7540
rect 6104 7500 10548 7528
rect 2464 7432 3096 7460
rect 3237 7463 3295 7469
rect 2464 7420 2470 7432
rect 3237 7429 3249 7463
rect 3283 7429 3295 7463
rect 3237 7423 3295 7429
rect 1443 7395 1501 7401
rect 1443 7361 1455 7395
rect 1489 7392 1501 7395
rect 2958 7392 2964 7404
rect 1489 7364 2964 7392
rect 1489 7361 1501 7364
rect 1443 7355 1501 7361
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 3252 7392 3280 7423
rect 4019 7395 4077 7401
rect 3252 7374 3746 7392
rect 3252 7364 3914 7374
rect 3718 7346 3914 7364
rect 4019 7361 4031 7395
rect 4065 7392 4077 7395
rect 6104 7392 6132 7500
rect 10520 7472 10548 7500
rect 10980 7500 13452 7528
rect 10502 7420 10508 7472
rect 10560 7420 10566 7472
rect 4065 7364 6132 7392
rect 4065 7361 4077 7364
rect 4019 7355 4077 7361
rect 6546 7352 6552 7404
rect 6604 7401 6610 7404
rect 6604 7395 6653 7401
rect 6604 7361 6607 7395
rect 6641 7361 6653 7395
rect 6604 7355 6653 7361
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 7742 7392 7748 7404
rect 6871 7364 7748 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 6604 7352 6610 7355
rect 7742 7352 7748 7364
rect 7800 7352 7806 7404
rect 8662 7392 8668 7404
rect 8404 7364 8668 7392
rect 937 7327 995 7333
rect 937 7293 949 7327
rect 983 7324 995 7327
rect 1210 7324 1216 7336
rect 983 7296 1216 7324
rect 983 7293 995 7296
rect 937 7287 995 7293
rect 1210 7284 1216 7296
rect 1268 7284 1274 7336
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 2682 7324 2688 7336
rect 1719 7296 2688 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 2682 7284 2688 7296
rect 2740 7284 2746 7336
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 3344 7296 3433 7324
rect 3344 7200 3372 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 3510 7284 3516 7336
rect 3568 7284 3574 7336
rect 3886 7324 3914 7346
rect 4249 7327 4307 7333
rect 4249 7324 4261 7327
rect 3886 7296 4261 7324
rect 4249 7293 4261 7296
rect 4295 7293 4307 7327
rect 4249 7287 4307 7293
rect 5258 7284 5264 7336
rect 5316 7324 5322 7336
rect 5905 7327 5963 7333
rect 5905 7324 5917 7327
rect 5316 7296 5917 7324
rect 5316 7284 5322 7296
rect 5736 7268 5764 7296
rect 5905 7293 5917 7296
rect 5951 7293 5963 7327
rect 5905 7287 5963 7293
rect 6089 7327 6147 7333
rect 6089 7293 6101 7327
rect 6135 7293 6147 7327
rect 6089 7287 6147 7293
rect 5718 7216 5724 7268
rect 5776 7216 5782 7268
rect 1394 7148 1400 7200
rect 1452 7197 1458 7200
rect 1452 7188 1461 7197
rect 1452 7160 1497 7188
rect 1452 7151 1461 7160
rect 1452 7148 1458 7151
rect 2774 7148 2780 7200
rect 2832 7148 2838 7200
rect 3326 7148 3332 7200
rect 3384 7148 3390 7200
rect 3970 7148 3976 7200
rect 4028 7197 4034 7200
rect 4028 7188 4037 7197
rect 6104 7188 6132 7287
rect 6178 7284 6184 7336
rect 6236 7324 6242 7336
rect 8404 7333 8432 7364
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 8754 7352 8760 7404
rect 8812 7392 8818 7404
rect 9033 7395 9091 7401
rect 9033 7392 9045 7395
rect 8812 7364 9045 7392
rect 8812 7352 8818 7364
rect 9033 7361 9045 7364
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 9539 7395 9597 7401
rect 9539 7361 9551 7395
rect 9585 7392 9597 7395
rect 10980 7392 11008 7500
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 13722 7488 13728 7540
rect 13780 7528 13786 7540
rect 18325 7531 18383 7537
rect 13780 7500 15424 7528
rect 13780 7488 13786 7500
rect 9585 7364 11008 7392
rect 11241 7395 11299 7401
rect 9585 7361 9597 7364
rect 9539 7355 9597 7361
rect 11241 7361 11253 7395
rect 11287 7392 11299 7395
rect 11422 7392 11428 7404
rect 11287 7364 11428 7392
rect 11287 7361 11299 7364
rect 11241 7355 11299 7361
rect 11422 7352 11428 7364
rect 11480 7352 11486 7404
rect 11747 7395 11805 7401
rect 11747 7361 11759 7395
rect 11793 7392 11805 7395
rect 12342 7392 12348 7404
rect 11793 7364 12348 7392
rect 11793 7361 11805 7364
rect 11747 7355 11805 7361
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 12492 7364 13952 7392
rect 12492 7352 12498 7364
rect 13924 7336 13952 7364
rect 14366 7352 14372 7404
rect 14424 7392 14430 7404
rect 14424 7364 14469 7392
rect 14424 7352 14430 7364
rect 14642 7352 14648 7404
rect 14700 7352 14706 7404
rect 15396 7392 15424 7500
rect 18325 7497 18337 7531
rect 18371 7528 18383 7531
rect 19794 7528 19800 7540
rect 18371 7500 19800 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 20530 7488 20536 7540
rect 20588 7488 20594 7540
rect 23382 7528 23388 7540
rect 21100 7500 23388 7528
rect 17954 7420 17960 7472
rect 18012 7420 18018 7472
rect 16580 7393 16638 7399
rect 15396 7364 16252 7392
rect 9398 7333 9404 7336
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 6236 7296 8217 7324
rect 6236 7284 6242 7296
rect 8205 7293 8217 7296
rect 8251 7293 8263 7327
rect 8205 7287 8263 7293
rect 8389 7327 8447 7333
rect 8389 7293 8401 7327
rect 8435 7293 8447 7327
rect 9360 7327 9404 7333
rect 9360 7324 9372 7327
rect 8389 7287 8447 7293
rect 9140 7296 9372 7324
rect 7558 7216 7564 7268
rect 7616 7256 7622 7268
rect 8404 7256 8432 7287
rect 7616 7228 8432 7256
rect 8665 7259 8723 7265
rect 7616 7216 7622 7228
rect 8665 7225 8677 7259
rect 8711 7256 8723 7259
rect 8938 7256 8944 7268
rect 8711 7228 8944 7256
rect 8711 7225 8723 7228
rect 8665 7219 8723 7225
rect 8938 7216 8944 7228
rect 8996 7256 9002 7268
rect 9140 7256 9168 7296
rect 9360 7293 9372 7296
rect 9360 7287 9404 7293
rect 9398 7284 9404 7287
rect 9456 7284 9462 7336
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7324 9827 7327
rect 10594 7324 10600 7336
rect 9815 7296 10600 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 10594 7284 10600 7296
rect 10652 7284 10658 7336
rect 11977 7327 12035 7333
rect 11977 7293 11989 7327
rect 12023 7324 12035 7327
rect 12710 7324 12716 7336
rect 12023 7296 12716 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 13078 7284 13084 7336
rect 13136 7284 13142 7336
rect 13817 7327 13875 7333
rect 13817 7293 13829 7327
rect 13863 7293 13875 7327
rect 13817 7287 13875 7293
rect 13096 7256 13124 7284
rect 8996 7228 9168 7256
rect 13004 7228 13124 7256
rect 13832 7256 13860 7287
rect 13906 7284 13912 7336
rect 13964 7284 13970 7336
rect 14734 7284 14740 7336
rect 14792 7324 14798 7336
rect 15102 7324 15108 7336
rect 14792 7296 15108 7324
rect 14792 7284 14798 7296
rect 15102 7284 15108 7296
rect 15160 7324 15166 7336
rect 16117 7327 16175 7333
rect 16117 7324 16129 7327
rect 15160 7296 16129 7324
rect 15160 7284 15166 7296
rect 16117 7293 16129 7296
rect 16163 7293 16175 7327
rect 16224 7324 16252 7364
rect 16580 7359 16592 7393
rect 16626 7392 16638 7393
rect 16666 7392 16672 7404
rect 16626 7364 16672 7392
rect 16626 7359 16638 7364
rect 16580 7353 16638 7359
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 17034 7352 17040 7404
rect 17092 7392 17098 7404
rect 18693 7395 18751 7401
rect 17092 7364 18552 7392
rect 17092 7352 17098 7364
rect 18524 7333 18552 7364
rect 18693 7361 18705 7395
rect 18739 7392 18751 7395
rect 18966 7392 18972 7404
rect 18739 7364 18972 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 18966 7352 18972 7364
rect 19024 7352 19030 7404
rect 19199 7395 19257 7401
rect 19199 7361 19211 7395
rect 19245 7392 19257 7395
rect 19429 7395 19487 7401
rect 19245 7364 19380 7392
rect 19245 7361 19257 7364
rect 19199 7355 19257 7361
rect 16853 7327 16911 7333
rect 16853 7324 16865 7327
rect 16224 7296 16865 7324
rect 16117 7287 16175 7293
rect 16853 7293 16865 7296
rect 16899 7293 16911 7327
rect 16853 7287 16911 7293
rect 18509 7327 18567 7333
rect 18509 7293 18521 7327
rect 18555 7324 18567 7327
rect 18598 7324 18604 7336
rect 18555 7296 18604 7324
rect 18555 7293 18567 7296
rect 18509 7287 18567 7293
rect 18598 7284 18604 7296
rect 18656 7284 18662 7336
rect 19352 7324 19380 7364
rect 19429 7361 19441 7395
rect 19475 7392 19487 7395
rect 20548 7392 20576 7488
rect 19475 7364 20576 7392
rect 19475 7361 19487 7364
rect 19429 7355 19487 7361
rect 20990 7324 20996 7336
rect 19352 7296 20996 7324
rect 20990 7284 20996 7296
rect 21048 7324 21054 7336
rect 21100 7333 21128 7500
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 23477 7531 23535 7537
rect 23477 7497 23489 7531
rect 23523 7528 23535 7531
rect 24026 7528 24032 7540
rect 23523 7500 24032 7528
rect 23523 7497 23535 7500
rect 23477 7491 23535 7497
rect 24026 7488 24032 7500
rect 24084 7488 24090 7540
rect 25314 7488 25320 7540
rect 25372 7488 25378 7540
rect 25869 7531 25927 7537
rect 25869 7497 25881 7531
rect 25915 7528 25927 7531
rect 26878 7528 26884 7540
rect 25915 7500 26884 7528
rect 25915 7497 25927 7500
rect 25869 7491 25927 7497
rect 26878 7488 26884 7500
rect 26936 7488 26942 7540
rect 27890 7488 27896 7540
rect 27948 7528 27954 7540
rect 28258 7528 28264 7540
rect 27948 7500 28264 7528
rect 27948 7488 27954 7500
rect 28258 7488 28264 7500
rect 28316 7488 28322 7540
rect 21634 7352 21640 7404
rect 21692 7392 21698 7404
rect 21780 7395 21838 7401
rect 21780 7392 21792 7395
rect 21692 7364 21792 7392
rect 21692 7352 21698 7364
rect 21780 7361 21792 7364
rect 21826 7361 21838 7395
rect 21780 7355 21838 7361
rect 21959 7395 22017 7401
rect 21959 7361 21971 7395
rect 22005 7392 22017 7395
rect 22005 7364 23796 7392
rect 22005 7361 22017 7364
rect 21959 7355 22017 7361
rect 21085 7327 21143 7333
rect 21085 7324 21097 7327
rect 21048 7296 21097 7324
rect 21048 7284 21054 7296
rect 21085 7293 21097 7296
rect 21131 7293 21143 7327
rect 21085 7287 21143 7293
rect 21450 7284 21456 7336
rect 21508 7284 21514 7336
rect 22186 7284 22192 7336
rect 22244 7284 22250 7336
rect 13998 7256 14004 7268
rect 13832 7228 14004 7256
rect 8996 7216 9002 7228
rect 6362 7188 6368 7200
rect 4028 7160 4073 7188
rect 6104 7160 6368 7188
rect 4028 7151 4037 7160
rect 4028 7148 4034 7151
rect 6362 7148 6368 7160
rect 6420 7148 6426 7200
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 6555 7191 6613 7197
rect 6555 7188 6567 7191
rect 6512 7160 6567 7188
rect 6512 7148 6518 7160
rect 6555 7157 6567 7160
rect 6601 7157 6613 7191
rect 6555 7151 6613 7157
rect 6730 7148 6736 7200
rect 6788 7188 6794 7200
rect 9858 7188 9864 7200
rect 6788 7160 9864 7188
rect 6788 7148 6794 7160
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 10870 7148 10876 7200
rect 10928 7148 10934 7200
rect 11707 7191 11765 7197
rect 11707 7157 11719 7191
rect 11753 7188 11765 7191
rect 12434 7188 12440 7200
rect 11753 7160 12440 7188
rect 11753 7157 11765 7160
rect 11707 7151 11765 7157
rect 12434 7148 12440 7160
rect 12492 7188 12498 7200
rect 13004 7188 13032 7228
rect 13998 7216 14004 7228
rect 14056 7216 14062 7268
rect 12492 7160 13032 7188
rect 12492 7148 12498 7160
rect 13078 7148 13084 7200
rect 13136 7148 13142 7200
rect 13633 7191 13691 7197
rect 13633 7157 13645 7191
rect 13679 7188 13691 7191
rect 14274 7188 14280 7200
rect 13679 7160 14280 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 14375 7191 14433 7197
rect 14375 7157 14387 7191
rect 14421 7188 14433 7191
rect 14550 7188 14556 7200
rect 14421 7160 14556 7188
rect 14421 7157 14433 7160
rect 14375 7151 14433 7157
rect 14550 7148 14556 7160
rect 14608 7148 14614 7200
rect 15286 7148 15292 7200
rect 15344 7188 15350 7200
rect 15749 7191 15807 7197
rect 15749 7188 15761 7191
rect 15344 7160 15761 7188
rect 15344 7148 15350 7160
rect 15749 7157 15761 7160
rect 15795 7157 15807 7191
rect 15749 7151 15807 7157
rect 16390 7148 16396 7200
rect 16448 7188 16454 7200
rect 16583 7191 16641 7197
rect 16583 7188 16595 7191
rect 16448 7160 16595 7188
rect 16448 7148 16454 7160
rect 16583 7157 16595 7160
rect 16629 7157 16641 7191
rect 16583 7151 16641 7157
rect 18782 7148 18788 7200
rect 18840 7188 18846 7200
rect 19159 7191 19217 7197
rect 19159 7188 19171 7191
rect 18840 7160 19171 7188
rect 18840 7148 18846 7160
rect 19159 7157 19171 7160
rect 19205 7157 19217 7191
rect 19159 7151 19217 7157
rect 19886 7148 19892 7200
rect 19944 7188 19950 7200
rect 20533 7191 20591 7197
rect 20533 7188 20545 7191
rect 19944 7160 20545 7188
rect 19944 7148 19950 7160
rect 20533 7157 20545 7160
rect 20579 7157 20591 7191
rect 21468 7188 21496 7284
rect 22646 7188 22652 7200
rect 21468 7160 22652 7188
rect 20533 7151 20591 7157
rect 22646 7148 22652 7160
rect 22704 7148 22710 7200
rect 23768 7188 23796 7364
rect 23842 7352 23848 7404
rect 23900 7352 23906 7404
rect 24118 7352 24124 7404
rect 24176 7352 24182 7404
rect 24351 7395 24409 7401
rect 24351 7361 24363 7395
rect 24397 7392 24409 7395
rect 25332 7392 25360 7488
rect 28902 7420 28908 7472
rect 28960 7460 28966 7472
rect 29273 7463 29331 7469
rect 29273 7460 29285 7463
rect 28960 7432 29285 7460
rect 28960 7420 28966 7432
rect 29273 7429 29285 7432
rect 29319 7429 29331 7463
rect 29273 7423 29331 7429
rect 29454 7420 29460 7472
rect 29512 7460 29518 7472
rect 29512 7432 29776 7460
rect 29512 7420 29518 7432
rect 28350 7392 28356 7404
rect 24397 7364 25360 7392
rect 26528 7377 28356 7392
rect 24397 7361 24409 7364
rect 24351 7355 24409 7361
rect 24136 7324 24164 7352
rect 26528 7346 26561 7377
rect 26549 7343 26561 7346
rect 26595 7364 28356 7377
rect 26595 7343 26607 7364
rect 28350 7352 28356 7364
rect 28408 7352 28414 7404
rect 28994 7352 29000 7404
rect 29052 7352 29058 7404
rect 26549 7337 26607 7343
rect 24581 7327 24639 7333
rect 24581 7324 24593 7327
rect 24136 7296 24593 7324
rect 24581 7293 24593 7296
rect 24627 7293 24639 7327
rect 24581 7287 24639 7293
rect 25314 7284 25320 7336
rect 25372 7324 25378 7336
rect 26050 7324 26056 7336
rect 25372 7296 26056 7324
rect 25372 7284 25378 7296
rect 26050 7284 26056 7296
rect 26108 7284 26114 7336
rect 26786 7284 26792 7336
rect 26844 7284 26850 7336
rect 29012 7324 29040 7352
rect 29748 7333 29776 7432
rect 29181 7327 29239 7333
rect 29181 7324 29193 7327
rect 29012 7296 29193 7324
rect 29181 7293 29193 7296
rect 29227 7293 29239 7327
rect 29181 7287 29239 7293
rect 29457 7327 29515 7333
rect 29457 7293 29469 7327
rect 29503 7293 29515 7327
rect 29457 7287 29515 7293
rect 29733 7327 29791 7333
rect 29733 7293 29745 7327
rect 29779 7293 29791 7327
rect 29733 7287 29791 7293
rect 28353 7259 28411 7265
rect 28353 7256 28365 7259
rect 27448 7228 28365 7256
rect 24118 7188 24124 7200
rect 23768 7160 24124 7188
rect 24118 7148 24124 7160
rect 24176 7148 24182 7200
rect 24302 7148 24308 7200
rect 24360 7197 24366 7200
rect 24360 7188 24369 7197
rect 24360 7160 24405 7188
rect 24360 7151 24369 7160
rect 24360 7148 24366 7151
rect 24486 7148 24492 7200
rect 24544 7188 24550 7200
rect 25866 7188 25872 7200
rect 24544 7160 25872 7188
rect 24544 7148 24550 7160
rect 25866 7148 25872 7160
rect 25924 7188 25930 7200
rect 26519 7191 26577 7197
rect 26519 7188 26531 7191
rect 25924 7160 26531 7188
rect 25924 7148 25930 7160
rect 26519 7157 26531 7160
rect 26565 7188 26577 7191
rect 26878 7188 26884 7200
rect 26565 7160 26884 7188
rect 26565 7157 26577 7160
rect 26519 7151 26577 7157
rect 26878 7148 26884 7160
rect 26936 7148 26942 7200
rect 27246 7148 27252 7200
rect 27304 7188 27310 7200
rect 27448 7188 27476 7228
rect 28353 7225 28365 7228
rect 28399 7225 28411 7259
rect 29472 7256 29500 7287
rect 28353 7219 28411 7225
rect 29196 7228 29500 7256
rect 29196 7200 29224 7228
rect 27304 7160 27476 7188
rect 27304 7148 27310 7160
rect 27890 7148 27896 7200
rect 27948 7148 27954 7200
rect 28258 7148 28264 7200
rect 28316 7188 28322 7200
rect 28445 7191 28503 7197
rect 28445 7188 28457 7191
rect 28316 7160 28457 7188
rect 28316 7148 28322 7160
rect 28445 7157 28457 7160
rect 28491 7157 28503 7191
rect 28445 7151 28503 7157
rect 28534 7148 28540 7200
rect 28592 7188 28598 7200
rect 28997 7191 29055 7197
rect 28997 7188 29009 7191
rect 28592 7160 29009 7188
rect 28592 7148 28598 7160
rect 28997 7157 29009 7160
rect 29043 7157 29055 7191
rect 28997 7151 29055 7157
rect 29178 7148 29184 7200
rect 29236 7148 29242 7200
rect 29270 7148 29276 7200
rect 29328 7188 29334 7200
rect 29549 7191 29607 7197
rect 29549 7188 29561 7191
rect 29328 7160 29561 7188
rect 29328 7148 29334 7160
rect 29549 7157 29561 7160
rect 29595 7157 29607 7191
rect 29549 7151 29607 7157
rect 552 7098 31072 7120
rect 552 7046 7988 7098
rect 8040 7046 8052 7098
rect 8104 7046 8116 7098
rect 8168 7046 8180 7098
rect 8232 7046 8244 7098
rect 8296 7046 15578 7098
rect 15630 7046 15642 7098
rect 15694 7046 15706 7098
rect 15758 7046 15770 7098
rect 15822 7046 15834 7098
rect 15886 7046 23168 7098
rect 23220 7046 23232 7098
rect 23284 7046 23296 7098
rect 23348 7046 23360 7098
rect 23412 7046 23424 7098
rect 23476 7046 30758 7098
rect 30810 7046 30822 7098
rect 30874 7046 30886 7098
rect 30938 7046 30950 7098
rect 31002 7046 31014 7098
rect 31066 7046 31072 7098
rect 552 7024 31072 7046
rect 1394 6944 1400 6996
rect 1452 6984 1458 6996
rect 1587 6987 1645 6993
rect 1587 6984 1599 6987
rect 1452 6956 1599 6984
rect 1452 6944 1458 6956
rect 1587 6953 1599 6956
rect 1633 6984 1645 6987
rect 1633 6956 2544 6984
rect 1633 6953 1645 6956
rect 1587 6947 1645 6953
rect 2516 6916 2544 6956
rect 2682 6944 2688 6996
rect 2740 6984 2746 6996
rect 2740 6956 4752 6984
rect 2740 6944 2746 6956
rect 3237 6919 3295 6925
rect 2516 6888 3188 6916
rect 1029 6851 1087 6857
rect 1029 6817 1041 6851
rect 1075 6817 1087 6851
rect 1029 6811 1087 6817
rect 1121 6851 1179 6857
rect 1121 6817 1133 6851
rect 1167 6848 1179 6851
rect 1210 6848 1216 6860
rect 1167 6820 1216 6848
rect 1167 6817 1179 6820
rect 1121 6811 1179 6817
rect 1044 6712 1072 6811
rect 1210 6808 1216 6820
rect 1268 6808 1274 6860
rect 3160 6848 3188 6888
rect 3237 6885 3249 6919
rect 3283 6916 3295 6919
rect 3418 6916 3424 6928
rect 3283 6888 3424 6916
rect 3283 6885 3295 6888
rect 3237 6879 3295 6885
rect 3418 6876 3424 6888
rect 3476 6876 3482 6928
rect 4724 6916 4752 6956
rect 5810 6944 5816 6996
rect 5868 6944 5874 6996
rect 6089 6987 6147 6993
rect 6089 6953 6101 6987
rect 6135 6953 6147 6987
rect 6089 6947 6147 6953
rect 6104 6916 6132 6947
rect 6454 6944 6460 6996
rect 6512 6984 6518 6996
rect 6923 6987 6981 6993
rect 6923 6984 6935 6987
rect 6512 6956 6935 6984
rect 6512 6944 6518 6956
rect 6923 6953 6935 6956
rect 6969 6984 6981 6987
rect 9131 6987 9189 6993
rect 9131 6984 9143 6987
rect 6969 6956 9143 6984
rect 6969 6953 6981 6956
rect 6923 6947 6981 6953
rect 9131 6953 9143 6956
rect 9177 6984 9189 6987
rect 9398 6984 9404 6996
rect 9177 6956 9404 6984
rect 9177 6953 9189 6956
rect 9131 6947 9189 6953
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 10502 6944 10508 6996
rect 10560 6944 10566 6996
rect 11241 6987 11299 6993
rect 11241 6984 11253 6987
rect 10980 6956 11253 6984
rect 4724 6888 6132 6916
rect 10778 6876 10784 6928
rect 10836 6916 10842 6928
rect 10980 6916 11008 6956
rect 11241 6953 11253 6956
rect 11287 6953 11299 6987
rect 11241 6947 11299 6953
rect 11974 6944 11980 6996
rect 12032 6944 12038 6996
rect 12894 6984 12900 6996
rect 12176 6956 12900 6984
rect 11992 6916 12020 6944
rect 10836 6888 11008 6916
rect 11440 6888 12020 6916
rect 10836 6876 10842 6888
rect 3694 6857 3700 6860
rect 3656 6851 3700 6857
rect 3656 6848 3668 6851
rect 3160 6820 3668 6848
rect 3656 6817 3668 6820
rect 3656 6811 3700 6817
rect 3694 6808 3700 6811
rect 3752 6808 3758 6860
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6848 4123 6851
rect 5166 6848 5172 6860
rect 4111 6820 5172 6848
rect 4111 6817 4123 6820
rect 4065 6811 4123 6817
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 5442 6808 5448 6860
rect 5500 6808 5506 6860
rect 5718 6808 5724 6860
rect 5776 6848 5782 6860
rect 5997 6851 6055 6857
rect 5997 6848 6009 6851
rect 5776 6820 6009 6848
rect 5776 6808 5782 6820
rect 5997 6817 6009 6820
rect 6043 6848 6055 6851
rect 6178 6848 6184 6860
rect 6043 6820 6184 6848
rect 6043 6817 6055 6820
rect 5997 6811 6055 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6817 6331 6851
rect 6273 6811 6331 6817
rect 1627 6783 1685 6789
rect 1627 6749 1639 6783
rect 1673 6780 1685 6783
rect 1762 6780 1768 6792
rect 1673 6752 1768 6780
rect 1673 6749 1685 6752
rect 1627 6743 1685 6749
rect 1762 6740 1768 6752
rect 1820 6740 1826 6792
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6780 1915 6783
rect 3329 6783 3387 6789
rect 1903 6752 2774 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 1118 6712 1124 6724
rect 1044 6684 1124 6712
rect 1118 6672 1124 6684
rect 1176 6672 1182 6724
rect 845 6647 903 6653
rect 845 6613 857 6647
rect 891 6644 903 6647
rect 1486 6644 1492 6656
rect 891 6616 1492 6644
rect 891 6613 903 6616
rect 845 6607 903 6613
rect 1486 6604 1492 6616
rect 1544 6604 1550 6656
rect 2746 6644 2774 6752
rect 3329 6749 3341 6783
rect 3375 6780 3387 6783
rect 3510 6780 3516 6792
rect 3375 6752 3516 6780
rect 3375 6749 3387 6752
rect 3329 6743 3387 6749
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 3835 6783 3893 6789
rect 3835 6749 3847 6783
rect 3881 6780 3893 6783
rect 6288 6780 6316 6811
rect 6362 6808 6368 6860
rect 6420 6848 6426 6860
rect 6457 6851 6515 6857
rect 6457 6848 6469 6851
rect 6420 6820 6469 6848
rect 6420 6808 6426 6820
rect 6457 6817 6469 6820
rect 6503 6848 6515 6851
rect 6503 6820 7144 6848
rect 6503 6817 6515 6820
rect 6457 6811 6515 6817
rect 6730 6780 6736 6792
rect 3881 6752 6224 6780
rect 6288 6752 6736 6780
rect 3881 6749 3893 6752
rect 3835 6743 3893 6749
rect 5994 6644 6000 6656
rect 2746 6616 6000 6644
rect 5994 6604 6000 6616
rect 6052 6604 6058 6656
rect 6196 6644 6224 6752
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 7006 6791 7012 6792
rect 6963 6785 7012 6791
rect 6963 6751 6975 6785
rect 7009 6751 7012 6785
rect 6963 6745 7012 6751
rect 7006 6740 7012 6745
rect 7064 6740 7070 6792
rect 7116 6780 7144 6820
rect 7190 6808 7196 6860
rect 7248 6808 7254 6860
rect 8665 6851 8723 6857
rect 8665 6817 8677 6851
rect 8711 6848 8723 6851
rect 8754 6848 8760 6860
rect 8711 6820 8760 6848
rect 8711 6817 8723 6820
rect 8665 6811 8723 6817
rect 8680 6780 8708 6811
rect 8754 6808 8760 6820
rect 8812 6808 8818 6860
rect 9401 6851 9459 6857
rect 9401 6817 9413 6851
rect 9447 6848 9459 6851
rect 9490 6848 9496 6860
rect 9447 6820 9496 6848
rect 9447 6817 9459 6820
rect 9401 6811 9459 6817
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 11146 6808 11152 6860
rect 11204 6808 11210 6860
rect 11440 6857 11468 6888
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6817 11483 6851
rect 11425 6811 11483 6817
rect 11514 6808 11520 6860
rect 11572 6808 11578 6860
rect 11606 6808 11612 6860
rect 11664 6848 11670 6860
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11664 6820 11989 6848
rect 11664 6808 11670 6820
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 7116 6752 8708 6780
rect 9171 6783 9229 6789
rect 9171 6749 9183 6783
rect 9217 6780 9229 6783
rect 11992 6780 12020 6811
rect 12066 6808 12072 6860
rect 12124 6808 12130 6860
rect 12176 6780 12204 6956
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 14642 6944 14648 6996
rect 14700 6984 14706 6996
rect 15013 6987 15071 6993
rect 15013 6984 15025 6987
rect 14700 6956 15025 6984
rect 14700 6944 14706 6956
rect 15013 6953 15025 6956
rect 15059 6953 15071 6987
rect 15013 6947 15071 6953
rect 15102 6944 15108 6996
rect 15160 6984 15166 6996
rect 16298 6984 16304 6996
rect 15160 6956 16304 6984
rect 15160 6944 15166 6956
rect 16298 6944 16304 6956
rect 16356 6944 16362 6996
rect 16390 6944 16396 6996
rect 16448 6944 16454 6996
rect 18966 6984 18972 6996
rect 18616 6956 18972 6984
rect 14550 6876 14556 6928
rect 14608 6916 14614 6928
rect 14918 6916 14924 6928
rect 14608 6888 14924 6916
rect 14608 6876 14614 6888
rect 14918 6876 14924 6888
rect 14976 6916 14982 6928
rect 16408 6916 16436 6944
rect 14976 6888 16436 6916
rect 14976 6876 14982 6888
rect 12434 6857 12440 6860
rect 12396 6851 12440 6857
rect 12396 6817 12408 6851
rect 12396 6811 12440 6817
rect 12434 6808 12440 6811
rect 12492 6808 12498 6860
rect 12805 6851 12863 6857
rect 12805 6817 12817 6851
rect 12851 6848 12863 6851
rect 13170 6848 13176 6860
rect 12851 6820 13176 6848
rect 12851 6817 12863 6820
rect 12805 6811 12863 6817
rect 13170 6808 13176 6820
rect 13228 6808 13234 6860
rect 13262 6808 13268 6860
rect 13320 6848 13326 6860
rect 14277 6851 14335 6857
rect 14277 6848 14289 6851
rect 13320 6820 14289 6848
rect 13320 6808 13326 6820
rect 14277 6817 14289 6820
rect 14323 6817 14335 6851
rect 14277 6811 14335 6817
rect 15197 6851 15255 6857
rect 15197 6817 15209 6851
rect 15243 6817 15255 6851
rect 15197 6811 15255 6817
rect 15289 6852 15347 6857
rect 15289 6851 15516 6852
rect 15289 6817 15301 6851
rect 15335 6824 15516 6851
rect 15335 6817 15347 6824
rect 15289 6811 15347 6817
rect 9217 6752 11928 6780
rect 11992 6752 12204 6780
rect 12532 6785 12590 6791
rect 9217 6749 9229 6752
rect 9171 6743 9229 6749
rect 8294 6672 8300 6724
rect 8352 6672 8358 6724
rect 10594 6672 10600 6724
rect 10652 6712 10658 6724
rect 10965 6715 11023 6721
rect 10965 6712 10977 6715
rect 10652 6684 10977 6712
rect 10652 6672 10658 6684
rect 10965 6681 10977 6684
rect 11011 6681 11023 6715
rect 10965 6675 11023 6681
rect 11054 6672 11060 6724
rect 11112 6712 11118 6724
rect 11793 6715 11851 6721
rect 11793 6712 11805 6715
rect 11112 6684 11805 6712
rect 11112 6672 11118 6684
rect 11793 6681 11805 6684
rect 11839 6681 11851 6715
rect 11793 6675 11851 6681
rect 7926 6644 7932 6656
rect 6196 6616 7932 6644
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 8386 6604 8392 6656
rect 8444 6644 8450 6656
rect 11606 6644 11612 6656
rect 8444 6616 11612 6644
rect 8444 6604 8450 6616
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 11698 6604 11704 6656
rect 11756 6604 11762 6656
rect 11900 6644 11928 6752
rect 12532 6751 12544 6785
rect 12578 6780 12590 6785
rect 12618 6780 12624 6792
rect 12578 6752 12624 6780
rect 12578 6751 12590 6752
rect 12532 6745 12590 6751
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 13446 6740 13452 6792
rect 13504 6780 13510 6792
rect 15212 6780 15240 6811
rect 13504 6752 15240 6780
rect 15488 6780 15516 6824
rect 15746 6808 15752 6860
rect 15804 6808 15810 6860
rect 15930 6808 15936 6860
rect 15988 6808 15994 6860
rect 16298 6808 16304 6860
rect 16356 6808 16362 6860
rect 16482 6808 16488 6860
rect 16540 6808 16546 6860
rect 18616 6857 18644 6956
rect 18966 6944 18972 6956
rect 19024 6944 19030 6996
rect 20625 6987 20683 6993
rect 20625 6953 20637 6987
rect 20671 6984 20683 6987
rect 21082 6984 21088 6996
rect 20671 6956 21088 6984
rect 20671 6953 20683 6956
rect 20625 6947 20683 6953
rect 21082 6944 21088 6956
rect 21140 6944 21146 6996
rect 21269 6987 21327 6993
rect 21269 6953 21281 6987
rect 21315 6984 21327 6987
rect 21542 6984 21548 6996
rect 21315 6956 21548 6984
rect 21315 6953 21327 6956
rect 21269 6947 21327 6953
rect 21542 6944 21548 6956
rect 21600 6944 21606 6996
rect 23934 6944 23940 6996
rect 23992 6944 23998 6996
rect 24118 6944 24124 6996
rect 24176 6984 24182 6996
rect 26421 6987 26479 6993
rect 24176 6956 25544 6984
rect 24176 6944 24182 6956
rect 22002 6916 22008 6928
rect 21744 6888 22008 6916
rect 21744 6860 21772 6888
rect 22002 6876 22008 6888
rect 22060 6876 22066 6928
rect 24026 6916 24032 6928
rect 23860 6888 24032 6916
rect 18601 6851 18659 6857
rect 17052 6820 18276 6848
rect 15948 6780 15976 6808
rect 15488 6752 15976 6780
rect 16393 6783 16451 6789
rect 13504 6740 13510 6752
rect 16393 6749 16405 6783
rect 16439 6780 16451 6783
rect 16500 6780 16528 6808
rect 16758 6789 16764 6792
rect 16439 6752 16528 6780
rect 16720 6783 16764 6789
rect 16439 6749 16451 6752
rect 16393 6743 16451 6749
rect 16720 6749 16732 6783
rect 16720 6743 16764 6749
rect 13998 6672 14004 6724
rect 14056 6712 14062 6724
rect 15473 6715 15531 6721
rect 15473 6712 15485 6715
rect 14056 6684 15485 6712
rect 14056 6672 14062 6684
rect 15473 6681 15485 6684
rect 15519 6681 15531 6715
rect 16408 6712 16436 6743
rect 16758 6740 16764 6743
rect 16816 6740 16822 6792
rect 16899 6783 16957 6789
rect 16899 6749 16911 6783
rect 16945 6780 16957 6783
rect 17052 6780 17080 6820
rect 18248 6792 18276 6820
rect 18601 6817 18613 6851
rect 18647 6817 18659 6851
rect 20714 6848 20720 6860
rect 18601 6811 18659 6817
rect 19214 6820 20720 6848
rect 16945 6752 17080 6780
rect 16945 6749 16957 6752
rect 16899 6743 16957 6749
rect 17126 6740 17132 6792
rect 17184 6740 17190 6792
rect 18230 6740 18236 6792
rect 18288 6740 18294 6792
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 18928 6783 18986 6789
rect 18928 6780 18940 6783
rect 18840 6752 18940 6780
rect 18840 6740 18846 6752
rect 18928 6749 18940 6752
rect 18974 6749 18986 6783
rect 18928 6743 18986 6749
rect 19107 6785 19165 6791
rect 19107 6751 19119 6785
rect 19153 6780 19165 6785
rect 19214 6780 19242 6820
rect 20714 6808 20720 6820
rect 20772 6808 20778 6860
rect 21085 6851 21143 6857
rect 21085 6817 21097 6851
rect 21131 6848 21143 6851
rect 21453 6851 21511 6857
rect 21131 6820 21404 6848
rect 21131 6817 21143 6820
rect 21085 6811 21143 6817
rect 21376 6792 21404 6820
rect 21453 6817 21465 6851
rect 21499 6817 21511 6851
rect 21453 6811 21511 6817
rect 19153 6752 19242 6780
rect 19337 6783 19395 6789
rect 19153 6751 19165 6752
rect 19107 6745 19165 6751
rect 19337 6749 19349 6783
rect 19383 6780 19395 6783
rect 20530 6780 20536 6792
rect 19383 6752 20536 6780
rect 19383 6749 19395 6752
rect 19337 6743 19395 6749
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 21358 6740 21364 6792
rect 21416 6740 21422 6792
rect 21468 6780 21496 6811
rect 21726 6808 21732 6860
rect 21784 6808 21790 6860
rect 22240 6851 22298 6857
rect 22240 6817 22252 6851
rect 22286 6848 22298 6851
rect 22286 6820 22600 6848
rect 22286 6817 22298 6820
rect 22240 6811 22298 6817
rect 21818 6780 21824 6792
rect 21468 6752 21824 6780
rect 21818 6740 21824 6752
rect 21876 6740 21882 6792
rect 21910 6740 21916 6792
rect 21968 6740 21974 6792
rect 22370 6740 22376 6792
rect 22428 6780 22434 6792
rect 22572 6780 22600 6820
rect 22646 6808 22652 6860
rect 22704 6808 22710 6860
rect 23014 6808 23020 6860
rect 23072 6848 23078 6860
rect 23860 6848 23888 6888
rect 24026 6876 24032 6888
rect 24084 6916 24090 6928
rect 25516 6916 25544 6956
rect 26421 6953 26433 6987
rect 26467 6984 26479 6987
rect 26786 6984 26792 6996
rect 26467 6956 26792 6984
rect 26467 6953 26479 6956
rect 26421 6947 26479 6953
rect 26786 6944 26792 6956
rect 26844 6944 26850 6996
rect 27982 6944 27988 6996
rect 28040 6984 28046 6996
rect 28083 6987 28141 6993
rect 28083 6984 28095 6987
rect 28040 6956 28095 6984
rect 28040 6944 28046 6956
rect 28083 6953 28095 6956
rect 28129 6953 28141 6987
rect 28083 6947 28141 6953
rect 27614 6916 27620 6928
rect 24084 6876 24118 6916
rect 25516 6888 27620 6916
rect 27614 6876 27620 6888
rect 27672 6876 27678 6928
rect 23072 6820 23888 6848
rect 24090 6872 24118 6876
rect 24090 6857 24164 6872
rect 24486 6857 24492 6860
rect 24090 6851 24179 6857
rect 24090 6844 24133 6851
rect 23072 6808 23078 6820
rect 24121 6817 24133 6844
rect 24167 6817 24179 6851
rect 24448 6851 24492 6857
rect 24448 6848 24460 6851
rect 24121 6811 24179 6817
rect 24366 6820 24460 6848
rect 24366 6780 24394 6820
rect 24448 6817 24460 6820
rect 24448 6811 24492 6817
rect 24486 6808 24492 6811
rect 24544 6808 24550 6860
rect 24857 6851 24915 6857
rect 24857 6817 24869 6851
rect 24903 6848 24915 6851
rect 25590 6848 25596 6860
rect 24903 6820 25596 6848
rect 24903 6817 24915 6820
rect 24857 6811 24915 6817
rect 25590 6808 25596 6820
rect 25648 6808 25654 6860
rect 25958 6808 25964 6860
rect 26016 6848 26022 6860
rect 26510 6848 26516 6860
rect 26016 6820 26516 6848
rect 26016 6808 26022 6820
rect 26510 6808 26516 6820
rect 26568 6848 26574 6860
rect 26605 6851 26663 6857
rect 26605 6848 26617 6851
rect 26568 6820 26617 6848
rect 26568 6808 26574 6820
rect 26605 6817 26617 6820
rect 26651 6817 26663 6851
rect 26605 6811 26663 6817
rect 27157 6851 27215 6857
rect 27157 6817 27169 6851
rect 27203 6817 27215 6851
rect 27157 6811 27215 6817
rect 28353 6851 28411 6857
rect 28353 6817 28365 6851
rect 28399 6848 28411 6851
rect 29638 6848 29644 6860
rect 28399 6820 29644 6848
rect 28399 6817 28411 6820
rect 28353 6811 28411 6817
rect 24670 6789 24676 6792
rect 22428 6752 22473 6780
rect 22572 6752 24026 6780
rect 22428 6740 22434 6752
rect 21634 6712 21640 6724
rect 15473 6675 15531 6681
rect 15856 6684 16436 6712
rect 20824 6684 21640 6712
rect 13909 6647 13967 6653
rect 13909 6644 13921 6647
rect 11900 6616 13921 6644
rect 13909 6613 13921 6616
rect 13955 6613 13967 6647
rect 13909 6607 13967 6613
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 15856 6644 15884 6684
rect 14608 6616 15884 6644
rect 14608 6604 14614 6616
rect 15930 6604 15936 6656
rect 15988 6604 15994 6656
rect 16114 6604 16120 6656
rect 16172 6604 16178 6656
rect 18417 6647 18475 6653
rect 18417 6613 18429 6647
rect 18463 6644 18475 6647
rect 20824 6644 20852 6684
rect 21634 6672 21640 6684
rect 21692 6672 21698 6724
rect 23998 6712 24026 6752
rect 24136 6752 24394 6780
rect 24627 6783 24676 6789
rect 24136 6712 24164 6752
rect 24627 6749 24639 6783
rect 24673 6749 24676 6783
rect 24627 6743 24676 6749
rect 24670 6740 24676 6743
rect 24728 6740 24734 6792
rect 26050 6740 26056 6792
rect 26108 6780 26114 6792
rect 27172 6780 27200 6811
rect 29638 6808 29644 6820
rect 29696 6808 29702 6860
rect 29733 6851 29791 6857
rect 29733 6817 29745 6851
rect 29779 6848 29791 6851
rect 30650 6848 30656 6860
rect 29779 6820 30656 6848
rect 29779 6817 29791 6820
rect 29733 6811 29791 6817
rect 30650 6808 30656 6820
rect 30708 6808 30714 6860
rect 27522 6780 27528 6792
rect 26108 6752 27528 6780
rect 26108 6740 26114 6752
rect 27522 6740 27528 6752
rect 27580 6740 27586 6792
rect 27617 6783 27675 6789
rect 27617 6749 27629 6783
rect 27663 6780 27675 6783
rect 27798 6780 27804 6792
rect 27663 6752 27804 6780
rect 27663 6749 27675 6752
rect 27617 6743 27675 6749
rect 27798 6740 27804 6752
rect 27856 6740 27862 6792
rect 28074 6740 28080 6792
rect 28132 6780 28138 6792
rect 28132 6752 28177 6780
rect 28132 6740 28138 6752
rect 29270 6740 29276 6792
rect 29328 6740 29334 6792
rect 23998 6684 24164 6712
rect 25866 6672 25872 6724
rect 25924 6712 25930 6724
rect 25924 6684 27384 6712
rect 25924 6672 25930 6684
rect 18463 6616 20852 6644
rect 20901 6647 20959 6653
rect 18463 6613 18475 6616
rect 18417 6607 18475 6613
rect 20901 6613 20913 6647
rect 20947 6644 20959 6647
rect 21082 6644 21088 6656
rect 20947 6616 21088 6644
rect 20947 6613 20959 6616
rect 20901 6607 20959 6613
rect 21082 6604 21088 6616
rect 21140 6604 21146 6656
rect 21545 6647 21603 6653
rect 21545 6613 21557 6647
rect 21591 6644 21603 6647
rect 22186 6644 22192 6656
rect 21591 6616 22192 6644
rect 21591 6613 21603 6616
rect 21545 6607 21603 6613
rect 22186 6604 22192 6616
rect 22244 6604 22250 6656
rect 22830 6604 22836 6656
rect 22888 6644 22894 6656
rect 25961 6647 26019 6653
rect 25961 6644 25973 6647
rect 22888 6616 25973 6644
rect 22888 6604 22894 6616
rect 25961 6613 25973 6616
rect 26007 6613 26019 6647
rect 25961 6607 26019 6613
rect 26234 6604 26240 6656
rect 26292 6644 26298 6656
rect 26510 6644 26516 6656
rect 26292 6616 26516 6644
rect 26292 6604 26298 6616
rect 26510 6604 26516 6616
rect 26568 6644 26574 6656
rect 27249 6647 27307 6653
rect 27249 6644 27261 6647
rect 26568 6616 27261 6644
rect 26568 6604 26574 6616
rect 27249 6613 27261 6616
rect 27295 6613 27307 6647
rect 27356 6644 27384 6684
rect 29288 6644 29316 6740
rect 27356 6616 29316 6644
rect 27249 6607 27307 6613
rect 552 6554 30912 6576
rect 552 6502 4193 6554
rect 4245 6502 4257 6554
rect 4309 6502 4321 6554
rect 4373 6502 4385 6554
rect 4437 6502 4449 6554
rect 4501 6502 11783 6554
rect 11835 6502 11847 6554
rect 11899 6502 11911 6554
rect 11963 6502 11975 6554
rect 12027 6502 12039 6554
rect 12091 6502 19373 6554
rect 19425 6502 19437 6554
rect 19489 6502 19501 6554
rect 19553 6502 19565 6554
rect 19617 6502 19629 6554
rect 19681 6502 26963 6554
rect 27015 6502 27027 6554
rect 27079 6502 27091 6554
rect 27143 6502 27155 6554
rect 27207 6502 27219 6554
rect 27271 6502 30912 6554
rect 552 6480 30912 6502
rect 5442 6440 5448 6452
rect 2746 6412 5448 6440
rect 1443 6307 1501 6313
rect 1443 6273 1455 6307
rect 1489 6304 1501 6307
rect 2746 6304 2774 6412
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 6362 6440 6368 6452
rect 6104 6412 6368 6440
rect 5813 6375 5871 6381
rect 5813 6341 5825 6375
rect 5859 6341 5871 6375
rect 5813 6335 5871 6341
rect 1489 6276 2774 6304
rect 3053 6307 3111 6313
rect 1489 6273 1501 6276
rect 1443 6267 1501 6273
rect 3053 6273 3065 6307
rect 3099 6304 3111 6307
rect 3835 6307 3893 6313
rect 3099 6276 3740 6304
rect 3099 6273 3111 6276
rect 3053 6267 3111 6273
rect 934 6196 940 6248
rect 992 6196 998 6248
rect 1670 6196 1676 6248
rect 1728 6196 1734 6248
rect 3329 6239 3387 6245
rect 3329 6205 3341 6239
rect 3375 6236 3387 6239
rect 3418 6236 3424 6248
rect 3375 6208 3424 6236
rect 3375 6205 3387 6208
rect 3329 6199 3387 6205
rect 3418 6196 3424 6208
rect 3476 6196 3482 6248
rect 3712 6236 3740 6276
rect 3835 6273 3847 6307
rect 3881 6304 3893 6307
rect 3970 6304 3976 6316
rect 3881 6276 3976 6304
rect 3881 6273 3893 6276
rect 3835 6267 3893 6273
rect 3970 6264 3976 6276
rect 4028 6264 4034 6316
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6304 4123 6307
rect 5828 6304 5856 6335
rect 6104 6313 6132 6412
rect 6362 6400 6368 6412
rect 6420 6400 6426 6452
rect 6638 6400 6644 6452
rect 6696 6440 6702 6452
rect 6696 6412 7512 6440
rect 6696 6400 6702 6412
rect 7484 6372 7512 6412
rect 7926 6400 7932 6452
rect 7984 6400 7990 6452
rect 8294 6400 8300 6452
rect 8352 6400 8358 6452
rect 8941 6443 8999 6449
rect 8941 6409 8953 6443
rect 8987 6440 8999 6443
rect 9674 6440 9680 6452
rect 8987 6412 9680 6440
rect 8987 6409 8999 6412
rect 8941 6403 8999 6409
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 9858 6400 9864 6452
rect 9916 6440 9922 6452
rect 11057 6443 11115 6449
rect 11057 6440 11069 6443
rect 9916 6412 11069 6440
rect 9916 6400 9922 6412
rect 11057 6409 11069 6412
rect 11103 6409 11115 6443
rect 11057 6403 11115 6409
rect 11238 6400 11244 6452
rect 11296 6440 11302 6452
rect 12066 6440 12072 6452
rect 11296 6412 12072 6440
rect 11296 6400 11302 6412
rect 12066 6400 12072 6412
rect 12124 6400 12130 6452
rect 12621 6443 12679 6449
rect 12621 6409 12633 6443
rect 12667 6440 12679 6443
rect 12710 6440 12716 6452
rect 12667 6412 12716 6440
rect 12667 6409 12679 6412
rect 12621 6403 12679 6409
rect 12710 6400 12716 6412
rect 12768 6400 12774 6452
rect 12986 6400 12992 6452
rect 13044 6440 13050 6452
rect 13081 6443 13139 6449
rect 13081 6440 13093 6443
rect 13044 6412 13093 6440
rect 13044 6400 13050 6412
rect 13081 6409 13093 6412
rect 13127 6409 13139 6443
rect 13081 6403 13139 6409
rect 13173 6443 13231 6449
rect 13173 6409 13185 6443
rect 13219 6440 13231 6443
rect 13630 6440 13636 6452
rect 13219 6412 13636 6440
rect 13219 6409 13231 6412
rect 13173 6403 13231 6409
rect 13630 6400 13636 6412
rect 13688 6400 13694 6452
rect 13722 6400 13728 6452
rect 13780 6400 13786 6452
rect 14458 6400 14464 6452
rect 14516 6440 14522 6452
rect 16393 6443 16451 6449
rect 16393 6440 16405 6443
rect 14516 6412 16405 6440
rect 14516 6400 14522 6412
rect 16393 6409 16405 6412
rect 16439 6409 16451 6443
rect 16393 6403 16451 6409
rect 18325 6443 18383 6449
rect 18325 6409 18337 6443
rect 18371 6440 18383 6443
rect 19058 6440 19064 6452
rect 18371 6412 19064 6440
rect 18371 6409 18383 6412
rect 18325 6403 18383 6409
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 20806 6440 20812 6452
rect 19904 6412 20812 6440
rect 8312 6372 8340 6400
rect 7484 6344 8340 6372
rect 10778 6332 10784 6384
rect 10836 6332 10842 6384
rect 11793 6375 11851 6381
rect 11793 6341 11805 6375
rect 11839 6372 11851 6375
rect 14366 6372 14372 6384
rect 11839 6344 14372 6372
rect 11839 6341 11851 6344
rect 11793 6335 11851 6341
rect 14366 6332 14372 6344
rect 14424 6332 14430 6384
rect 6454 6313 6460 6316
rect 4111 6276 5856 6304
rect 6089 6307 6147 6313
rect 4111 6273 4123 6276
rect 4065 6267 4123 6273
rect 6089 6273 6101 6307
rect 6135 6273 6147 6307
rect 6089 6267 6147 6273
rect 6416 6307 6460 6313
rect 6416 6273 6428 6307
rect 6416 6267 6460 6273
rect 6454 6264 6460 6267
rect 6512 6264 6518 6316
rect 6638 6311 6644 6316
rect 6595 6305 6644 6311
rect 6595 6271 6607 6305
rect 6641 6271 6644 6305
rect 6595 6265 6644 6271
rect 6638 6264 6644 6265
rect 6696 6264 6702 6316
rect 6822 6264 6828 6316
rect 6880 6264 6886 6316
rect 7466 6264 7472 6316
rect 7524 6264 7530 6316
rect 8754 6264 8760 6316
rect 8812 6304 8818 6316
rect 9217 6307 9275 6313
rect 9217 6304 9229 6307
rect 8812 6276 9229 6304
rect 8812 6264 8818 6276
rect 9217 6273 9229 6276
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 9398 6264 9404 6316
rect 9456 6304 9462 6316
rect 9544 6307 9602 6313
rect 9544 6304 9556 6307
rect 9456 6276 9556 6304
rect 9456 6264 9462 6276
rect 9544 6273 9556 6276
rect 9590 6273 9602 6307
rect 9544 6267 9602 6273
rect 9723 6307 9781 6313
rect 9723 6273 9735 6307
rect 9769 6304 9781 6307
rect 9953 6307 10011 6313
rect 9769 6276 9904 6304
rect 9769 6273 9781 6276
rect 9723 6267 9781 6273
rect 4798 6236 4804 6248
rect 3712 6208 4804 6236
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 5534 6196 5540 6248
rect 5592 6236 5598 6248
rect 5721 6239 5779 6245
rect 5721 6236 5733 6239
rect 5592 6208 5733 6236
rect 5592 6196 5598 6208
rect 5721 6205 5733 6208
rect 5767 6205 5779 6239
rect 5721 6199 5779 6205
rect 5997 6239 6055 6245
rect 5997 6205 6009 6239
rect 6043 6236 6055 6239
rect 7098 6236 7104 6248
rect 6043 6208 7104 6236
rect 6043 6205 6055 6208
rect 5997 6199 6055 6205
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 7484 6236 7512 6264
rect 8386 6236 8392 6248
rect 7484 6208 8392 6236
rect 8386 6196 8392 6208
rect 8444 6196 8450 6248
rect 8846 6196 8852 6248
rect 8904 6196 8910 6248
rect 9122 6196 9128 6248
rect 9180 6196 9186 6248
rect 9876 6236 9904 6276
rect 9953 6273 9965 6307
rect 9999 6304 10011 6307
rect 10796 6304 10824 6332
rect 13446 6304 13452 6316
rect 9999 6276 10824 6304
rect 11716 6276 13452 6304
rect 9999 6273 10011 6276
rect 9953 6267 10011 6273
rect 10226 6236 10232 6248
rect 9876 6208 10232 6236
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 11422 6196 11428 6248
rect 11480 6236 11486 6248
rect 11716 6245 11744 6276
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 11480 6208 11713 6236
rect 11480 6196 11486 6208
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 11977 6239 12035 6245
rect 11977 6205 11989 6239
rect 12023 6236 12035 6239
rect 12066 6236 12072 6248
rect 12023 6208 12072 6236
rect 12023 6205 12035 6208
rect 11977 6199 12035 6205
rect 12066 6196 12072 6208
rect 12124 6196 12130 6248
rect 12158 6196 12164 6248
rect 12216 6236 12222 6248
rect 12544 6245 12572 6276
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 14274 6264 14280 6316
rect 14332 6304 14338 6316
rect 14734 6304 14740 6316
rect 14332 6276 14504 6304
rect 14332 6264 14338 6276
rect 12802 6245 12808 6248
rect 12253 6239 12311 6245
rect 12253 6236 12265 6239
rect 12216 6208 12265 6236
rect 12216 6196 12222 6208
rect 12253 6205 12265 6208
rect 12299 6205 12311 6239
rect 12253 6199 12311 6205
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6205 12587 6239
rect 12797 6236 12808 6245
rect 12529 6199 12587 6205
rect 12636 6208 12808 6236
rect 8864 6168 8892 6196
rect 7484 6140 9352 6168
rect 1394 6060 1400 6112
rect 1452 6109 1458 6112
rect 1452 6100 1461 6109
rect 3234 6100 3240 6112
rect 1452 6072 3240 6100
rect 1452 6063 1461 6072
rect 1452 6060 1458 6063
rect 3234 6060 3240 6072
rect 3292 6100 3298 6112
rect 3418 6100 3424 6112
rect 3292 6072 3424 6100
rect 3292 6060 3298 6072
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 3694 6060 3700 6112
rect 3752 6100 3758 6112
rect 3795 6103 3853 6109
rect 3795 6100 3807 6103
rect 3752 6072 3807 6100
rect 3752 6060 3758 6072
rect 3795 6069 3807 6072
rect 3841 6069 3853 6103
rect 3795 6063 3853 6069
rect 5166 6060 5172 6112
rect 5224 6060 5230 6112
rect 5537 6103 5595 6109
rect 5537 6069 5549 6103
rect 5583 6100 5595 6103
rect 5626 6100 5632 6112
rect 5583 6072 5632 6100
rect 5583 6069 5595 6072
rect 5537 6063 5595 6069
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 5810 6060 5816 6112
rect 5868 6100 5874 6112
rect 6362 6100 6368 6112
rect 5868 6072 6368 6100
rect 5868 6060 5874 6072
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 7484 6100 7512 6140
rect 6788 6072 7512 6100
rect 6788 6060 6794 6072
rect 8570 6060 8576 6112
rect 8628 6060 8634 6112
rect 8665 6103 8723 6109
rect 8665 6069 8677 6103
rect 8711 6100 8723 6103
rect 9214 6100 9220 6112
rect 8711 6072 9220 6100
rect 8711 6069 8723 6072
rect 8665 6063 8723 6069
rect 9214 6060 9220 6072
rect 9272 6060 9278 6112
rect 9324 6100 9352 6140
rect 11054 6128 11060 6180
rect 11112 6168 11118 6180
rect 12268 6168 12296 6199
rect 12636 6168 12664 6208
rect 12797 6199 12808 6208
rect 12802 6196 12808 6199
rect 12860 6196 12866 6248
rect 12894 6196 12900 6248
rect 12952 6196 12958 6248
rect 13354 6196 13360 6248
rect 13412 6196 13418 6248
rect 13909 6239 13967 6245
rect 13909 6205 13921 6239
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 11112 6140 12664 6168
rect 11112 6128 11118 6140
rect 13630 6128 13636 6180
rect 13688 6168 13694 6180
rect 13924 6168 13952 6199
rect 14090 6196 14096 6248
rect 14148 6196 14154 6248
rect 14476 6168 14504 6276
rect 14568 6276 14740 6304
rect 14568 6245 14596 6276
rect 14660 6274 14694 6276
rect 14734 6264 14740 6276
rect 14792 6264 14798 6316
rect 14918 6313 14924 6316
rect 14880 6307 14924 6313
rect 14880 6273 14892 6307
rect 14880 6267 14924 6273
rect 14918 6264 14924 6267
rect 14976 6264 14982 6316
rect 15059 6307 15117 6313
rect 15059 6273 15071 6307
rect 15105 6304 15117 6307
rect 15378 6304 15384 6316
rect 15105 6276 15384 6304
rect 15105 6273 15117 6276
rect 15059 6267 15117 6273
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 17865 6307 17923 6313
rect 17512 6276 17724 6304
rect 14553 6239 14611 6245
rect 14553 6205 14565 6239
rect 14599 6205 14611 6239
rect 15289 6239 15347 6245
rect 15289 6236 15301 6239
rect 14666 6232 15301 6236
rect 14553 6199 14611 6205
rect 14660 6208 15301 6232
rect 14660 6204 14694 6208
rect 15289 6205 15301 6208
rect 15335 6205 15347 6239
rect 14660 6168 14688 6204
rect 15289 6199 15347 6205
rect 16761 6239 16819 6245
rect 16761 6205 16773 6239
rect 16807 6236 16819 6239
rect 16850 6236 16856 6248
rect 16807 6208 16856 6236
rect 16807 6205 16819 6208
rect 16761 6199 16819 6205
rect 16850 6196 16856 6208
rect 16908 6236 16914 6248
rect 17512 6245 17540 6276
rect 17497 6239 17555 6245
rect 16908 6208 17448 6236
rect 16908 6196 16914 6208
rect 13688 6140 13860 6168
rect 13924 6140 14418 6168
rect 14476 6140 14688 6168
rect 13688 6128 13694 6140
rect 9490 6100 9496 6112
rect 9324 6072 9496 6100
rect 9490 6060 9496 6072
rect 9548 6060 9554 6112
rect 11514 6060 11520 6112
rect 11572 6060 11578 6112
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 11974 6100 11980 6112
rect 11848 6072 11980 6100
rect 11848 6060 11854 6072
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12069 6103 12127 6109
rect 12069 6069 12081 6103
rect 12115 6100 12127 6103
rect 12250 6100 12256 6112
rect 12115 6072 12256 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12250 6060 12256 6072
rect 12308 6060 12314 6112
rect 12345 6103 12403 6109
rect 12345 6069 12357 6103
rect 12391 6100 12403 6103
rect 13354 6100 13360 6112
rect 12391 6072 13360 6100
rect 12391 6069 12403 6072
rect 12345 6063 12403 6069
rect 13354 6060 13360 6072
rect 13412 6060 13418 6112
rect 13832 6100 13860 6140
rect 14185 6103 14243 6109
rect 14185 6100 14197 6103
rect 13832 6072 14197 6100
rect 14185 6069 14197 6072
rect 14231 6069 14243 6103
rect 14390 6100 14418 6140
rect 16666 6128 16672 6180
rect 16724 6168 16730 6180
rect 17037 6171 17095 6177
rect 17037 6168 17049 6171
rect 16724 6140 17049 6168
rect 16724 6128 16730 6140
rect 17037 6137 17049 6140
rect 17083 6137 17095 6171
rect 17420 6168 17448 6208
rect 17497 6205 17509 6239
rect 17543 6205 17555 6239
rect 17497 6199 17555 6205
rect 17589 6239 17647 6245
rect 17589 6205 17601 6239
rect 17635 6205 17647 6239
rect 17696 6236 17724 6276
rect 17865 6273 17877 6307
rect 17911 6304 17923 6307
rect 18782 6304 18788 6316
rect 17911 6276 18788 6304
rect 17911 6273 17923 6276
rect 17865 6267 17923 6273
rect 18782 6264 18788 6276
rect 18840 6264 18846 6316
rect 19904 6313 19932 6412
rect 20806 6400 20812 6412
rect 20864 6400 20870 6452
rect 21082 6400 21088 6452
rect 21140 6440 21146 6452
rect 21140 6412 21496 6440
rect 21140 6400 21146 6412
rect 21468 6372 21496 6412
rect 21634 6400 21640 6452
rect 21692 6440 21698 6452
rect 21692 6412 25452 6440
rect 21692 6400 21698 6412
rect 21468 6344 23520 6372
rect 19889 6307 19947 6313
rect 19168 6276 19748 6304
rect 17696 6208 18184 6236
rect 17589 6199 17647 6205
rect 17604 6168 17632 6199
rect 18156 6180 18184 6208
rect 18506 6196 18512 6248
rect 18564 6196 18570 6248
rect 19168 6245 19196 6276
rect 19720 6245 19748 6276
rect 19889 6273 19901 6307
rect 19935 6273 19947 6307
rect 19889 6267 19947 6273
rect 20395 6307 20453 6313
rect 20395 6273 20407 6307
rect 20441 6304 20453 6307
rect 20441 6276 20760 6304
rect 20441 6273 20453 6276
rect 20395 6267 20453 6273
rect 20732 6248 20760 6276
rect 21910 6264 21916 6316
rect 21968 6304 21974 6316
rect 23014 6304 23020 6316
rect 21968 6276 23020 6304
rect 21968 6264 21974 6276
rect 23014 6264 23020 6276
rect 23072 6264 23078 6316
rect 23382 6264 23388 6316
rect 23440 6264 23446 6316
rect 23492 6304 23520 6344
rect 24210 6304 24216 6316
rect 23492 6276 24216 6304
rect 24210 6264 24216 6276
rect 24268 6264 24274 6316
rect 24535 6307 24593 6313
rect 24535 6273 24547 6307
rect 24581 6304 24593 6307
rect 25424 6304 25452 6412
rect 27614 6400 27620 6452
rect 27672 6440 27678 6452
rect 28537 6443 28595 6449
rect 28537 6440 28549 6443
rect 27672 6412 28549 6440
rect 27672 6400 27678 6412
rect 28537 6409 28549 6412
rect 28583 6409 28595 6443
rect 28537 6403 28595 6409
rect 28166 6332 28172 6384
rect 28224 6372 28230 6384
rect 28224 6344 28994 6372
rect 28224 6332 28230 6344
rect 27160 6305 27218 6311
rect 24581 6276 25176 6304
rect 25424 6302 27016 6304
rect 27160 6302 27172 6305
rect 25424 6276 27172 6302
rect 24581 6273 24593 6276
rect 24535 6267 24593 6273
rect 20254 6245 20260 6248
rect 18877 6239 18935 6245
rect 18877 6205 18889 6239
rect 18923 6205 18935 6239
rect 18877 6199 18935 6205
rect 19153 6239 19211 6245
rect 19153 6205 19165 6239
rect 19199 6205 19211 6239
rect 19153 6199 19211 6205
rect 19429 6239 19487 6245
rect 19429 6205 19441 6239
rect 19475 6236 19487 6239
rect 19705 6239 19763 6245
rect 19475 6208 19509 6236
rect 19475 6205 19487 6208
rect 19429 6199 19487 6205
rect 19705 6205 19717 6239
rect 19751 6236 19763 6239
rect 20216 6239 20260 6245
rect 19751 6208 20024 6236
rect 19751 6205 19763 6208
rect 19705 6199 19763 6205
rect 17862 6168 17868 6180
rect 17420 6140 17868 6168
rect 17037 6131 17095 6137
rect 17862 6128 17868 6140
rect 17920 6128 17926 6180
rect 18138 6128 18144 6180
rect 18196 6128 18202 6180
rect 18892 6168 18920 6199
rect 19444 6168 19472 6199
rect 19996 6180 20024 6208
rect 20216 6205 20228 6239
rect 20216 6199 20260 6205
rect 20254 6196 20260 6199
rect 20312 6196 20318 6248
rect 20622 6196 20628 6248
rect 20680 6196 20686 6248
rect 20714 6196 20720 6248
rect 20772 6196 20778 6248
rect 22281 6239 22339 6245
rect 22281 6205 22293 6239
rect 22327 6236 22339 6239
rect 22327 6208 22416 6236
rect 22327 6205 22339 6208
rect 22281 6199 22339 6205
rect 18892 6140 19656 6168
rect 15378 6100 15384 6112
rect 14390 6072 15384 6100
rect 14185 6063 14243 6069
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 17310 6060 17316 6112
rect 17368 6060 17374 6112
rect 18414 6060 18420 6112
rect 18472 6100 18478 6112
rect 18693 6103 18751 6109
rect 18693 6100 18705 6103
rect 18472 6072 18705 6100
rect 18472 6060 18478 6072
rect 18693 6069 18705 6072
rect 18739 6069 18751 6103
rect 18693 6063 18751 6069
rect 18966 6060 18972 6112
rect 19024 6060 19030 6112
rect 19058 6060 19064 6112
rect 19116 6100 19122 6112
rect 19245 6103 19303 6109
rect 19245 6100 19257 6103
rect 19116 6072 19257 6100
rect 19116 6060 19122 6072
rect 19245 6069 19257 6072
rect 19291 6069 19303 6103
rect 19245 6063 19303 6069
rect 19518 6060 19524 6112
rect 19576 6060 19582 6112
rect 19628 6100 19656 6140
rect 19978 6128 19984 6180
rect 20036 6128 20042 6180
rect 21634 6128 21640 6180
rect 21692 6168 21698 6180
rect 21818 6168 21824 6180
rect 21692 6140 21824 6168
rect 21692 6128 21698 6140
rect 21818 6128 21824 6140
rect 21876 6168 21882 6180
rect 22388 6168 22416 6208
rect 22554 6196 22560 6248
rect 22612 6196 22618 6248
rect 22738 6196 22744 6248
rect 22796 6196 22802 6248
rect 23566 6196 23572 6248
rect 23624 6196 23630 6248
rect 24029 6239 24087 6245
rect 24029 6205 24041 6239
rect 24075 6205 24087 6239
rect 24029 6199 24087 6205
rect 23584 6168 23612 6196
rect 24044 6168 24072 6199
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 25148 6236 25176 6276
rect 26988 6274 27172 6276
rect 27160 6271 27172 6274
rect 27206 6271 27218 6305
rect 27160 6265 27218 6271
rect 27433 6307 27491 6313
rect 27433 6273 27445 6307
rect 27479 6304 27491 6307
rect 28534 6304 28540 6316
rect 27479 6276 28540 6304
rect 27479 6273 27491 6276
rect 27433 6267 27491 6273
rect 28534 6264 28540 6276
rect 28592 6264 28598 6316
rect 25148 6208 25636 6236
rect 25608 6180 25636 6208
rect 26050 6196 26056 6248
rect 26108 6236 26114 6248
rect 26602 6236 26608 6248
rect 26108 6208 26608 6236
rect 26108 6196 26114 6208
rect 26602 6196 26608 6208
rect 26660 6236 26666 6248
rect 26697 6239 26755 6245
rect 26697 6236 26709 6239
rect 26660 6208 26709 6236
rect 26660 6196 26666 6208
rect 26697 6205 26709 6208
rect 26743 6205 26755 6239
rect 28626 6236 28632 6248
rect 26697 6199 26755 6205
rect 26804 6208 28632 6236
rect 21876 6140 23612 6168
rect 23860 6140 24072 6168
rect 21876 6128 21882 6140
rect 21652 6100 21680 6128
rect 23860 6112 23888 6140
rect 25590 6128 25596 6180
rect 25648 6128 25654 6180
rect 26145 6171 26203 6177
rect 26145 6137 26157 6171
rect 26191 6168 26203 6171
rect 26418 6168 26424 6180
rect 26191 6140 26424 6168
rect 26191 6137 26203 6140
rect 26145 6131 26203 6137
rect 26418 6128 26424 6140
rect 26476 6128 26482 6180
rect 19628 6072 21680 6100
rect 21910 6060 21916 6112
rect 21968 6060 21974 6112
rect 22094 6060 22100 6112
rect 22152 6060 22158 6112
rect 22373 6103 22431 6109
rect 22373 6069 22385 6103
rect 22419 6100 22431 6103
rect 22554 6100 22560 6112
rect 22419 6072 22560 6100
rect 22419 6069 22431 6072
rect 22373 6063 22431 6069
rect 22554 6060 22560 6072
rect 22612 6060 22618 6112
rect 23842 6060 23848 6112
rect 23900 6060 23906 6112
rect 24486 6060 24492 6112
rect 24544 6109 24550 6112
rect 24544 6063 24553 6109
rect 24544 6060 24550 6063
rect 24670 6060 24676 6112
rect 24728 6100 24734 6112
rect 26804 6100 26832 6208
rect 28626 6196 28632 6208
rect 28684 6196 28690 6248
rect 28966 6236 28994 6344
rect 29181 6239 29239 6245
rect 29181 6236 29193 6239
rect 28966 6208 29193 6236
rect 29181 6205 29193 6208
rect 29227 6205 29239 6239
rect 29181 6199 29239 6205
rect 24728 6072 26832 6100
rect 24728 6060 24734 6072
rect 26970 6060 26976 6112
rect 27028 6100 27034 6112
rect 27154 6100 27160 6112
rect 27212 6109 27218 6112
rect 27028 6072 27160 6100
rect 27028 6060 27034 6072
rect 27154 6060 27160 6072
rect 27212 6063 27221 6109
rect 27212 6060 27218 6063
rect 27338 6060 27344 6112
rect 27396 6100 27402 6112
rect 27798 6100 27804 6112
rect 27396 6072 27804 6100
rect 27396 6060 27402 6072
rect 27798 6060 27804 6072
rect 27856 6060 27862 6112
rect 28997 6103 29055 6109
rect 28997 6069 29009 6103
rect 29043 6100 29055 6103
rect 29270 6100 29276 6112
rect 29043 6072 29276 6100
rect 29043 6069 29055 6072
rect 28997 6063 29055 6069
rect 29270 6060 29276 6072
rect 29328 6060 29334 6112
rect 552 6010 31072 6032
rect 552 5958 7988 6010
rect 8040 5958 8052 6010
rect 8104 5958 8116 6010
rect 8168 5958 8180 6010
rect 8232 5958 8244 6010
rect 8296 5958 15578 6010
rect 15630 5958 15642 6010
rect 15694 5958 15706 6010
rect 15758 5958 15770 6010
rect 15822 5958 15834 6010
rect 15886 5958 23168 6010
rect 23220 5958 23232 6010
rect 23284 5958 23296 6010
rect 23348 5958 23360 6010
rect 23412 5958 23424 6010
rect 23476 5958 30758 6010
rect 30810 5958 30822 6010
rect 30874 5958 30886 6010
rect 30938 5958 30950 6010
rect 31002 5958 31014 6010
rect 31066 5958 31072 6010
rect 552 5936 31072 5958
rect 845 5899 903 5905
rect 845 5865 857 5899
rect 891 5896 903 5899
rect 1946 5896 1952 5908
rect 891 5868 1952 5896
rect 891 5865 903 5868
rect 845 5859 903 5865
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 5166 5896 5172 5908
rect 2746 5868 5172 5896
rect 1026 5720 1032 5772
rect 1084 5720 1090 5772
rect 1394 5720 1400 5772
rect 1452 5760 1458 5772
rect 1632 5763 1690 5769
rect 1632 5760 1644 5763
rect 1452 5732 1644 5760
rect 1452 5720 1458 5732
rect 1632 5729 1644 5732
rect 1678 5729 1690 5763
rect 2746 5760 2774 5868
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 5350 5856 5356 5908
rect 5408 5896 5414 5908
rect 7193 5899 7251 5905
rect 7193 5896 7205 5899
rect 5408 5868 7205 5896
rect 5408 5856 5414 5868
rect 7193 5865 7205 5868
rect 7239 5865 7251 5899
rect 7193 5859 7251 5865
rect 8303 5899 8361 5905
rect 8303 5865 8315 5899
rect 8349 5896 8361 5899
rect 8478 5896 8484 5908
rect 8349 5868 8484 5896
rect 8349 5865 8361 5868
rect 8303 5859 8361 5865
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 8662 5856 8668 5908
rect 8720 5896 8726 5908
rect 8720 5868 10732 5896
rect 8720 5856 8726 5868
rect 10704 5840 10732 5868
rect 10778 5856 10784 5908
rect 10836 5856 10842 5908
rect 11057 5899 11115 5905
rect 11057 5865 11069 5899
rect 11103 5896 11115 5899
rect 11103 5868 11744 5896
rect 11103 5865 11115 5868
rect 11057 5859 11115 5865
rect 6086 5788 6092 5840
rect 6144 5788 6150 5840
rect 6656 5800 7696 5828
rect 6656 5772 6684 5800
rect 7668 5772 7696 5800
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 9824 5800 10640 5828
rect 9824 5788 9830 5800
rect 1632 5723 1690 5729
rect 1964 5732 2774 5760
rect 1801 5713 1859 5719
rect 934 5652 940 5704
rect 992 5692 998 5704
rect 1305 5695 1363 5701
rect 1305 5692 1317 5695
rect 992 5664 1317 5692
rect 992 5652 998 5664
rect 1305 5661 1317 5664
rect 1351 5661 1363 5695
rect 1801 5679 1813 5713
rect 1847 5692 1859 5713
rect 1964 5692 1992 5732
rect 3602 5720 3608 5772
rect 3660 5760 3666 5772
rect 3840 5763 3898 5769
rect 3840 5760 3852 5763
rect 3660 5732 3852 5760
rect 3660 5720 3666 5732
rect 3840 5729 3852 5732
rect 3886 5760 3898 5763
rect 4522 5760 4528 5772
rect 3886 5732 4528 5760
rect 3886 5729 3898 5732
rect 3840 5723 3898 5729
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 5534 5720 5540 5772
rect 5592 5720 5598 5772
rect 5810 5720 5816 5772
rect 5868 5720 5874 5772
rect 6178 5720 6184 5772
rect 6236 5760 6242 5772
rect 6549 5763 6607 5769
rect 6549 5760 6561 5763
rect 6236 5732 6561 5760
rect 6236 5720 6242 5732
rect 6549 5729 6561 5732
rect 6595 5760 6607 5763
rect 6638 5760 6644 5772
rect 6595 5732 6644 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 6825 5763 6883 5769
rect 6825 5729 6837 5763
rect 6871 5729 6883 5763
rect 6825 5723 6883 5729
rect 1847 5679 1992 5692
rect 1801 5673 1992 5679
rect 1816 5664 1992 5673
rect 1305 5655 1363 5661
rect 2038 5652 2044 5704
rect 2096 5652 2102 5704
rect 2866 5652 2872 5704
rect 2924 5692 2930 5704
rect 3513 5695 3571 5701
rect 3513 5692 3525 5695
rect 2924 5664 3525 5692
rect 2924 5652 2930 5664
rect 3513 5661 3525 5664
rect 3559 5692 3571 5695
rect 3694 5692 3700 5704
rect 3559 5664 3700 5692
rect 3559 5661 3571 5664
rect 3513 5655 3571 5661
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 4062 5701 4068 5704
rect 4019 5695 4068 5701
rect 4019 5661 4031 5695
rect 4065 5661 4068 5695
rect 4019 5655 4068 5661
rect 4062 5652 4068 5655
rect 4120 5652 4126 5704
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 4706 5692 4712 5704
rect 4295 5664 4712 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 5552 5692 5580 5720
rect 6840 5692 6868 5723
rect 7098 5720 7104 5772
rect 7156 5720 7162 5772
rect 7377 5763 7435 5769
rect 7377 5760 7389 5763
rect 7208 5732 7389 5760
rect 7208 5704 7236 5732
rect 7377 5729 7389 5732
rect 7423 5729 7435 5763
rect 7377 5723 7435 5729
rect 7650 5720 7656 5772
rect 7708 5720 7714 5772
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 8573 5763 8631 5769
rect 8573 5760 8585 5763
rect 7800 5732 8585 5760
rect 7800 5720 7806 5732
rect 8573 5729 8585 5732
rect 8619 5729 8631 5763
rect 8573 5723 8631 5729
rect 10229 5763 10287 5769
rect 10229 5729 10241 5763
rect 10275 5729 10287 5763
rect 10229 5723 10287 5729
rect 5552 5664 6868 5692
rect 5442 5584 5448 5636
rect 5500 5624 5506 5636
rect 6641 5627 6699 5633
rect 6641 5624 6653 5627
rect 5500 5596 6653 5624
rect 5500 5584 5506 5596
rect 6641 5593 6653 5596
rect 6687 5593 6699 5627
rect 6840 5624 6868 5664
rect 7190 5652 7196 5704
rect 7248 5652 7254 5704
rect 7834 5652 7840 5704
rect 7892 5652 7898 5704
rect 8386 5701 8392 5704
rect 8343 5695 8392 5701
rect 8343 5661 8355 5695
rect 8389 5661 8392 5695
rect 8343 5655 8392 5661
rect 8386 5652 8392 5655
rect 8444 5652 8450 5704
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5692 10011 5695
rect 10134 5692 10140 5704
rect 9999 5664 10140 5692
rect 9999 5661 10011 5664
rect 9953 5655 10011 5661
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 10244 5692 10272 5723
rect 10502 5720 10508 5772
rect 10560 5720 10566 5772
rect 10612 5769 10640 5800
rect 10686 5788 10692 5840
rect 10744 5788 10750 5840
rect 10597 5763 10655 5769
rect 10597 5729 10609 5763
rect 10643 5760 10655 5763
rect 10778 5760 10784 5772
rect 10643 5732 10784 5760
rect 10643 5729 10655 5732
rect 10597 5723 10655 5729
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 11054 5720 11060 5772
rect 11112 5720 11118 5772
rect 11238 5720 11244 5772
rect 11296 5720 11302 5772
rect 11517 5763 11575 5769
rect 11517 5760 11529 5763
rect 11348 5732 11529 5760
rect 11072 5692 11100 5720
rect 11348 5692 11376 5732
rect 11517 5729 11529 5732
rect 11563 5729 11575 5763
rect 11517 5723 11575 5729
rect 11606 5720 11612 5772
rect 11664 5720 11670 5772
rect 11716 5760 11744 5868
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 12075 5899 12133 5905
rect 12075 5896 12087 5899
rect 12032 5868 12087 5896
rect 12032 5856 12038 5868
rect 12075 5865 12087 5868
rect 12121 5865 12133 5899
rect 12075 5859 12133 5865
rect 12250 5856 12256 5908
rect 12308 5896 12314 5908
rect 13906 5896 13912 5908
rect 12308 5868 13912 5896
rect 12308 5856 12314 5868
rect 13906 5856 13912 5868
rect 13964 5856 13970 5908
rect 20530 5856 20536 5908
rect 20588 5856 20594 5908
rect 20622 5856 20628 5908
rect 20680 5896 20686 5908
rect 20809 5899 20867 5905
rect 20809 5896 20821 5899
rect 20680 5868 20821 5896
rect 20680 5856 20686 5868
rect 20809 5865 20821 5868
rect 20855 5865 20867 5899
rect 20809 5859 20867 5865
rect 21910 5856 21916 5908
rect 21968 5856 21974 5908
rect 24486 5856 24492 5908
rect 24544 5896 24550 5908
rect 24587 5899 24645 5905
rect 24587 5896 24599 5899
rect 24544 5868 24599 5896
rect 24544 5856 24550 5868
rect 24587 5865 24599 5868
rect 24633 5865 24645 5899
rect 24587 5859 24645 5865
rect 26694 5856 26700 5908
rect 26752 5896 26758 5908
rect 26752 5868 27292 5896
rect 26752 5856 26758 5868
rect 19978 5788 19984 5840
rect 20036 5828 20042 5840
rect 20036 5800 21772 5828
rect 20036 5788 20042 5800
rect 12345 5763 12403 5769
rect 12345 5760 12357 5763
rect 11716 5732 12357 5760
rect 12345 5729 12357 5732
rect 12391 5729 12403 5763
rect 12345 5723 12403 5729
rect 13725 5763 13783 5769
rect 13725 5729 13737 5763
rect 13771 5760 13783 5763
rect 13771 5732 14323 5760
rect 13771 5729 13783 5732
rect 13725 5723 13783 5729
rect 12072 5695 12130 5701
rect 12072 5692 12084 5695
rect 10244 5664 11376 5692
rect 11440 5664 12084 5692
rect 6840 5596 7880 5624
rect 6641 5587 6699 5593
rect 1486 5516 1492 5568
rect 1544 5556 1550 5568
rect 2038 5556 2044 5568
rect 1544 5528 2044 5556
rect 1544 5516 1550 5528
rect 2038 5516 2044 5528
rect 2096 5516 2102 5568
rect 3329 5559 3387 5565
rect 3329 5525 3341 5559
rect 3375 5556 3387 5559
rect 3970 5556 3976 5568
rect 3375 5528 3976 5556
rect 3375 5525 3387 5528
rect 3329 5519 3387 5525
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 5534 5516 5540 5568
rect 5592 5516 5598 5568
rect 6365 5559 6423 5565
rect 6365 5525 6377 5559
rect 6411 5556 6423 5559
rect 6546 5556 6552 5568
rect 6411 5528 6552 5556
rect 6411 5525 6423 5528
rect 6365 5519 6423 5525
rect 6546 5516 6552 5528
rect 6604 5516 6610 5568
rect 6730 5516 6736 5568
rect 6788 5556 6794 5568
rect 6917 5559 6975 5565
rect 6917 5556 6929 5559
rect 6788 5528 6929 5556
rect 6788 5516 6794 5528
rect 6917 5525 6929 5528
rect 6963 5525 6975 5559
rect 6917 5519 6975 5525
rect 7466 5516 7472 5568
rect 7524 5516 7530 5568
rect 7852 5556 7880 5596
rect 9490 5584 9496 5636
rect 9548 5624 9554 5636
rect 10502 5624 10508 5636
rect 9548 5596 10508 5624
rect 9548 5584 9554 5596
rect 10502 5584 10508 5596
rect 10560 5584 10566 5636
rect 11238 5584 11244 5636
rect 11296 5624 11302 5636
rect 11440 5624 11468 5664
rect 12072 5661 12084 5664
rect 12118 5661 12130 5695
rect 12072 5655 12130 5661
rect 13814 5652 13820 5704
rect 13872 5652 13878 5704
rect 14182 5701 14188 5704
rect 14144 5695 14188 5701
rect 14144 5661 14156 5695
rect 14144 5655 14188 5661
rect 14182 5652 14188 5655
rect 14240 5652 14246 5704
rect 14295 5703 14323 5732
rect 14366 5720 14372 5772
rect 14424 5760 14430 5772
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 14424 5732 14565 5760
rect 14424 5720 14430 5732
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 16444 5763 16502 5769
rect 16444 5729 16456 5763
rect 16490 5760 16502 5763
rect 16666 5760 16672 5772
rect 16490 5732 16672 5760
rect 16490 5729 16502 5732
rect 16444 5723 16502 5729
rect 16666 5720 16672 5732
rect 16724 5720 16730 5772
rect 16853 5763 16911 5769
rect 16853 5729 16865 5763
rect 16899 5760 16911 5763
rect 17310 5760 17316 5772
rect 16899 5732 17316 5760
rect 16899 5729 16911 5732
rect 16853 5723 16911 5729
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 18138 5720 18144 5772
rect 18196 5760 18202 5772
rect 19061 5763 19119 5769
rect 18196 5732 18920 5760
rect 18196 5720 18202 5732
rect 18524 5704 18552 5732
rect 14280 5697 14338 5703
rect 14280 5663 14292 5697
rect 14326 5663 14338 5697
rect 14280 5657 14338 5663
rect 15930 5652 15936 5704
rect 15988 5692 15994 5704
rect 16117 5695 16175 5701
rect 16117 5692 16129 5695
rect 15988 5664 16129 5692
rect 15988 5652 15994 5664
rect 16117 5661 16129 5664
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 16574 5652 16580 5704
rect 16632 5652 16638 5704
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5661 18383 5695
rect 18325 5655 18383 5661
rect 11296 5596 11468 5624
rect 11296 5584 11302 5596
rect 8662 5556 8668 5568
rect 7852 5528 8668 5556
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 10042 5516 10048 5568
rect 10100 5516 10106 5568
rect 10321 5559 10379 5565
rect 10321 5525 10333 5559
rect 10367 5556 10379 5559
rect 10962 5556 10968 5568
rect 10367 5528 10968 5556
rect 10367 5525 10379 5528
rect 10321 5519 10379 5525
rect 10962 5516 10968 5528
rect 11020 5516 11026 5568
rect 11333 5559 11391 5565
rect 11333 5525 11345 5559
rect 11379 5556 11391 5559
rect 12250 5556 12256 5568
rect 11379 5528 12256 5556
rect 11379 5525 11391 5528
rect 11333 5519 11391 5525
rect 12250 5516 12256 5528
rect 12308 5516 12314 5568
rect 15841 5559 15899 5565
rect 15841 5525 15853 5559
rect 15887 5556 15899 5559
rect 16758 5556 16764 5568
rect 15887 5528 16764 5556
rect 15887 5525 15899 5528
rect 15841 5519 15899 5525
rect 16758 5516 16764 5528
rect 16816 5516 16822 5568
rect 18138 5516 18144 5568
rect 18196 5516 18202 5568
rect 18340 5556 18368 5655
rect 18506 5652 18512 5704
rect 18564 5652 18570 5704
rect 18690 5701 18696 5704
rect 18652 5695 18696 5701
rect 18652 5661 18664 5695
rect 18652 5655 18696 5661
rect 18690 5652 18696 5655
rect 18748 5652 18754 5704
rect 18782 5652 18788 5704
rect 18840 5652 18846 5704
rect 18892 5692 18920 5732
rect 19061 5729 19073 5763
rect 19107 5760 19119 5763
rect 19518 5760 19524 5772
rect 19107 5732 19524 5760
rect 19107 5729 19119 5732
rect 19061 5723 19119 5729
rect 19518 5720 19524 5732
rect 19576 5720 19582 5772
rect 20732 5769 20760 5800
rect 20717 5763 20775 5769
rect 20717 5729 20729 5763
rect 20763 5729 20775 5763
rect 20717 5723 20775 5729
rect 20993 5763 21051 5769
rect 20993 5729 21005 5763
rect 21039 5729 21051 5763
rect 20993 5723 21051 5729
rect 21453 5763 21511 5769
rect 21453 5729 21465 5763
rect 21499 5760 21511 5763
rect 21634 5760 21640 5772
rect 21499 5732 21640 5760
rect 21499 5729 21511 5732
rect 21453 5723 21511 5729
rect 21008 5692 21036 5723
rect 21634 5720 21640 5732
rect 21692 5720 21698 5772
rect 21744 5769 21772 5800
rect 21729 5763 21787 5769
rect 21729 5729 21741 5763
rect 21775 5760 21787 5763
rect 21818 5760 21824 5772
rect 21775 5732 21824 5760
rect 21775 5729 21787 5732
rect 21729 5723 21787 5729
rect 21818 5720 21824 5732
rect 21876 5720 21882 5772
rect 21928 5760 21956 5856
rect 26050 5788 26056 5840
rect 26108 5828 26114 5840
rect 26326 5828 26332 5840
rect 26108 5800 26332 5828
rect 26108 5788 26114 5800
rect 26326 5788 26332 5800
rect 26384 5828 26390 5840
rect 27062 5828 27068 5840
rect 26384 5800 27068 5828
rect 26384 5788 26390 5800
rect 22296 5760 22419 5764
rect 21928 5736 22419 5760
rect 21928 5732 22324 5736
rect 18892 5664 21772 5692
rect 21269 5627 21327 5633
rect 21269 5593 21281 5627
rect 21315 5624 21327 5627
rect 21634 5624 21640 5636
rect 21315 5596 21640 5624
rect 21315 5593 21327 5596
rect 21269 5587 21327 5593
rect 21634 5584 21640 5596
rect 21692 5584 21698 5636
rect 18598 5556 18604 5568
rect 18340 5528 18604 5556
rect 18598 5516 18604 5528
rect 18656 5516 18662 5568
rect 20346 5516 20352 5568
rect 20404 5516 20410 5568
rect 21082 5516 21088 5568
rect 21140 5556 21146 5568
rect 21545 5559 21603 5565
rect 21545 5556 21557 5559
rect 21140 5528 21557 5556
rect 21140 5516 21146 5528
rect 21545 5525 21557 5528
rect 21591 5525 21603 5559
rect 21744 5556 21772 5664
rect 21910 5652 21916 5704
rect 21968 5652 21974 5704
rect 22278 5701 22284 5704
rect 22240 5695 22284 5701
rect 22240 5661 22252 5695
rect 22240 5655 22284 5661
rect 22278 5652 22284 5655
rect 22336 5652 22342 5704
rect 22391 5703 22419 5736
rect 22554 5720 22560 5772
rect 22612 5760 22618 5772
rect 26896 5769 26924 5800
rect 27062 5788 27068 5800
rect 27120 5788 27126 5840
rect 22649 5763 22707 5769
rect 22649 5760 22661 5763
rect 22612 5732 22661 5760
rect 22612 5720 22618 5732
rect 22649 5729 22661 5732
rect 22695 5729 22707 5763
rect 22649 5723 22707 5729
rect 24029 5763 24087 5769
rect 24029 5729 24041 5763
rect 24075 5760 24087 5763
rect 26605 5763 26663 5769
rect 24075 5732 24624 5760
rect 24075 5729 24087 5732
rect 24029 5723 24087 5729
rect 22376 5697 22434 5703
rect 22376 5663 22388 5697
rect 22422 5663 22434 5697
rect 22376 5657 22434 5663
rect 23842 5652 23848 5704
rect 23900 5692 23906 5704
rect 24596 5701 24624 5732
rect 26605 5729 26617 5763
rect 26651 5729 26663 5763
rect 26605 5723 26663 5729
rect 26881 5763 26939 5769
rect 26881 5729 26893 5763
rect 26927 5729 26939 5763
rect 26881 5723 26939 5729
rect 24121 5695 24179 5701
rect 24121 5692 24133 5695
rect 23900 5664 24133 5692
rect 23900 5652 23906 5664
rect 24121 5661 24133 5664
rect 24167 5661 24179 5695
rect 24121 5655 24179 5661
rect 24584 5695 24642 5701
rect 24584 5661 24596 5695
rect 24630 5661 24642 5695
rect 24584 5655 24642 5661
rect 24854 5652 24860 5704
rect 24912 5652 24918 5704
rect 25866 5652 25872 5704
rect 25924 5692 25930 5704
rect 26142 5692 26148 5704
rect 25924 5664 26148 5692
rect 25924 5652 25930 5664
rect 26142 5652 26148 5664
rect 26200 5692 26206 5704
rect 26620 5692 26648 5723
rect 26970 5720 26976 5772
rect 27028 5760 27034 5772
rect 27157 5763 27215 5769
rect 27157 5760 27169 5763
rect 27028 5732 27169 5760
rect 27028 5720 27034 5732
rect 27157 5729 27169 5732
rect 27203 5729 27215 5763
rect 27264 5760 27292 5868
rect 27522 5856 27528 5908
rect 27580 5856 27586 5908
rect 27991 5899 28049 5905
rect 27991 5896 28003 5899
rect 27632 5868 28003 5896
rect 27540 5769 27568 5856
rect 27433 5763 27491 5769
rect 27433 5760 27445 5763
rect 27264 5732 27445 5760
rect 27157 5723 27215 5729
rect 27433 5729 27445 5732
rect 27479 5729 27491 5763
rect 27433 5723 27491 5729
rect 27533 5763 27591 5769
rect 27533 5729 27545 5763
rect 27579 5729 27591 5763
rect 27533 5723 27591 5729
rect 26200 5664 26648 5692
rect 26200 5652 26206 5664
rect 27338 5652 27344 5704
rect 27396 5692 27402 5704
rect 27632 5694 27660 5868
rect 27991 5865 28003 5868
rect 28037 5865 28049 5899
rect 27991 5859 28049 5865
rect 29362 5856 29368 5908
rect 29420 5856 29426 5908
rect 27798 5720 27804 5772
rect 27856 5760 27862 5772
rect 28261 5763 28319 5769
rect 28261 5760 28273 5763
rect 27856 5732 28273 5760
rect 27856 5720 27862 5732
rect 28261 5729 28273 5732
rect 28307 5729 28319 5763
rect 28261 5723 28319 5729
rect 27540 5692 27660 5694
rect 27396 5666 27660 5692
rect 28031 5695 28089 5701
rect 27396 5664 27568 5666
rect 27396 5652 27402 5664
rect 28031 5661 28043 5695
rect 28077 5692 28089 5695
rect 28166 5692 28172 5704
rect 28077 5664 28172 5692
rect 28077 5661 28089 5664
rect 28031 5655 28089 5661
rect 28166 5652 28172 5664
rect 28224 5652 28230 5704
rect 26421 5627 26479 5633
rect 26421 5593 26433 5627
rect 26467 5624 26479 5627
rect 26786 5624 26792 5636
rect 26467 5596 26792 5624
rect 26467 5593 26479 5596
rect 26421 5587 26479 5593
rect 26786 5584 26792 5596
rect 26844 5584 26850 5636
rect 22462 5556 22468 5568
rect 21744 5528 22468 5556
rect 21545 5519 21603 5525
rect 22462 5516 22468 5528
rect 22520 5516 22526 5568
rect 26142 5516 26148 5568
rect 26200 5516 26206 5568
rect 26694 5516 26700 5568
rect 26752 5516 26758 5568
rect 26878 5516 26884 5568
rect 26936 5556 26942 5568
rect 26973 5559 27031 5565
rect 26973 5556 26985 5559
rect 26936 5528 26985 5556
rect 26936 5516 26942 5528
rect 26973 5525 26985 5528
rect 27019 5525 27031 5559
rect 26973 5519 27031 5525
rect 27249 5559 27307 5565
rect 27249 5525 27261 5559
rect 27295 5556 27307 5559
rect 28166 5556 28172 5568
rect 27295 5528 28172 5556
rect 27295 5525 27307 5528
rect 27249 5519 27307 5525
rect 28166 5516 28172 5528
rect 28224 5516 28230 5568
rect 552 5466 30912 5488
rect 552 5414 4193 5466
rect 4245 5414 4257 5466
rect 4309 5414 4321 5466
rect 4373 5414 4385 5466
rect 4437 5414 4449 5466
rect 4501 5414 11783 5466
rect 11835 5414 11847 5466
rect 11899 5414 11911 5466
rect 11963 5414 11975 5466
rect 12027 5414 12039 5466
rect 12091 5414 19373 5466
rect 19425 5414 19437 5466
rect 19489 5414 19501 5466
rect 19553 5414 19565 5466
rect 19617 5414 19629 5466
rect 19681 5414 26963 5466
rect 27015 5414 27027 5466
rect 27079 5414 27091 5466
rect 27143 5414 27155 5466
rect 27207 5414 27219 5466
rect 27271 5414 30912 5466
rect 552 5392 30912 5414
rect 2961 5355 3019 5361
rect 2961 5321 2973 5355
rect 3007 5352 3019 5355
rect 4062 5352 4068 5364
rect 3007 5324 4068 5352
rect 3007 5321 3019 5324
rect 2961 5315 3019 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 7466 5352 7472 5364
rect 4212 5324 7472 5352
rect 4212 5312 4218 5324
rect 7466 5312 7472 5324
rect 7524 5312 7530 5364
rect 9490 5352 9496 5364
rect 8772 5324 9496 5352
rect 3510 5244 3516 5296
rect 3568 5244 3574 5296
rect 8665 5287 8723 5293
rect 8665 5284 8677 5287
rect 7760 5256 8677 5284
rect 1673 5219 1731 5225
rect 1448 5207 1624 5216
rect 1433 5201 1624 5207
rect 1433 5167 1445 5201
rect 1479 5188 1624 5201
rect 1479 5167 1491 5188
rect 1433 5161 1491 5167
rect 934 5108 940 5160
rect 992 5108 998 5160
rect 1596 5148 1624 5188
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 4062 5216 4068 5228
rect 1719 5188 4068 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 4387 5219 4445 5225
rect 4387 5185 4399 5219
rect 4433 5216 4445 5219
rect 5718 5216 5724 5228
rect 4433 5188 5724 5216
rect 4433 5185 4445 5188
rect 4387 5179 4445 5185
rect 5718 5176 5724 5188
rect 5776 5176 5782 5228
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5216 6055 5219
rect 6552 5219 6610 5225
rect 6552 5216 6564 5219
rect 6043 5188 6564 5216
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 6552 5185 6564 5188
rect 6598 5185 6610 5219
rect 6552 5179 6610 5185
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 7760 5216 7788 5256
rect 8665 5253 8677 5256
rect 8711 5253 8723 5287
rect 8665 5247 8723 5253
rect 8772 5216 8800 5324
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 10686 5312 10692 5364
rect 10744 5352 10750 5364
rect 13265 5355 13323 5361
rect 10744 5324 12664 5352
rect 10744 5312 10750 5324
rect 12636 5284 12664 5324
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13906 5352 13912 5364
rect 13311 5324 13912 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 13906 5312 13912 5324
rect 13964 5312 13970 5364
rect 15749 5355 15807 5361
rect 15749 5321 15761 5355
rect 15795 5352 15807 5355
rect 16574 5352 16580 5364
rect 15795 5324 16580 5352
rect 15795 5321 15807 5324
rect 15749 5315 15807 5321
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17184 5324 20668 5352
rect 17184 5312 17190 5324
rect 13630 5284 13636 5296
rect 12636 5256 13636 5284
rect 13630 5244 13636 5256
rect 13688 5244 13694 5296
rect 20640 5284 20668 5324
rect 20714 5312 20720 5364
rect 20772 5312 20778 5364
rect 20824 5324 25268 5352
rect 20824 5284 20852 5324
rect 20640 5256 20852 5284
rect 23109 5287 23167 5293
rect 23109 5253 23121 5287
rect 23155 5284 23167 5287
rect 23474 5284 23480 5296
rect 23155 5256 23480 5284
rect 23155 5253 23167 5256
rect 23109 5247 23167 5253
rect 23474 5244 23480 5256
rect 23532 5244 23538 5296
rect 25240 5284 25268 5324
rect 25590 5312 25596 5364
rect 25648 5352 25654 5364
rect 25685 5355 25743 5361
rect 25685 5352 25697 5355
rect 25648 5324 25697 5352
rect 25648 5312 25654 5324
rect 25685 5321 25697 5324
rect 25731 5321 25743 5355
rect 29457 5355 29515 5361
rect 29457 5352 29469 5355
rect 25685 5315 25743 5321
rect 25792 5324 29469 5352
rect 25792 5284 25820 5324
rect 29457 5321 29469 5324
rect 29503 5321 29515 5355
rect 29457 5315 29515 5321
rect 25240 5256 25820 5284
rect 25958 5244 25964 5296
rect 26016 5244 26022 5296
rect 26602 5244 26608 5296
rect 26660 5284 26666 5296
rect 26660 5256 26740 5284
rect 26660 5244 26666 5256
rect 9496 5219 9554 5225
rect 9496 5216 9508 5219
rect 6871 5188 7788 5216
rect 8588 5188 8800 5216
rect 9419 5214 9508 5216
rect 9283 5188 9508 5214
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 1596 5120 3832 5148
rect 2958 5040 2964 5092
rect 3016 5080 3022 5092
rect 3234 5080 3240 5092
rect 3016 5052 3240 5080
rect 3016 5040 3022 5052
rect 3234 5040 3240 5052
rect 3292 5080 3298 5092
rect 3329 5083 3387 5089
rect 3329 5080 3341 5083
rect 3292 5052 3341 5080
rect 3292 5040 3298 5052
rect 3329 5049 3341 5052
rect 3375 5049 3387 5083
rect 3329 5043 3387 5049
rect 1394 4972 1400 5024
rect 1452 5021 1458 5024
rect 1452 5012 1461 5021
rect 1452 4984 1497 5012
rect 1452 4975 1461 4984
rect 1452 4972 1458 4975
rect 2038 4972 2044 5024
rect 2096 5012 2102 5024
rect 2314 5012 2320 5024
rect 2096 4984 2320 5012
rect 2096 4972 2102 4984
rect 2314 4972 2320 4984
rect 2372 4972 2378 5024
rect 3804 5012 3832 5120
rect 3878 5108 3884 5160
rect 3936 5108 3942 5160
rect 4154 5108 4160 5160
rect 4212 5157 4218 5160
rect 4212 5151 4266 5157
rect 4212 5117 4220 5151
rect 4254 5117 4266 5151
rect 4212 5111 4266 5117
rect 4617 5151 4675 5157
rect 4617 5117 4629 5151
rect 4663 5148 4675 5151
rect 5442 5148 5448 5160
rect 4663 5120 5448 5148
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 4212 5108 4218 5111
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 5902 5108 5908 5160
rect 5960 5108 5966 5160
rect 6089 5151 6147 5157
rect 6089 5117 6101 5151
rect 6135 5117 6147 5151
rect 6089 5111 6147 5117
rect 6416 5151 6474 5157
rect 6416 5117 6428 5151
rect 6462 5148 6474 5151
rect 8478 5148 8484 5160
rect 6462 5120 8484 5148
rect 6462 5117 6474 5120
rect 6416 5111 6474 5117
rect 5920 5012 5948 5108
rect 3804 4984 5948 5012
rect 6104 5012 6132 5111
rect 8478 5108 8484 5120
rect 8536 5108 8542 5160
rect 8588 5157 8616 5188
rect 9283 5186 9447 5188
rect 8573 5151 8631 5157
rect 8573 5117 8585 5151
rect 8619 5117 8631 5151
rect 8573 5111 8631 5117
rect 8662 5108 8668 5160
rect 8720 5148 8726 5160
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 8720 5120 8861 5148
rect 8720 5108 8726 5120
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 8938 5108 8944 5160
rect 8996 5148 9002 5160
rect 9033 5151 9091 5157
rect 9033 5148 9045 5151
rect 8996 5120 9045 5148
rect 8996 5108 9002 5120
rect 9033 5117 9045 5120
rect 9079 5117 9091 5151
rect 9283 5148 9311 5186
rect 9496 5185 9508 5188
rect 9542 5185 9554 5219
rect 9496 5179 9554 5185
rect 9674 5176 9680 5228
rect 9732 5216 9738 5228
rect 9769 5219 9827 5225
rect 9769 5216 9781 5219
rect 9732 5188 9781 5216
rect 9732 5176 9738 5188
rect 9769 5185 9781 5188
rect 9815 5185 9827 5219
rect 9769 5179 9827 5185
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 11704 5219 11762 5225
rect 11704 5216 11716 5219
rect 11195 5188 11716 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11704 5185 11716 5188
rect 11750 5185 11762 5219
rect 11704 5179 11762 5185
rect 13354 5176 13360 5228
rect 13412 5216 13418 5228
rect 13412 5188 13852 5216
rect 13412 5176 13418 5188
rect 9033 5111 9091 5117
rect 9146 5120 9311 5148
rect 9360 5151 9418 5157
rect 8205 5083 8263 5089
rect 8205 5049 8217 5083
rect 8251 5080 8263 5083
rect 9146 5080 9174 5120
rect 9360 5117 9372 5151
rect 9406 5148 9418 5151
rect 9582 5148 9588 5160
rect 9406 5120 9588 5148
rect 9406 5117 9418 5120
rect 9360 5111 9418 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 11241 5151 11299 5157
rect 11241 5117 11253 5151
rect 11287 5148 11299 5151
rect 11330 5148 11336 5160
rect 11287 5120 11336 5148
rect 11287 5117 11299 5120
rect 11241 5111 11299 5117
rect 11330 5108 11336 5120
rect 11388 5108 11394 5160
rect 11514 5108 11520 5160
rect 11572 5148 11578 5160
rect 11977 5151 12035 5157
rect 11977 5148 11989 5151
rect 11572 5120 11989 5148
rect 11572 5108 11578 5120
rect 11977 5117 11989 5120
rect 12023 5117 12035 5151
rect 11977 5111 12035 5117
rect 13725 5151 13783 5157
rect 13725 5117 13737 5151
rect 13771 5117 13783 5151
rect 13824 5148 13852 5188
rect 13906 5176 13912 5228
rect 13964 5216 13970 5228
rect 14188 5219 14246 5225
rect 14188 5216 14200 5219
rect 13964 5188 14200 5216
rect 13964 5176 13970 5188
rect 14188 5185 14200 5188
rect 14234 5185 14246 5219
rect 14188 5179 14246 5185
rect 16114 5176 16120 5228
rect 16172 5216 16178 5228
rect 16396 5219 16454 5225
rect 16396 5216 16408 5219
rect 16172 5188 16408 5216
rect 16172 5176 16178 5188
rect 16396 5185 16408 5188
rect 16442 5185 16454 5219
rect 16396 5179 16454 5185
rect 18138 5176 18144 5228
rect 18196 5216 18202 5228
rect 19156 5219 19214 5225
rect 19156 5216 19168 5219
rect 18196 5188 19168 5216
rect 18196 5176 18202 5188
rect 19156 5185 19168 5188
rect 19202 5185 19214 5219
rect 19156 5179 19214 5185
rect 20254 5176 20260 5228
rect 20312 5216 20318 5228
rect 21228 5219 21286 5225
rect 21228 5216 21240 5219
rect 20312 5188 21240 5216
rect 20312 5176 20318 5188
rect 21228 5185 21240 5188
rect 21274 5185 21286 5219
rect 21380 5201 21438 5207
rect 21380 5198 21392 5201
rect 21228 5179 21286 5185
rect 21376 5167 21392 5198
rect 21426 5167 21438 5201
rect 21634 5176 21640 5228
rect 21692 5176 21698 5228
rect 21928 5188 23428 5216
rect 21376 5161 21438 5167
rect 14461 5151 14519 5157
rect 14461 5148 14473 5151
rect 13824 5120 14473 5148
rect 13725 5111 13783 5117
rect 14461 5117 14473 5120
rect 14507 5117 14519 5151
rect 14461 5111 14519 5117
rect 8251 5052 9174 5080
rect 13740 5080 13768 5111
rect 15930 5108 15936 5160
rect 15988 5108 15994 5160
rect 16669 5151 16727 5157
rect 16669 5117 16681 5151
rect 16715 5148 16727 5151
rect 18414 5148 18420 5160
rect 16715 5120 18420 5148
rect 16715 5117 16727 5120
rect 16669 5111 16727 5117
rect 18414 5108 18420 5120
rect 18472 5108 18478 5160
rect 18506 5108 18512 5160
rect 18564 5108 18570 5160
rect 18598 5108 18604 5160
rect 18656 5148 18662 5160
rect 18693 5151 18751 5157
rect 18693 5148 18705 5151
rect 18656 5120 18705 5148
rect 18656 5108 18662 5120
rect 18693 5117 18705 5120
rect 18739 5117 18751 5151
rect 19429 5151 19487 5157
rect 19429 5148 19441 5151
rect 18693 5111 18751 5117
rect 18803 5120 19441 5148
rect 13814 5080 13820 5092
rect 13740 5052 13820 5080
rect 8251 5049 8263 5052
rect 8205 5043 8263 5049
rect 13814 5040 13820 5052
rect 13872 5040 13878 5092
rect 18046 5040 18052 5092
rect 18104 5040 18110 5092
rect 18803 5080 18831 5120
rect 19429 5117 19441 5120
rect 19475 5117 19487 5151
rect 19429 5111 19487 5117
rect 20806 5108 20812 5160
rect 20864 5148 20870 5160
rect 20901 5151 20959 5157
rect 20901 5148 20913 5151
rect 20864 5120 20913 5148
rect 20864 5108 20870 5120
rect 20901 5117 20913 5120
rect 20947 5117 20959 5151
rect 21376 5148 21404 5161
rect 21928 5160 21956 5188
rect 20901 5111 20959 5117
rect 21008 5120 21404 5148
rect 21008 5080 21036 5120
rect 21910 5108 21916 5160
rect 21968 5108 21974 5160
rect 22002 5108 22008 5160
rect 22060 5148 22066 5160
rect 22060 5120 23060 5148
rect 22060 5108 22066 5120
rect 23032 5080 23060 5120
rect 23290 5108 23296 5160
rect 23348 5108 23354 5160
rect 23400 5148 23428 5188
rect 23566 5176 23572 5228
rect 23624 5216 23630 5228
rect 24308 5219 24366 5225
rect 24308 5216 24320 5219
rect 23624 5188 24320 5216
rect 23624 5176 23630 5188
rect 24308 5185 24320 5188
rect 24354 5185 24366 5219
rect 24308 5179 24366 5185
rect 25038 5176 25044 5228
rect 25096 5216 25102 5228
rect 25976 5216 26004 5244
rect 26712 5225 26740 5256
rect 28994 5244 29000 5296
rect 29052 5284 29058 5296
rect 31202 5284 31208 5296
rect 29052 5256 31208 5284
rect 29052 5244 29058 5256
rect 25096 5188 26004 5216
rect 26697 5219 26755 5225
rect 25096 5176 25102 5188
rect 26697 5185 26709 5219
rect 26743 5185 26755 5219
rect 27890 5216 27896 5228
rect 26697 5179 26755 5185
rect 27172 5201 27896 5216
rect 27172 5170 27205 5201
rect 27193 5167 27205 5170
rect 27239 5188 27896 5201
rect 27239 5167 27251 5188
rect 27890 5176 27896 5188
rect 27948 5176 27954 5228
rect 27193 5161 27251 5167
rect 23658 5148 23664 5160
rect 23400 5120 23664 5148
rect 23658 5108 23664 5120
rect 23716 5148 23722 5160
rect 23845 5151 23903 5157
rect 23845 5148 23857 5151
rect 23716 5120 23857 5148
rect 23716 5108 23722 5120
rect 23845 5117 23857 5120
rect 23891 5117 23903 5151
rect 24581 5151 24639 5157
rect 24581 5148 24593 5151
rect 23845 5111 23903 5117
rect 23952 5120 24593 5148
rect 23106 5080 23112 5092
rect 18340 5052 18831 5080
rect 20824 5052 21036 5080
rect 22296 5052 22968 5080
rect 23032 5052 23112 5080
rect 6362 5012 6368 5024
rect 6104 4984 6368 5012
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 8389 5015 8447 5021
rect 8389 5012 8401 5015
rect 6880 4984 8401 5012
rect 6880 4972 6886 4984
rect 8389 4981 8401 4984
rect 8435 4981 8447 5015
rect 8389 4975 8447 4981
rect 9030 4972 9036 5024
rect 9088 5012 9094 5024
rect 11514 5012 11520 5024
rect 9088 4984 11520 5012
rect 9088 4972 9094 4984
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 11698 4972 11704 5024
rect 11756 5021 11762 5024
rect 11756 5012 11765 5021
rect 11756 4984 11801 5012
rect 11756 4975 11765 4984
rect 11756 4972 11762 4975
rect 14182 4972 14188 5024
rect 14240 5021 14246 5024
rect 14240 5012 14249 5021
rect 16399 5015 16457 5021
rect 14240 4984 14285 5012
rect 14240 4975 14249 4984
rect 16399 4981 16411 5015
rect 16445 5012 16457 5015
rect 16666 5012 16672 5024
rect 16445 4984 16672 5012
rect 16445 4981 16457 4984
rect 16399 4975 16457 4981
rect 14240 4972 14246 4975
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 18340 5021 18368 5052
rect 20824 5024 20852 5052
rect 22296 5024 22324 5052
rect 18325 5015 18383 5021
rect 18325 4981 18337 5015
rect 18371 4981 18383 5015
rect 18325 4975 18383 4981
rect 18690 4972 18696 5024
rect 18748 5012 18754 5024
rect 19159 5015 19217 5021
rect 19159 5012 19171 5015
rect 18748 4984 19171 5012
rect 18748 4972 18754 4984
rect 19159 4981 19171 4984
rect 19205 4981 19217 5015
rect 19159 4975 19217 4981
rect 20806 4972 20812 5024
rect 20864 4972 20870 5024
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 21634 5012 21640 5024
rect 20956 4984 21640 5012
rect 20956 4972 20962 4984
rect 21634 4972 21640 4984
rect 21692 4972 21698 5024
rect 22278 4972 22284 5024
rect 22336 4972 22342 5024
rect 22646 4972 22652 5024
rect 22704 5012 22710 5024
rect 22741 5015 22799 5021
rect 22741 5012 22753 5015
rect 22704 4984 22753 5012
rect 22704 4972 22710 4984
rect 22741 4981 22753 4984
rect 22787 4981 22799 5015
rect 22940 5012 22968 5052
rect 23106 5040 23112 5052
rect 23164 5040 23170 5092
rect 23474 5040 23480 5092
rect 23532 5080 23538 5092
rect 23952 5080 23980 5120
rect 24581 5117 24593 5120
rect 24627 5117 24639 5151
rect 24581 5111 24639 5117
rect 25314 5108 25320 5160
rect 25372 5148 25378 5160
rect 25866 5148 25872 5160
rect 25372 5120 25872 5148
rect 25372 5108 25378 5120
rect 25866 5108 25872 5120
rect 25924 5108 25930 5160
rect 27430 5108 27436 5160
rect 27488 5108 27494 5160
rect 29196 5157 29224 5256
rect 31202 5244 31208 5256
rect 31260 5244 31266 5296
rect 29181 5151 29239 5157
rect 29181 5117 29193 5151
rect 29227 5117 29239 5151
rect 29181 5111 29239 5117
rect 29273 5151 29331 5157
rect 29273 5117 29285 5151
rect 29319 5148 29331 5151
rect 29914 5148 29920 5160
rect 29319 5120 29920 5148
rect 29319 5117 29331 5120
rect 29273 5111 29331 5117
rect 23532 5052 23980 5080
rect 23532 5040 23538 5052
rect 29086 5040 29092 5092
rect 29144 5080 29150 5092
rect 29288 5080 29316 5111
rect 29914 5108 29920 5120
rect 29972 5108 29978 5160
rect 29144 5052 29316 5080
rect 29144 5040 29150 5052
rect 24311 5015 24369 5021
rect 24311 5012 24323 5015
rect 22940 4984 24323 5012
rect 22741 4975 22799 4981
rect 24311 4981 24323 4984
rect 24357 4981 24369 5015
rect 24311 4975 24369 4981
rect 27163 5015 27221 5021
rect 27163 4981 27175 5015
rect 27209 5012 27221 5015
rect 27338 5012 27344 5024
rect 27209 4984 27344 5012
rect 27209 4981 27221 4984
rect 27163 4975 27221 4981
rect 27338 4972 27344 4984
rect 27396 4972 27402 5024
rect 27430 4972 27436 5024
rect 27488 5012 27494 5024
rect 28537 5015 28595 5021
rect 28537 5012 28549 5015
rect 27488 4984 28549 5012
rect 27488 4972 27494 4984
rect 28537 4981 28549 4984
rect 28583 4981 28595 5015
rect 28537 4975 28595 4981
rect 28994 4972 29000 5024
rect 29052 4972 29058 5024
rect 552 4922 31072 4944
rect 552 4870 7988 4922
rect 8040 4870 8052 4922
rect 8104 4870 8116 4922
rect 8168 4870 8180 4922
rect 8232 4870 8244 4922
rect 8296 4870 15578 4922
rect 15630 4870 15642 4922
rect 15694 4870 15706 4922
rect 15758 4870 15770 4922
rect 15822 4870 15834 4922
rect 15886 4870 23168 4922
rect 23220 4870 23232 4922
rect 23284 4870 23296 4922
rect 23348 4870 23360 4922
rect 23412 4870 23424 4922
rect 23476 4870 30758 4922
rect 30810 4870 30822 4922
rect 30874 4870 30886 4922
rect 30938 4870 30950 4922
rect 31002 4870 31014 4922
rect 31066 4870 31072 4922
rect 552 4848 31072 4870
rect 845 4811 903 4817
rect 845 4777 857 4811
rect 891 4808 903 4811
rect 1854 4808 1860 4820
rect 891 4780 1860 4808
rect 891 4777 903 4780
rect 845 4771 903 4777
rect 1854 4768 1860 4780
rect 1912 4768 1918 4820
rect 3142 4768 3148 4820
rect 3200 4768 3206 4820
rect 3979 4811 4037 4817
rect 3979 4777 3991 4811
rect 4025 4808 4037 4811
rect 4522 4808 4528 4820
rect 4025 4780 4528 4808
rect 4025 4777 4037 4780
rect 3979 4771 4037 4777
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 7650 4768 7656 4820
rect 7708 4768 7714 4820
rect 7929 4811 7987 4817
rect 7929 4777 7941 4811
rect 7975 4808 7987 4811
rect 8386 4808 8392 4820
rect 7975 4780 8392 4808
rect 7975 4777 7987 4780
rect 7929 4771 7987 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 9131 4811 9189 4817
rect 9131 4777 9143 4811
rect 9177 4808 9189 4811
rect 9490 4808 9496 4820
rect 9177 4780 9496 4808
rect 9177 4777 9189 4780
rect 9131 4771 9189 4777
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 10689 4811 10747 4817
rect 10689 4777 10701 4811
rect 10735 4808 10747 4811
rect 11238 4808 11244 4820
rect 10735 4780 11244 4808
rect 10735 4777 10747 4780
rect 10689 4771 10747 4777
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 11422 4768 11428 4820
rect 11480 4768 11486 4820
rect 11698 4768 11704 4820
rect 11756 4808 11762 4820
rect 12075 4811 12133 4817
rect 12075 4808 12087 4811
rect 11756 4780 12087 4808
rect 11756 4768 11762 4780
rect 12075 4777 12087 4780
rect 12121 4777 12133 4811
rect 12075 4771 12133 4777
rect 14182 4768 14188 4820
rect 14240 4808 14246 4820
rect 14283 4811 14341 4817
rect 14283 4808 14295 4811
rect 14240 4780 14295 4808
rect 14240 4768 14246 4780
rect 14283 4777 14295 4780
rect 14329 4777 14341 4811
rect 14283 4771 14341 4777
rect 18046 4768 18052 4820
rect 18104 4768 18110 4820
rect 18141 4811 18199 4817
rect 18141 4777 18153 4811
rect 18187 4808 18199 4811
rect 18782 4808 18788 4820
rect 18187 4780 18788 4808
rect 18187 4777 18199 4780
rect 18141 4771 18199 4777
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 20349 4811 20407 4817
rect 20349 4777 20361 4811
rect 20395 4808 20407 4811
rect 20806 4808 20812 4820
rect 20395 4780 20812 4808
rect 20395 4777 20407 4780
rect 20349 4771 20407 4777
rect 20806 4768 20812 4780
rect 20864 4768 20870 4820
rect 20898 4768 20904 4820
rect 20956 4768 20962 4820
rect 21726 4768 21732 4820
rect 21784 4768 21790 4820
rect 22094 4768 22100 4820
rect 22152 4768 22158 4820
rect 22278 4768 22284 4820
rect 22336 4808 22342 4820
rect 22471 4811 22529 4817
rect 22471 4808 22483 4811
rect 22336 4780 22483 4808
rect 22336 4768 22342 4780
rect 22471 4777 22483 4780
rect 22517 4777 22529 4811
rect 22471 4771 22529 4777
rect 24213 4811 24271 4817
rect 24213 4777 24225 4811
rect 24259 4808 24271 4811
rect 24670 4808 24676 4820
rect 24259 4780 24676 4808
rect 24259 4777 24271 4780
rect 24213 4771 24271 4777
rect 24670 4768 24676 4780
rect 24728 4768 24734 4820
rect 24762 4768 24768 4820
rect 24820 4768 24826 4820
rect 26050 4808 26056 4820
rect 24964 4780 26056 4808
rect 1029 4675 1087 4681
rect 1029 4672 1041 4675
rect 860 4644 1041 4672
rect 860 4468 888 4644
rect 1029 4641 1041 4644
rect 1075 4641 1087 4675
rect 1029 4635 1087 4641
rect 1394 4632 1400 4684
rect 1452 4681 1458 4684
rect 1452 4675 1506 4681
rect 1452 4641 1460 4675
rect 1494 4641 1506 4675
rect 1452 4635 1506 4641
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 1903 4644 3464 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 1452 4632 1458 4635
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1121 4607 1179 4613
rect 1121 4604 1133 4607
rect 992 4576 1133 4604
rect 992 4564 998 4576
rect 1121 4573 1133 4576
rect 1167 4573 1179 4607
rect 1121 4567 1179 4573
rect 1627 4607 1685 4613
rect 1627 4573 1639 4607
rect 1673 4604 1685 4607
rect 1964 4604 2268 4606
rect 2774 4604 2780 4616
rect 1673 4578 2780 4604
rect 1673 4576 1992 4578
rect 2240 4576 2780 4578
rect 1673 4573 1685 4576
rect 1627 4567 1685 4573
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 3234 4468 3240 4480
rect 860 4440 3240 4468
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 3436 4468 3464 4644
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 5994 4672 6000 4684
rect 4212 4644 6000 4672
rect 4212 4632 4218 4644
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 6178 4632 6184 4684
rect 6236 4681 6242 4684
rect 6236 4675 6290 4681
rect 6236 4641 6244 4675
rect 6278 4641 6290 4675
rect 6236 4635 6290 4641
rect 6236 4632 6242 4635
rect 6546 4632 6552 4684
rect 6604 4672 6610 4684
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 6604 4644 6653 4672
rect 6604 4632 6610 4644
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 6641 4635 6699 4641
rect 6914 4632 6920 4684
rect 6972 4632 6978 4684
rect 7668 4672 7696 4768
rect 8297 4675 8355 4681
rect 8297 4672 8309 4675
rect 7668 4644 8309 4672
rect 8297 4641 8309 4644
rect 8343 4641 8355 4675
rect 8297 4635 8355 4641
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4672 8631 4675
rect 9030 4672 9036 4684
rect 8619 4644 9036 4672
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4604 3571 4607
rect 3786 4604 3792 4616
rect 3559 4576 3792 4604
rect 3559 4573 3571 4576
rect 3513 4567 3571 4573
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 3970 4564 3976 4616
rect 4028 4604 4034 4616
rect 4249 4607 4307 4613
rect 4028 4576 4073 4604
rect 4028 4564 4034 4576
rect 4249 4573 4261 4607
rect 4295 4604 4307 4607
rect 5810 4604 5816 4616
rect 4295 4576 5816 4604
rect 4295 4573 4307 4576
rect 4249 4567 4307 4573
rect 5810 4564 5816 4576
rect 5868 4564 5874 4616
rect 5902 4564 5908 4616
rect 5960 4564 5966 4616
rect 6411 4607 6469 4613
rect 6411 4573 6423 4607
rect 6457 4604 6469 4607
rect 6932 4604 6960 4632
rect 6457 4576 6960 4604
rect 6457 4573 6469 4576
rect 6411 4567 6469 4573
rect 7742 4564 7748 4616
rect 7800 4604 7806 4616
rect 7800 4576 8156 4604
rect 7800 4564 7806 4576
rect 8128 4545 8156 4576
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 8588 4604 8616 4635
rect 9030 4632 9036 4644
rect 9088 4632 9094 4684
rect 9674 4672 9680 4684
rect 9324 4644 9680 4672
rect 8260 4576 8616 4604
rect 8665 4607 8723 4613
rect 8260 4564 8266 4576
rect 8665 4573 8677 4607
rect 8711 4604 8723 4607
rect 8938 4604 8944 4616
rect 8711 4576 8944 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 8938 4564 8944 4576
rect 8996 4564 9002 4616
rect 9171 4607 9229 4613
rect 9171 4573 9183 4607
rect 9217 4604 9229 4607
rect 9324 4604 9352 4644
rect 9674 4632 9680 4644
rect 9732 4632 9738 4684
rect 11149 4675 11207 4681
rect 11149 4641 11161 4675
rect 11195 4672 11207 4675
rect 11440 4672 11468 4768
rect 15933 4743 15991 4749
rect 15933 4709 15945 4743
rect 15979 4740 15991 4743
rect 16114 4740 16120 4752
rect 15979 4712 16120 4740
rect 15979 4709 15991 4712
rect 15933 4703 15991 4709
rect 16114 4700 16120 4712
rect 16172 4700 16178 4752
rect 11195 4644 11468 4672
rect 11195 4641 11207 4644
rect 11149 4635 11207 4641
rect 9217 4576 9352 4604
rect 9401 4607 9459 4613
rect 9217 4573 9229 4576
rect 9171 4567 9229 4573
rect 9401 4573 9413 4607
rect 9447 4604 9459 4607
rect 9447 4576 11008 4604
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 10980 4545 11008 4576
rect 8113 4539 8171 4545
rect 5460 4508 5948 4536
rect 5460 4468 5488 4508
rect 3436 4440 5488 4468
rect 5534 4428 5540 4480
rect 5592 4428 5598 4480
rect 5920 4468 5948 4508
rect 8113 4505 8125 4539
rect 8159 4505 8171 4539
rect 10965 4539 11023 4545
rect 8113 4499 8171 4505
rect 8312 4508 8708 4536
rect 6822 4468 6828 4480
rect 5920 4440 6828 4468
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 7098 4428 7104 4480
rect 7156 4468 7162 4480
rect 8312 4468 8340 4508
rect 7156 4440 8340 4468
rect 7156 4428 7162 4440
rect 8386 4428 8392 4480
rect 8444 4428 8450 4480
rect 8680 4468 8708 4508
rect 10965 4505 10977 4539
rect 11011 4505 11023 4539
rect 10965 4499 11023 4505
rect 11164 4468 11192 4635
rect 11514 4632 11520 4684
rect 11572 4632 11578 4684
rect 12250 4632 12256 4684
rect 12308 4672 12314 4684
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 12308 4644 12357 4672
rect 12308 4632 12314 4644
rect 12345 4641 12357 4644
rect 12391 4641 12403 4675
rect 12345 4635 12403 4641
rect 12434 4632 12440 4684
rect 12492 4632 12498 4684
rect 13725 4675 13783 4681
rect 13725 4641 13737 4675
rect 13771 4672 13783 4675
rect 13771 4644 14323 4672
rect 13771 4641 13783 4644
rect 13725 4635 13783 4641
rect 11330 4564 11336 4616
rect 11388 4604 11394 4616
rect 11606 4604 11612 4616
rect 11388 4576 11612 4604
rect 11388 4564 11394 4576
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 12158 4613 12164 4616
rect 12115 4607 12164 4613
rect 12115 4573 12127 4607
rect 12161 4573 12164 4607
rect 12115 4567 12164 4573
rect 12158 4564 12164 4567
rect 12216 4564 12222 4616
rect 12452 4604 12480 4632
rect 12452 4576 13768 4604
rect 11514 4496 11520 4548
rect 11572 4496 11578 4548
rect 8680 4440 11192 4468
rect 11330 4428 11336 4480
rect 11388 4428 11394 4480
rect 11532 4468 11560 4496
rect 12802 4468 12808 4480
rect 11532 4440 12808 4468
rect 12802 4428 12808 4440
rect 12860 4428 12866 4480
rect 13740 4468 13768 4576
rect 13814 4564 13820 4616
rect 13872 4564 13878 4616
rect 14295 4615 14323 4644
rect 16758 4632 16764 4684
rect 16816 4632 16822 4684
rect 18064 4672 18092 4768
rect 18064 4644 18828 4672
rect 14280 4609 14338 4615
rect 14280 4575 14292 4609
rect 14326 4575 14338 4609
rect 14280 4569 14338 4575
rect 14366 4564 14372 4616
rect 14424 4604 14430 4616
rect 14553 4607 14611 4613
rect 14553 4604 14565 4607
rect 14424 4576 14565 4604
rect 14424 4564 14430 4576
rect 14553 4573 14565 4576
rect 14599 4573 14611 4607
rect 14553 4567 14611 4573
rect 16114 4564 16120 4616
rect 16172 4564 16178 4616
rect 16482 4613 16488 4616
rect 16444 4607 16488 4613
rect 16444 4573 16456 4607
rect 16444 4567 16488 4573
rect 16482 4564 16488 4567
rect 16540 4564 16546 4616
rect 16623 4607 16681 4613
rect 16623 4573 16635 4607
rect 16669 4604 16681 4607
rect 16776 4604 16804 4632
rect 18800 4631 18828 4644
rect 19058 4632 19064 4684
rect 19116 4632 19122 4684
rect 20438 4632 20444 4684
rect 20496 4672 20502 4684
rect 20717 4675 20775 4681
rect 20717 4672 20729 4675
rect 20496 4644 20729 4672
rect 20496 4632 20502 4644
rect 20717 4641 20729 4644
rect 20763 4672 20775 4675
rect 20916 4672 20944 4768
rect 21744 4740 21772 4768
rect 21008 4712 21772 4740
rect 21008 4684 21036 4712
rect 20763 4644 20944 4672
rect 20763 4641 20775 4644
rect 20717 4635 20775 4641
rect 20990 4632 20996 4684
rect 21048 4632 21054 4684
rect 21453 4675 21511 4681
rect 21453 4641 21465 4675
rect 21499 4672 21511 4675
rect 21634 4672 21640 4684
rect 21499 4644 21640 4672
rect 21499 4641 21511 4644
rect 21453 4635 21511 4641
rect 21634 4632 21640 4644
rect 21692 4632 21698 4684
rect 21744 4681 21772 4712
rect 21729 4675 21787 4681
rect 21729 4641 21741 4675
rect 21775 4641 21787 4675
rect 21729 4635 21787 4641
rect 21910 4632 21916 4684
rect 21968 4672 21974 4684
rect 22005 4675 22063 4681
rect 22005 4672 22017 4675
rect 21968 4644 22017 4672
rect 21968 4632 21974 4644
rect 22005 4641 22017 4644
rect 22051 4641 22063 4675
rect 22112 4672 22140 4768
rect 24964 4740 24992 4780
rect 26050 4768 26056 4780
rect 26108 4768 26114 4820
rect 26605 4811 26663 4817
rect 26605 4808 26617 4811
rect 26160 4780 26617 4808
rect 24688 4712 24992 4740
rect 24688 4681 24716 4712
rect 25038 4700 25044 4752
rect 25096 4700 25102 4752
rect 25590 4700 25596 4752
rect 25648 4740 25654 4752
rect 26160 4740 26188 4780
rect 26605 4777 26617 4780
rect 26651 4777 26663 4811
rect 26605 4771 26663 4777
rect 27246 4768 27252 4820
rect 27304 4768 27310 4820
rect 27338 4768 27344 4820
rect 27396 4808 27402 4820
rect 28258 4808 28264 4820
rect 28316 4817 28322 4820
rect 27396 4780 28264 4808
rect 27396 4768 27402 4780
rect 28258 4768 28264 4780
rect 28316 4771 28325 4817
rect 28316 4768 28322 4771
rect 25648 4712 26188 4740
rect 26252 4712 27108 4740
rect 25648 4700 25654 4712
rect 22296 4672 22508 4676
rect 24397 4675 24455 4681
rect 22112 4648 22784 4672
rect 22112 4644 22324 4648
rect 22480 4644 22784 4648
rect 22005 4635 22063 4641
rect 18800 4625 18862 4631
rect 16669 4576 16804 4604
rect 16853 4607 16911 4613
rect 16669 4573 16681 4576
rect 16623 4567 16681 4573
rect 16853 4573 16865 4607
rect 16899 4604 16911 4607
rect 18325 4607 18383 4613
rect 16899 4576 17908 4604
rect 16899 4573 16911 4576
rect 16853 4567 16911 4573
rect 14366 4468 14372 4480
rect 13740 4440 14372 4468
rect 14366 4428 14372 4440
rect 14424 4428 14430 4480
rect 17880 4468 17908 4576
rect 18325 4573 18337 4607
rect 18371 4604 18383 4607
rect 18506 4604 18512 4616
rect 18371 4576 18512 4604
rect 18371 4573 18383 4576
rect 18325 4567 18383 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 18690 4613 18696 4616
rect 18652 4607 18696 4613
rect 18652 4573 18664 4607
rect 18652 4567 18696 4573
rect 18690 4564 18696 4567
rect 18748 4564 18754 4616
rect 18800 4594 18816 4625
rect 18804 4591 18816 4594
rect 18850 4591 18862 4625
rect 18804 4585 18862 4591
rect 19150 4564 19156 4616
rect 19208 4604 19214 4616
rect 22370 4604 22376 4616
rect 19208 4576 22376 4604
rect 19208 4564 19214 4576
rect 22370 4564 22376 4576
rect 22428 4564 22434 4616
rect 22511 4607 22569 4613
rect 22511 4573 22523 4607
rect 22557 4604 22569 4607
rect 22646 4604 22652 4616
rect 22557 4576 22652 4604
rect 22557 4573 22569 4576
rect 22511 4567 22569 4573
rect 22646 4564 22652 4576
rect 22704 4564 22710 4616
rect 22756 4613 22784 4644
rect 24397 4641 24409 4675
rect 24443 4641 24455 4675
rect 24397 4635 24455 4641
rect 24673 4675 24731 4681
rect 24673 4641 24685 4675
rect 24719 4641 24731 4675
rect 24673 4635 24731 4641
rect 24949 4675 25007 4681
rect 24949 4641 24961 4675
rect 24995 4672 25007 4675
rect 25056 4672 25084 4700
rect 24995 4644 25084 4672
rect 24995 4641 25007 4644
rect 24949 4635 25007 4641
rect 22741 4607 22799 4613
rect 22741 4573 22753 4607
rect 22787 4573 22799 4607
rect 24412 4604 24440 4635
rect 25130 4632 25136 4684
rect 25188 4672 25194 4684
rect 25225 4675 25283 4681
rect 25225 4672 25237 4675
rect 25188 4644 25237 4672
rect 25188 4632 25194 4644
rect 25225 4641 25237 4644
rect 25271 4641 25283 4675
rect 25225 4635 25283 4641
rect 25501 4675 25559 4681
rect 25501 4641 25513 4675
rect 25547 4672 25559 4675
rect 26252 4672 26280 4712
rect 25547 4644 26280 4672
rect 26421 4675 26479 4681
rect 25547 4641 25559 4644
rect 25501 4635 25559 4641
rect 26421 4641 26433 4675
rect 26467 4672 26479 4675
rect 26602 4672 26608 4684
rect 26467 4644 26608 4672
rect 26467 4641 26479 4644
rect 26421 4635 26479 4641
rect 26602 4632 26608 4644
rect 26660 4632 26666 4684
rect 27080 4681 27108 4712
rect 27430 4700 27436 4752
rect 27488 4700 27494 4752
rect 27706 4700 27712 4752
rect 27764 4740 27770 4752
rect 27764 4712 27936 4740
rect 27764 4700 27770 4712
rect 27065 4675 27123 4681
rect 27065 4641 27077 4675
rect 27111 4672 27123 4675
rect 27338 4672 27344 4684
rect 27111 4644 27344 4672
rect 27111 4641 27123 4644
rect 27065 4635 27123 4641
rect 27338 4632 27344 4644
rect 27396 4632 27402 4684
rect 25314 4604 25320 4616
rect 24412 4576 25320 4604
rect 22741 4567 22799 4573
rect 25314 4564 25320 4576
rect 25372 4564 25378 4616
rect 25406 4564 25412 4616
rect 25464 4604 25470 4616
rect 27448 4604 27476 4700
rect 27522 4632 27528 4684
rect 27580 4672 27586 4684
rect 27801 4675 27859 4681
rect 27801 4672 27813 4675
rect 27580 4644 27813 4672
rect 27580 4632 27586 4644
rect 27801 4641 27813 4644
rect 27847 4641 27859 4675
rect 27801 4635 27859 4641
rect 25464 4576 27476 4604
rect 27908 4604 27936 4712
rect 28537 4675 28595 4681
rect 28537 4641 28549 4675
rect 28583 4672 28595 4675
rect 28902 4672 28908 4684
rect 28583 4644 28908 4672
rect 28583 4641 28595 4644
rect 28537 4635 28595 4641
rect 28902 4632 28908 4644
rect 28960 4632 28966 4684
rect 28264 4607 28322 4613
rect 28264 4604 28276 4607
rect 27908 4576 28276 4604
rect 25464 4564 25470 4576
rect 28264 4573 28276 4576
rect 28310 4573 28322 4607
rect 28264 4567 28322 4573
rect 20533 4539 20591 4545
rect 20533 4536 20545 4539
rect 19720 4508 20545 4536
rect 18966 4468 18972 4480
rect 17880 4440 18972 4468
rect 18966 4428 18972 4440
rect 19024 4428 19030 4480
rect 19058 4428 19064 4480
rect 19116 4468 19122 4480
rect 19720 4468 19748 4508
rect 20533 4505 20545 4508
rect 20579 4505 20591 4539
rect 20533 4499 20591 4505
rect 21269 4539 21327 4545
rect 21269 4505 21281 4539
rect 21315 4536 21327 4539
rect 21818 4536 21824 4548
rect 21315 4508 21824 4536
rect 21315 4505 21327 4508
rect 21269 4499 21327 4505
rect 21818 4496 21824 4508
rect 21876 4496 21882 4548
rect 27246 4536 27252 4548
rect 23955 4508 27252 4536
rect 19116 4440 19748 4468
rect 19116 4428 19122 4440
rect 20070 4428 20076 4480
rect 20128 4468 20134 4480
rect 20809 4471 20867 4477
rect 20809 4468 20821 4471
rect 20128 4440 20821 4468
rect 20128 4428 20134 4440
rect 20809 4437 20821 4440
rect 20855 4437 20867 4471
rect 20809 4431 20867 4437
rect 21542 4428 21548 4480
rect 21600 4428 21606 4480
rect 21634 4428 21640 4480
rect 21692 4468 21698 4480
rect 23955 4468 23983 4508
rect 27246 4496 27252 4508
rect 27304 4496 27310 4548
rect 29641 4539 29699 4545
rect 29641 4505 29653 4539
rect 29687 4505 29699 4539
rect 29641 4499 29699 4505
rect 21692 4440 23983 4468
rect 24029 4471 24087 4477
rect 21692 4428 21698 4440
rect 24029 4437 24041 4471
rect 24075 4468 24087 4471
rect 24302 4468 24308 4480
rect 24075 4440 24308 4468
rect 24075 4437 24087 4440
rect 24029 4431 24087 4437
rect 24302 4428 24308 4440
rect 24360 4428 24366 4480
rect 24489 4471 24547 4477
rect 24489 4437 24501 4471
rect 24535 4468 24547 4471
rect 24670 4468 24676 4480
rect 24535 4440 24676 4468
rect 24535 4437 24547 4440
rect 24489 4431 24547 4437
rect 24670 4428 24676 4440
rect 24728 4428 24734 4480
rect 25038 4428 25044 4480
rect 25096 4428 25102 4480
rect 25314 4428 25320 4480
rect 25372 4428 25378 4480
rect 25498 4428 25504 4480
rect 25556 4468 25562 4480
rect 29656 4468 29684 4499
rect 25556 4440 29684 4468
rect 25556 4428 25562 4440
rect 552 4378 30912 4400
rect 552 4326 4193 4378
rect 4245 4326 4257 4378
rect 4309 4326 4321 4378
rect 4373 4326 4385 4378
rect 4437 4326 4449 4378
rect 4501 4326 11783 4378
rect 11835 4326 11847 4378
rect 11899 4326 11911 4378
rect 11963 4326 11975 4378
rect 12027 4326 12039 4378
rect 12091 4326 19373 4378
rect 19425 4326 19437 4378
rect 19489 4326 19501 4378
rect 19553 4326 19565 4378
rect 19617 4326 19629 4378
rect 19681 4326 26963 4378
rect 27015 4326 27027 4378
rect 27079 4326 27091 4378
rect 27143 4326 27155 4378
rect 27207 4326 27219 4378
rect 27271 4326 30912 4378
rect 552 4304 30912 4326
rect 2746 4236 5120 4264
rect 2406 4156 2412 4208
rect 2464 4196 2470 4208
rect 2746 4196 2774 4236
rect 2464 4168 2774 4196
rect 5092 4196 5120 4236
rect 5718 4224 5724 4276
rect 5776 4224 5782 4276
rect 8386 4264 8392 4276
rect 5828 4236 8392 4264
rect 5828 4196 5856 4236
rect 8386 4224 8392 4236
rect 8444 4224 8450 4276
rect 11885 4267 11943 4273
rect 9646 4236 11284 4264
rect 5092 4168 5856 4196
rect 2464 4156 2470 4168
rect 7650 4156 7656 4208
rect 7708 4196 7714 4208
rect 8570 4196 8576 4208
rect 7708 4168 8576 4196
rect 7708 4156 7714 4168
rect 8570 4156 8576 4168
rect 8628 4156 8634 4208
rect 9646 4196 9674 4236
rect 9858 4196 9864 4208
rect 8680 4168 9674 4196
rect 9728 4168 9864 4196
rect 3050 4128 3056 4140
rect 1448 4119 3056 4128
rect 1433 4113 3056 4119
rect 1433 4079 1445 4113
rect 1479 4100 3056 4113
rect 1479 4079 1491 4100
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 4203 4131 4261 4137
rect 3252 4100 4067 4128
rect 1433 4073 1491 4079
rect 934 4020 940 4072
rect 992 4020 998 4072
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4060 1731 4063
rect 1946 4060 1952 4072
rect 1719 4032 1952 4060
rect 1719 4029 1731 4032
rect 1673 4023 1731 4029
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 2498 4020 2504 4072
rect 2556 4060 2562 4072
rect 3252 4060 3280 4100
rect 2556 4032 3280 4060
rect 2556 4020 2562 4032
rect 3326 4020 3332 4072
rect 3384 4060 3390 4072
rect 3602 4060 3608 4072
rect 3384 4032 3608 4060
rect 3384 4020 3390 4032
rect 3602 4020 3608 4032
rect 3660 4020 3666 4072
rect 3697 4063 3755 4069
rect 3697 4029 3709 4063
rect 3743 4060 3755 4063
rect 3786 4060 3792 4072
rect 3743 4032 3792 4060
rect 3743 4029 3755 4032
rect 3697 4023 3755 4029
rect 3786 4020 3792 4032
rect 3844 4020 3850 4072
rect 4039 4069 4067 4100
rect 4203 4097 4215 4131
rect 4249 4128 4261 4131
rect 4798 4128 4804 4140
rect 4249 4100 4804 4128
rect 4249 4097 4261 4100
rect 4203 4091 4261 4097
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 5534 4088 5540 4140
rect 5592 4128 5598 4140
rect 6368 4131 6426 4137
rect 6368 4128 6380 4131
rect 5592 4100 6380 4128
rect 5592 4088 5598 4100
rect 6368 4097 6380 4100
rect 6414 4097 6426 4131
rect 6368 4091 6426 4097
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 6730 4128 6736 4140
rect 6687 4100 6736 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 6730 4088 6736 4100
rect 6788 4088 6794 4140
rect 8680 4128 8708 4168
rect 6840 4100 8708 4128
rect 4024 4063 4082 4069
rect 4024 4029 4036 4063
rect 4070 4060 4082 4063
rect 4338 4060 4344 4072
rect 4070 4032 4344 4060
rect 4070 4029 4082 4032
rect 4024 4023 4082 4029
rect 4338 4020 4344 4032
rect 4396 4020 4402 4072
rect 4433 4063 4491 4069
rect 4433 4029 4445 4063
rect 4479 4060 4491 4063
rect 5626 4060 5632 4072
rect 4479 4032 5632 4060
rect 4479 4029 4491 4032
rect 4433 4023 4491 4029
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 5902 4020 5908 4072
rect 5960 4020 5966 4072
rect 5994 4020 6000 4072
rect 6052 4060 6058 4072
rect 6232 4063 6290 4069
rect 6232 4060 6244 4063
rect 6052 4032 6244 4060
rect 6052 4020 6058 4032
rect 6232 4029 6244 4032
rect 6278 4060 6290 4063
rect 6840 4060 6868 4100
rect 9030 4088 9036 4140
rect 9088 4128 9094 4140
rect 9728 4128 9756 4168
rect 9858 4156 9864 4168
rect 9916 4156 9922 4208
rect 11256 4196 11284 4236
rect 11885 4233 11897 4267
rect 11931 4264 11943 4267
rect 12158 4264 12164 4276
rect 11931 4236 12164 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 13265 4267 13323 4273
rect 13265 4233 13277 4267
rect 13311 4264 13323 4267
rect 13814 4264 13820 4276
rect 13311 4236 13820 4264
rect 13311 4233 13323 4236
rect 13265 4227 13323 4233
rect 13814 4224 13820 4236
rect 13872 4224 13878 4276
rect 15102 4264 15108 4276
rect 13924 4236 15108 4264
rect 13924 4196 13952 4236
rect 15102 4224 15108 4236
rect 15160 4224 15166 4276
rect 16209 4267 16267 4273
rect 16209 4233 16221 4267
rect 16255 4264 16267 4267
rect 16298 4264 16304 4276
rect 16255 4236 16304 4264
rect 16255 4233 16267 4236
rect 16209 4227 16267 4233
rect 16298 4224 16304 4236
rect 16356 4224 16362 4276
rect 18138 4224 18144 4276
rect 18196 4264 18202 4276
rect 21634 4264 21640 4276
rect 18196 4236 21640 4264
rect 18196 4224 18202 4236
rect 21634 4224 21640 4236
rect 21692 4224 21698 4276
rect 21726 4224 21732 4276
rect 21784 4224 21790 4276
rect 23106 4224 23112 4276
rect 23164 4264 23170 4276
rect 25130 4264 25136 4276
rect 23164 4236 25136 4264
rect 23164 4224 23170 4236
rect 25130 4224 25136 4236
rect 25188 4224 25194 4276
rect 27338 4224 27344 4276
rect 27396 4264 27402 4276
rect 29086 4264 29092 4276
rect 27396 4236 29092 4264
rect 27396 4224 27402 4236
rect 29086 4224 29092 4236
rect 29144 4224 29150 4276
rect 11256 4168 13952 4196
rect 14182 4156 14188 4208
rect 14240 4156 14246 4208
rect 18230 4156 18236 4208
rect 18288 4156 18294 4208
rect 21744 4196 21772 4224
rect 21744 4168 23428 4196
rect 9088 4100 9260 4128
rect 9088 4088 9094 4100
rect 6278 4032 6868 4060
rect 6278 4029 6290 4032
rect 6232 4023 6290 4029
rect 6914 4020 6920 4072
rect 6972 4060 6978 4072
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 6972 4032 8493 4060
rect 6972 4020 6978 4032
rect 8481 4029 8493 4032
rect 8527 4060 8539 4063
rect 8662 4060 8668 4072
rect 8527 4032 8668 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 9232 4069 9260 4100
rect 9692 4100 9756 4128
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4029 9275 4063
rect 9217 4023 9275 4029
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4060 9551 4063
rect 9692 4060 9720 4100
rect 10042 4088 10048 4140
rect 10100 4088 10106 4140
rect 10134 4088 10140 4140
rect 10192 4128 10198 4140
rect 10324 4131 10382 4137
rect 10324 4128 10336 4131
rect 10192 4100 10336 4128
rect 10192 4088 10198 4100
rect 10324 4097 10336 4100
rect 10370 4097 10382 4131
rect 10324 4091 10382 4097
rect 10502 4088 10508 4140
rect 10560 4128 10566 4140
rect 11514 4128 11520 4140
rect 10560 4100 11520 4128
rect 10560 4088 10566 4100
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 11698 4088 11704 4140
rect 11756 4128 11762 4140
rect 12253 4131 12311 4137
rect 12253 4128 12265 4131
rect 11756 4100 12265 4128
rect 11756 4088 11762 4100
rect 12253 4097 12265 4100
rect 12299 4097 12311 4131
rect 13262 4128 13268 4140
rect 12253 4091 12311 4097
rect 12406 4100 13268 4128
rect 9769 4063 9827 4069
rect 9769 4060 9781 4063
rect 9539 4032 9781 4060
rect 9539 4029 9551 4032
rect 9493 4023 9551 4029
rect 9769 4029 9781 4032
rect 9815 4029 9827 4063
rect 9769 4023 9827 4029
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4029 9919 4063
rect 10060 4060 10088 4088
rect 10597 4063 10655 4069
rect 10597 4060 10609 4063
rect 10060 4032 10609 4060
rect 9861 4023 9919 4029
rect 10597 4029 10609 4032
rect 10643 4029 10655 4063
rect 12069 4063 12127 4069
rect 12069 4060 12081 4063
rect 10597 4023 10655 4029
rect 11348 4032 12081 4060
rect 5258 3952 5264 4004
rect 5316 3992 5322 4004
rect 5442 3992 5448 4004
rect 5316 3964 5448 3992
rect 5316 3952 5322 3964
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 9876 3992 9904 4023
rect 9950 3992 9956 4004
rect 9508 3964 9720 3992
rect 9876 3964 9956 3992
rect 9508 3936 9536 3964
rect 1394 3884 1400 3936
rect 1452 3933 1458 3936
rect 1452 3924 1461 3933
rect 1452 3896 1497 3924
rect 1452 3887 1461 3896
rect 1452 3884 1458 3887
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 2682 3924 2688 3936
rect 1636 3896 2688 3924
rect 1636 3884 1642 3896
rect 2682 3884 2688 3896
rect 2740 3884 2746 3936
rect 2774 3884 2780 3936
rect 2832 3884 2838 3936
rect 3421 3927 3479 3933
rect 3421 3893 3433 3927
rect 3467 3924 3479 3927
rect 6178 3924 6184 3936
rect 3467 3896 6184 3924
rect 3467 3893 3479 3896
rect 3421 3887 3479 3893
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 7742 3884 7748 3936
rect 7800 3884 7806 3936
rect 8570 3884 8576 3936
rect 8628 3884 8634 3936
rect 9030 3884 9036 3936
rect 9088 3884 9094 3936
rect 9306 3884 9312 3936
rect 9364 3884 9370 3936
rect 9490 3884 9496 3936
rect 9548 3884 9554 3936
rect 9582 3884 9588 3936
rect 9640 3884 9646 3936
rect 9692 3924 9720 3964
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 10327 3927 10385 3933
rect 10327 3924 10339 3927
rect 9692 3896 10339 3924
rect 10327 3893 10339 3896
rect 10373 3893 10385 3927
rect 10327 3887 10385 3893
rect 10686 3884 10692 3936
rect 10744 3924 10750 3936
rect 11348 3924 11376 4032
rect 12069 4029 12081 4032
rect 12115 4060 12127 4063
rect 12406 4060 12434 4100
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 13909 4131 13967 4137
rect 13909 4097 13921 4131
rect 13955 4128 13967 4131
rect 14200 4128 14228 4156
rect 16758 4128 16764 4140
rect 13955 4100 14228 4128
rect 14660 4113 16764 4128
rect 13955 4097 13967 4100
rect 13909 4091 13967 4097
rect 14660 4082 14693 4113
rect 14681 4079 14693 4082
rect 14727 4100 16764 4113
rect 14727 4079 14739 4100
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 17129 4131 17187 4137
rect 16904 4119 17080 4128
rect 16889 4113 17080 4119
rect 14681 4073 14739 4079
rect 16889 4079 16901 4113
rect 16935 4100 17080 4113
rect 16935 4079 16947 4100
rect 16889 4073 16947 4079
rect 12115 4032 12434 4060
rect 12115 4029 12127 4032
rect 12069 4023 12127 4029
rect 12802 4020 12808 4072
rect 12860 4020 12866 4072
rect 13630 4020 13636 4072
rect 13688 4020 13694 4072
rect 13998 4020 14004 4072
rect 14056 4060 14062 4072
rect 14185 4063 14243 4069
rect 14185 4060 14197 4063
rect 14056 4032 14197 4060
rect 14056 4020 14062 4032
rect 14185 4029 14197 4032
rect 14231 4060 14243 4063
rect 14550 4060 14556 4072
rect 14231 4032 14556 4060
rect 14231 4029 14243 4032
rect 14185 4023 14243 4029
rect 14550 4020 14556 4032
rect 14608 4020 14614 4072
rect 14918 4020 14924 4072
rect 14976 4020 14982 4072
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 16393 4063 16451 4069
rect 16393 4060 16405 4063
rect 16264 4032 16405 4060
rect 16264 4020 16270 4032
rect 16393 4029 16405 4032
rect 16439 4029 16451 4063
rect 17052 4060 17080 4100
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 18046 4128 18052 4140
rect 17175 4100 18052 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 18690 4088 18696 4140
rect 18748 4128 18754 4140
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 18748 4100 19441 4128
rect 18748 4088 18754 4100
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 19429 4091 19487 4097
rect 20346 4088 20352 4140
rect 20404 4128 20410 4140
rect 20444 4131 20502 4137
rect 20444 4128 20456 4131
rect 20404 4100 20456 4128
rect 20404 4088 20410 4100
rect 20444 4097 20456 4100
rect 20490 4097 20502 4131
rect 20444 4091 20502 4097
rect 20530 4088 20536 4140
rect 20588 4088 20594 4140
rect 20717 4131 20775 4137
rect 20717 4097 20729 4131
rect 20763 4128 20775 4131
rect 21082 4128 21088 4140
rect 20763 4100 21088 4128
rect 20763 4097 20775 4100
rect 20717 4091 20775 4097
rect 21082 4088 21088 4100
rect 21140 4088 21146 4140
rect 17052 4032 18920 4060
rect 16393 4023 16451 4029
rect 12989 3995 13047 4001
rect 12989 3961 13001 3995
rect 13035 3992 13047 3995
rect 14274 3992 14280 4004
rect 13035 3964 14280 3992
rect 13035 3961 13047 3964
rect 12989 3955 13047 3961
rect 14274 3952 14280 3964
rect 14332 3952 14338 4004
rect 18506 3952 18512 4004
rect 18564 3992 18570 4004
rect 18782 3992 18788 4004
rect 18564 3964 18788 3992
rect 18564 3952 18570 3964
rect 18782 3952 18788 3964
rect 18840 3952 18846 4004
rect 18892 3992 18920 4032
rect 19242 4020 19248 4072
rect 19300 4020 19306 4072
rect 19981 4063 20039 4069
rect 19981 4029 19993 4063
rect 20027 4060 20039 4063
rect 20548 4060 20576 4088
rect 20027 4032 20576 4060
rect 20027 4029 20039 4032
rect 19981 4023 20039 4029
rect 22370 4020 22376 4072
rect 22428 4020 22434 4072
rect 23106 4020 23112 4072
rect 23164 4020 23170 4072
rect 23400 4069 23428 4168
rect 23842 4088 23848 4140
rect 23900 4128 23906 4140
rect 24029 4131 24087 4137
rect 24029 4128 24041 4131
rect 23900 4100 24041 4128
rect 23900 4088 23906 4100
rect 24029 4097 24041 4100
rect 24075 4097 24087 4131
rect 24029 4091 24087 4097
rect 24302 4088 24308 4140
rect 24360 4128 24366 4140
rect 24492 4131 24550 4137
rect 24492 4128 24504 4131
rect 24360 4100 24504 4128
rect 24360 4088 24366 4100
rect 24492 4097 24504 4100
rect 24538 4097 24550 4131
rect 24492 4091 24550 4097
rect 24670 4088 24676 4140
rect 24728 4128 24734 4140
rect 24765 4131 24823 4137
rect 24765 4128 24777 4131
rect 24728 4100 24777 4128
rect 24728 4088 24734 4100
rect 24765 4097 24777 4100
rect 24811 4097 24823 4131
rect 24765 4091 24823 4097
rect 26142 4088 26148 4140
rect 26200 4128 26206 4140
rect 26700 4131 26758 4137
rect 26700 4128 26712 4131
rect 26200 4100 26712 4128
rect 26200 4088 26206 4100
rect 26700 4097 26712 4100
rect 26746 4097 26758 4131
rect 26700 4091 26758 4097
rect 26786 4088 26792 4140
rect 26844 4128 26850 4140
rect 26973 4131 27031 4137
rect 26973 4128 26985 4131
rect 26844 4100 26985 4128
rect 26844 4088 26850 4100
rect 26973 4097 26985 4100
rect 27019 4097 27031 4131
rect 26973 4091 27031 4097
rect 23385 4063 23443 4069
rect 23385 4029 23397 4063
rect 23431 4029 23443 4063
rect 23385 4023 23443 4029
rect 26234 4020 26240 4072
rect 26292 4060 26298 4072
rect 27338 4060 27344 4072
rect 26292 4032 27344 4060
rect 26292 4020 26298 4032
rect 27338 4020 27344 4032
rect 27396 4020 27402 4072
rect 19702 3992 19708 4004
rect 18892 3964 19708 3992
rect 19702 3952 19708 3964
rect 19760 3952 19766 4004
rect 22094 3952 22100 4004
rect 22152 3952 22158 4004
rect 22278 3952 22284 4004
rect 22336 3992 22342 4004
rect 22646 3992 22652 4004
rect 22336 3964 22652 3992
rect 22336 3952 22342 3964
rect 22646 3952 22652 3964
rect 22704 3952 22710 4004
rect 24118 3992 24124 4004
rect 22940 3964 24124 3992
rect 10744 3896 11376 3924
rect 10744 3884 10750 3896
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 12434 3924 12440 3936
rect 11480 3896 12440 3924
rect 11480 3884 11486 3896
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 12621 3927 12679 3933
rect 12621 3893 12633 3927
rect 12667 3924 12679 3927
rect 14458 3924 14464 3936
rect 12667 3896 14464 3924
rect 12667 3893 12679 3896
rect 12621 3887 12679 3893
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 14651 3927 14709 3933
rect 14651 3893 14663 3927
rect 14697 3924 14709 3927
rect 14826 3924 14832 3936
rect 14697 3896 14832 3924
rect 14697 3893 14709 3896
rect 14651 3887 14709 3893
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 16666 3884 16672 3936
rect 16724 3924 16730 3936
rect 16859 3927 16917 3933
rect 16859 3924 16871 3927
rect 16724 3896 16871 3924
rect 16724 3884 16730 3896
rect 16859 3893 16871 3896
rect 16905 3893 16917 3927
rect 16859 3887 16917 3893
rect 17862 3884 17868 3936
rect 17920 3924 17926 3936
rect 18877 3927 18935 3933
rect 18877 3924 18889 3927
rect 17920 3896 18889 3924
rect 17920 3884 17926 3896
rect 18877 3893 18889 3896
rect 18923 3893 18935 3927
rect 18877 3887 18935 3893
rect 20254 3884 20260 3936
rect 20312 3924 20318 3936
rect 22940 3933 22968 3964
rect 24118 3952 24124 3964
rect 24176 3952 24182 4004
rect 20447 3927 20505 3933
rect 20447 3924 20459 3927
rect 20312 3896 20459 3924
rect 20312 3884 20318 3896
rect 20447 3893 20459 3896
rect 20493 3893 20505 3927
rect 20447 3887 20505 3893
rect 22925 3927 22983 3933
rect 22925 3893 22937 3927
rect 22971 3893 22983 3927
rect 22925 3887 22983 3893
rect 23201 3927 23259 3933
rect 23201 3893 23213 3927
rect 23247 3924 23259 3927
rect 24394 3924 24400 3936
rect 23247 3896 24400 3924
rect 23247 3893 23259 3896
rect 23201 3887 23259 3893
rect 24394 3884 24400 3896
rect 24452 3884 24458 3936
rect 24486 3884 24492 3936
rect 24544 3933 24550 3936
rect 24544 3924 24553 3933
rect 24544 3896 24589 3924
rect 24544 3887 24553 3896
rect 24544 3884 24550 3887
rect 26050 3884 26056 3936
rect 26108 3884 26114 3936
rect 26694 3884 26700 3936
rect 26752 3933 26758 3936
rect 26752 3887 26761 3933
rect 26752 3884 26758 3887
rect 28074 3884 28080 3936
rect 28132 3884 28138 3936
rect 552 3834 31072 3856
rect 552 3782 7988 3834
rect 8040 3782 8052 3834
rect 8104 3782 8116 3834
rect 8168 3782 8180 3834
rect 8232 3782 8244 3834
rect 8296 3782 15578 3834
rect 15630 3782 15642 3834
rect 15694 3782 15706 3834
rect 15758 3782 15770 3834
rect 15822 3782 15834 3834
rect 15886 3782 23168 3834
rect 23220 3782 23232 3834
rect 23284 3782 23296 3834
rect 23348 3782 23360 3834
rect 23412 3782 23424 3834
rect 23476 3782 30758 3834
rect 30810 3782 30822 3834
rect 30874 3782 30886 3834
rect 30938 3782 30950 3834
rect 31002 3782 31014 3834
rect 31066 3782 31072 3834
rect 552 3760 31072 3782
rect 845 3723 903 3729
rect 845 3689 857 3723
rect 891 3720 903 3723
rect 1578 3720 1584 3732
rect 891 3692 1256 3720
rect 891 3689 903 3692
rect 845 3683 903 3689
rect 1029 3587 1087 3593
rect 1029 3553 1041 3587
rect 1075 3553 1087 3587
rect 1029 3547 1087 3553
rect 1044 3380 1072 3547
rect 1228 3516 1256 3692
rect 1320 3692 1584 3720
rect 1320 3593 1348 3692
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 1762 3680 1768 3732
rect 1820 3729 1826 3732
rect 1820 3720 1829 3729
rect 2498 3720 2504 3732
rect 1820 3692 2504 3720
rect 1820 3683 1829 3692
rect 1820 3680 1826 3683
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 2774 3720 2780 3732
rect 2746 3680 2780 3720
rect 2832 3680 2838 3732
rect 3786 3680 3792 3732
rect 3844 3720 3850 3732
rect 3979 3723 4037 3729
rect 3979 3720 3991 3723
rect 3844 3692 3991 3720
rect 3844 3680 3850 3692
rect 3979 3689 3991 3692
rect 4025 3689 4037 3723
rect 3979 3683 4037 3689
rect 4338 3680 4344 3732
rect 4396 3720 4402 3732
rect 5074 3720 5080 3732
rect 4396 3692 5080 3720
rect 4396 3680 4402 3692
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 5810 3680 5816 3732
rect 5868 3680 5874 3732
rect 5902 3680 5908 3732
rect 5960 3720 5966 3732
rect 6270 3720 6276 3732
rect 5960 3692 6276 3720
rect 5960 3680 5966 3692
rect 6270 3680 6276 3692
rect 6328 3720 6334 3732
rect 6641 3723 6699 3729
rect 6641 3720 6653 3723
rect 6328 3692 6653 3720
rect 6328 3680 6334 3692
rect 6641 3689 6653 3692
rect 6687 3720 6699 3723
rect 6914 3720 6920 3732
rect 6687 3692 6920 3720
rect 6687 3689 6699 3692
rect 6641 3683 6699 3689
rect 6914 3680 6920 3692
rect 6972 3680 6978 3732
rect 8303 3723 8361 3729
rect 8303 3720 8315 3723
rect 7576 3692 8315 3720
rect 1305 3587 1363 3593
rect 1305 3553 1317 3587
rect 1351 3553 1363 3587
rect 2746 3584 2774 3680
rect 7576 3664 7604 3692
rect 8303 3689 8315 3692
rect 8349 3720 8361 3723
rect 8478 3720 8484 3732
rect 8349 3692 8484 3720
rect 8349 3689 8361 3692
rect 8303 3683 8361 3689
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 9674 3680 9680 3732
rect 9732 3680 9738 3732
rect 9858 3680 9864 3732
rect 9916 3680 9922 3732
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 11149 3723 11207 3729
rect 11149 3720 11161 3723
rect 10008 3692 11161 3720
rect 10008 3680 10014 3692
rect 11149 3689 11161 3692
rect 11195 3689 11207 3723
rect 11149 3683 11207 3689
rect 11698 3680 11704 3732
rect 11756 3720 11762 3732
rect 12075 3723 12133 3729
rect 12075 3720 12087 3723
rect 11756 3692 12087 3720
rect 11756 3680 11762 3692
rect 12075 3689 12087 3692
rect 12121 3689 12133 3723
rect 12075 3683 12133 3689
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 14090 3720 14096 3732
rect 12492 3692 14096 3720
rect 12492 3680 12498 3692
rect 14090 3680 14096 3692
rect 14148 3680 14154 3732
rect 14182 3680 14188 3732
rect 14240 3720 14246 3732
rect 14283 3723 14341 3729
rect 14283 3720 14295 3723
rect 14240 3692 14295 3720
rect 14240 3680 14246 3692
rect 14283 3689 14295 3692
rect 14329 3689 14341 3723
rect 14283 3683 14341 3689
rect 16574 3680 16580 3732
rect 16632 3729 16638 3732
rect 16632 3720 16641 3729
rect 16632 3692 16677 3720
rect 16632 3683 16641 3692
rect 16632 3680 16638 3683
rect 16758 3680 16764 3732
rect 16816 3720 16822 3732
rect 20162 3720 20168 3732
rect 16816 3692 20168 3720
rect 16816 3680 16822 3692
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 20254 3680 20260 3732
rect 20312 3720 20318 3732
rect 21266 3720 21272 3732
rect 20312 3692 21272 3720
rect 20312 3680 20318 3692
rect 21266 3680 21272 3692
rect 21324 3720 21330 3732
rect 21735 3723 21793 3729
rect 21735 3720 21747 3723
rect 21324 3692 21747 3720
rect 21324 3680 21330 3692
rect 21735 3689 21747 3692
rect 21781 3689 21793 3723
rect 21735 3683 21793 3689
rect 22094 3680 22100 3732
rect 22152 3720 22158 3732
rect 23566 3720 23572 3732
rect 22152 3692 23572 3720
rect 22152 3680 22158 3692
rect 23566 3680 23572 3692
rect 23624 3680 23630 3732
rect 23750 3680 23756 3732
rect 23808 3720 23814 3732
rect 23808 3692 26004 3720
rect 23808 3680 23814 3692
rect 4982 3612 4988 3664
rect 5040 3652 5046 3664
rect 5040 3624 6040 3652
rect 5040 3612 5046 3624
rect 1305 3547 1363 3553
rect 1964 3556 2774 3584
rect 1801 3537 1859 3543
rect 1486 3516 1492 3528
rect 1228 3488 1492 3516
rect 1486 3476 1492 3488
rect 1544 3476 1550 3528
rect 1801 3503 1813 3537
rect 1847 3516 1859 3537
rect 1964 3516 1992 3556
rect 2866 3544 2872 3596
rect 2924 3584 2930 3596
rect 3510 3584 3516 3596
rect 2924 3556 3516 3584
rect 2924 3544 2930 3556
rect 3510 3544 3516 3556
rect 3568 3544 3574 3596
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3584 4307 3587
rect 5350 3584 5356 3596
rect 4295 3556 5356 3584
rect 4295 3553 4307 3556
rect 4249 3547 4307 3553
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 6012 3593 6040 3624
rect 6454 3612 6460 3664
rect 6512 3652 6518 3664
rect 6512 3624 7328 3652
rect 6512 3612 6518 3624
rect 5997 3587 6055 3593
rect 5997 3553 6009 3587
rect 6043 3553 6055 3587
rect 5997 3547 6055 3553
rect 6362 3544 6368 3596
rect 6420 3584 6426 3596
rect 6420 3556 6868 3584
rect 6420 3544 6426 3556
rect 1847 3503 1992 3516
rect 1801 3497 1992 3503
rect 1816 3488 1992 3497
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3516 2099 3519
rect 2406 3516 2412 3528
rect 2087 3488 2412 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 2406 3476 2412 3488
rect 2464 3476 2470 3528
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 3976 3521 4034 3527
rect 3976 3518 3988 3521
rect 3850 3516 3988 3518
rect 3467 3490 3988 3516
rect 3467 3488 3878 3490
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 3976 3487 3988 3490
rect 4022 3487 4034 3521
rect 3976 3481 4034 3487
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3516 5687 3519
rect 6730 3516 6736 3528
rect 5675 3488 6736 3516
rect 5675 3485 5687 3488
rect 5629 3479 5687 3485
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 6840 3516 6868 3556
rect 7098 3544 7104 3596
rect 7156 3584 7162 3596
rect 7300 3593 7328 3624
rect 7558 3612 7564 3664
rect 7616 3612 7622 3664
rect 7742 3612 7748 3664
rect 7800 3612 7806 3664
rect 9876 3652 9904 3680
rect 11422 3652 11428 3664
rect 9876 3624 10824 3652
rect 7193 3587 7251 3593
rect 7193 3584 7205 3587
rect 7156 3556 7205 3584
rect 7156 3544 7162 3556
rect 7193 3553 7205 3556
rect 7239 3553 7251 3587
rect 7193 3547 7251 3553
rect 7285 3587 7343 3593
rect 7285 3553 7297 3587
rect 7331 3553 7343 3587
rect 7760 3584 7788 3612
rect 7760 3556 8064 3584
rect 7285 3547 7343 3553
rect 7834 3516 7840 3528
rect 6840 3488 7840 3516
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 8036 3516 8064 3556
rect 9030 3544 9036 3596
rect 9088 3584 9094 3596
rect 9950 3584 9956 3596
rect 9088 3556 9956 3584
rect 9088 3544 9094 3556
rect 9950 3544 9956 3556
rect 10008 3544 10014 3596
rect 10045 3587 10103 3593
rect 10045 3553 10057 3587
rect 10091 3584 10103 3587
rect 10686 3584 10692 3596
rect 10091 3556 10692 3584
rect 10091 3553 10103 3556
rect 10045 3547 10103 3553
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 10796 3593 10824 3624
rect 10980 3624 11428 3652
rect 10781 3587 10839 3593
rect 10781 3553 10793 3587
rect 10827 3553 10839 3587
rect 10781 3547 10839 3553
rect 8300 3519 8358 3525
rect 8300 3516 8312 3519
rect 8036 3488 8312 3516
rect 8300 3485 8312 3488
rect 8346 3485 8358 3519
rect 8300 3479 8358 3485
rect 8386 3476 8392 3528
rect 8444 3516 8450 3528
rect 8573 3519 8631 3525
rect 8573 3516 8585 3519
rect 8444 3488 8585 3516
rect 8444 3476 8450 3488
rect 8573 3485 8585 3488
rect 8619 3485 8631 3519
rect 8573 3479 8631 3485
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 10229 3519 10287 3525
rect 10229 3516 10241 3519
rect 9548 3488 10241 3516
rect 9548 3476 9554 3488
rect 10229 3485 10241 3488
rect 10275 3485 10287 3519
rect 10980 3516 11008 3624
rect 11422 3612 11428 3624
rect 11480 3612 11486 3664
rect 11057 3587 11115 3593
rect 11057 3553 11069 3587
rect 11103 3553 11115 3587
rect 11057 3547 11115 3553
rect 10229 3479 10287 3485
rect 10520 3488 11008 3516
rect 11072 3516 11100 3547
rect 11330 3544 11336 3596
rect 11388 3584 11394 3596
rect 12345 3587 12403 3593
rect 12345 3584 12357 3587
rect 11388 3556 12357 3584
rect 11388 3544 11394 3556
rect 12345 3553 12357 3556
rect 12391 3553 12403 3587
rect 12345 3547 12403 3553
rect 13725 3587 13783 3593
rect 13725 3553 13737 3587
rect 13771 3584 13783 3587
rect 13771 3556 14323 3584
rect 13771 3553 13783 3556
rect 13725 3547 13783 3553
rect 11606 3516 11612 3528
rect 11072 3488 11612 3516
rect 7190 3448 7196 3460
rect 6380 3420 7196 3448
rect 3694 3380 3700 3392
rect 1044 3352 3700 3380
rect 3694 3340 3700 3352
rect 3752 3340 3758 3392
rect 3786 3340 3792 3392
rect 3844 3380 3850 3392
rect 6380 3380 6408 3420
rect 7190 3408 7196 3420
rect 7248 3408 7254 3460
rect 3844 3352 6408 3380
rect 7009 3383 7067 3389
rect 3844 3340 3850 3352
rect 7009 3349 7021 3383
rect 7055 3380 7067 3383
rect 8386 3380 8392 3392
rect 7055 3352 8392 3380
rect 7055 3349 7067 3352
rect 7009 3343 7067 3349
rect 8386 3340 8392 3352
rect 8444 3340 8450 3392
rect 8478 3340 8484 3392
rect 8536 3380 8542 3392
rect 10520 3380 10548 3488
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 12158 3525 12164 3528
rect 12115 3519 12164 3525
rect 12115 3485 12127 3519
rect 12161 3485 12164 3519
rect 12115 3479 12164 3485
rect 12158 3476 12164 3479
rect 12216 3476 12222 3528
rect 13814 3476 13820 3528
rect 13872 3476 13878 3528
rect 14295 3527 14323 3556
rect 14458 3544 14464 3596
rect 14516 3584 14522 3596
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 14516 3556 14565 3584
rect 14516 3544 14522 3556
rect 14553 3553 14565 3556
rect 14599 3553 14611 3587
rect 14553 3547 14611 3553
rect 15933 3587 15991 3593
rect 15933 3553 15945 3587
rect 15979 3584 15991 3587
rect 18233 3587 18291 3593
rect 15979 3556 16623 3584
rect 15979 3553 15991 3556
rect 15933 3547 15991 3553
rect 14280 3521 14338 3527
rect 14280 3487 14292 3521
rect 14326 3487 14338 3521
rect 14280 3481 14338 3487
rect 14366 3476 14372 3528
rect 14424 3516 14430 3528
rect 16114 3516 16120 3528
rect 14424 3488 16120 3516
rect 14424 3476 14430 3488
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 16595 3527 16623 3556
rect 18233 3553 18245 3587
rect 18279 3584 18291 3587
rect 18279 3556 18831 3584
rect 18279 3553 18291 3556
rect 18233 3547 18291 3553
rect 16580 3521 16638 3527
rect 16580 3487 16592 3521
rect 16626 3487 16638 3521
rect 16580 3481 16638 3487
rect 16850 3476 16856 3528
rect 16908 3476 16914 3528
rect 18690 3525 18696 3528
rect 18325 3519 18383 3525
rect 18325 3485 18337 3519
rect 18371 3485 18383 3519
rect 18325 3479 18383 3485
rect 18652 3519 18696 3525
rect 18652 3485 18664 3519
rect 18652 3479 18696 3485
rect 10612 3420 11560 3448
rect 10612 3389 10640 3420
rect 8536 3352 10548 3380
rect 10597 3383 10655 3389
rect 8536 3340 8542 3352
rect 10597 3349 10609 3383
rect 10643 3349 10655 3383
rect 11532 3380 11560 3420
rect 14274 3380 14280 3392
rect 11532 3352 14280 3380
rect 10597 3343 10655 3349
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 16132 3380 16160 3476
rect 17862 3408 17868 3460
rect 17920 3408 17926 3460
rect 17880 3380 17908 3408
rect 16132 3352 17908 3380
rect 18340 3380 18368 3479
rect 18690 3476 18696 3479
rect 18748 3476 18754 3528
rect 18803 3527 18831 3556
rect 19058 3544 19064 3596
rect 19116 3544 19122 3596
rect 20625 3587 20683 3593
rect 20625 3553 20637 3587
rect 20671 3584 20683 3587
rect 20714 3584 20720 3596
rect 20671 3556 20720 3584
rect 20671 3553 20683 3556
rect 20625 3547 20683 3553
rect 20714 3544 20720 3556
rect 20772 3584 20778 3596
rect 20898 3584 20904 3596
rect 20772 3556 20904 3584
rect 20772 3544 20778 3556
rect 20898 3544 20904 3556
rect 20956 3584 20962 3596
rect 21269 3587 21327 3593
rect 21269 3584 21281 3587
rect 20956 3556 21281 3584
rect 20956 3544 20962 3556
rect 21269 3553 21281 3556
rect 21315 3553 21327 3587
rect 21269 3547 21327 3553
rect 21818 3544 21824 3596
rect 21876 3584 21882 3596
rect 22005 3587 22063 3593
rect 22005 3584 22017 3587
rect 21876 3556 22017 3584
rect 21876 3544 21882 3556
rect 22005 3553 22017 3556
rect 22051 3553 22063 3587
rect 22005 3547 22063 3553
rect 23385 3587 23443 3593
rect 23385 3553 23397 3587
rect 23431 3584 23443 3587
rect 23431 3556 23983 3584
rect 23431 3553 23443 3556
rect 23385 3547 23443 3553
rect 21732 3537 21790 3543
rect 18788 3521 18846 3527
rect 18788 3487 18800 3521
rect 18834 3487 18846 3521
rect 18788 3481 18846 3487
rect 20441 3519 20499 3525
rect 20441 3485 20453 3519
rect 20487 3516 20499 3519
rect 21732 3516 21744 3537
rect 20487 3503 21744 3516
rect 21778 3503 21790 3537
rect 20487 3497 21790 3503
rect 23477 3519 23535 3525
rect 20487 3488 21775 3497
rect 20487 3485 20499 3488
rect 20441 3479 20499 3485
rect 23477 3485 23489 3519
rect 23523 3518 23535 3519
rect 23523 3516 23612 3518
rect 23658 3516 23664 3528
rect 23523 3490 23664 3516
rect 23523 3485 23535 3490
rect 23584 3488 23664 3490
rect 23477 3479 23535 3485
rect 23658 3476 23664 3488
rect 23716 3476 23722 3528
rect 23842 3525 23848 3528
rect 23804 3519 23848 3525
rect 23804 3485 23816 3519
rect 23804 3479 23848 3485
rect 23842 3476 23848 3479
rect 23900 3476 23906 3528
rect 23955 3527 23983 3556
rect 24118 3544 24124 3596
rect 24176 3584 24182 3596
rect 24213 3587 24271 3593
rect 24213 3584 24225 3587
rect 24176 3556 24225 3584
rect 24176 3544 24182 3556
rect 24213 3553 24225 3556
rect 24259 3553 24271 3587
rect 24213 3547 24271 3553
rect 24486 3544 24492 3596
rect 24544 3544 24550 3596
rect 25406 3544 25412 3596
rect 25464 3584 25470 3596
rect 25685 3587 25743 3593
rect 25685 3584 25697 3587
rect 25464 3556 25697 3584
rect 25464 3544 25470 3556
rect 25685 3553 25697 3556
rect 25731 3584 25743 3587
rect 25774 3584 25780 3596
rect 25731 3556 25780 3584
rect 25731 3553 25743 3556
rect 25685 3547 25743 3553
rect 25774 3544 25780 3556
rect 25832 3544 25838 3596
rect 23940 3521 23998 3527
rect 23940 3487 23952 3521
rect 23986 3487 23998 3521
rect 24504 3516 24532 3544
rect 25869 3519 25927 3525
rect 25869 3516 25881 3519
rect 24504 3488 25881 3516
rect 23940 3481 23998 3487
rect 25869 3485 25881 3488
rect 25915 3485 25927 3519
rect 25869 3479 25927 3485
rect 18598 3380 18604 3392
rect 18340 3352 18604 3380
rect 18598 3340 18604 3352
rect 18656 3380 18662 3392
rect 18782 3380 18788 3392
rect 18656 3352 18788 3380
rect 18656 3340 18662 3352
rect 18782 3340 18788 3352
rect 18840 3380 18846 3392
rect 20717 3383 20775 3389
rect 20717 3380 20729 3383
rect 18840 3352 20729 3380
rect 18840 3340 18846 3352
rect 20717 3349 20729 3352
rect 20763 3349 20775 3383
rect 20717 3343 20775 3349
rect 24670 3340 24676 3392
rect 24728 3380 24734 3392
rect 25317 3383 25375 3389
rect 25317 3380 25329 3383
rect 24728 3352 25329 3380
rect 24728 3340 24734 3352
rect 25317 3349 25329 3352
rect 25363 3349 25375 3383
rect 25976 3380 26004 3692
rect 26528 3692 27292 3720
rect 26528 3664 26556 3692
rect 26510 3612 26516 3664
rect 26568 3612 26574 3664
rect 26694 3612 26700 3664
rect 26752 3652 26758 3664
rect 27264 3661 27292 3692
rect 27338 3680 27344 3732
rect 27396 3680 27402 3732
rect 27522 3680 27528 3732
rect 27580 3680 27586 3732
rect 28258 3680 28264 3732
rect 28316 3720 28322 3732
rect 28359 3723 28417 3729
rect 28359 3720 28371 3723
rect 28316 3692 28371 3720
rect 28316 3680 28322 3692
rect 28359 3689 28371 3692
rect 28405 3689 28417 3723
rect 28359 3683 28417 3689
rect 26881 3655 26939 3661
rect 26881 3652 26893 3655
rect 26752 3624 26893 3652
rect 26752 3612 26758 3624
rect 26881 3621 26893 3624
rect 26927 3621 26939 3655
rect 26881 3615 26939 3621
rect 27249 3655 27307 3661
rect 27249 3621 27261 3655
rect 27295 3652 27307 3655
rect 27430 3652 27436 3664
rect 27295 3624 27436 3652
rect 27295 3621 27307 3624
rect 27249 3615 27307 3621
rect 27430 3612 27436 3624
rect 27488 3612 27494 3664
rect 26142 3544 26148 3596
rect 26200 3584 26206 3596
rect 26605 3587 26663 3593
rect 26605 3584 26617 3587
rect 26200 3556 26617 3584
rect 26200 3544 26206 3556
rect 26605 3553 26617 3556
rect 26651 3553 26663 3587
rect 27540 3584 27568 3680
rect 27893 3587 27951 3593
rect 27893 3584 27905 3587
rect 27540 3556 27905 3584
rect 26605 3547 26663 3553
rect 27893 3553 27905 3556
rect 27939 3553 27951 3587
rect 27893 3547 27951 3553
rect 28629 3587 28687 3593
rect 28629 3553 28641 3587
rect 28675 3584 28687 3587
rect 29822 3584 29828 3596
rect 28675 3556 29828 3584
rect 28675 3553 28687 3556
rect 28629 3547 28687 3553
rect 29822 3544 29828 3556
rect 29880 3544 29886 3596
rect 28350 3476 28356 3528
rect 28408 3476 28414 3528
rect 29733 3451 29791 3457
rect 29733 3417 29745 3451
rect 29779 3417 29791 3451
rect 29733 3411 29791 3417
rect 29748 3380 29776 3411
rect 25976 3352 29776 3380
rect 25317 3343 25375 3349
rect 552 3290 30912 3312
rect 552 3238 4193 3290
rect 4245 3238 4257 3290
rect 4309 3238 4321 3290
rect 4373 3238 4385 3290
rect 4437 3238 4449 3290
rect 4501 3238 11783 3290
rect 11835 3238 11847 3290
rect 11899 3238 11911 3290
rect 11963 3238 11975 3290
rect 12027 3238 12039 3290
rect 12091 3238 19373 3290
rect 19425 3238 19437 3290
rect 19489 3238 19501 3290
rect 19553 3238 19565 3290
rect 19617 3238 19629 3290
rect 19681 3238 26963 3290
rect 27015 3238 27027 3290
rect 27079 3238 27091 3290
rect 27143 3238 27155 3290
rect 27207 3238 27219 3290
rect 27271 3238 30912 3290
rect 552 3216 30912 3238
rect 2682 3136 2688 3188
rect 2740 3176 2746 3188
rect 3421 3179 3479 3185
rect 3421 3176 3433 3179
rect 2740 3148 3433 3176
rect 2740 3136 2746 3148
rect 3421 3145 3433 3148
rect 3467 3145 3479 3179
rect 3421 3139 3479 3145
rect 3605 3179 3663 3185
rect 3605 3145 3617 3179
rect 3651 3176 3663 3179
rect 3786 3176 3792 3188
rect 3651 3148 3792 3176
rect 3651 3145 3663 3148
rect 3605 3139 3663 3145
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 5626 3176 5632 3188
rect 3896 3148 5632 3176
rect 2961 3111 3019 3117
rect 2961 3077 2973 3111
rect 3007 3108 3019 3111
rect 3896 3108 3924 3148
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 8478 3176 8484 3188
rect 6104 3148 8484 3176
rect 6104 3108 6132 3148
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 9582 3136 9588 3188
rect 9640 3176 9646 3188
rect 11790 3176 11796 3188
rect 9640 3148 11796 3176
rect 9640 3136 9646 3148
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 16850 3136 16856 3188
rect 16908 3176 16914 3188
rect 18141 3179 18199 3185
rect 18141 3176 18153 3179
rect 16908 3148 18153 3176
rect 16908 3136 16914 3148
rect 18141 3145 18153 3148
rect 18187 3145 18199 3179
rect 19242 3176 19248 3188
rect 18141 3139 18199 3145
rect 18248 3148 19248 3176
rect 3007 3080 3924 3108
rect 5368 3080 6132 3108
rect 3007 3077 3019 3080
rect 2961 3071 3019 3077
rect 1443 3043 1501 3049
rect 1443 3009 1455 3043
rect 1489 3040 1501 3043
rect 3142 3040 3148 3052
rect 1489 3012 3148 3040
rect 1489 3009 1501 3012
rect 1443 3003 1501 3009
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 3234 3000 3240 3052
rect 3292 3040 3298 3052
rect 3292 3012 3832 3040
rect 3292 3000 3298 3012
rect 937 2975 995 2981
rect 937 2941 949 2975
rect 983 2972 995 2975
rect 1578 2972 1584 2984
rect 983 2944 1584 2972
rect 983 2941 995 2944
rect 937 2935 995 2941
rect 1578 2932 1584 2944
rect 1636 2932 1642 2984
rect 3804 2981 3832 3012
rect 3878 3000 3884 3052
rect 3936 3000 3942 3052
rect 4430 3047 4436 3052
rect 4387 3041 4436 3047
rect 4387 3007 4399 3041
rect 4433 3007 4436 3041
rect 4387 3001 4436 3007
rect 4430 3000 4436 3001
rect 4488 3000 4494 3052
rect 4522 3000 4528 3052
rect 4580 3040 4586 3052
rect 4617 3043 4675 3049
rect 4617 3040 4629 3043
rect 4580 3012 4629 3040
rect 4580 3000 4586 3012
rect 4617 3009 4629 3012
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2972 1731 2975
rect 3789 2975 3847 2981
rect 1719 2944 2774 2972
rect 1719 2941 1731 2944
rect 1673 2935 1731 2941
rect 2746 2904 2774 2944
rect 3789 2941 3801 2975
rect 3835 2941 3847 2975
rect 5258 2972 5264 2984
rect 3789 2935 3847 2941
rect 3896 2944 5264 2972
rect 3510 2904 3516 2916
rect 2746 2876 3516 2904
rect 3510 2864 3516 2876
rect 3568 2904 3574 2916
rect 3896 2904 3924 2944
rect 5258 2932 5264 2944
rect 5316 2932 5322 2984
rect 3568 2876 3924 2904
rect 3568 2864 3574 2876
rect 1403 2839 1461 2845
rect 1403 2805 1415 2839
rect 1449 2836 1461 2839
rect 1762 2836 1768 2848
rect 1449 2808 1768 2836
rect 1449 2805 1461 2808
rect 1403 2799 1461 2805
rect 1762 2796 1768 2808
rect 1820 2796 1826 2848
rect 4347 2839 4405 2845
rect 4347 2805 4359 2839
rect 4393 2836 4405 2839
rect 5368 2836 5396 3080
rect 7834 3068 7840 3120
rect 7892 3108 7898 3120
rect 8665 3111 8723 3117
rect 8665 3108 8677 3111
rect 7892 3080 8677 3108
rect 7892 3068 7898 3080
rect 8665 3077 8677 3080
rect 8711 3077 8723 3111
rect 8665 3071 8723 3077
rect 17954 3068 17960 3120
rect 18012 3108 18018 3120
rect 18248 3108 18276 3148
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 20714 3136 20720 3188
rect 20772 3176 20778 3188
rect 20772 3148 22324 3176
rect 20772 3136 20778 3148
rect 18012 3080 18276 3108
rect 18012 3068 18018 3080
rect 6086 3000 6092 3052
rect 6144 3040 6150 3052
rect 6362 3040 6368 3052
rect 6144 3012 6368 3040
rect 6144 3000 6150 3012
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 6638 3047 6644 3052
rect 6595 3041 6644 3047
rect 6595 3007 6607 3041
rect 6641 3007 6644 3041
rect 6595 3001 6644 3007
rect 6638 3000 6644 3001
rect 6696 3000 6702 3052
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3040 8263 3043
rect 9496 3043 9554 3049
rect 9496 3040 9508 3043
rect 8251 3012 9508 3040
rect 8251 3009 8263 3012
rect 8205 3003 8263 3009
rect 9496 3009 9508 3012
rect 9542 3009 9554 3043
rect 9496 3003 9554 3009
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 11704 3043 11762 3049
rect 11704 3040 11716 3043
rect 11195 3012 11716 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 11704 3009 11716 3012
rect 11750 3009 11762 3043
rect 11704 3003 11762 3009
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 11848 3012 11989 3040
rect 11848 3000 11854 3012
rect 11977 3009 11989 3012
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 13357 3043 13415 3049
rect 13357 3009 13369 3043
rect 13403 3040 13415 3043
rect 14188 3043 14246 3049
rect 14188 3040 14200 3043
rect 13403 3012 14200 3040
rect 13403 3009 13415 3012
rect 13357 3003 13415 3009
rect 14188 3009 14200 3012
rect 14234 3009 14246 3043
rect 14188 3003 14246 3009
rect 14274 3000 14280 3052
rect 14332 3040 14338 3052
rect 14461 3043 14519 3049
rect 14461 3040 14473 3043
rect 14332 3012 14473 3040
rect 14332 3000 14338 3012
rect 14461 3009 14473 3012
rect 14507 3009 14519 3043
rect 14461 3003 14519 3009
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3040 15899 3043
rect 16396 3043 16454 3049
rect 16396 3040 16408 3043
rect 15887 3012 16408 3040
rect 15887 3009 15899 3012
rect 15841 3003 15899 3009
rect 16396 3009 16408 3012
rect 16442 3009 16454 3043
rect 16396 3003 16454 3009
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3040 18107 3043
rect 19156 3043 19214 3049
rect 19156 3040 19168 3043
rect 18095 3012 19168 3040
rect 18095 3009 18107 3012
rect 18049 3003 18107 3009
rect 19156 3009 19168 3012
rect 19202 3009 19214 3043
rect 19156 3003 19214 3009
rect 19429 3043 19487 3049
rect 19429 3009 19441 3043
rect 19475 3040 19487 3043
rect 20070 3040 20076 3052
rect 19475 3012 20076 3040
rect 19475 3009 19487 3012
rect 19429 3003 19487 3009
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 21364 3043 21422 3049
rect 21364 3040 21376 3043
rect 20855 3012 21376 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 21364 3009 21376 3012
rect 21410 3009 21422 3043
rect 21364 3003 21422 3009
rect 21542 3000 21548 3052
rect 21600 3040 21606 3052
rect 21637 3043 21695 3049
rect 21637 3040 21649 3043
rect 21600 3012 21649 3040
rect 21600 3000 21606 3012
rect 21637 3009 21649 3012
rect 21683 3009 21695 3043
rect 21637 3003 21695 3009
rect 5442 2932 5448 2984
rect 5500 2972 5506 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 5500 2944 6837 2972
rect 5500 2932 5506 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2972 8539 2975
rect 9030 2972 9036 2984
rect 8527 2944 9036 2972
rect 8527 2941 8539 2944
rect 8481 2935 8539 2941
rect 9030 2932 9036 2944
rect 9088 2932 9094 2984
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 9769 2975 9827 2981
rect 9769 2972 9781 2975
rect 9364 2944 9781 2972
rect 9364 2932 9370 2944
rect 9769 2941 9781 2944
rect 9815 2941 9827 2975
rect 9769 2935 9827 2941
rect 11238 2932 11244 2984
rect 11296 2972 11302 2984
rect 11606 2972 11612 2984
rect 11296 2944 11612 2972
rect 11296 2932 11302 2944
rect 11606 2932 11612 2944
rect 11664 2932 11670 2984
rect 13725 2975 13783 2981
rect 13725 2941 13737 2975
rect 13771 2972 13783 2975
rect 13814 2972 13820 2984
rect 13771 2944 13820 2972
rect 13771 2941 13783 2944
rect 13725 2935 13783 2941
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 15933 2975 15991 2981
rect 15933 2941 15945 2975
rect 15979 2972 15991 2975
rect 16022 2972 16028 2984
rect 15979 2944 16028 2972
rect 15979 2941 15991 2944
rect 15933 2935 15991 2941
rect 16022 2932 16028 2944
rect 16080 2932 16086 2984
rect 16669 2975 16727 2981
rect 16669 2941 16681 2975
rect 16715 2972 16727 2975
rect 17954 2972 17960 2984
rect 16715 2944 17960 2972
rect 16715 2941 16727 2944
rect 16669 2935 16727 2941
rect 17954 2932 17960 2944
rect 18012 2932 18018 2984
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2941 18383 2975
rect 18325 2935 18383 2941
rect 5994 2864 6000 2916
rect 6052 2864 6058 2916
rect 18340 2904 18368 2935
rect 18598 2932 18604 2984
rect 18656 2972 18662 2984
rect 18693 2975 18751 2981
rect 18693 2972 18705 2975
rect 18656 2944 18705 2972
rect 18656 2932 18662 2944
rect 18693 2941 18705 2944
rect 18739 2941 18751 2975
rect 20438 2972 20444 2984
rect 18693 2935 18751 2941
rect 18806 2944 20444 2972
rect 18806 2904 18834 2944
rect 20438 2932 20444 2944
rect 20496 2932 20502 2984
rect 20898 2932 20904 2984
rect 20956 2972 20962 2984
rect 21726 2972 21732 2984
rect 20956 2944 21732 2972
rect 20956 2932 20962 2944
rect 21726 2932 21732 2944
rect 21784 2932 21790 2984
rect 22296 2972 22324 3148
rect 22370 3136 22376 3188
rect 22428 3176 22434 3188
rect 25406 3176 25412 3188
rect 22428 3148 25412 3176
rect 22428 3136 22434 3148
rect 25406 3136 25412 3148
rect 25464 3136 25470 3188
rect 26050 3136 26056 3188
rect 26108 3136 26114 3188
rect 26160 3148 28580 3176
rect 22646 3068 22652 3120
rect 22704 3108 22710 3120
rect 23842 3108 23848 3120
rect 22704 3080 23848 3108
rect 22704 3068 22710 3080
rect 23842 3068 23848 3080
rect 23900 3068 23906 3120
rect 25685 3111 25743 3117
rect 25685 3077 25697 3111
rect 25731 3077 25743 3111
rect 25685 3071 25743 3077
rect 23017 3043 23075 3049
rect 23017 3009 23029 3043
rect 23063 3040 23075 3043
rect 24308 3043 24366 3049
rect 24308 3040 24320 3043
rect 23063 3012 24320 3040
rect 23063 3009 23075 3012
rect 23017 3003 23075 3009
rect 24308 3009 24320 3012
rect 24354 3009 24366 3043
rect 24308 3003 24366 3009
rect 24394 3000 24400 3052
rect 24452 3040 24458 3052
rect 24581 3043 24639 3049
rect 24581 3040 24593 3043
rect 24452 3012 24593 3040
rect 24452 3000 24458 3012
rect 24581 3009 24593 3012
rect 24627 3009 24639 3043
rect 24581 3003 24639 3009
rect 24762 3000 24768 3052
rect 24820 3040 24826 3052
rect 25700 3040 25728 3071
rect 24820 3012 25728 3040
rect 26068 3040 26096 3136
rect 26160 3120 26188 3148
rect 26142 3068 26148 3120
rect 26200 3068 26206 3120
rect 28552 3108 28580 3148
rect 28626 3136 28632 3188
rect 28684 3136 28690 3188
rect 29454 3136 29460 3188
rect 29512 3176 29518 3188
rect 29730 3176 29736 3188
rect 29512 3148 29736 3176
rect 29512 3136 29518 3148
rect 29730 3136 29736 3148
rect 29788 3136 29794 3188
rect 28552 3080 29316 3108
rect 26700 3043 26758 3049
rect 26700 3040 26712 3043
rect 26068 3012 26712 3040
rect 24820 3000 24826 3012
rect 26700 3009 26712 3012
rect 26746 3009 26758 3043
rect 26700 3003 26758 3009
rect 26786 3000 26792 3052
rect 26844 3040 26850 3052
rect 26973 3043 27031 3049
rect 26973 3040 26985 3043
rect 26844 3012 26985 3040
rect 26844 3000 26850 3012
rect 26973 3009 26985 3012
rect 27019 3009 27031 3043
rect 26973 3003 27031 3009
rect 27614 3000 27620 3052
rect 27672 3040 27678 3052
rect 29181 3043 29239 3049
rect 29181 3040 29193 3043
rect 27672 3012 29193 3040
rect 27672 3000 27678 3012
rect 29181 3009 29193 3012
rect 29227 3009 29239 3043
rect 29181 3003 29239 3009
rect 23201 2975 23259 2981
rect 22296 2944 23152 2972
rect 23124 2904 23152 2944
rect 23201 2941 23213 2975
rect 23247 2972 23259 2975
rect 23658 2972 23664 2984
rect 23247 2944 23664 2972
rect 23247 2941 23259 2944
rect 23201 2935 23259 2941
rect 23658 2932 23664 2944
rect 23716 2972 23722 2984
rect 23845 2975 23903 2981
rect 23845 2972 23857 2975
rect 23716 2944 23857 2972
rect 23716 2932 23722 2944
rect 23845 2941 23857 2944
rect 23891 2941 23903 2975
rect 25682 2972 25688 2984
rect 23845 2935 23903 2941
rect 23955 2944 25688 2972
rect 23955 2904 23983 2944
rect 25682 2932 25688 2944
rect 25740 2972 25746 2984
rect 26142 2972 26148 2984
rect 25740 2944 26148 2972
rect 25740 2932 25746 2944
rect 26142 2932 26148 2944
rect 26200 2932 26206 2984
rect 26234 2932 26240 2984
rect 26292 2932 26298 2984
rect 26602 2932 26608 2984
rect 26660 2972 26666 2984
rect 28258 2972 28264 2984
rect 26660 2944 28264 2972
rect 26660 2932 26666 2944
rect 28258 2932 28264 2944
rect 28316 2972 28322 2984
rect 28445 2975 28503 2981
rect 28445 2972 28457 2975
rect 28316 2944 28457 2972
rect 28316 2932 28322 2944
rect 28445 2941 28457 2944
rect 28491 2941 28503 2975
rect 28445 2935 28503 2941
rect 28997 2975 29055 2981
rect 28997 2941 29009 2975
rect 29043 2972 29055 2975
rect 29288 2972 29316 3080
rect 29043 2944 29316 2972
rect 29043 2941 29055 2944
rect 28997 2935 29055 2941
rect 18340 2876 18834 2904
rect 22664 2876 22876 2904
rect 23124 2876 23983 2904
rect 4393 2808 5396 2836
rect 6555 2839 6613 2845
rect 4393 2805 4405 2808
rect 4347 2799 4405 2805
rect 6555 2805 6567 2839
rect 6601 2836 6613 2839
rect 6822 2836 6828 2848
rect 6601 2808 6828 2836
rect 6601 2805 6613 2808
rect 6555 2799 6613 2805
rect 6822 2796 6828 2808
rect 6880 2836 6886 2848
rect 7558 2836 7564 2848
rect 6880 2808 7564 2836
rect 6880 2796 6886 2808
rect 7558 2796 7564 2808
rect 7616 2796 7622 2848
rect 9122 2796 9128 2848
rect 9180 2836 9186 2848
rect 9490 2836 9496 2848
rect 9548 2845 9554 2848
rect 9180 2808 9496 2836
rect 9180 2796 9186 2808
rect 9490 2796 9496 2808
rect 9548 2799 9557 2845
rect 9548 2796 9554 2799
rect 11698 2796 11704 2848
rect 11756 2845 11762 2848
rect 11756 2836 11765 2845
rect 11756 2808 11801 2836
rect 11756 2799 11765 2808
rect 11756 2796 11762 2799
rect 14182 2796 14188 2848
rect 14240 2845 14246 2848
rect 14240 2836 14249 2845
rect 14240 2808 14285 2836
rect 14240 2799 14249 2808
rect 14240 2796 14246 2799
rect 15378 2796 15384 2848
rect 15436 2836 15442 2848
rect 16298 2836 16304 2848
rect 15436 2808 16304 2836
rect 15436 2796 15442 2808
rect 16298 2796 16304 2808
rect 16356 2796 16362 2848
rect 16399 2839 16457 2845
rect 16399 2805 16411 2839
rect 16445 2836 16457 2839
rect 16574 2836 16580 2848
rect 16445 2808 16580 2836
rect 16445 2805 16457 2808
rect 16399 2799 16457 2805
rect 16574 2796 16580 2808
rect 16632 2796 16638 2848
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 19159 2839 19217 2845
rect 19159 2836 19171 2839
rect 18748 2808 19171 2836
rect 18748 2796 18754 2808
rect 19159 2805 19171 2808
rect 19205 2805 19217 2839
rect 19159 2799 19217 2805
rect 21266 2796 21272 2848
rect 21324 2836 21330 2848
rect 21367 2839 21425 2845
rect 21367 2836 21379 2839
rect 21324 2808 21379 2836
rect 21324 2796 21330 2808
rect 21367 2805 21379 2808
rect 21413 2805 21425 2839
rect 21367 2799 21425 2805
rect 21726 2796 21732 2848
rect 21784 2836 21790 2848
rect 22664 2836 22692 2876
rect 21784 2808 22692 2836
rect 22848 2836 22876 2876
rect 23293 2839 23351 2845
rect 23293 2836 23305 2839
rect 22848 2808 23305 2836
rect 21784 2796 21790 2808
rect 23293 2805 23305 2808
rect 23339 2805 23351 2839
rect 23293 2799 23351 2805
rect 23842 2796 23848 2848
rect 23900 2836 23906 2848
rect 24118 2836 24124 2848
rect 23900 2808 24124 2836
rect 23900 2796 23906 2808
rect 24118 2796 24124 2808
rect 24176 2836 24182 2848
rect 24311 2839 24369 2845
rect 24311 2836 24323 2839
rect 24176 2808 24323 2836
rect 24176 2796 24182 2808
rect 24311 2805 24323 2808
rect 24357 2805 24369 2839
rect 24311 2799 24369 2805
rect 26694 2796 26700 2848
rect 26752 2845 26758 2848
rect 26752 2836 26761 2845
rect 26752 2808 26797 2836
rect 26752 2799 26761 2808
rect 26752 2796 26758 2799
rect 27338 2796 27344 2848
rect 27396 2836 27402 2848
rect 28077 2839 28135 2845
rect 28077 2836 28089 2839
rect 27396 2808 28089 2836
rect 27396 2796 27402 2808
rect 28077 2805 28089 2808
rect 28123 2805 28135 2839
rect 28077 2799 28135 2805
rect 552 2746 31072 2768
rect 552 2694 7988 2746
rect 8040 2694 8052 2746
rect 8104 2694 8116 2746
rect 8168 2694 8180 2746
rect 8232 2694 8244 2746
rect 8296 2694 15578 2746
rect 15630 2694 15642 2746
rect 15694 2694 15706 2746
rect 15758 2694 15770 2746
rect 15822 2694 15834 2746
rect 15886 2694 23168 2746
rect 23220 2694 23232 2746
rect 23284 2694 23296 2746
rect 23348 2694 23360 2746
rect 23412 2694 23424 2746
rect 23476 2694 30758 2746
rect 30810 2694 30822 2746
rect 30874 2694 30886 2746
rect 30938 2694 30950 2746
rect 31002 2694 31014 2746
rect 31066 2694 31072 2746
rect 552 2672 31072 2694
rect 845 2635 903 2641
rect 845 2601 857 2635
rect 891 2632 903 2635
rect 891 2604 1440 2632
rect 891 2601 903 2604
rect 845 2595 903 2601
rect 934 2524 940 2576
rect 992 2564 998 2576
rect 992 2536 1348 2564
rect 992 2524 998 2536
rect 1029 2499 1087 2505
rect 1029 2465 1041 2499
rect 1075 2496 1087 2499
rect 1118 2496 1124 2508
rect 1075 2468 1124 2496
rect 1075 2465 1087 2468
rect 1029 2459 1087 2465
rect 1118 2456 1124 2468
rect 1176 2456 1182 2508
rect 1320 2505 1348 2536
rect 1305 2499 1363 2505
rect 1305 2465 1317 2499
rect 1351 2465 1363 2499
rect 1412 2496 1440 2604
rect 1762 2592 1768 2644
rect 1820 2641 1826 2644
rect 1820 2595 1829 2641
rect 1820 2592 1826 2595
rect 3142 2592 3148 2644
rect 3200 2592 3206 2644
rect 4706 2632 4712 2644
rect 3252 2604 4712 2632
rect 1670 2496 1676 2508
rect 1412 2468 1676 2496
rect 1305 2459 1363 2465
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 2314 2496 2320 2508
rect 1826 2468 2320 2496
rect 1826 2439 1854 2468
rect 2314 2456 2320 2468
rect 2372 2456 2378 2508
rect 1811 2433 1869 2439
rect 1811 2399 1823 2433
rect 1857 2399 1869 2433
rect 1811 2393 1869 2399
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2428 2099 2431
rect 3252 2428 3280 2604
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 5994 2592 6000 2644
rect 6052 2632 6058 2644
rect 6822 2632 6828 2644
rect 6052 2604 6500 2632
rect 6052 2592 6058 2604
rect 5902 2564 5908 2576
rect 5736 2536 5908 2564
rect 3326 2456 3332 2508
rect 3384 2496 3390 2508
rect 3513 2499 3571 2505
rect 3513 2496 3525 2499
rect 3384 2468 3525 2496
rect 3384 2456 3390 2468
rect 3513 2465 3525 2468
rect 3559 2465 3571 2499
rect 3513 2459 3571 2465
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 4522 2496 4528 2508
rect 4295 2468 4528 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 4522 2456 4528 2468
rect 4580 2456 4586 2508
rect 4706 2456 4712 2508
rect 4764 2496 4770 2508
rect 5736 2496 5764 2536
rect 5902 2524 5908 2536
rect 5960 2564 5966 2576
rect 6089 2567 6147 2573
rect 6089 2564 6101 2567
rect 5960 2536 6101 2564
rect 5960 2524 5966 2536
rect 6089 2533 6101 2536
rect 6135 2533 6147 2567
rect 6089 2527 6147 2533
rect 6472 2508 6500 2604
rect 6570 2604 6828 2632
rect 4764 2468 5764 2496
rect 4764 2456 4770 2468
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 6362 2496 6368 2508
rect 5868 2468 6368 2496
rect 5868 2456 5874 2468
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 6454 2456 6460 2508
rect 6512 2456 6518 2508
rect 3840 2431 3898 2437
rect 3840 2428 3852 2431
rect 2087 2400 3280 2428
rect 3528 2400 3852 2428
rect 2087 2397 2099 2400
rect 2041 2391 2099 2397
rect 3528 2292 3556 2400
rect 3840 2397 3852 2400
rect 3886 2397 3898 2431
rect 3840 2391 3898 2397
rect 3970 2388 3976 2440
rect 4028 2388 4034 2440
rect 6570 2428 6598 2604
rect 6822 2592 6828 2604
rect 6880 2632 6886 2644
rect 6923 2635 6981 2641
rect 6923 2632 6935 2635
rect 6880 2604 6935 2632
rect 6880 2592 6886 2604
rect 6923 2601 6935 2604
rect 6969 2601 6981 2635
rect 6923 2595 6981 2601
rect 9122 2592 9128 2644
rect 9180 2641 9186 2644
rect 9180 2632 9189 2641
rect 9180 2604 9225 2632
rect 9180 2595 9189 2604
rect 9180 2592 9186 2595
rect 11238 2592 11244 2644
rect 11296 2592 11302 2644
rect 11698 2592 11704 2644
rect 11756 2632 11762 2644
rect 12075 2635 12133 2641
rect 12075 2632 12087 2635
rect 11756 2604 12087 2632
rect 11756 2592 11762 2604
rect 12075 2601 12087 2604
rect 12121 2601 12133 2635
rect 12075 2595 12133 2601
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 13722 2632 13728 2644
rect 12492 2604 13728 2632
rect 12492 2592 12498 2604
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 14182 2592 14188 2644
rect 14240 2632 14246 2644
rect 14283 2635 14341 2641
rect 14283 2632 14295 2635
rect 14240 2604 14295 2632
rect 14240 2592 14246 2604
rect 14283 2601 14295 2604
rect 14329 2601 14341 2635
rect 14283 2595 14341 2601
rect 16574 2592 16580 2644
rect 16632 2641 16638 2644
rect 16632 2632 16641 2641
rect 16632 2604 16677 2632
rect 16632 2595 16641 2604
rect 16632 2592 16638 2595
rect 18230 2592 18236 2644
rect 18288 2632 18294 2644
rect 20990 2632 20996 2644
rect 18288 2604 20996 2632
rect 18288 2592 18294 2604
rect 20990 2592 20996 2604
rect 21048 2592 21054 2644
rect 21266 2592 21272 2644
rect 21324 2632 21330 2644
rect 21735 2635 21793 2641
rect 21735 2632 21747 2635
rect 21324 2604 21747 2632
rect 21324 2592 21330 2604
rect 21735 2601 21747 2604
rect 21781 2601 21793 2635
rect 26694 2632 26700 2644
rect 21735 2595 21793 2601
rect 23492 2604 26700 2632
rect 20441 2567 20499 2573
rect 20441 2533 20453 2567
rect 20487 2564 20499 2567
rect 20487 2536 21407 2564
rect 20487 2533 20499 2536
rect 20441 2527 20499 2533
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 6788 2468 6963 2496
rect 6788 2456 6794 2468
rect 6935 2439 6963 2468
rect 7190 2456 7196 2508
rect 7248 2456 7254 2508
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 8619 2468 9168 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 4908 2400 6598 2428
rect 6920 2433 6978 2439
rect 9140 2437 9168 2468
rect 9306 2456 9312 2508
rect 9364 2496 9370 2508
rect 9401 2499 9459 2505
rect 9401 2496 9413 2499
rect 9364 2468 9413 2496
rect 9364 2456 9370 2468
rect 9401 2465 9413 2468
rect 9447 2465 9459 2499
rect 9401 2459 9459 2465
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2496 11207 2499
rect 11882 2496 11888 2508
rect 11195 2468 11888 2496
rect 11195 2465 11207 2468
rect 11149 2459 11207 2465
rect 11882 2456 11888 2468
rect 11940 2456 11946 2508
rect 15933 2499 15991 2505
rect 11992 2468 12388 2496
rect 4908 2292 4936 2400
rect 6920 2399 6932 2433
rect 6966 2399 6978 2433
rect 6920 2393 6978 2399
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 9128 2431 9186 2437
rect 9128 2397 9140 2431
rect 9174 2397 9186 2431
rect 9128 2391 9186 2397
rect 5626 2320 5632 2372
rect 5684 2360 5690 2372
rect 6362 2360 6368 2372
rect 5684 2332 6368 2360
rect 5684 2320 5690 2332
rect 6362 2320 6368 2332
rect 6420 2320 6426 2372
rect 3528 2264 4936 2292
rect 5537 2295 5595 2301
rect 5537 2261 5549 2295
rect 5583 2292 5595 2295
rect 7282 2292 7288 2304
rect 5583 2264 7288 2292
rect 5583 2261 5595 2264
rect 5537 2255 5595 2261
rect 7282 2252 7288 2264
rect 7340 2252 7346 2304
rect 8680 2292 8708 2391
rect 11238 2388 11244 2440
rect 11296 2428 11302 2440
rect 11606 2428 11612 2440
rect 11296 2400 11612 2428
rect 11296 2388 11302 2400
rect 11606 2388 11612 2400
rect 11664 2388 11670 2440
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 11992 2428 12020 2468
rect 12158 2437 12164 2440
rect 11848 2400 12020 2428
rect 12115 2431 12164 2437
rect 11848 2388 11854 2400
rect 12115 2397 12127 2431
rect 12161 2397 12164 2431
rect 12115 2391 12164 2397
rect 12158 2388 12164 2391
rect 12216 2388 12222 2440
rect 12360 2437 12388 2468
rect 13096 2468 14596 2496
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 9030 2292 9036 2304
rect 8680 2264 9036 2292
rect 9030 2252 9036 2264
rect 9088 2252 9094 2304
rect 10689 2295 10747 2301
rect 10689 2261 10701 2295
rect 10735 2292 10747 2295
rect 11974 2292 11980 2304
rect 10735 2264 11980 2292
rect 10735 2261 10747 2264
rect 10689 2255 10747 2261
rect 11974 2252 11980 2264
rect 12032 2252 12038 2304
rect 12342 2252 12348 2304
rect 12400 2292 12406 2304
rect 13096 2292 13124 2468
rect 13722 2388 13728 2440
rect 13780 2428 13786 2440
rect 13817 2431 13875 2437
rect 13817 2428 13829 2431
rect 13780 2400 13829 2428
rect 13780 2388 13786 2400
rect 13817 2397 13829 2400
rect 13863 2397 13875 2431
rect 13817 2391 13875 2397
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 14568 2437 14596 2468
rect 15933 2465 15945 2499
rect 15979 2496 15991 2499
rect 18233 2499 18291 2505
rect 15979 2468 16620 2496
rect 15979 2465 15991 2468
rect 15933 2459 15991 2465
rect 14280 2431 14338 2437
rect 14280 2428 14292 2431
rect 14148 2400 14292 2428
rect 14148 2388 14154 2400
rect 14280 2397 14292 2400
rect 14326 2397 14338 2431
rect 14280 2391 14338 2397
rect 14553 2431 14611 2437
rect 14553 2397 14565 2431
rect 14599 2397 14611 2431
rect 14553 2391 14611 2397
rect 16022 2388 16028 2440
rect 16080 2428 16086 2440
rect 16592 2437 16620 2468
rect 18233 2465 18245 2499
rect 18279 2496 18291 2499
rect 18279 2468 18828 2496
rect 18279 2465 18291 2468
rect 18233 2459 18291 2465
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 16080 2400 16129 2428
rect 16080 2388 16086 2400
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 16580 2431 16638 2437
rect 16580 2397 16592 2431
rect 16626 2397 16638 2431
rect 16580 2391 16638 2397
rect 16853 2431 16911 2437
rect 16853 2397 16865 2431
rect 16899 2428 16911 2431
rect 17770 2428 17776 2440
rect 16899 2400 17776 2428
rect 16899 2397 16911 2400
rect 16853 2391 16911 2397
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 18325 2431 18383 2437
rect 18325 2397 18337 2431
rect 18371 2428 18383 2431
rect 18506 2428 18512 2440
rect 18371 2400 18512 2428
rect 18371 2397 18383 2400
rect 18325 2391 18383 2397
rect 18506 2388 18512 2400
rect 18564 2388 18570 2440
rect 18690 2437 18696 2440
rect 18652 2431 18696 2437
rect 18652 2397 18664 2431
rect 18652 2391 18696 2397
rect 18690 2388 18696 2391
rect 18748 2388 18754 2440
rect 18800 2437 18828 2468
rect 19150 2456 19156 2508
rect 19208 2496 19214 2508
rect 20530 2496 20536 2508
rect 19208 2468 20536 2496
rect 19208 2456 19214 2468
rect 20530 2456 20536 2468
rect 20588 2456 20594 2508
rect 20806 2456 20812 2508
rect 20864 2496 20870 2508
rect 21269 2499 21327 2505
rect 21269 2496 21281 2499
rect 20864 2468 21281 2496
rect 20864 2456 20870 2468
rect 21269 2465 21281 2468
rect 21315 2465 21327 2499
rect 21379 2496 21407 2536
rect 23492 2496 23520 2604
rect 26694 2592 26700 2604
rect 26752 2632 26758 2644
rect 26887 2635 26945 2641
rect 26887 2632 26899 2635
rect 26752 2604 26899 2632
rect 26752 2592 26758 2604
rect 26887 2601 26899 2604
rect 26933 2601 26945 2635
rect 26887 2595 26945 2601
rect 28810 2592 28816 2644
rect 28868 2592 28874 2644
rect 29362 2592 29368 2644
rect 29420 2592 29426 2644
rect 23658 2524 23664 2576
rect 23716 2564 23722 2576
rect 23937 2567 23995 2573
rect 23937 2564 23949 2567
rect 23716 2536 23949 2564
rect 23716 2524 23722 2536
rect 23937 2533 23949 2536
rect 23983 2533 23995 2567
rect 23937 2527 23995 2533
rect 26418 2524 26424 2576
rect 26476 2524 26482 2576
rect 29086 2564 29092 2576
rect 28644 2536 29092 2564
rect 21379 2468 21680 2496
rect 21269 2459 21327 2465
rect 18788 2431 18846 2437
rect 18788 2397 18800 2431
rect 18834 2397 18846 2431
rect 18788 2391 18846 2397
rect 19061 2431 19119 2437
rect 19061 2397 19073 2431
rect 19107 2428 19119 2431
rect 20717 2431 20775 2437
rect 19107 2400 20668 2428
rect 19107 2397 19119 2400
rect 19061 2391 19119 2397
rect 13170 2320 13176 2372
rect 13228 2360 13234 2372
rect 20640 2360 20668 2400
rect 20717 2397 20729 2431
rect 20763 2428 20775 2431
rect 21174 2428 21180 2440
rect 20763 2400 21180 2428
rect 20763 2397 20775 2400
rect 20717 2391 20775 2397
rect 21174 2388 21180 2400
rect 21232 2388 21238 2440
rect 21652 2428 21680 2468
rect 21928 2468 23520 2496
rect 23569 2499 23627 2505
rect 21928 2440 21956 2468
rect 23569 2465 23581 2499
rect 23615 2496 23627 2499
rect 23750 2496 23756 2508
rect 23615 2468 23756 2496
rect 23615 2465 23627 2468
rect 23569 2459 23627 2465
rect 23750 2456 23756 2468
rect 23808 2496 23814 2508
rect 24026 2496 24032 2508
rect 23808 2468 24032 2496
rect 23808 2456 23814 2468
rect 24026 2456 24032 2468
rect 24084 2496 24090 2508
rect 24121 2499 24179 2505
rect 24121 2496 24133 2499
rect 24084 2468 24133 2496
rect 24084 2456 24090 2468
rect 24121 2465 24133 2468
rect 24167 2465 24179 2499
rect 24121 2459 24179 2465
rect 21732 2431 21790 2437
rect 21732 2428 21744 2431
rect 21652 2400 21744 2428
rect 21732 2397 21744 2400
rect 21778 2397 21790 2431
rect 21732 2391 21790 2397
rect 21910 2388 21916 2440
rect 21968 2388 21974 2440
rect 22002 2388 22008 2440
rect 22060 2388 22066 2440
rect 24136 2428 24164 2459
rect 24854 2456 24860 2508
rect 24912 2456 24918 2508
rect 26436 2496 26464 2524
rect 26436 2468 26740 2496
rect 24617 2449 24675 2455
rect 24617 2446 24629 2449
rect 24302 2428 24308 2440
rect 24136 2400 24308 2428
rect 24302 2388 24308 2400
rect 24360 2388 24366 2440
rect 24486 2437 24492 2440
rect 24448 2431 24492 2437
rect 24448 2397 24460 2431
rect 24448 2391 24492 2397
rect 24486 2388 24492 2391
rect 24544 2388 24550 2440
rect 24596 2415 24629 2446
rect 24663 2440 24675 2449
rect 24663 2415 24676 2440
rect 24596 2400 24676 2415
rect 24670 2388 24676 2400
rect 24728 2388 24734 2440
rect 25682 2388 25688 2440
rect 25740 2428 25746 2440
rect 26234 2428 26240 2440
rect 25740 2400 26240 2428
rect 25740 2388 25746 2400
rect 26234 2388 26240 2400
rect 26292 2428 26298 2440
rect 26421 2431 26479 2437
rect 26421 2428 26433 2431
rect 26292 2400 26433 2428
rect 26292 2388 26298 2400
rect 26421 2397 26433 2400
rect 26467 2397 26479 2431
rect 26712 2428 26740 2468
rect 27062 2456 27068 2508
rect 27120 2496 27126 2508
rect 28644 2505 28672 2536
rect 29086 2524 29092 2536
rect 29144 2564 29150 2576
rect 29454 2564 29460 2576
rect 29144 2536 29460 2564
rect 29144 2524 29150 2536
rect 29454 2524 29460 2536
rect 29512 2524 29518 2576
rect 27157 2499 27215 2505
rect 27157 2496 27169 2499
rect 27120 2468 27169 2496
rect 27120 2456 27126 2468
rect 27157 2465 27169 2468
rect 27203 2465 27215 2499
rect 28629 2499 28687 2505
rect 28629 2496 28641 2499
rect 27157 2459 27215 2465
rect 27264 2468 28641 2496
rect 26884 2431 26942 2437
rect 26884 2428 26896 2431
rect 26712 2400 26896 2428
rect 26421 2391 26479 2397
rect 26884 2397 26896 2400
rect 26930 2397 26942 2431
rect 26884 2391 26942 2397
rect 26970 2388 26976 2440
rect 27028 2428 27034 2440
rect 27264 2428 27292 2468
rect 28629 2465 28641 2468
rect 28675 2465 28687 2499
rect 28629 2459 28687 2465
rect 28810 2456 28816 2508
rect 28868 2496 28874 2508
rect 28905 2499 28963 2505
rect 28905 2496 28917 2499
rect 28868 2468 28917 2496
rect 28868 2456 28874 2468
rect 28905 2465 28917 2468
rect 28951 2465 28963 2499
rect 28905 2459 28963 2465
rect 29181 2499 29239 2505
rect 29181 2465 29193 2499
rect 29227 2496 29239 2499
rect 29730 2496 29736 2508
rect 29227 2468 29736 2496
rect 29227 2465 29239 2468
rect 29181 2459 29239 2465
rect 29730 2456 29736 2468
rect 29788 2456 29794 2508
rect 29546 2428 29552 2440
rect 27028 2400 27292 2428
rect 28092 2400 29552 2428
rect 27028 2388 27034 2400
rect 21266 2360 21272 2372
rect 13228 2332 13860 2360
rect 20640 2332 21272 2360
rect 13228 2320 13234 2332
rect 12400 2264 13124 2292
rect 13633 2295 13691 2301
rect 12400 2252 12406 2264
rect 13633 2261 13645 2295
rect 13679 2292 13691 2295
rect 13722 2292 13728 2304
rect 13679 2264 13728 2292
rect 13679 2261 13691 2264
rect 13633 2255 13691 2261
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 13832 2292 13860 2332
rect 21266 2320 21272 2332
rect 21324 2320 21330 2372
rect 23474 2360 23480 2372
rect 22940 2332 23480 2360
rect 16666 2292 16672 2304
rect 13832 2264 16672 2292
rect 16666 2252 16672 2264
rect 16724 2292 16730 2304
rect 19242 2292 19248 2304
rect 16724 2264 19248 2292
rect 16724 2252 16730 2264
rect 19242 2252 19248 2264
rect 19300 2292 19306 2304
rect 20622 2292 20628 2304
rect 19300 2264 20628 2292
rect 19300 2252 19306 2264
rect 20622 2252 20628 2264
rect 20680 2252 20686 2304
rect 20990 2252 20996 2304
rect 21048 2292 21054 2304
rect 22940 2292 22968 2332
rect 23474 2320 23480 2332
rect 23532 2320 23538 2372
rect 21048 2264 22968 2292
rect 21048 2252 21054 2264
rect 23014 2252 23020 2304
rect 23072 2292 23078 2304
rect 23109 2295 23167 2301
rect 23109 2292 23121 2295
rect 23072 2264 23121 2292
rect 23072 2252 23078 2264
rect 23109 2261 23121 2264
rect 23155 2261 23167 2295
rect 23109 2255 23167 2261
rect 24302 2252 24308 2304
rect 24360 2292 24366 2304
rect 25961 2295 26019 2301
rect 25961 2292 25973 2295
rect 24360 2264 25973 2292
rect 24360 2252 24366 2264
rect 25961 2261 25973 2264
rect 26007 2261 26019 2295
rect 25961 2255 26019 2261
rect 26602 2252 26608 2304
rect 26660 2292 26666 2304
rect 28092 2292 28120 2400
rect 29546 2388 29552 2400
rect 29604 2388 29610 2440
rect 29086 2320 29092 2372
rect 29144 2320 29150 2372
rect 26660 2264 28120 2292
rect 26660 2252 26666 2264
rect 28258 2252 28264 2304
rect 28316 2252 28322 2304
rect 552 2202 30912 2224
rect 552 2150 4193 2202
rect 4245 2150 4257 2202
rect 4309 2150 4321 2202
rect 4373 2150 4385 2202
rect 4437 2150 4449 2202
rect 4501 2150 11783 2202
rect 11835 2150 11847 2202
rect 11899 2150 11911 2202
rect 11963 2150 11975 2202
rect 12027 2150 12039 2202
rect 12091 2150 19373 2202
rect 19425 2150 19437 2202
rect 19489 2150 19501 2202
rect 19553 2150 19565 2202
rect 19617 2150 19629 2202
rect 19681 2150 26963 2202
rect 27015 2150 27027 2202
rect 27079 2150 27091 2202
rect 27143 2150 27155 2202
rect 27207 2150 27219 2202
rect 27271 2150 30912 2202
rect 552 2128 30912 2150
rect 1302 2088 1308 2100
rect 952 2060 1308 2088
rect 952 1961 980 2060
rect 1302 2048 1308 2060
rect 1360 2088 1366 2100
rect 2866 2088 2872 2100
rect 1360 2060 2872 2088
rect 1360 2048 1366 2060
rect 2866 2048 2872 2060
rect 2924 2048 2930 2100
rect 2961 2091 3019 2097
rect 2961 2057 2973 2091
rect 3007 2088 3019 2091
rect 3970 2088 3976 2100
rect 3007 2060 3976 2088
rect 3007 2057 3019 2060
rect 2961 2051 3019 2057
rect 3970 2048 3976 2060
rect 4028 2048 4034 2100
rect 4614 2048 4620 2100
rect 4672 2088 4678 2100
rect 5353 2091 5411 2097
rect 5353 2088 5365 2091
rect 4672 2060 5365 2088
rect 4672 2048 4678 2060
rect 5353 2057 5365 2060
rect 5399 2057 5411 2091
rect 5353 2051 5411 2057
rect 6638 2048 6644 2100
rect 6696 2088 6702 2100
rect 7745 2091 7803 2097
rect 7745 2088 7757 2091
rect 6696 2060 7757 2088
rect 6696 2048 6702 2060
rect 7745 2057 7757 2060
rect 7791 2057 7803 2091
rect 7745 2051 7803 2057
rect 8757 2091 8815 2097
rect 8757 2057 8769 2091
rect 8803 2088 8815 2091
rect 8846 2088 8852 2100
rect 8803 2060 8852 2088
rect 8803 2057 8815 2060
rect 8757 2051 8815 2057
rect 8846 2048 8852 2060
rect 8904 2048 8910 2100
rect 10962 2048 10968 2100
rect 11020 2088 11026 2100
rect 11974 2088 11980 2100
rect 11020 2060 11980 2088
rect 11020 2048 11026 2060
rect 11974 2048 11980 2060
rect 12032 2048 12038 2100
rect 12066 2048 12072 2100
rect 12124 2088 12130 2100
rect 13170 2088 13176 2100
rect 12124 2060 13176 2088
rect 12124 2048 12130 2060
rect 13170 2048 13176 2060
rect 13228 2048 13234 2100
rect 13265 2091 13323 2097
rect 13265 2057 13277 2091
rect 13311 2088 13323 2091
rect 14090 2088 14096 2100
rect 13311 2060 14096 2088
rect 13311 2057 13323 2060
rect 13265 2051 13323 2057
rect 14090 2048 14096 2060
rect 14148 2048 14154 2100
rect 14550 2048 14556 2100
rect 14608 2088 14614 2100
rect 14608 2060 17908 2088
rect 14608 2048 14614 2060
rect 3237 2023 3295 2029
rect 3237 1989 3249 2023
rect 3283 2020 3295 2023
rect 3418 2020 3424 2032
rect 3283 1992 3424 2020
rect 3283 1989 3295 1992
rect 3237 1983 3295 1989
rect 3418 1980 3424 1992
rect 3476 1980 3482 2032
rect 17880 2020 17908 2060
rect 17954 2048 17960 2100
rect 18012 2088 18018 2100
rect 18049 2091 18107 2097
rect 18049 2088 18061 2091
rect 18012 2060 18061 2088
rect 18012 2048 18018 2060
rect 18049 2057 18061 2060
rect 18095 2057 18107 2091
rect 21450 2088 21456 2100
rect 18049 2051 18107 2057
rect 18248 2060 21456 2088
rect 18248 2020 18276 2060
rect 21450 2048 21456 2060
rect 21508 2048 21514 2100
rect 22002 2048 22008 2100
rect 22060 2088 22066 2100
rect 23845 2091 23903 2097
rect 23845 2088 23857 2091
rect 22060 2060 23857 2088
rect 22060 2048 22066 2060
rect 23845 2057 23857 2060
rect 23891 2057 23903 2091
rect 23845 2051 23903 2057
rect 23952 2060 26280 2088
rect 17880 1992 18276 2020
rect 18325 2023 18383 2029
rect 18325 1989 18337 2023
rect 18371 1989 18383 2023
rect 18325 1983 18383 1989
rect 937 1955 995 1961
rect 937 1921 949 1955
rect 983 1921 995 1955
rect 937 1915 995 1921
rect 1443 1955 1501 1961
rect 1443 1921 1455 1955
rect 1489 1921 1501 1955
rect 1443 1915 1501 1921
rect 1673 1955 1731 1961
rect 1673 1921 1685 1955
rect 1719 1952 1731 1955
rect 2590 1952 2596 1964
rect 1719 1924 2596 1952
rect 1719 1921 1731 1924
rect 1673 1915 1731 1921
rect 1458 1884 1486 1915
rect 2590 1912 2596 1924
rect 2648 1912 2654 1964
rect 3694 1952 3700 1964
rect 3436 1924 3700 1952
rect 2130 1884 2136 1896
rect 1458 1856 2136 1884
rect 2130 1844 2136 1856
rect 2188 1844 2194 1896
rect 3326 1844 3332 1896
rect 3384 1844 3390 1896
rect 3436 1893 3464 1924
rect 3694 1912 3700 1924
rect 3752 1912 3758 1964
rect 4062 1959 4068 1964
rect 4019 1953 4068 1959
rect 4019 1919 4031 1953
rect 4065 1919 4068 1953
rect 4019 1913 4068 1919
rect 4062 1912 4068 1913
rect 4120 1912 4126 1964
rect 4246 1912 4252 1964
rect 4304 1912 4310 1964
rect 5905 1955 5963 1961
rect 5905 1921 5917 1955
rect 5951 1952 5963 1955
rect 6270 1952 6276 1964
rect 5951 1924 6276 1952
rect 5951 1921 5963 1924
rect 5905 1915 5963 1921
rect 6270 1912 6276 1924
rect 6328 1912 6334 1964
rect 6362 1912 6368 1964
rect 6420 1912 6426 1964
rect 9030 1912 9036 1964
rect 9088 1912 9094 1964
rect 9214 1912 9220 1964
rect 9272 1952 9278 1964
rect 9360 1955 9418 1961
rect 9360 1952 9372 1955
rect 9272 1924 9372 1952
rect 9272 1912 9278 1924
rect 9360 1921 9372 1924
rect 9406 1921 9418 1955
rect 9360 1915 9418 1921
rect 9490 1912 9496 1964
rect 9548 1952 9554 1964
rect 11149 1955 11207 1961
rect 9548 1924 9593 1952
rect 9548 1912 9554 1924
rect 11149 1921 11161 1955
rect 11195 1952 11207 1955
rect 11704 1955 11762 1961
rect 11704 1952 11716 1955
rect 11195 1924 11716 1952
rect 11195 1921 11207 1924
rect 11149 1915 11207 1921
rect 11704 1921 11716 1924
rect 11750 1921 11762 1955
rect 11704 1915 11762 1921
rect 11790 1912 11796 1964
rect 11848 1912 11854 1964
rect 11974 1912 11980 1964
rect 12032 1912 12038 1964
rect 13630 1912 13636 1964
rect 13688 1912 13694 1964
rect 13998 1961 14004 1964
rect 13960 1955 14004 1961
rect 13960 1921 13972 1955
rect 13960 1915 14004 1921
rect 13998 1912 14004 1915
rect 14056 1912 14062 1964
rect 14112 1955 14170 1961
rect 14112 1921 14124 1955
rect 14158 1952 14170 1955
rect 15749 1955 15807 1961
rect 14158 1924 14228 1952
rect 14158 1921 14170 1924
rect 14112 1915 14170 1921
rect 3421 1887 3479 1893
rect 3421 1853 3433 1887
rect 3467 1853 3479 1887
rect 3421 1847 3479 1853
rect 3513 1887 3571 1893
rect 3513 1853 3525 1887
rect 3559 1853 3571 1887
rect 3513 1847 3571 1853
rect 3344 1816 3372 1844
rect 3528 1816 3556 1847
rect 3786 1844 3792 1896
rect 3844 1893 3850 1896
rect 3844 1887 3898 1893
rect 3844 1853 3852 1887
rect 3886 1853 3898 1887
rect 3844 1847 3898 1853
rect 3844 1844 3850 1847
rect 6178 1844 6184 1896
rect 6236 1884 6242 1896
rect 6641 1887 6699 1893
rect 6641 1884 6653 1887
rect 6236 1856 6653 1884
rect 6236 1844 6242 1856
rect 6641 1853 6653 1856
rect 6687 1853 6699 1887
rect 6641 1847 6699 1853
rect 8478 1844 8484 1896
rect 8536 1844 8542 1896
rect 9766 1844 9772 1896
rect 9824 1844 9830 1896
rect 11238 1844 11244 1896
rect 11296 1844 11302 1896
rect 11568 1887 11626 1893
rect 11568 1853 11580 1887
rect 11614 1884 11626 1887
rect 11808 1884 11836 1912
rect 14200 1884 14228 1924
rect 15749 1921 15761 1955
rect 15795 1952 15807 1955
rect 16304 1955 16362 1961
rect 16304 1952 16316 1955
rect 15795 1924 16316 1952
rect 15795 1921 15807 1924
rect 15749 1915 15807 1921
rect 16304 1921 16316 1924
rect 16350 1921 16362 1955
rect 16304 1915 16362 1921
rect 16577 1955 16635 1961
rect 16577 1921 16589 1955
rect 16623 1952 16635 1955
rect 18340 1952 18368 1983
rect 18506 1980 18512 2032
rect 18564 1980 18570 2032
rect 23109 2023 23167 2029
rect 23109 1989 23121 2023
rect 23155 1989 23167 2023
rect 23109 1983 23167 1989
rect 16623 1924 18368 1952
rect 18524 1952 18552 1980
rect 18693 1955 18751 1961
rect 18693 1952 18705 1955
rect 18524 1924 18705 1952
rect 16623 1921 16635 1924
rect 16577 1915 16635 1921
rect 18693 1921 18705 1924
rect 18739 1921 18751 1955
rect 18693 1915 18751 1921
rect 19150 1912 19156 1964
rect 19208 1952 19214 1964
rect 20809 1955 20867 1961
rect 19208 1924 19253 1952
rect 19208 1912 19214 1924
rect 20809 1921 20821 1955
rect 20855 1952 20867 1955
rect 21364 1955 21422 1961
rect 21364 1952 21376 1955
rect 20855 1924 21376 1952
rect 20855 1921 20867 1924
rect 20809 1915 20867 1921
rect 21364 1921 21376 1924
rect 21410 1921 21422 1955
rect 21364 1915 21422 1921
rect 21450 1912 21456 1964
rect 21508 1912 21514 1964
rect 21637 1955 21695 1961
rect 21637 1921 21649 1955
rect 21683 1952 21695 1955
rect 23124 1952 23152 1983
rect 23474 1980 23480 2032
rect 23532 2020 23538 2032
rect 23952 2020 23980 2060
rect 23532 1992 23980 2020
rect 23532 1980 23538 1992
rect 21683 1924 23152 1952
rect 23216 1950 23980 1952
rect 24044 1950 24532 1952
rect 23216 1924 24532 1950
rect 21683 1921 21695 1924
rect 21637 1915 21695 1921
rect 11614 1856 11836 1884
rect 13648 1880 14044 1884
rect 14108 1880 14228 1884
rect 13648 1856 14228 1880
rect 11614 1853 11626 1856
rect 11568 1847 11626 1853
rect 3344 1788 3556 1816
rect 13648 1760 13676 1856
rect 14016 1852 14136 1856
rect 14366 1844 14372 1896
rect 14424 1844 14430 1896
rect 15841 1887 15899 1893
rect 15841 1853 15853 1887
rect 15887 1884 15899 1887
rect 15930 1884 15936 1896
rect 15887 1856 15936 1884
rect 15887 1853 15899 1856
rect 15841 1847 15899 1853
rect 15930 1844 15936 1856
rect 15988 1844 15994 1896
rect 18230 1844 18236 1896
rect 18288 1844 18294 1896
rect 18322 1844 18328 1896
rect 18380 1884 18386 1896
rect 18509 1887 18567 1893
rect 18509 1884 18521 1887
rect 18380 1856 18521 1884
rect 18380 1844 18386 1856
rect 18509 1853 18521 1856
rect 18555 1853 18567 1887
rect 18509 1847 18567 1853
rect 17954 1776 17960 1828
rect 18012 1776 18018 1828
rect 1403 1751 1461 1757
rect 1403 1717 1415 1751
rect 1449 1748 1461 1751
rect 1762 1748 1768 1760
rect 1449 1720 1768 1748
rect 1449 1717 1461 1720
rect 1403 1711 1461 1717
rect 1762 1708 1768 1720
rect 1820 1748 1826 1760
rect 4706 1748 4712 1760
rect 1820 1720 4712 1748
rect 1820 1708 1826 1720
rect 4706 1708 4712 1720
rect 4764 1748 4770 1760
rect 6371 1751 6429 1757
rect 6371 1748 6383 1751
rect 4764 1720 6383 1748
rect 4764 1708 4770 1720
rect 6371 1717 6383 1720
rect 6417 1717 6429 1751
rect 6371 1711 6429 1717
rect 6546 1708 6552 1760
rect 6604 1748 6610 1760
rect 12066 1748 12072 1760
rect 6604 1720 12072 1748
rect 6604 1708 6610 1720
rect 12066 1708 12072 1720
rect 12124 1708 12130 1760
rect 13630 1708 13636 1760
rect 13688 1708 13694 1760
rect 16307 1751 16365 1757
rect 16307 1717 16319 1751
rect 16353 1748 16365 1751
rect 16574 1748 16580 1760
rect 16353 1720 16580 1748
rect 16353 1717 16365 1720
rect 16307 1711 16365 1717
rect 16574 1708 16580 1720
rect 16632 1708 16638 1760
rect 18524 1748 18552 1847
rect 18966 1844 18972 1896
rect 19024 1893 19030 1896
rect 19024 1887 19078 1893
rect 19024 1853 19032 1887
rect 19066 1853 19078 1887
rect 19024 1847 19078 1853
rect 19024 1844 19030 1847
rect 19426 1844 19432 1896
rect 19484 1844 19490 1896
rect 20901 1887 20959 1893
rect 20901 1853 20913 1887
rect 20947 1853 20959 1887
rect 21468 1884 21496 1912
rect 22738 1884 22744 1896
rect 21468 1856 22744 1884
rect 20901 1847 20959 1853
rect 20714 1776 20720 1828
rect 20772 1776 20778 1828
rect 20806 1776 20812 1828
rect 20864 1816 20870 1828
rect 20916 1816 20944 1847
rect 22738 1844 22744 1856
rect 22796 1844 22802 1896
rect 22922 1844 22928 1896
rect 22980 1884 22986 1896
rect 23216 1884 23244 1924
rect 23952 1922 24072 1924
rect 22980 1856 23244 1884
rect 22980 1844 22986 1856
rect 23290 1844 23296 1896
rect 23348 1844 23354 1896
rect 23474 1844 23480 1896
rect 23532 1884 23538 1896
rect 23569 1887 23627 1893
rect 23569 1884 23581 1887
rect 23532 1856 23581 1884
rect 23532 1844 23538 1856
rect 23569 1853 23581 1856
rect 23615 1853 23627 1887
rect 23569 1847 23627 1853
rect 24029 1887 24087 1893
rect 24029 1853 24041 1887
rect 24075 1853 24087 1887
rect 24029 1847 24087 1853
rect 24305 1887 24363 1893
rect 24305 1853 24317 1887
rect 24351 1884 24363 1887
rect 24394 1884 24400 1896
rect 24351 1856 24400 1884
rect 24351 1853 24363 1856
rect 24305 1847 24363 1853
rect 20864 1788 20944 1816
rect 23017 1819 23075 1825
rect 20864 1776 20870 1788
rect 23017 1785 23029 1819
rect 23063 1816 23075 1819
rect 23934 1816 23940 1828
rect 23063 1788 23940 1816
rect 23063 1785 23075 1788
rect 23017 1779 23075 1785
rect 23934 1776 23940 1788
rect 23992 1776 23998 1828
rect 19058 1748 19064 1760
rect 18524 1720 19064 1748
rect 19058 1708 19064 1720
rect 19116 1708 19122 1760
rect 19242 1708 19248 1760
rect 19300 1748 19306 1760
rect 20732 1748 20760 1776
rect 19300 1720 20760 1748
rect 19300 1708 19306 1720
rect 21174 1708 21180 1760
rect 21232 1748 21238 1760
rect 21367 1751 21425 1757
rect 21367 1748 21379 1751
rect 21232 1720 21379 1748
rect 21232 1708 21238 1720
rect 21367 1717 21379 1720
rect 21413 1717 21425 1751
rect 21367 1711 21425 1717
rect 22830 1708 22836 1760
rect 22888 1748 22894 1760
rect 23385 1751 23443 1757
rect 23385 1748 23397 1751
rect 22888 1720 23397 1748
rect 22888 1708 22894 1720
rect 23385 1717 23397 1720
rect 23431 1717 23443 1751
rect 23385 1711 23443 1717
rect 23658 1708 23664 1760
rect 23716 1748 23722 1760
rect 24044 1748 24072 1847
rect 24394 1844 24400 1856
rect 24452 1844 24458 1896
rect 24504 1884 24532 1924
rect 24762 1912 24768 1964
rect 24820 1912 24826 1964
rect 25038 1912 25044 1964
rect 25096 1912 25102 1964
rect 26252 1884 26280 2060
rect 26326 2048 26332 2100
rect 26384 2048 26390 2100
rect 27430 2088 27436 2100
rect 26715 2060 27436 2088
rect 26715 1961 26743 2060
rect 27430 2048 27436 2060
rect 27488 2048 27494 2100
rect 27890 2048 27896 2100
rect 27948 2088 27954 2100
rect 28626 2088 28632 2100
rect 27948 2060 28632 2088
rect 27948 2048 27954 2060
rect 28626 2048 28632 2060
rect 28684 2048 28690 2100
rect 28718 2048 28724 2100
rect 28776 2048 28782 2100
rect 29178 1980 29184 2032
rect 29236 1980 29242 2032
rect 26697 1955 26755 1961
rect 26697 1921 26709 1955
rect 26743 1921 26755 1955
rect 26697 1915 26755 1921
rect 27203 1955 27261 1961
rect 27203 1921 27215 1955
rect 27249 1952 27261 1955
rect 27338 1952 27344 1964
rect 27249 1924 27344 1952
rect 27249 1921 27261 1924
rect 27203 1915 27261 1921
rect 27338 1912 27344 1924
rect 27396 1912 27402 1964
rect 27433 1955 27491 1961
rect 27433 1921 27445 1955
rect 27479 1952 27491 1955
rect 29270 1952 29276 1964
rect 27479 1924 29276 1952
rect 27479 1921 27491 1924
rect 27433 1915 27491 1921
rect 29270 1912 29276 1924
rect 29328 1912 29334 1964
rect 26970 1884 26976 1896
rect 24504 1856 25728 1884
rect 26252 1856 26976 1884
rect 23716 1720 24072 1748
rect 23716 1708 23722 1720
rect 24210 1708 24216 1760
rect 24268 1748 24274 1760
rect 24578 1748 24584 1760
rect 24268 1720 24584 1748
rect 24268 1708 24274 1720
rect 24578 1708 24584 1720
rect 24636 1748 24642 1760
rect 24771 1751 24829 1757
rect 24771 1748 24783 1751
rect 24636 1720 24783 1748
rect 24636 1708 24642 1720
rect 24771 1717 24783 1720
rect 24817 1717 24829 1751
rect 25700 1748 25728 1856
rect 26970 1844 26976 1856
rect 27028 1844 27034 1896
rect 27798 1844 27804 1896
rect 27856 1884 27862 1896
rect 28902 1884 28908 1896
rect 27856 1856 28908 1884
rect 27856 1844 27862 1856
rect 28902 1844 28908 1856
rect 28960 1844 28966 1896
rect 28997 1887 29055 1893
rect 28997 1853 29009 1887
rect 29043 1884 29055 1887
rect 30006 1884 30012 1896
rect 29043 1856 30012 1884
rect 29043 1853 29055 1856
rect 28997 1847 29055 1853
rect 27062 1748 27068 1760
rect 25700 1720 27068 1748
rect 24771 1711 24829 1717
rect 27062 1708 27068 1720
rect 27120 1708 27126 1760
rect 27163 1751 27221 1757
rect 27163 1717 27175 1751
rect 27209 1748 27221 1751
rect 27522 1748 27528 1760
rect 27209 1720 27528 1748
rect 27209 1717 27221 1720
rect 27163 1711 27221 1717
rect 27522 1708 27528 1720
rect 27580 1708 27586 1760
rect 27706 1708 27712 1760
rect 27764 1748 27770 1760
rect 28810 1748 28816 1760
rect 27764 1720 28816 1748
rect 27764 1708 27770 1720
rect 28810 1708 28816 1720
rect 28868 1748 28874 1760
rect 29012 1748 29040 1847
rect 30006 1844 30012 1856
rect 30064 1844 30070 1896
rect 28868 1720 29040 1748
rect 28868 1708 28874 1720
rect 552 1658 31072 1680
rect 552 1606 7988 1658
rect 8040 1606 8052 1658
rect 8104 1606 8116 1658
rect 8168 1606 8180 1658
rect 8232 1606 8244 1658
rect 8296 1606 15578 1658
rect 15630 1606 15642 1658
rect 15694 1606 15706 1658
rect 15758 1606 15770 1658
rect 15822 1606 15834 1658
rect 15886 1606 23168 1658
rect 23220 1606 23232 1658
rect 23284 1606 23296 1658
rect 23348 1606 23360 1658
rect 23412 1606 23424 1658
rect 23476 1606 30758 1658
rect 30810 1606 30822 1658
rect 30874 1606 30886 1658
rect 30938 1606 30950 1658
rect 31002 1606 31014 1658
rect 31066 1606 31072 1658
rect 552 1584 31072 1606
rect 1762 1504 1768 1556
rect 1820 1553 1826 1556
rect 1820 1507 1829 1553
rect 1820 1504 1826 1507
rect 3786 1504 3792 1556
rect 3844 1544 3850 1556
rect 3979 1547 4037 1553
rect 3979 1544 3991 1547
rect 3844 1516 3991 1544
rect 3844 1504 3850 1516
rect 3979 1513 3991 1516
rect 4025 1544 4037 1547
rect 4614 1544 4620 1556
rect 4025 1516 4620 1544
rect 4025 1513 4037 1516
rect 3979 1507 4037 1513
rect 4614 1504 4620 1516
rect 4672 1504 4678 1556
rect 5534 1504 5540 1556
rect 5592 1504 5598 1556
rect 6822 1504 6828 1556
rect 6880 1544 6886 1556
rect 6923 1547 6981 1553
rect 6923 1544 6935 1547
rect 6880 1516 6935 1544
rect 6880 1504 6886 1516
rect 6923 1513 6935 1516
rect 6969 1513 6981 1547
rect 9030 1544 9036 1556
rect 6923 1507 6981 1513
rect 8680 1516 9036 1544
rect 5074 1436 5080 1488
rect 5132 1476 5138 1488
rect 6089 1479 6147 1485
rect 6089 1476 6101 1479
rect 5132 1448 6101 1476
rect 5132 1436 5138 1448
rect 6089 1445 6101 1448
rect 6135 1445 6147 1479
rect 6089 1439 6147 1445
rect 8680 1420 8708 1516
rect 9030 1504 9036 1516
rect 9088 1504 9094 1556
rect 11333 1547 11391 1553
rect 11333 1513 11345 1547
rect 11379 1513 11391 1547
rect 11333 1507 11391 1513
rect 11348 1476 11376 1507
rect 11698 1504 11704 1556
rect 11756 1544 11762 1556
rect 12075 1547 12133 1553
rect 12075 1544 12087 1547
rect 11756 1516 12087 1544
rect 11756 1504 11762 1516
rect 12075 1513 12087 1516
rect 12121 1513 12133 1547
rect 12075 1507 12133 1513
rect 12250 1504 12256 1556
rect 12308 1544 12314 1556
rect 12308 1516 13584 1544
rect 12308 1504 12314 1516
rect 13556 1476 13584 1516
rect 13630 1504 13636 1556
rect 13688 1504 13694 1556
rect 14090 1504 14096 1556
rect 14148 1544 14154 1556
rect 14283 1547 14341 1553
rect 14283 1544 14295 1547
rect 14148 1516 14295 1544
rect 14148 1504 14154 1516
rect 14283 1513 14295 1516
rect 14329 1513 14341 1547
rect 14283 1507 14341 1513
rect 16574 1504 16580 1556
rect 16632 1553 16638 1556
rect 16632 1544 16641 1553
rect 16632 1516 16677 1544
rect 16632 1507 16641 1516
rect 16632 1504 16638 1507
rect 18690 1504 18696 1556
rect 18748 1544 18754 1556
rect 18791 1547 18849 1553
rect 18791 1544 18803 1547
rect 18748 1516 18803 1544
rect 18748 1504 18754 1516
rect 18791 1513 18803 1516
rect 18837 1513 18849 1547
rect 18791 1507 18849 1513
rect 19426 1504 19432 1556
rect 19484 1544 19490 1556
rect 20533 1547 20591 1553
rect 20533 1544 20545 1547
rect 19484 1516 20545 1544
rect 19484 1504 19490 1516
rect 20533 1513 20545 1516
rect 20579 1513 20591 1547
rect 20533 1507 20591 1513
rect 21174 1504 21180 1556
rect 21232 1544 21238 1556
rect 21735 1547 21793 1553
rect 21735 1544 21747 1547
rect 21232 1516 21747 1544
rect 21232 1504 21238 1516
rect 21735 1513 21747 1516
rect 21781 1513 21793 1547
rect 21735 1507 21793 1513
rect 22738 1504 22744 1556
rect 22796 1544 22802 1556
rect 24486 1544 24492 1556
rect 22796 1516 24492 1544
rect 22796 1504 22802 1516
rect 24486 1504 24492 1516
rect 24544 1504 24550 1556
rect 26421 1547 26479 1553
rect 26421 1544 26433 1547
rect 24872 1516 26433 1544
rect 20441 1479 20499 1485
rect 11348 1448 11750 1476
rect 13556 1448 13952 1476
rect 1210 1368 1216 1420
rect 1268 1368 1274 1420
rect 1302 1368 1308 1420
rect 1360 1368 1366 1420
rect 1946 1408 1952 1420
rect 1826 1380 1952 1408
rect 1826 1351 1854 1380
rect 1946 1368 1952 1380
rect 2004 1368 2010 1420
rect 3421 1411 3479 1417
rect 3421 1377 3433 1411
rect 3467 1408 3479 1411
rect 3467 1380 5764 1408
rect 3467 1377 3479 1380
rect 3421 1371 3479 1377
rect 1811 1345 1869 1351
rect 1811 1311 1823 1345
rect 1857 1311 1869 1345
rect 1811 1305 1869 1311
rect 2038 1300 2044 1352
rect 2096 1300 2102 1352
rect 3326 1300 3332 1352
rect 3384 1340 3390 1352
rect 3513 1343 3571 1349
rect 3513 1340 3525 1343
rect 3384 1312 3525 1340
rect 3384 1300 3390 1312
rect 3513 1309 3525 1312
rect 3559 1340 3571 1343
rect 3878 1340 3884 1352
rect 3559 1312 3884 1340
rect 3559 1309 3571 1312
rect 3513 1303 3571 1309
rect 3878 1300 3884 1312
rect 3936 1300 3942 1352
rect 4062 1349 4068 1352
rect 4019 1343 4068 1349
rect 4019 1309 4031 1343
rect 4065 1309 4068 1343
rect 4019 1303 4068 1309
rect 4062 1300 4068 1303
rect 4120 1300 4126 1352
rect 4249 1343 4307 1349
rect 4249 1309 4261 1343
rect 4295 1340 4307 1343
rect 5350 1340 5356 1352
rect 4295 1312 5356 1340
rect 4295 1309 4307 1312
rect 4249 1303 4307 1309
rect 5350 1300 5356 1312
rect 5408 1300 5414 1352
rect 5736 1340 5764 1380
rect 5810 1368 5816 1420
rect 5868 1368 5874 1420
rect 6454 1368 6460 1420
rect 6512 1368 6518 1420
rect 8662 1368 8668 1420
rect 8720 1368 8726 1420
rect 9490 1408 9496 1420
rect 8864 1380 9496 1408
rect 6920 1361 6978 1367
rect 6920 1340 6932 1361
rect 5736 1327 6932 1340
rect 6966 1327 6978 1361
rect 5736 1321 6978 1327
rect 7193 1343 7251 1349
rect 5736 1312 6960 1321
rect 7193 1309 7205 1343
rect 7239 1340 7251 1343
rect 8573 1343 8631 1349
rect 7239 1312 7880 1340
rect 7239 1309 7251 1312
rect 7193 1303 7251 1309
rect 1029 1207 1087 1213
rect 1029 1173 1041 1207
rect 1075 1204 1087 1207
rect 7852 1204 7880 1312
rect 8573 1309 8585 1343
rect 8619 1340 8631 1343
rect 8864 1340 8892 1380
rect 9490 1368 9496 1380
rect 9548 1368 9554 1420
rect 11146 1368 11152 1420
rect 11204 1408 11210 1420
rect 11241 1411 11299 1417
rect 11241 1408 11253 1411
rect 11204 1380 11253 1408
rect 11204 1368 11210 1380
rect 11241 1377 11253 1380
rect 11287 1377 11299 1411
rect 11241 1371 11299 1377
rect 11514 1368 11520 1420
rect 11572 1368 11578 1420
rect 11606 1368 11612 1420
rect 11664 1368 11670 1420
rect 11722 1408 11750 1448
rect 12250 1408 12256 1420
rect 11722 1380 12256 1408
rect 12250 1368 12256 1380
rect 12308 1368 12314 1420
rect 13538 1368 13544 1420
rect 13596 1408 13602 1420
rect 13924 1408 13952 1448
rect 20441 1445 20453 1479
rect 20487 1476 20499 1479
rect 20487 1448 21404 1476
rect 20487 1445 20499 1448
rect 20441 1439 20499 1445
rect 15933 1411 15991 1417
rect 13596 1380 13676 1408
rect 13924 1380 14596 1408
rect 13596 1368 13602 1380
rect 9030 1349 9036 1352
rect 8619 1312 8892 1340
rect 8992 1343 9036 1349
rect 8619 1309 8631 1312
rect 8573 1303 8631 1309
rect 8992 1309 9004 1343
rect 8992 1303 9036 1309
rect 9030 1300 9036 1303
rect 9088 1300 9094 1352
rect 9214 1349 9220 1352
rect 9171 1343 9220 1349
rect 9171 1309 9183 1343
rect 9217 1309 9220 1343
rect 9171 1303 9220 1309
rect 9214 1300 9220 1303
rect 9272 1300 9278 1352
rect 9306 1300 9312 1352
rect 9364 1340 9370 1352
rect 9401 1343 9459 1349
rect 9401 1340 9413 1343
rect 9364 1312 9413 1340
rect 9364 1300 9370 1312
rect 9401 1309 9413 1312
rect 9447 1309 9459 1343
rect 9401 1303 9459 1309
rect 10781 1343 10839 1349
rect 10781 1309 10793 1343
rect 10827 1340 10839 1343
rect 12072 1343 12130 1349
rect 12072 1340 12084 1343
rect 10827 1312 12084 1340
rect 10827 1309 10839 1312
rect 10781 1303 10839 1309
rect 12072 1309 12084 1312
rect 12118 1309 12130 1343
rect 12072 1303 12130 1309
rect 12158 1300 12164 1352
rect 12216 1340 12222 1352
rect 12345 1343 12403 1349
rect 12345 1340 12357 1343
rect 12216 1312 12357 1340
rect 12216 1300 12222 1312
rect 12345 1309 12357 1312
rect 12391 1309 12403 1343
rect 13648 1340 13676 1380
rect 13817 1343 13875 1349
rect 13817 1342 13829 1343
rect 13740 1340 13829 1342
rect 13648 1314 13829 1340
rect 13648 1312 13768 1314
rect 12345 1303 12403 1309
rect 13817 1309 13829 1314
rect 13863 1309 13875 1343
rect 13817 1303 13875 1309
rect 13998 1300 14004 1352
rect 14056 1340 14062 1352
rect 14568 1349 14596 1380
rect 15933 1377 15945 1411
rect 15979 1408 15991 1411
rect 18233 1411 18291 1417
rect 15979 1380 16620 1408
rect 15979 1377 15991 1380
rect 15933 1371 15991 1377
rect 14280 1343 14338 1349
rect 14280 1340 14292 1343
rect 14056 1312 14292 1340
rect 14056 1300 14062 1312
rect 14280 1309 14292 1312
rect 14326 1309 14338 1343
rect 14280 1303 14338 1309
rect 14553 1343 14611 1349
rect 14553 1309 14565 1343
rect 14599 1309 14611 1343
rect 14553 1303 14611 1309
rect 16022 1300 16028 1352
rect 16080 1340 16086 1352
rect 16592 1349 16620 1380
rect 18233 1377 18245 1411
rect 18279 1408 18291 1411
rect 18279 1380 18828 1408
rect 18279 1377 18291 1380
rect 18233 1371 18291 1377
rect 16117 1343 16175 1349
rect 16117 1340 16129 1343
rect 16080 1312 16129 1340
rect 16080 1300 16086 1312
rect 16117 1309 16129 1312
rect 16163 1309 16175 1343
rect 16117 1303 16175 1309
rect 16580 1343 16638 1349
rect 16580 1309 16592 1343
rect 16626 1309 16638 1343
rect 16580 1303 16638 1309
rect 16850 1300 16856 1352
rect 16908 1300 16914 1352
rect 18325 1343 18383 1349
rect 18325 1309 18337 1343
rect 18371 1340 18383 1343
rect 18506 1340 18512 1352
rect 18371 1312 18512 1340
rect 18371 1309 18383 1312
rect 18325 1303 18383 1309
rect 18506 1300 18512 1312
rect 18564 1300 18570 1352
rect 18800 1349 18828 1380
rect 20714 1368 20720 1420
rect 20772 1368 20778 1420
rect 20806 1368 20812 1420
rect 20864 1408 20870 1420
rect 20864 1380 20944 1408
rect 20864 1368 20870 1380
rect 18788 1343 18846 1349
rect 18788 1309 18800 1343
rect 18834 1309 18846 1343
rect 18788 1303 18846 1309
rect 19061 1343 19119 1349
rect 19061 1309 19073 1343
rect 19107 1340 19119 1343
rect 20916 1340 20944 1380
rect 20990 1368 20996 1420
rect 21048 1368 21054 1420
rect 21269 1343 21327 1349
rect 21269 1340 21281 1343
rect 19107 1312 20852 1340
rect 20916 1312 21281 1340
rect 19107 1309 19119 1312
rect 19061 1303 19119 1309
rect 20824 1281 20852 1312
rect 21269 1309 21281 1312
rect 21315 1309 21327 1343
rect 21376 1340 21404 1448
rect 23385 1411 23443 1417
rect 23385 1377 23397 1411
rect 23431 1408 23443 1411
rect 23566 1408 23572 1420
rect 23431 1380 23572 1408
rect 23431 1377 23443 1380
rect 23385 1371 23443 1377
rect 23566 1368 23572 1380
rect 23624 1368 23630 1420
rect 23804 1411 23862 1417
rect 23804 1377 23816 1411
rect 23850 1408 23862 1411
rect 24026 1408 24032 1420
rect 23850 1380 24032 1408
rect 23850 1377 23862 1380
rect 23804 1371 23862 1377
rect 24026 1368 24032 1380
rect 24084 1368 24090 1420
rect 24872 1408 24900 1516
rect 26421 1513 26433 1516
rect 26467 1513 26479 1547
rect 26421 1507 26479 1513
rect 27157 1547 27215 1553
rect 27157 1513 27169 1547
rect 27203 1513 27215 1547
rect 27157 1507 27215 1513
rect 27172 1476 27200 1507
rect 27246 1504 27252 1556
rect 27304 1544 27310 1556
rect 27433 1547 27491 1553
rect 27433 1544 27445 1547
rect 27304 1516 27445 1544
rect 27304 1504 27310 1516
rect 27433 1513 27445 1516
rect 27479 1513 27491 1547
rect 27433 1507 27491 1513
rect 27522 1504 27528 1556
rect 27580 1544 27586 1556
rect 27991 1547 28049 1553
rect 27991 1544 28003 1547
rect 27580 1516 28003 1544
rect 27580 1504 27586 1516
rect 27991 1513 28003 1516
rect 28037 1513 28049 1547
rect 27991 1507 28049 1513
rect 28626 1504 28632 1556
rect 28684 1544 28690 1556
rect 29365 1547 29423 1553
rect 29365 1544 29377 1547
rect 28684 1516 29377 1544
rect 28684 1504 28690 1516
rect 29365 1513 29377 1516
rect 29411 1513 29423 1547
rect 29365 1507 29423 1513
rect 24228 1380 24900 1408
rect 24964 1448 27200 1476
rect 27264 1448 27660 1476
rect 21732 1343 21790 1349
rect 21732 1340 21744 1343
rect 21376 1312 21744 1340
rect 21269 1303 21327 1309
rect 21732 1309 21744 1312
rect 21778 1309 21790 1343
rect 21732 1303 21790 1309
rect 22005 1343 22063 1349
rect 22005 1309 22017 1343
rect 22051 1340 22063 1343
rect 22830 1340 22836 1352
rect 22051 1312 22836 1340
rect 22051 1309 22063 1312
rect 22005 1303 22063 1309
rect 22830 1300 22836 1312
rect 22888 1300 22894 1352
rect 23474 1300 23480 1352
rect 23532 1300 23538 1352
rect 23934 1300 23940 1352
rect 23992 1340 23998 1352
rect 24228 1349 24256 1380
rect 24213 1343 24271 1349
rect 23992 1312 24037 1340
rect 23992 1300 23998 1312
rect 24213 1309 24225 1343
rect 24259 1309 24271 1343
rect 24213 1303 24271 1309
rect 24578 1300 24584 1352
rect 24636 1340 24642 1352
rect 24964 1340 24992 1448
rect 25590 1368 25596 1420
rect 25648 1368 25654 1420
rect 25682 1368 25688 1420
rect 25740 1408 25746 1420
rect 25777 1411 25835 1417
rect 25777 1408 25789 1411
rect 25740 1380 25789 1408
rect 25740 1368 25746 1380
rect 25777 1377 25789 1380
rect 25823 1377 25835 1411
rect 25777 1371 25835 1377
rect 26602 1368 26608 1420
rect 26660 1368 26666 1420
rect 26881 1411 26939 1417
rect 26881 1377 26893 1411
rect 26927 1377 26939 1411
rect 26881 1371 26939 1377
rect 24636 1312 24992 1340
rect 26896 1340 26924 1371
rect 26970 1368 26976 1420
rect 27028 1368 27034 1420
rect 27264 1417 27292 1448
rect 27249 1411 27307 1417
rect 27249 1408 27261 1411
rect 27080 1380 27261 1408
rect 27080 1340 27108 1380
rect 27249 1377 27261 1380
rect 27295 1377 27307 1411
rect 27249 1371 27307 1377
rect 27430 1368 27436 1420
rect 27488 1408 27494 1420
rect 27525 1411 27583 1417
rect 27525 1408 27537 1411
rect 27488 1380 27537 1408
rect 27488 1368 27494 1380
rect 27525 1377 27537 1380
rect 27571 1377 27583 1411
rect 27632 1408 27660 1448
rect 27798 1408 27804 1420
rect 27632 1380 27804 1408
rect 27525 1371 27583 1377
rect 27798 1368 27804 1380
rect 27856 1368 27862 1420
rect 29730 1368 29736 1420
rect 29788 1368 29794 1420
rect 28021 1361 28079 1367
rect 28021 1358 28033 1361
rect 27706 1340 27712 1352
rect 26896 1312 27108 1340
rect 27540 1312 27712 1340
rect 24636 1300 24642 1312
rect 20809 1275 20867 1281
rect 20809 1241 20821 1275
rect 20855 1241 20867 1275
rect 20809 1235 20867 1241
rect 1075 1176 7880 1204
rect 1075 1173 1087 1176
rect 1029 1167 1087 1173
rect 8018 1164 8024 1216
rect 8076 1204 8082 1216
rect 9766 1204 9772 1216
rect 8076 1176 9772 1204
rect 8076 1164 8082 1176
rect 9766 1164 9772 1176
rect 9824 1164 9830 1216
rect 11057 1207 11115 1213
rect 11057 1173 11069 1207
rect 11103 1204 11115 1207
rect 12342 1204 12348 1216
rect 11103 1176 12348 1204
rect 11103 1173 11115 1176
rect 11057 1167 11115 1173
rect 12342 1164 12348 1176
rect 12400 1164 12406 1216
rect 14274 1164 14280 1216
rect 14332 1204 14338 1216
rect 19426 1204 19432 1216
rect 14332 1176 19432 1204
rect 14332 1164 14338 1176
rect 19426 1164 19432 1176
rect 19484 1164 19490 1216
rect 21910 1164 21916 1216
rect 21968 1204 21974 1216
rect 23492 1204 23520 1300
rect 26326 1232 26332 1284
rect 26384 1272 26390 1284
rect 27540 1272 27568 1312
rect 27706 1300 27712 1312
rect 27764 1300 27770 1352
rect 28000 1327 28033 1358
rect 28067 1352 28079 1361
rect 28067 1327 28080 1352
rect 28000 1312 28080 1327
rect 28074 1300 28080 1312
rect 28132 1300 28138 1352
rect 28166 1300 28172 1352
rect 28224 1340 28230 1352
rect 28261 1343 28319 1349
rect 28261 1340 28273 1343
rect 28224 1312 28273 1340
rect 28224 1300 28230 1312
rect 28261 1309 28273 1312
rect 28307 1309 28319 1343
rect 28261 1303 28319 1309
rect 26384 1244 27568 1272
rect 26384 1232 26390 1244
rect 23842 1204 23848 1216
rect 21968 1176 23848 1204
rect 21968 1164 21974 1176
rect 23842 1164 23848 1176
rect 23900 1164 23906 1216
rect 24394 1164 24400 1216
rect 24452 1204 24458 1216
rect 25869 1207 25927 1213
rect 25869 1204 25881 1207
rect 24452 1176 25881 1204
rect 24452 1164 24458 1176
rect 25869 1173 25881 1176
rect 25915 1173 25927 1207
rect 25869 1167 25927 1173
rect 26694 1164 26700 1216
rect 26752 1164 26758 1216
rect 26878 1164 26884 1216
rect 26936 1204 26942 1216
rect 29822 1204 29828 1216
rect 26936 1176 29828 1204
rect 26936 1164 26942 1176
rect 29822 1164 29828 1176
rect 29880 1164 29886 1216
rect 29914 1164 29920 1216
rect 29972 1164 29978 1216
rect 552 1114 30912 1136
rect 552 1062 4193 1114
rect 4245 1062 4257 1114
rect 4309 1062 4321 1114
rect 4373 1062 4385 1114
rect 4437 1062 4449 1114
rect 4501 1062 11783 1114
rect 11835 1062 11847 1114
rect 11899 1062 11911 1114
rect 11963 1062 11975 1114
rect 12027 1062 12039 1114
rect 12091 1062 19373 1114
rect 19425 1062 19437 1114
rect 19489 1062 19501 1114
rect 19553 1062 19565 1114
rect 19617 1062 19629 1114
rect 19681 1062 26963 1114
rect 27015 1062 27027 1114
rect 27079 1062 27091 1114
rect 27143 1062 27155 1114
rect 27207 1062 27219 1114
rect 27271 1062 30912 1114
rect 552 1040 30912 1062
rect 3326 1000 3332 1012
rect 952 972 3332 1000
rect 952 873 980 972
rect 3326 960 3332 972
rect 3384 960 3390 1012
rect 3510 960 3516 1012
rect 3568 960 3574 1012
rect 3881 1003 3939 1009
rect 3881 969 3893 1003
rect 3927 1000 3939 1003
rect 4798 1000 4804 1012
rect 3927 972 4804 1000
rect 3927 969 3939 972
rect 3881 963 3939 969
rect 4798 960 4804 972
rect 4856 960 4862 1012
rect 4982 960 4988 1012
rect 5040 960 5046 1012
rect 5169 1003 5227 1009
rect 5169 969 5181 1003
rect 5215 1000 5227 1003
rect 5258 1000 5264 1012
rect 5215 972 5264 1000
rect 5215 969 5227 972
rect 5169 963 5227 969
rect 5258 960 5264 972
rect 5316 960 5322 1012
rect 5445 1003 5503 1009
rect 5445 969 5457 1003
rect 5491 1000 5503 1003
rect 8113 1003 8171 1009
rect 5491 972 7512 1000
rect 5491 969 5503 972
rect 5445 963 5503 969
rect 937 867 995 873
rect 1486 871 1492 876
rect 937 833 949 867
rect 983 833 995 867
rect 937 827 995 833
rect 1443 865 1492 871
rect 1443 831 1455 865
rect 1489 831 1492 865
rect 1443 825 1492 831
rect 1486 824 1492 825
rect 1544 824 1550 876
rect 3053 867 3111 873
rect 3053 833 3065 867
rect 3099 864 3111 867
rect 5000 864 5028 960
rect 7484 932 7512 972
rect 8113 969 8125 1003
rect 8159 1000 8171 1003
rect 9214 1000 9220 1012
rect 8159 972 9220 1000
rect 8159 969 8171 972
rect 8113 963 8171 969
rect 9214 960 9220 972
rect 9272 960 9278 1012
rect 10962 960 10968 1012
rect 11020 960 11026 1012
rect 13541 1003 13599 1009
rect 11256 972 13492 1000
rect 8294 932 8300 944
rect 7484 904 8300 932
rect 8294 892 8300 904
rect 8352 892 8358 944
rect 3099 836 5028 864
rect 3099 833 3111 836
rect 3053 827 3111 833
rect 5166 824 5172 876
rect 5224 864 5230 876
rect 6089 867 6147 873
rect 5224 836 5672 864
rect 5224 824 5230 836
rect 5644 808 5672 836
rect 6089 833 6101 867
rect 6135 864 6147 867
rect 6454 864 6460 876
rect 6135 836 6460 864
rect 6135 833 6147 836
rect 6089 827 6147 833
rect 6454 824 6460 836
rect 6512 824 6518 876
rect 6638 873 6644 876
rect 6595 867 6644 873
rect 6595 833 6607 867
rect 6641 833 6644 867
rect 6595 827 6644 833
rect 6638 824 6644 827
rect 6696 824 6702 876
rect 6730 824 6736 876
rect 6788 864 6794 876
rect 6825 867 6883 873
rect 6825 864 6837 867
rect 6788 836 6837 864
rect 6788 824 6794 836
rect 6825 833 6837 836
rect 6871 833 6883 867
rect 6825 827 6883 833
rect 7282 824 7288 876
rect 7340 864 7346 876
rect 7340 836 8294 864
rect 7340 824 7346 836
rect 1673 799 1731 805
rect 1673 765 1685 799
rect 1719 796 1731 799
rect 1719 768 2774 796
rect 1719 765 1731 768
rect 1673 759 1731 765
rect 2746 728 2774 768
rect 3602 756 3608 808
rect 3660 796 3666 808
rect 5353 799 5411 805
rect 5353 796 5365 799
rect 3660 768 5365 796
rect 3660 756 3666 768
rect 5353 765 5365 768
rect 5399 765 5411 799
rect 5353 759 5411 765
rect 5626 756 5632 808
rect 5684 756 5690 808
rect 5994 756 6000 808
rect 6052 756 6058 808
rect 8018 796 8024 808
rect 6196 768 8024 796
rect 2746 700 4292 728
rect 4264 672 4292 700
rect 1403 663 1461 669
rect 1403 629 1415 663
rect 1449 660 1461 663
rect 3786 660 3792 672
rect 1449 632 3792 660
rect 1449 629 1461 632
rect 1403 623 1461 629
rect 3786 620 3792 632
rect 3844 620 3850 672
rect 4246 620 4252 672
rect 4304 620 4310 672
rect 5813 663 5871 669
rect 5813 629 5825 663
rect 5859 660 5871 663
rect 6196 660 6224 768
rect 8018 756 8024 768
rect 8076 756 8082 808
rect 8266 728 8294 836
rect 8662 824 8668 876
rect 8720 824 8726 876
rect 9030 873 9036 876
rect 8992 867 9036 873
rect 8992 833 9004 867
rect 8992 827 9036 833
rect 9030 824 9036 827
rect 9088 824 9094 876
rect 9128 867 9186 873
rect 9128 833 9140 867
rect 9174 833 9186 867
rect 9128 827 9186 833
rect 8570 756 8576 808
rect 8628 756 8634 808
rect 8680 792 9076 796
rect 9143 792 9171 827
rect 9398 824 9404 876
rect 9456 824 9462 876
rect 11256 873 11284 972
rect 13464 932 13492 972
rect 13541 969 13553 1003
rect 13587 1000 13599 1003
rect 14366 1000 14372 1012
rect 13587 972 14372 1000
rect 13587 969 13599 972
rect 13541 963 13599 969
rect 14366 960 14372 972
rect 14424 960 14430 1012
rect 16117 1003 16175 1009
rect 16117 969 16129 1003
rect 16163 1000 16175 1003
rect 16850 1000 16856 1012
rect 16163 972 16856 1000
rect 16163 969 16175 972
rect 16117 963 16175 969
rect 16850 960 16856 972
rect 16908 960 16914 1012
rect 17770 960 17776 1012
rect 17828 1000 17834 1012
rect 18693 1003 18751 1009
rect 18693 1000 18705 1003
rect 17828 972 18705 1000
rect 17828 960 17834 972
rect 18693 969 18705 972
rect 18739 969 18751 1003
rect 20714 1000 20720 1012
rect 18693 963 18751 969
rect 18800 972 20720 1000
rect 13464 904 13860 932
rect 11790 873 11796 876
rect 11241 867 11299 873
rect 11241 833 11253 867
rect 11287 833 11299 867
rect 11241 827 11299 833
rect 11747 867 11796 873
rect 11747 833 11759 867
rect 11793 833 11796 867
rect 11747 827 11796 833
rect 11790 824 11796 827
rect 11848 824 11854 876
rect 13630 864 13636 876
rect 12176 836 13636 864
rect 12176 812 12204 836
rect 13630 824 13636 836
rect 13688 824 13694 876
rect 11146 796 11152 808
rect 8680 768 9171 792
rect 8680 728 8708 768
rect 9048 764 9171 768
rect 10244 768 11152 796
rect 10244 740 10272 768
rect 11146 756 11152 768
rect 11204 756 11210 808
rect 11882 796 11888 808
rect 11256 768 11888 796
rect 8266 700 8708 728
rect 10226 688 10232 740
rect 10284 688 10290 740
rect 11256 728 11284 768
rect 11882 756 11888 768
rect 11940 756 11946 808
rect 11977 799 12035 805
rect 11977 765 11989 799
rect 12023 796 12035 799
rect 12130 796 12204 812
rect 13832 808 13860 904
rect 18230 892 18236 944
rect 18288 892 18294 944
rect 14274 824 14280 876
rect 14332 873 14338 876
rect 14332 867 14381 873
rect 14332 833 14335 867
rect 14369 833 14381 867
rect 16899 867 16957 873
rect 14332 827 14381 833
rect 14476 836 16528 864
rect 14332 824 14338 827
rect 12023 784 12204 796
rect 12023 768 12158 784
rect 12023 765 12035 768
rect 11977 759 12035 765
rect 12986 756 12992 808
rect 13044 796 13050 808
rect 13725 799 13783 805
rect 13725 796 13737 799
rect 13044 768 13737 796
rect 13044 756 13050 768
rect 13725 765 13737 768
rect 13771 765 13783 799
rect 13725 759 13783 765
rect 13814 756 13820 808
rect 13872 756 13878 808
rect 14144 799 14202 805
rect 14144 796 14156 799
rect 13924 768 14156 796
rect 13924 728 13952 768
rect 14144 765 14156 768
rect 14190 796 14202 799
rect 14476 796 14504 836
rect 14190 768 14504 796
rect 14190 765 14202 768
rect 14144 759 14202 765
rect 14550 756 14556 808
rect 14608 756 14614 808
rect 15378 756 15384 808
rect 15436 796 15442 808
rect 16301 799 16359 805
rect 16301 796 16313 799
rect 15436 768 16313 796
rect 15436 756 15442 768
rect 16301 765 16313 768
rect 16347 765 16359 799
rect 16301 759 16359 765
rect 16393 799 16451 805
rect 16393 765 16405 799
rect 16439 765 16451 799
rect 16500 796 16528 836
rect 16899 833 16911 867
rect 16945 864 16957 867
rect 18800 864 18828 972
rect 20714 960 20720 972
rect 20772 960 20778 1012
rect 20824 972 23428 1000
rect 18874 892 18880 944
rect 18932 932 18938 944
rect 18932 904 19012 932
rect 18932 892 18938 904
rect 18984 873 19012 904
rect 16945 836 18828 864
rect 18969 867 19027 873
rect 16945 833 16957 836
rect 16899 827 16957 833
rect 18969 833 18981 867
rect 19015 833 19027 867
rect 18969 827 19027 833
rect 19150 824 19156 876
rect 19208 824 19214 876
rect 19334 873 19340 876
rect 19296 867 19340 873
rect 19296 833 19308 867
rect 19296 827 19340 833
rect 19334 824 19340 827
rect 19392 824 19398 876
rect 19518 871 19524 876
rect 19475 865 19524 871
rect 19475 831 19487 865
rect 19521 831 19524 865
rect 19475 825 19524 831
rect 19518 824 19524 825
rect 19576 824 19582 876
rect 19705 867 19763 873
rect 19705 833 19717 867
rect 19751 864 19763 867
rect 20714 864 20720 876
rect 19751 836 20720 864
rect 19751 833 19763 836
rect 19705 827 19763 833
rect 20714 824 20720 836
rect 20772 824 20778 876
rect 16720 799 16778 805
rect 16720 796 16732 799
rect 16500 768 16732 796
rect 16393 759 16451 765
rect 16720 765 16732 768
rect 16766 796 16778 799
rect 17034 796 17040 808
rect 16766 768 17040 796
rect 16766 765 16778 768
rect 16720 759 16778 765
rect 10336 700 11284 728
rect 13004 700 13952 728
rect 16408 728 16436 759
rect 17034 756 17040 768
rect 17092 756 17098 808
rect 17126 756 17132 808
rect 17184 756 17190 808
rect 18877 799 18935 805
rect 18877 765 18889 799
rect 18923 772 18935 799
rect 19168 796 19196 824
rect 20824 796 20852 972
rect 21266 892 21272 944
rect 21324 892 21330 944
rect 23400 932 23428 972
rect 23474 960 23480 1012
rect 23532 1000 23538 1012
rect 23569 1003 23627 1009
rect 23569 1000 23581 1003
rect 23532 972 23581 1000
rect 23532 960 23538 972
rect 23569 969 23581 972
rect 23615 969 23627 1003
rect 24578 1000 24584 1012
rect 23569 963 23627 969
rect 23676 972 24584 1000
rect 23676 932 23704 972
rect 24578 960 24584 972
rect 24636 960 24642 1012
rect 25682 960 25688 1012
rect 25740 960 25746 1012
rect 26694 1000 26700 1012
rect 26160 972 26700 1000
rect 23400 904 23704 932
rect 26053 935 26111 941
rect 26053 901 26065 935
rect 26099 901 26111 935
rect 26053 895 26111 901
rect 21545 867 21603 873
rect 21545 833 21557 867
rect 21591 864 21603 867
rect 21910 864 21916 876
rect 21591 836 21916 864
rect 21591 833 21603 836
rect 21545 827 21603 833
rect 21910 824 21916 836
rect 21968 824 21974 876
rect 22051 867 22109 873
rect 22051 833 22063 867
rect 22097 864 22109 867
rect 23014 864 23020 876
rect 22097 836 23020 864
rect 22097 833 22109 836
rect 22051 827 22109 833
rect 23014 824 23020 836
rect 23072 824 23078 876
rect 23566 824 23572 876
rect 23624 864 23630 876
rect 24308 867 24366 873
rect 24308 864 24320 867
rect 23624 836 24320 864
rect 23624 824 23630 836
rect 24308 833 24320 836
rect 24354 833 24366 867
rect 24308 827 24366 833
rect 24581 867 24639 873
rect 24581 833 24593 867
rect 24627 864 24639 867
rect 26068 864 26096 895
rect 24627 836 26096 864
rect 24627 833 24639 836
rect 24581 827 24639 833
rect 18923 765 19104 772
rect 19168 768 20852 796
rect 21453 799 21511 805
rect 18877 759 19104 765
rect 21453 765 21465 799
rect 21499 796 21511 799
rect 22186 796 22192 808
rect 21499 768 22192 796
rect 21499 765 21511 768
rect 21453 759 21511 765
rect 18892 744 19104 759
rect 16408 700 16528 728
rect 5859 632 6224 660
rect 6555 663 6613 669
rect 5859 629 5871 632
rect 5813 623 5871 629
rect 6555 629 6567 663
rect 6601 660 6613 663
rect 6822 660 6828 672
rect 6601 632 6828 660
rect 6601 629 6613 632
rect 6555 623 6613 629
rect 6822 620 6828 632
rect 6880 620 6886 672
rect 8389 663 8447 669
rect 8389 629 8401 663
rect 8435 660 8447 663
rect 10336 660 10364 700
rect 8435 632 10364 660
rect 10689 663 10747 669
rect 8435 629 8447 632
rect 8389 623 8447 629
rect 10689 629 10701 663
rect 10735 660 10747 663
rect 11606 660 11612 672
rect 10735 632 11612 660
rect 10735 629 10747 632
rect 10689 623 10747 629
rect 11606 620 11612 632
rect 11664 620 11670 672
rect 11707 663 11765 669
rect 11707 629 11719 663
rect 11753 660 11765 663
rect 13004 660 13032 700
rect 16500 672 16528 700
rect 11753 632 13032 660
rect 11753 629 11765 632
rect 11707 623 11765 629
rect 13078 620 13084 672
rect 13136 620 13142 672
rect 14458 620 14464 672
rect 14516 660 14522 672
rect 15657 663 15715 669
rect 15657 660 15669 663
rect 14516 632 15669 660
rect 14516 620 14522 632
rect 15657 629 15669 632
rect 15703 629 15715 663
rect 15657 623 15715 629
rect 16482 620 16488 672
rect 16540 620 16546 672
rect 19076 660 19104 744
rect 21358 728 21364 740
rect 20364 700 21364 728
rect 20364 660 20392 700
rect 21358 688 21364 700
rect 21416 728 21422 740
rect 21468 728 21496 759
rect 22186 756 22192 768
rect 22244 756 22250 808
rect 22281 799 22339 805
rect 22281 765 22293 799
rect 22327 796 22339 799
rect 22327 768 23796 796
rect 22327 765 22339 768
rect 22281 759 22339 765
rect 21416 700 21496 728
rect 23768 728 23796 768
rect 23842 756 23848 808
rect 23900 756 23906 808
rect 26160 796 26188 972
rect 26694 960 26700 972
rect 26752 960 26758 1012
rect 28534 960 28540 1012
rect 28592 960 28598 1012
rect 29181 1003 29239 1009
rect 29181 1000 29193 1003
rect 29012 972 29193 1000
rect 29012 944 29040 972
rect 29181 969 29193 972
rect 29227 969 29239 1003
rect 29181 963 29239 969
rect 29454 960 29460 1012
rect 29512 960 29518 1012
rect 28994 892 29000 944
rect 29052 892 29058 944
rect 26878 864 26884 876
rect 26252 836 26884 864
rect 26252 805 26280 836
rect 26878 824 26884 836
rect 26936 824 26942 876
rect 27203 867 27261 873
rect 27203 833 27215 867
rect 27249 864 27261 867
rect 28258 864 28264 876
rect 27249 836 28264 864
rect 27249 833 27261 836
rect 27203 827 27261 833
rect 28258 824 28264 836
rect 28316 824 28322 876
rect 29086 864 29092 876
rect 28920 836 29092 864
rect 23952 768 26188 796
rect 26237 799 26295 805
rect 23952 728 23980 768
rect 26237 765 26249 799
rect 26283 765 26295 799
rect 26237 759 26295 765
rect 26326 756 26332 808
rect 26384 796 26390 808
rect 26421 799 26479 805
rect 26421 796 26433 799
rect 26384 768 26433 796
rect 26384 756 26390 768
rect 26421 765 26433 768
rect 26467 765 26479 799
rect 26421 759 26479 765
rect 26697 799 26755 805
rect 26697 765 26709 799
rect 26743 796 26755 799
rect 27338 796 27344 808
rect 26743 768 27344 796
rect 26743 765 26755 768
rect 26697 759 26755 765
rect 27338 756 27344 768
rect 27396 756 27402 808
rect 27433 799 27491 805
rect 27433 765 27445 799
rect 27479 796 27491 799
rect 28920 796 28948 836
rect 29086 824 29092 836
rect 29144 824 29150 876
rect 27479 768 28948 796
rect 28997 799 29055 805
rect 27479 765 27491 768
rect 27433 759 27491 765
rect 28997 765 29009 799
rect 29043 796 29055 799
rect 29362 796 29368 808
rect 29043 768 29368 796
rect 29043 765 29055 768
rect 28997 759 29055 765
rect 29362 756 29368 768
rect 29420 756 29426 808
rect 23768 700 23980 728
rect 21416 688 21422 700
rect 19076 632 20392 660
rect 20438 620 20444 672
rect 20496 660 20502 672
rect 20809 663 20867 669
rect 20809 660 20821 663
rect 20496 632 20821 660
rect 20496 620 20502 632
rect 20809 629 20821 632
rect 20855 629 20867 663
rect 20809 623 20867 629
rect 22002 620 22008 672
rect 22060 669 22066 672
rect 22060 623 22069 669
rect 22060 620 22066 623
rect 22186 620 22192 672
rect 22244 660 22250 672
rect 23658 660 23664 672
rect 22244 632 23664 660
rect 22244 620 22250 632
rect 23658 620 23664 632
rect 23716 620 23722 672
rect 23934 620 23940 672
rect 23992 660 23998 672
rect 24311 663 24369 669
rect 24311 660 24323 663
rect 23992 632 24323 660
rect 23992 620 23998 632
rect 24311 629 24323 632
rect 24357 629 24369 663
rect 24311 623 24369 629
rect 24486 620 24492 672
rect 24544 660 24550 672
rect 26605 663 26663 669
rect 26605 660 26617 663
rect 24544 632 26617 660
rect 24544 620 24550 632
rect 26605 629 26617 632
rect 26651 629 26663 663
rect 26605 623 26663 629
rect 27163 663 27221 669
rect 27163 629 27175 663
rect 27209 660 27221 663
rect 27522 660 27528 672
rect 27209 632 27528 660
rect 27209 629 27221 632
rect 27163 623 27221 629
rect 27522 620 27528 632
rect 27580 620 27586 672
rect 552 570 31072 592
rect 552 518 7988 570
rect 8040 518 8052 570
rect 8104 518 8116 570
rect 8168 518 8180 570
rect 8232 518 8244 570
rect 8296 518 15578 570
rect 15630 518 15642 570
rect 15694 518 15706 570
rect 15758 518 15770 570
rect 15822 518 15834 570
rect 15886 518 23168 570
rect 23220 518 23232 570
rect 23284 518 23296 570
rect 23348 518 23360 570
rect 23412 518 23424 570
rect 23476 518 30758 570
rect 30810 518 30822 570
rect 30874 518 30886 570
rect 30938 518 30950 570
rect 31002 518 31014 570
rect 31066 518 31072 570
rect 552 496 31072 518
rect 1486 416 1492 468
rect 1544 416 1550 468
rect 2038 416 2044 468
rect 2096 456 2102 468
rect 2096 428 2774 456
rect 2096 416 2102 428
rect 1504 184 1532 416
rect 2746 252 2774 428
rect 5626 416 5632 468
rect 5684 416 5690 468
rect 5994 416 6000 468
rect 6052 456 6058 468
rect 10226 456 10232 468
rect 6052 428 10232 456
rect 6052 416 6058 428
rect 10226 416 10232 428
rect 10284 416 10290 468
rect 14458 456 14464 468
rect 11164 428 14464 456
rect 5644 388 5672 416
rect 8570 388 8576 400
rect 5644 360 8576 388
rect 8570 348 8576 360
rect 8628 388 8634 400
rect 10778 388 10784 400
rect 8628 360 10784 388
rect 8628 348 8634 360
rect 10778 348 10784 360
rect 10836 348 10842 400
rect 3970 280 3976 332
rect 4028 320 4034 332
rect 11164 320 11192 428
rect 14458 416 14464 428
rect 14516 416 14522 468
rect 17126 416 17132 468
rect 17184 456 17190 468
rect 19150 456 19156 468
rect 17184 428 19156 456
rect 17184 416 17190 428
rect 19150 416 19156 428
rect 19208 416 19214 468
rect 19518 416 19524 468
rect 19576 456 19582 468
rect 22094 456 22100 468
rect 19576 428 22100 456
rect 19576 416 19582 428
rect 22094 416 22100 428
rect 22152 416 22158 468
rect 24302 416 24308 468
rect 24360 416 24366 468
rect 13630 348 13636 400
rect 13688 388 13694 400
rect 22922 388 22928 400
rect 13688 360 22928 388
rect 13688 348 13694 360
rect 22922 348 22928 360
rect 22980 348 22986 400
rect 12986 320 12992 332
rect 4028 292 11192 320
rect 12406 292 12992 320
rect 4028 280 4034 292
rect 7650 252 7656 264
rect 2746 224 7656 252
rect 7650 212 7656 224
rect 7708 212 7714 264
rect 10778 212 10784 264
rect 10836 252 10842 264
rect 12406 252 12434 292
rect 12986 280 12992 292
rect 13044 280 13050 332
rect 13078 280 13084 332
rect 13136 280 13142 332
rect 17034 280 17040 332
rect 17092 320 17098 332
rect 22094 320 22100 332
rect 17092 292 22100 320
rect 17092 280 17098 292
rect 22094 280 22100 292
rect 22152 280 22158 332
rect 22186 280 22192 332
rect 22244 320 22250 332
rect 24320 320 24348 416
rect 22244 292 24348 320
rect 22244 280 22250 292
rect 10836 224 12434 252
rect 10836 212 10842 224
rect 13096 184 13124 280
rect 1504 156 13124 184
rect 13814 144 13820 196
rect 13872 184 13878 196
rect 16482 184 16488 196
rect 13872 156 16488 184
rect 13872 144 13878 156
rect 16482 144 16488 156
rect 16540 184 16546 196
rect 23750 184 23756 196
rect 16540 156 23756 184
rect 16540 144 16546 156
rect 23750 144 23756 156
rect 23808 144 23814 196
rect 22094 76 22100 128
rect 22152 116 22158 128
rect 24210 116 24216 128
rect 22152 88 24216 116
rect 22152 76 22158 88
rect 24210 76 24216 88
rect 24268 76 24274 128
rect 3878 8 3884 60
rect 3936 48 3942 60
rect 16206 48 16212 60
rect 3936 20 16212 48
rect 3936 8 3942 20
rect 16206 8 16212 20
rect 16264 48 16270 60
rect 18874 48 18880 60
rect 16264 20 18880 48
rect 16264 8 16270 20
rect 18874 8 18880 20
rect 18932 8 18938 60
<< via1 >>
rect 8208 22244 8260 22296
rect 11152 22244 11204 22296
rect 12256 22244 12308 22296
rect 6460 22176 6512 22228
rect 10048 22176 10100 22228
rect 10968 22176 11020 22228
rect 11060 22176 11112 22228
rect 14464 22176 14516 22228
rect 6092 22108 6144 22160
rect 9404 22108 9456 22160
rect 9956 22040 10008 22092
rect 10416 22040 10468 22092
rect 14004 22040 14056 22092
rect 2136 21836 2188 21888
rect 6644 21904 6696 21956
rect 12072 21904 12124 21956
rect 12256 21904 12308 21956
rect 12716 21904 12768 21956
rect 24124 22244 24176 22296
rect 22468 22176 22520 22228
rect 25596 22176 25648 22228
rect 14280 22040 14332 22092
rect 19340 22040 19392 22092
rect 19708 22040 19760 22092
rect 19892 21972 19944 22024
rect 23756 22108 23808 22160
rect 21088 22040 21140 22092
rect 27988 22040 28040 22092
rect 20352 21904 20404 21956
rect 6920 21836 6972 21888
rect 10232 21836 10284 21888
rect 10324 21836 10376 21888
rect 12624 21836 12676 21888
rect 12808 21836 12860 21888
rect 14188 21836 14240 21888
rect 16856 21836 16908 21888
rect 18880 21836 18932 21888
rect 19248 21836 19300 21888
rect 22468 21972 22520 22024
rect 25412 21972 25464 22024
rect 21456 21904 21508 21956
rect 23664 21904 23716 21956
rect 23940 21904 23992 21956
rect 31300 21904 31352 21956
rect 20536 21836 20588 21888
rect 23572 21836 23624 21888
rect 24124 21836 24176 21888
rect 25688 21836 25740 21888
rect 4193 21734 4245 21786
rect 4257 21734 4309 21786
rect 4321 21734 4373 21786
rect 4385 21734 4437 21786
rect 4449 21734 4501 21786
rect 11783 21734 11835 21786
rect 11847 21734 11899 21786
rect 11911 21734 11963 21786
rect 11975 21734 12027 21786
rect 12039 21734 12091 21786
rect 19373 21734 19425 21786
rect 19437 21734 19489 21786
rect 19501 21734 19553 21786
rect 19565 21734 19617 21786
rect 19629 21734 19681 21786
rect 26963 21734 27015 21786
rect 27027 21734 27079 21786
rect 27091 21734 27143 21786
rect 27155 21734 27207 21786
rect 27219 21734 27271 21786
rect 2504 21632 2556 21684
rect 2872 21632 2924 21684
rect 2136 21471 2188 21480
rect 2136 21437 2145 21471
rect 2145 21437 2179 21471
rect 2179 21437 2188 21471
rect 2136 21428 2188 21437
rect 3056 21496 3108 21548
rect 3240 21471 3292 21480
rect 1400 21360 1452 21412
rect 2780 21360 2832 21412
rect 1492 21292 1544 21344
rect 3240 21437 3249 21471
rect 3249 21437 3283 21471
rect 3283 21437 3292 21471
rect 3240 21428 3292 21437
rect 3976 21471 4028 21480
rect 3976 21437 3985 21471
rect 3985 21437 4019 21471
rect 4019 21437 4028 21471
rect 3976 21428 4028 21437
rect 5632 21471 5684 21480
rect 5632 21437 5641 21471
rect 5641 21437 5675 21471
rect 5675 21437 5684 21471
rect 5632 21428 5684 21437
rect 3700 21335 3752 21344
rect 3700 21301 3715 21335
rect 3715 21301 3749 21335
rect 3749 21301 3752 21335
rect 3700 21292 3752 21301
rect 5080 21335 5132 21344
rect 5080 21301 5089 21335
rect 5089 21301 5123 21335
rect 5123 21301 5132 21335
rect 5080 21292 5132 21301
rect 6092 21564 6144 21616
rect 6460 21632 6512 21684
rect 6920 21675 6972 21684
rect 6920 21641 6929 21675
rect 6929 21641 6963 21675
rect 6963 21641 6972 21675
rect 6920 21632 6972 21641
rect 6920 21496 6972 21548
rect 8208 21607 8260 21616
rect 8208 21573 8217 21607
rect 8217 21573 8251 21607
rect 8251 21573 8260 21607
rect 8208 21564 8260 21573
rect 8576 21564 8628 21616
rect 9404 21632 9456 21684
rect 10324 21607 10376 21616
rect 10324 21573 10333 21607
rect 10333 21573 10367 21607
rect 10367 21573 10376 21607
rect 10324 21564 10376 21573
rect 7288 21428 7340 21480
rect 11428 21539 11480 21548
rect 11428 21505 11440 21539
rect 11440 21505 11474 21539
rect 11474 21505 11480 21539
rect 12716 21632 12768 21684
rect 12808 21675 12860 21684
rect 12808 21641 12817 21675
rect 12817 21641 12851 21675
rect 12851 21641 12860 21675
rect 12808 21632 12860 21641
rect 14556 21632 14608 21684
rect 17132 21632 17184 21684
rect 19064 21564 19116 21616
rect 21088 21632 21140 21684
rect 22376 21632 22428 21684
rect 11428 21496 11480 21505
rect 13820 21496 13872 21548
rect 8576 21471 8628 21480
rect 8576 21437 8585 21471
rect 8585 21437 8619 21471
rect 8619 21437 8628 21471
rect 8576 21428 8628 21437
rect 8852 21428 8904 21480
rect 10416 21428 10468 21480
rect 10692 21428 10744 21480
rect 10784 21471 10836 21480
rect 10784 21437 10793 21471
rect 10793 21437 10827 21471
rect 10827 21437 10836 21471
rect 10784 21428 10836 21437
rect 10876 21428 10928 21480
rect 11060 21428 11112 21480
rect 11244 21428 11296 21480
rect 11704 21471 11756 21480
rect 11704 21437 11713 21471
rect 11713 21437 11747 21471
rect 11747 21437 11756 21471
rect 11704 21428 11756 21437
rect 13360 21471 13412 21480
rect 13360 21437 13369 21471
rect 13369 21437 13403 21471
rect 13403 21437 13412 21471
rect 13360 21428 13412 21437
rect 14280 21471 14332 21480
rect 14280 21437 14289 21471
rect 14289 21437 14323 21471
rect 14323 21437 14332 21471
rect 14280 21428 14332 21437
rect 14556 21471 14608 21480
rect 14556 21437 14565 21471
rect 14565 21437 14599 21471
rect 14599 21437 14608 21471
rect 14556 21428 14608 21437
rect 14648 21428 14700 21480
rect 16856 21539 16908 21548
rect 16856 21505 16865 21539
rect 16865 21505 16899 21539
rect 16899 21505 16908 21539
rect 16856 21496 16908 21505
rect 19248 21496 19300 21548
rect 19616 21496 19668 21548
rect 6644 21403 6696 21412
rect 6644 21369 6653 21403
rect 6653 21369 6687 21403
rect 6687 21369 6696 21403
rect 6644 21360 6696 21369
rect 8484 21360 8536 21412
rect 9312 21360 9364 21412
rect 16396 21360 16448 21412
rect 8300 21292 8352 21344
rect 8668 21292 8720 21344
rect 11336 21292 11388 21344
rect 11612 21292 11664 21344
rect 12348 21292 12400 21344
rect 13728 21335 13780 21344
rect 13728 21301 13737 21335
rect 13737 21301 13771 21335
rect 13771 21301 13780 21335
rect 13728 21292 13780 21301
rect 16120 21335 16172 21344
rect 16120 21301 16129 21335
rect 16129 21301 16163 21335
rect 16163 21301 16172 21335
rect 16120 21292 16172 21301
rect 18788 21428 18840 21480
rect 18880 21471 18932 21480
rect 18880 21437 18889 21471
rect 18889 21437 18923 21471
rect 18923 21437 18932 21471
rect 18880 21428 18932 21437
rect 16764 21403 16816 21412
rect 16764 21369 16773 21403
rect 16773 21369 16807 21403
rect 16807 21369 16816 21403
rect 16764 21360 16816 21369
rect 20720 21428 20772 21480
rect 18972 21292 19024 21344
rect 20536 21292 20588 21344
rect 21272 21292 21324 21344
rect 21456 21539 21508 21548
rect 21456 21505 21465 21539
rect 21465 21505 21499 21539
rect 21499 21505 21508 21539
rect 21456 21496 21508 21505
rect 22008 21496 22060 21548
rect 22468 21539 22520 21548
rect 22468 21505 22477 21539
rect 22477 21505 22511 21539
rect 22511 21505 22520 21539
rect 22468 21496 22520 21505
rect 22192 21471 22244 21480
rect 22192 21437 22201 21471
rect 22201 21437 22235 21471
rect 22235 21437 22244 21471
rect 22192 21428 22244 21437
rect 22284 21471 22336 21480
rect 22284 21437 22318 21471
rect 22318 21437 22336 21471
rect 22284 21428 22336 21437
rect 23204 21471 23256 21480
rect 23204 21437 23213 21471
rect 23213 21437 23247 21471
rect 23247 21437 23256 21471
rect 23204 21428 23256 21437
rect 23572 21471 23624 21480
rect 23572 21437 23581 21471
rect 23581 21437 23615 21471
rect 23615 21437 23624 21471
rect 23572 21428 23624 21437
rect 23940 21564 23992 21616
rect 25504 21564 25556 21616
rect 29000 21564 29052 21616
rect 24492 21539 24544 21548
rect 24492 21505 24501 21539
rect 24501 21505 24535 21539
rect 24535 21505 24544 21539
rect 24492 21496 24544 21505
rect 24584 21496 24636 21548
rect 25412 21496 25464 21548
rect 25780 21496 25832 21548
rect 23940 21428 23992 21480
rect 22744 21292 22796 21344
rect 22928 21292 22980 21344
rect 23020 21292 23072 21344
rect 24768 21471 24820 21480
rect 24768 21437 24777 21471
rect 24777 21437 24811 21471
rect 24811 21437 24820 21471
rect 24768 21428 24820 21437
rect 25688 21428 25740 21480
rect 27804 21428 27856 21480
rect 28356 21496 28408 21548
rect 25044 21292 25096 21344
rect 25688 21292 25740 21344
rect 28080 21360 28132 21412
rect 30380 21428 30432 21480
rect 30564 21471 30616 21480
rect 30564 21437 30573 21471
rect 30573 21437 30607 21471
rect 30607 21437 30616 21471
rect 30564 21428 30616 21437
rect 27436 21292 27488 21344
rect 28448 21292 28500 21344
rect 30288 21360 30340 21412
rect 29736 21335 29788 21344
rect 29736 21301 29745 21335
rect 29745 21301 29779 21335
rect 29779 21301 29788 21335
rect 29736 21292 29788 21301
rect 30104 21292 30156 21344
rect 7988 21190 8040 21242
rect 8052 21190 8104 21242
rect 8116 21190 8168 21242
rect 8180 21190 8232 21242
rect 8244 21190 8296 21242
rect 15578 21190 15630 21242
rect 15642 21190 15694 21242
rect 15706 21190 15758 21242
rect 15770 21190 15822 21242
rect 15834 21190 15886 21242
rect 23168 21190 23220 21242
rect 23232 21190 23284 21242
rect 23296 21190 23348 21242
rect 23360 21190 23412 21242
rect 23424 21190 23476 21242
rect 30758 21190 30810 21242
rect 30822 21190 30874 21242
rect 30886 21190 30938 21242
rect 30950 21190 31002 21242
rect 31014 21190 31066 21242
rect 848 21131 900 21140
rect 848 21097 857 21131
rect 857 21097 891 21131
rect 891 21097 900 21131
rect 848 21088 900 21097
rect 3700 21088 3752 21140
rect 6092 21088 6144 21140
rect 6644 21088 6696 21140
rect 5908 21020 5960 21072
rect 7840 21020 7892 21072
rect 1492 20884 1544 20936
rect 1768 20884 1820 20936
rect 1860 20927 1912 20936
rect 1860 20893 1869 20927
rect 1869 20893 1903 20927
rect 1903 20893 1912 20927
rect 1860 20884 1912 20893
rect 3240 20884 3292 20936
rect 3516 20884 3568 20936
rect 3700 20927 3752 20936
rect 3700 20893 3702 20927
rect 3702 20893 3752 20927
rect 3700 20884 3752 20893
rect 3792 20927 3844 20936
rect 3792 20893 3804 20927
rect 3804 20893 3838 20927
rect 3838 20893 3844 20927
rect 3792 20884 3844 20893
rect 4068 20927 4120 20936
rect 4068 20893 4077 20927
rect 4077 20893 4111 20927
rect 4111 20893 4120 20927
rect 4068 20884 4120 20893
rect 5816 20927 5868 20936
rect 5816 20893 5825 20927
rect 5825 20893 5859 20927
rect 5859 20893 5868 20927
rect 5816 20884 5868 20893
rect 7748 20952 7800 21004
rect 10968 21020 11020 21072
rect 8668 20952 8720 21004
rect 6552 20927 6604 20936
rect 6552 20893 6561 20927
rect 6561 20893 6595 20927
rect 6595 20893 6604 20927
rect 6552 20884 6604 20893
rect 5540 20748 5592 20800
rect 6460 20748 6512 20800
rect 7656 20748 7708 20800
rect 8760 20927 8812 20936
rect 8760 20893 8769 20927
rect 8769 20893 8803 20927
rect 8803 20893 8812 20927
rect 8760 20884 8812 20893
rect 8852 20884 8904 20936
rect 10508 20952 10560 21004
rect 8944 20748 8996 20800
rect 11060 20884 11112 20936
rect 11520 20927 11572 20936
rect 11520 20893 11522 20927
rect 11522 20893 11572 20927
rect 10876 20816 10928 20868
rect 11520 20884 11572 20893
rect 16120 21088 16172 21140
rect 17960 21088 18012 21140
rect 21272 21088 21324 21140
rect 22192 21088 22244 21140
rect 14004 21020 14056 21072
rect 14188 21020 14240 21072
rect 15568 21020 15620 21072
rect 13912 20952 13964 21004
rect 14372 20995 14424 21004
rect 14372 20961 14381 20995
rect 14381 20961 14415 20995
rect 14415 20961 14424 20995
rect 14372 20952 14424 20961
rect 15936 21020 15988 21072
rect 22836 21020 22888 21072
rect 25044 21020 25096 21072
rect 25872 21020 25924 21072
rect 13820 20884 13872 20936
rect 16212 20952 16264 21004
rect 11428 20748 11480 20800
rect 12256 20748 12308 20800
rect 16304 20884 16356 20936
rect 20628 20952 20680 21004
rect 14280 20816 14332 20868
rect 18880 20884 18932 20936
rect 16764 20748 16816 20800
rect 17224 20748 17276 20800
rect 19248 20927 19300 20936
rect 19248 20893 19257 20927
rect 19257 20893 19291 20927
rect 19291 20893 19300 20927
rect 23112 20952 23164 21004
rect 19248 20884 19300 20893
rect 21180 20884 21232 20936
rect 25136 20952 25188 21004
rect 22652 20748 22704 20800
rect 22744 20748 22796 20800
rect 24492 20748 24544 20800
rect 27436 20952 27488 21004
rect 26700 20927 26752 20936
rect 26700 20893 26709 20927
rect 26709 20893 26743 20927
rect 26743 20893 26752 20927
rect 26700 20884 26752 20893
rect 26792 20884 26844 20936
rect 26884 20884 26936 20936
rect 29460 20884 29512 20936
rect 29644 20884 29696 20936
rect 26884 20748 26936 20800
rect 4193 20646 4245 20698
rect 4257 20646 4309 20698
rect 4321 20646 4373 20698
rect 4385 20646 4437 20698
rect 4449 20646 4501 20698
rect 11783 20646 11835 20698
rect 11847 20646 11899 20698
rect 11911 20646 11963 20698
rect 11975 20646 12027 20698
rect 12039 20646 12091 20698
rect 19373 20646 19425 20698
rect 19437 20646 19489 20698
rect 19501 20646 19553 20698
rect 19565 20646 19617 20698
rect 19629 20646 19681 20698
rect 26963 20646 27015 20698
rect 27027 20646 27079 20698
rect 27091 20646 27143 20698
rect 27155 20646 27207 20698
rect 27219 20646 27271 20698
rect 1768 20544 1820 20596
rect 3240 20408 3292 20460
rect 1216 20340 1268 20392
rect 1676 20383 1728 20392
rect 1676 20349 1685 20383
rect 1685 20349 1719 20383
rect 1719 20349 1728 20383
rect 1676 20340 1728 20349
rect 2780 20340 2832 20392
rect 6644 20544 6696 20596
rect 6920 20544 6972 20596
rect 6000 20476 6052 20528
rect 7748 20476 7800 20528
rect 10508 20544 10560 20596
rect 10876 20544 10928 20596
rect 10968 20544 11020 20596
rect 14188 20544 14240 20596
rect 14372 20544 14424 20596
rect 15108 20544 15160 20596
rect 15200 20544 15252 20596
rect 16396 20544 16448 20596
rect 21364 20544 21416 20596
rect 21548 20544 21600 20596
rect 5080 20408 5132 20460
rect 6460 20451 6512 20460
rect 6460 20417 6462 20451
rect 6462 20417 6512 20451
rect 6460 20408 6512 20417
rect 4712 20340 4764 20392
rect 4896 20340 4948 20392
rect 5448 20340 5500 20392
rect 6828 20383 6880 20392
rect 6828 20349 6837 20383
rect 6837 20349 6871 20383
rect 6871 20349 6880 20383
rect 6828 20340 6880 20349
rect 7104 20340 7156 20392
rect 8392 20383 8444 20392
rect 8392 20349 8401 20383
rect 8401 20349 8435 20383
rect 8435 20349 8444 20383
rect 8392 20340 8444 20349
rect 3976 20272 4028 20324
rect 1400 20247 1452 20256
rect 1400 20213 1415 20247
rect 1415 20213 1449 20247
rect 1449 20213 1452 20247
rect 1400 20204 1452 20213
rect 1768 20204 1820 20256
rect 4252 20204 4304 20256
rect 4620 20204 4672 20256
rect 4896 20204 4948 20256
rect 9496 20340 9548 20392
rect 10232 20340 10284 20392
rect 10968 20340 11020 20392
rect 11244 20340 11296 20392
rect 8668 20204 8720 20256
rect 11612 20204 11664 20256
rect 13268 20204 13320 20256
rect 15936 20408 15988 20460
rect 19248 20451 19300 20460
rect 19248 20417 19257 20451
rect 19257 20417 19291 20451
rect 19291 20417 19300 20451
rect 19248 20408 19300 20417
rect 21180 20408 21232 20460
rect 27068 20544 27120 20596
rect 27436 20544 27488 20596
rect 29368 20544 29420 20596
rect 23112 20476 23164 20528
rect 14280 20383 14332 20392
rect 14280 20349 14296 20383
rect 14296 20349 14330 20383
rect 14330 20349 14332 20383
rect 14280 20340 14332 20349
rect 16396 20383 16448 20392
rect 16396 20349 16405 20383
rect 16405 20349 16439 20383
rect 16439 20349 16448 20383
rect 16396 20340 16448 20349
rect 20628 20340 20680 20392
rect 14832 20272 14884 20324
rect 16212 20272 16264 20324
rect 17960 20315 18012 20324
rect 17960 20281 17969 20315
rect 17969 20281 18003 20315
rect 18003 20281 18012 20315
rect 17960 20272 18012 20281
rect 15384 20204 15436 20256
rect 17500 20247 17552 20256
rect 17500 20213 17509 20247
rect 17509 20213 17543 20247
rect 17543 20213 17552 20247
rect 17500 20204 17552 20213
rect 18788 20315 18840 20324
rect 18788 20281 18797 20315
rect 18797 20281 18831 20315
rect 18831 20281 18840 20315
rect 18788 20272 18840 20281
rect 25136 20340 25188 20392
rect 25688 20340 25740 20392
rect 26424 20408 26476 20460
rect 26608 20408 26660 20460
rect 27068 20383 27120 20392
rect 18696 20204 18748 20256
rect 22008 20204 22060 20256
rect 23112 20272 23164 20324
rect 23480 20272 23532 20324
rect 24400 20272 24452 20324
rect 27068 20349 27070 20383
rect 27070 20349 27120 20383
rect 27068 20340 27120 20349
rect 26608 20272 26660 20324
rect 22468 20204 22520 20256
rect 24768 20204 24820 20256
rect 26240 20247 26292 20256
rect 26240 20213 26249 20247
rect 26249 20213 26283 20247
rect 26283 20213 26292 20247
rect 26240 20204 26292 20213
rect 26516 20204 26568 20256
rect 29092 20383 29144 20392
rect 29092 20349 29101 20383
rect 29101 20349 29135 20383
rect 29135 20349 29144 20383
rect 29092 20340 29144 20349
rect 29276 20383 29328 20392
rect 29276 20349 29285 20383
rect 29285 20349 29319 20383
rect 29319 20349 29328 20383
rect 29276 20340 29328 20349
rect 29368 20383 29420 20392
rect 29368 20349 29377 20383
rect 29377 20349 29411 20383
rect 29411 20349 29420 20383
rect 29368 20340 29420 20349
rect 29000 20204 29052 20256
rect 29828 20204 29880 20256
rect 30196 20204 30248 20256
rect 31208 20204 31260 20256
rect 7988 20102 8040 20154
rect 8052 20102 8104 20154
rect 8116 20102 8168 20154
rect 8180 20102 8232 20154
rect 8244 20102 8296 20154
rect 15578 20102 15630 20154
rect 15642 20102 15694 20154
rect 15706 20102 15758 20154
rect 15770 20102 15822 20154
rect 15834 20102 15886 20154
rect 23168 20102 23220 20154
rect 23232 20102 23284 20154
rect 23296 20102 23348 20154
rect 23360 20102 23412 20154
rect 23424 20102 23476 20154
rect 30758 20102 30810 20154
rect 30822 20102 30874 20154
rect 30886 20102 30938 20154
rect 30950 20102 31002 20154
rect 31014 20102 31066 20154
rect 1768 20000 1820 20052
rect 3792 20000 3844 20052
rect 4252 20000 4304 20052
rect 7840 20043 7892 20052
rect 7840 20009 7849 20043
rect 7849 20009 7883 20043
rect 7883 20009 7892 20043
rect 7840 20000 7892 20009
rect 9588 20000 9640 20052
rect 664 19864 716 19916
rect 1216 19864 1268 19916
rect 2872 19864 2924 19916
rect 1860 19839 1912 19848
rect 1860 19805 1869 19839
rect 1869 19805 1903 19839
rect 1903 19805 1912 19839
rect 1860 19796 1912 19805
rect 3516 19839 3568 19848
rect 3516 19805 3525 19839
rect 3525 19805 3559 19839
rect 3559 19805 3568 19839
rect 3516 19796 3568 19805
rect 3700 19796 3752 19848
rect 3884 19839 3936 19848
rect 3884 19805 3886 19839
rect 3886 19805 3936 19839
rect 3884 19796 3936 19805
rect 4712 19796 4764 19848
rect 5080 19796 5132 19848
rect 5172 19796 5224 19848
rect 5816 19839 5868 19848
rect 5816 19805 5825 19839
rect 5825 19805 5859 19839
rect 5859 19805 5868 19839
rect 5816 19796 5868 19805
rect 6184 19839 6236 19848
rect 6184 19805 6186 19839
rect 6186 19805 6236 19839
rect 6184 19796 6236 19805
rect 6920 19864 6972 19916
rect 8392 19932 8444 19984
rect 8208 19907 8260 19916
rect 8208 19873 8217 19907
rect 8217 19873 8251 19907
rect 8251 19873 8260 19907
rect 8208 19864 8260 19873
rect 6552 19839 6604 19848
rect 6552 19805 6561 19839
rect 6561 19805 6595 19839
rect 6595 19805 6604 19839
rect 6552 19796 6604 19805
rect 7656 19796 7708 19848
rect 8392 19839 8444 19848
rect 8392 19805 8401 19839
rect 8401 19805 8435 19839
rect 8435 19805 8444 19839
rect 8392 19796 8444 19805
rect 9036 19864 9088 19916
rect 11244 20000 11296 20052
rect 11520 20000 11572 20052
rect 13636 20000 13688 20052
rect 13912 20043 13964 20052
rect 13912 20009 13921 20043
rect 13921 20009 13955 20043
rect 13955 20009 13964 20043
rect 13912 20000 13964 20009
rect 14832 20000 14884 20052
rect 10876 19864 10928 19916
rect 11244 19886 11296 19938
rect 16580 20000 16632 20052
rect 22192 20000 22244 20052
rect 22836 20000 22888 20052
rect 8852 19839 8904 19848
rect 8852 19805 8854 19839
rect 8854 19805 8904 19839
rect 8852 19796 8904 19805
rect 8944 19839 8996 19848
rect 8944 19805 8956 19839
rect 8956 19805 8990 19839
rect 8990 19805 8996 19839
rect 8944 19796 8996 19805
rect 9220 19839 9272 19848
rect 9220 19805 9229 19839
rect 9229 19805 9263 19839
rect 9263 19805 9272 19839
rect 9220 19796 9272 19805
rect 848 19703 900 19712
rect 848 19669 857 19703
rect 857 19669 891 19703
rect 891 19669 900 19703
rect 848 19660 900 19669
rect 5448 19660 5500 19712
rect 7748 19660 7800 19712
rect 9956 19728 10008 19780
rect 8484 19660 8536 19712
rect 10324 19660 10376 19712
rect 11428 19796 11480 19848
rect 16028 19864 16080 19916
rect 16304 19907 16356 19916
rect 16304 19873 16313 19907
rect 16313 19873 16347 19907
rect 16347 19873 16356 19907
rect 16304 19864 16356 19873
rect 12256 19796 12308 19848
rect 12532 19839 12584 19848
rect 12532 19805 12544 19839
rect 12544 19805 12578 19839
rect 12578 19805 12584 19839
rect 12532 19796 12584 19805
rect 14188 19796 14240 19848
rect 14464 19796 14516 19848
rect 16212 19839 16264 19848
rect 16212 19805 16221 19839
rect 16221 19805 16255 19839
rect 16255 19805 16264 19839
rect 16212 19796 16264 19805
rect 17500 19864 17552 19916
rect 17960 19864 18012 19916
rect 18788 19864 18840 19916
rect 20628 19864 20680 19916
rect 21548 19907 21600 19916
rect 21548 19873 21557 19907
rect 21557 19873 21591 19907
rect 21591 19873 21600 19907
rect 21548 19864 21600 19873
rect 22744 19932 22796 19984
rect 23940 20000 23992 20052
rect 24768 20000 24820 20052
rect 26516 20000 26568 20052
rect 27804 20043 27856 20052
rect 27804 20009 27813 20043
rect 27813 20009 27847 20043
rect 27847 20009 27856 20043
rect 27804 20000 27856 20009
rect 30196 20043 30248 20052
rect 30196 20009 30205 20043
rect 30205 20009 30239 20043
rect 30239 20009 30248 20043
rect 30196 20000 30248 20009
rect 16948 19839 17000 19848
rect 16948 19805 16957 19839
rect 16957 19805 16991 19839
rect 16991 19805 17000 19839
rect 16948 19796 17000 19805
rect 20076 19796 20128 19848
rect 16672 19728 16724 19780
rect 20720 19728 20772 19780
rect 23572 19864 23624 19916
rect 22468 19839 22520 19848
rect 22468 19805 22477 19839
rect 22477 19805 22511 19839
rect 22511 19805 22520 19839
rect 22468 19796 22520 19805
rect 23112 19796 23164 19848
rect 23940 19864 23992 19916
rect 25136 19864 25188 19916
rect 24676 19839 24728 19848
rect 24676 19805 24685 19839
rect 24685 19805 24719 19839
rect 24719 19805 24728 19839
rect 24676 19796 24728 19805
rect 26792 19796 26844 19848
rect 27620 19796 27672 19848
rect 28540 19796 28592 19848
rect 29000 19796 29052 19848
rect 29552 19796 29604 19848
rect 14740 19660 14792 19712
rect 15200 19660 15252 19712
rect 15844 19703 15896 19712
rect 15844 19669 15853 19703
rect 15853 19669 15887 19703
rect 15887 19669 15896 19703
rect 15844 19660 15896 19669
rect 18604 19660 18656 19712
rect 19800 19660 19852 19712
rect 20444 19660 20496 19712
rect 22100 19660 22152 19712
rect 22468 19660 22520 19712
rect 26700 19660 26752 19712
rect 29184 19660 29236 19712
rect 30288 19660 30340 19712
rect 4193 19558 4245 19610
rect 4257 19558 4309 19610
rect 4321 19558 4373 19610
rect 4385 19558 4437 19610
rect 4449 19558 4501 19610
rect 11783 19558 11835 19610
rect 11847 19558 11899 19610
rect 11911 19558 11963 19610
rect 11975 19558 12027 19610
rect 12039 19558 12091 19610
rect 19373 19558 19425 19610
rect 19437 19558 19489 19610
rect 19501 19558 19553 19610
rect 19565 19558 19617 19610
rect 19629 19558 19681 19610
rect 26963 19558 27015 19610
rect 27027 19558 27079 19610
rect 27091 19558 27143 19610
rect 27155 19558 27207 19610
rect 27219 19558 27271 19610
rect 848 19456 900 19508
rect 2780 19320 2832 19372
rect 3976 19456 4028 19508
rect 3700 19388 3752 19440
rect 4252 19388 4304 19440
rect 4620 19456 4672 19508
rect 6184 19456 6236 19508
rect 7104 19499 7156 19508
rect 7104 19465 7113 19499
rect 7113 19465 7147 19499
rect 7147 19465 7156 19499
rect 7104 19456 7156 19465
rect 7564 19456 7616 19508
rect 8208 19456 8260 19508
rect 8668 19456 8720 19508
rect 8852 19456 8904 19508
rect 1216 19252 1268 19304
rect 2504 19252 2556 19304
rect 3056 19295 3108 19304
rect 3056 19261 3065 19295
rect 3065 19261 3099 19295
rect 3099 19261 3108 19295
rect 3056 19252 3108 19261
rect 3148 19252 3200 19304
rect 2964 19184 3016 19236
rect 3792 19252 3844 19304
rect 3884 19295 3936 19304
rect 3884 19261 3893 19295
rect 3893 19261 3927 19295
rect 3927 19261 3936 19295
rect 3884 19252 3936 19261
rect 4344 19252 4396 19304
rect 5080 19320 5132 19372
rect 5540 19320 5592 19372
rect 6460 19320 6512 19372
rect 6920 19320 6972 19372
rect 8208 19320 8260 19372
rect 6276 19252 6328 19304
rect 7656 19295 7708 19304
rect 7656 19261 7665 19295
rect 7665 19261 7699 19295
rect 7699 19261 7708 19295
rect 7656 19252 7708 19261
rect 7748 19252 7800 19304
rect 8576 19320 8628 19372
rect 4252 19227 4304 19236
rect 4252 19193 4261 19227
rect 4261 19193 4295 19227
rect 4295 19193 4304 19227
rect 4252 19184 4304 19193
rect 4620 19184 4672 19236
rect 4712 19184 4764 19236
rect 4804 19227 4856 19236
rect 4804 19193 4813 19227
rect 4813 19193 4847 19227
rect 4847 19193 4856 19227
rect 4804 19184 4856 19193
rect 4988 19184 5040 19236
rect 5356 19184 5408 19236
rect 1768 19116 1820 19168
rect 4068 19116 4120 19168
rect 4160 19116 4212 19168
rect 5908 19116 5960 19168
rect 6000 19116 6052 19168
rect 7472 19159 7524 19168
rect 7472 19125 7481 19159
rect 7481 19125 7515 19159
rect 7515 19125 7524 19159
rect 7472 19116 7524 19125
rect 7840 19227 7892 19236
rect 7840 19193 7849 19227
rect 7849 19193 7883 19227
rect 7883 19193 7892 19227
rect 7840 19184 7892 19193
rect 10232 19499 10284 19508
rect 10232 19465 10241 19499
rect 10241 19465 10275 19499
rect 10275 19465 10284 19499
rect 10232 19456 10284 19465
rect 10324 19456 10376 19508
rect 14648 19456 14700 19508
rect 15384 19499 15436 19508
rect 15384 19465 15393 19499
rect 15393 19465 15427 19499
rect 15427 19465 15436 19499
rect 15384 19456 15436 19465
rect 20076 19499 20128 19508
rect 20076 19465 20085 19499
rect 20085 19465 20119 19499
rect 20119 19465 20128 19499
rect 20076 19456 20128 19465
rect 20628 19456 20680 19508
rect 13268 19388 13320 19440
rect 10784 19320 10836 19372
rect 15844 19320 15896 19372
rect 10692 19295 10744 19304
rect 10692 19261 10701 19295
rect 10701 19261 10735 19295
rect 10735 19261 10744 19295
rect 10692 19252 10744 19261
rect 11152 19252 11204 19304
rect 11244 19295 11296 19304
rect 11244 19261 11253 19295
rect 11253 19261 11287 19295
rect 11287 19261 11296 19295
rect 11244 19252 11296 19261
rect 12256 19252 12308 19304
rect 13544 19295 13596 19304
rect 13544 19261 13553 19295
rect 13553 19261 13587 19295
rect 13587 19261 13596 19295
rect 13544 19252 13596 19261
rect 13636 19252 13688 19304
rect 14096 19252 14148 19304
rect 15936 19295 15988 19304
rect 15936 19261 15945 19295
rect 15945 19261 15979 19295
rect 15979 19261 15988 19295
rect 15936 19252 15988 19261
rect 16028 19252 16080 19304
rect 24676 19456 24728 19508
rect 22192 19388 22244 19440
rect 23664 19388 23716 19440
rect 18696 19363 18748 19372
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 8760 19116 8812 19168
rect 8852 19159 8904 19168
rect 8852 19125 8867 19159
rect 8867 19125 8901 19159
rect 8901 19125 8904 19159
rect 17040 19184 17092 19236
rect 17960 19227 18012 19236
rect 17960 19193 17969 19227
rect 17969 19193 18003 19227
rect 18003 19193 18012 19227
rect 17960 19184 18012 19193
rect 18236 19295 18288 19304
rect 18236 19261 18245 19295
rect 18245 19261 18279 19295
rect 18279 19261 18288 19295
rect 18236 19252 18288 19261
rect 18328 19252 18380 19304
rect 19248 19252 19300 19304
rect 20444 19295 20496 19304
rect 20444 19261 20453 19295
rect 20453 19261 20487 19295
rect 20487 19261 20496 19295
rect 20444 19252 20496 19261
rect 20720 19363 20772 19372
rect 20720 19329 20729 19363
rect 20729 19329 20763 19363
rect 20763 19329 20772 19363
rect 20720 19320 20772 19329
rect 21088 19320 21140 19372
rect 21916 19320 21968 19372
rect 22100 19320 22152 19372
rect 29368 19388 29420 19440
rect 29920 19320 29972 19372
rect 8852 19116 8904 19125
rect 11520 19116 11572 19168
rect 12440 19116 12492 19168
rect 14004 19116 14056 19168
rect 18512 19116 18564 19168
rect 21640 19116 21692 19168
rect 23572 19252 23624 19304
rect 22376 19184 22428 19236
rect 22744 19184 22796 19236
rect 22928 19184 22980 19236
rect 24032 19227 24084 19236
rect 24032 19193 24041 19227
rect 24041 19193 24075 19227
rect 24075 19193 24084 19227
rect 24032 19184 24084 19193
rect 24400 19252 24452 19304
rect 25596 19252 25648 19304
rect 26976 19252 27028 19304
rect 28540 19184 28592 19236
rect 24124 19159 24176 19168
rect 24124 19125 24133 19159
rect 24133 19125 24167 19159
rect 24167 19125 24176 19159
rect 24124 19116 24176 19125
rect 24492 19116 24544 19168
rect 24952 19159 25004 19168
rect 24952 19125 24967 19159
rect 24967 19125 25001 19159
rect 25001 19125 25004 19159
rect 24952 19116 25004 19125
rect 25320 19116 25372 19168
rect 29276 19252 29328 19304
rect 30656 19320 30708 19372
rect 29092 19227 29144 19236
rect 29092 19193 29101 19227
rect 29101 19193 29135 19227
rect 29135 19193 29144 19227
rect 29092 19184 29144 19193
rect 30012 19184 30064 19236
rect 30472 19184 30524 19236
rect 30288 19159 30340 19168
rect 30288 19125 30297 19159
rect 30297 19125 30331 19159
rect 30331 19125 30340 19159
rect 30288 19116 30340 19125
rect 7988 19014 8040 19066
rect 8052 19014 8104 19066
rect 8116 19014 8168 19066
rect 8180 19014 8232 19066
rect 8244 19014 8296 19066
rect 15578 19014 15630 19066
rect 15642 19014 15694 19066
rect 15706 19014 15758 19066
rect 15770 19014 15822 19066
rect 15834 19014 15886 19066
rect 23168 19014 23220 19066
rect 23232 19014 23284 19066
rect 23296 19014 23348 19066
rect 23360 19014 23412 19066
rect 23424 19014 23476 19066
rect 30758 19014 30810 19066
rect 30822 19014 30874 19066
rect 30886 19014 30938 19066
rect 30950 19014 31002 19066
rect 31014 19014 31066 19066
rect 1584 18912 1636 18964
rect 1308 18751 1360 18760
rect 1308 18717 1317 18751
rect 1317 18717 1351 18751
rect 1351 18717 1360 18751
rect 1308 18708 1360 18717
rect 1952 18708 2004 18760
rect 3700 18776 3752 18828
rect 3976 18776 4028 18828
rect 5540 18912 5592 18964
rect 5908 18912 5960 18964
rect 6184 18912 6236 18964
rect 7472 18912 7524 18964
rect 9864 18912 9916 18964
rect 13912 18912 13964 18964
rect 3424 18708 3476 18760
rect 4160 18708 4212 18760
rect 4896 18819 4948 18828
rect 4896 18785 4905 18819
rect 4905 18785 4939 18819
rect 4939 18785 4948 18819
rect 4896 18776 4948 18785
rect 3516 18640 3568 18692
rect 4344 18640 4396 18692
rect 4528 18640 4580 18692
rect 4620 18640 4672 18692
rect 4712 18683 4764 18692
rect 4712 18649 4721 18683
rect 4721 18649 4755 18683
rect 4755 18649 4764 18683
rect 4712 18640 4764 18649
rect 5448 18819 5500 18828
rect 5448 18785 5457 18819
rect 5457 18785 5491 18819
rect 5491 18785 5500 18819
rect 5448 18776 5500 18785
rect 1032 18615 1084 18624
rect 1032 18581 1041 18615
rect 1041 18581 1075 18615
rect 1075 18581 1084 18615
rect 1032 18572 1084 18581
rect 3332 18615 3384 18624
rect 3332 18581 3341 18615
rect 3341 18581 3375 18615
rect 3375 18581 3384 18615
rect 3332 18572 3384 18581
rect 3700 18615 3752 18624
rect 3700 18581 3709 18615
rect 3709 18581 3743 18615
rect 3743 18581 3752 18615
rect 3700 18572 3752 18581
rect 4804 18572 4856 18624
rect 8576 18844 8628 18896
rect 8668 18844 8720 18896
rect 5908 18819 5960 18828
rect 5908 18785 5917 18819
rect 5917 18785 5951 18819
rect 5951 18785 5960 18819
rect 5908 18776 5960 18785
rect 6460 18776 6512 18828
rect 10784 18887 10836 18896
rect 10784 18853 10793 18887
rect 10793 18853 10827 18887
rect 10827 18853 10836 18887
rect 10784 18844 10836 18853
rect 11612 18844 11664 18896
rect 16396 18912 16448 18964
rect 6184 18708 6236 18760
rect 6368 18753 6420 18760
rect 6368 18719 6380 18753
rect 6380 18719 6414 18753
rect 6414 18719 6420 18753
rect 6368 18708 6420 18719
rect 7472 18708 7524 18760
rect 7748 18708 7800 18760
rect 8300 18640 8352 18692
rect 8208 18572 8260 18624
rect 8484 18615 8536 18624
rect 8484 18581 8493 18615
rect 8493 18581 8527 18615
rect 8527 18581 8536 18615
rect 8484 18572 8536 18581
rect 8576 18572 8628 18624
rect 9404 18751 9456 18760
rect 9404 18717 9413 18751
rect 9413 18717 9447 18751
rect 9447 18717 9456 18751
rect 9404 18708 9456 18717
rect 9588 18708 9640 18760
rect 9496 18572 9548 18624
rect 10508 18708 10560 18760
rect 10232 18640 10284 18692
rect 10692 18640 10744 18692
rect 15292 18844 15344 18896
rect 16120 18844 16172 18896
rect 18420 18912 18472 18964
rect 18512 18844 18564 18896
rect 20720 18912 20772 18964
rect 22560 18844 22612 18896
rect 23020 18912 23072 18964
rect 24952 18912 25004 18964
rect 11244 18708 11296 18760
rect 11520 18708 11572 18760
rect 12164 18751 12216 18760
rect 12164 18717 12166 18751
rect 12166 18717 12216 18751
rect 12164 18708 12216 18717
rect 14188 18819 14240 18828
rect 14188 18785 14197 18819
rect 14197 18785 14231 18819
rect 14231 18785 14240 18819
rect 14188 18776 14240 18785
rect 14372 18776 14424 18828
rect 12900 18708 12952 18760
rect 15936 18776 15988 18828
rect 16304 18819 16356 18828
rect 16304 18785 16313 18819
rect 16313 18785 16347 18819
rect 16347 18785 16356 18819
rect 16304 18776 16356 18785
rect 16672 18776 16724 18828
rect 16948 18819 17000 18828
rect 16948 18785 16957 18819
rect 16957 18785 16991 18819
rect 16991 18785 17000 18819
rect 16948 18776 17000 18785
rect 15016 18708 15068 18760
rect 16396 18708 16448 18760
rect 20444 18776 20496 18828
rect 17684 18708 17736 18760
rect 16672 18640 16724 18692
rect 20352 18708 20404 18760
rect 21640 18776 21692 18828
rect 23940 18776 23992 18828
rect 26608 18819 26660 18828
rect 26608 18785 26617 18819
rect 26617 18785 26651 18819
rect 26651 18785 26660 18819
rect 26608 18776 26660 18785
rect 26700 18776 26752 18828
rect 20444 18640 20496 18692
rect 23848 18708 23900 18760
rect 22744 18640 22796 18692
rect 23480 18640 23532 18692
rect 11152 18572 11204 18624
rect 13820 18615 13872 18624
rect 13820 18581 13829 18615
rect 13829 18581 13863 18615
rect 13863 18581 13872 18615
rect 13820 18572 13872 18581
rect 18696 18572 18748 18624
rect 20720 18572 20772 18624
rect 22928 18572 22980 18624
rect 24308 18708 24360 18760
rect 24584 18751 24636 18760
rect 24584 18717 24596 18751
rect 24596 18717 24630 18751
rect 24630 18717 24636 18751
rect 24584 18708 24636 18717
rect 26424 18708 26476 18760
rect 29184 18776 29236 18828
rect 29368 18776 29420 18828
rect 29736 18776 29788 18828
rect 24400 18572 24452 18624
rect 26056 18640 26108 18692
rect 28264 18708 28316 18760
rect 30196 18776 30248 18828
rect 25964 18615 26016 18624
rect 25964 18581 25973 18615
rect 25973 18581 26007 18615
rect 26007 18581 26016 18615
rect 25964 18572 26016 18581
rect 26424 18615 26476 18624
rect 26424 18581 26433 18615
rect 26433 18581 26467 18615
rect 26467 18581 26476 18615
rect 26424 18572 26476 18581
rect 27712 18572 27764 18624
rect 29276 18572 29328 18624
rect 29736 18572 29788 18624
rect 30288 18615 30340 18624
rect 30288 18581 30297 18615
rect 30297 18581 30331 18615
rect 30331 18581 30340 18615
rect 30288 18572 30340 18581
rect 4193 18470 4245 18522
rect 4257 18470 4309 18522
rect 4321 18470 4373 18522
rect 4385 18470 4437 18522
rect 4449 18470 4501 18522
rect 11783 18470 11835 18522
rect 11847 18470 11899 18522
rect 11911 18470 11963 18522
rect 11975 18470 12027 18522
rect 12039 18470 12091 18522
rect 19373 18470 19425 18522
rect 19437 18470 19489 18522
rect 19501 18470 19553 18522
rect 19565 18470 19617 18522
rect 19629 18470 19681 18522
rect 26963 18470 27015 18522
rect 27027 18470 27079 18522
rect 27091 18470 27143 18522
rect 27155 18470 27207 18522
rect 27219 18470 27271 18522
rect 1216 18368 1268 18420
rect 2780 18411 2832 18420
rect 2780 18377 2789 18411
rect 2789 18377 2823 18411
rect 2823 18377 2832 18411
rect 2780 18368 2832 18377
rect 3424 18368 3476 18420
rect 3976 18368 4028 18420
rect 4804 18368 4856 18420
rect 5172 18368 5224 18420
rect 5264 18368 5316 18420
rect 5632 18368 5684 18420
rect 6736 18368 6788 18420
rect 6920 18368 6972 18420
rect 8852 18368 8904 18420
rect 9588 18368 9640 18420
rect 2964 18232 3016 18284
rect 5908 18300 5960 18352
rect 8484 18300 8536 18352
rect 3884 18232 3936 18284
rect 5540 18232 5592 18284
rect 5632 18232 5684 18284
rect 8300 18232 8352 18284
rect 9680 18232 9732 18284
rect 1216 18164 1268 18216
rect 2688 18164 2740 18216
rect 3516 18164 3568 18216
rect 3976 18207 4028 18216
rect 3976 18173 3985 18207
rect 3985 18173 4019 18207
rect 4019 18173 4028 18207
rect 3976 18164 4028 18173
rect 4068 18164 4120 18216
rect 6000 18207 6052 18216
rect 6000 18173 6009 18207
rect 6009 18173 6043 18207
rect 6043 18173 6052 18207
rect 6000 18164 6052 18173
rect 6092 18207 6144 18216
rect 6092 18173 6101 18207
rect 6101 18173 6135 18207
rect 6135 18173 6144 18207
rect 6092 18164 6144 18173
rect 8852 18207 8904 18216
rect 8852 18173 8854 18207
rect 8854 18173 8904 18207
rect 8852 18164 8904 18173
rect 9956 18164 10008 18216
rect 8576 18096 8628 18148
rect 12532 18411 12584 18420
rect 12532 18377 12541 18411
rect 12541 18377 12575 18411
rect 12575 18377 12584 18411
rect 12532 18368 12584 18377
rect 13084 18411 13136 18420
rect 13084 18377 13093 18411
rect 13093 18377 13127 18411
rect 13127 18377 13136 18411
rect 13084 18368 13136 18377
rect 13452 18368 13504 18420
rect 14188 18368 14240 18420
rect 16396 18368 16448 18420
rect 17684 18368 17736 18420
rect 11612 18232 11664 18284
rect 13728 18232 13780 18284
rect 1676 18028 1728 18080
rect 1768 18028 1820 18080
rect 6184 18028 6236 18080
rect 6736 18028 6788 18080
rect 7656 18028 7708 18080
rect 10048 18028 10100 18080
rect 10692 18028 10744 18080
rect 14372 18207 14424 18216
rect 14372 18173 14381 18207
rect 14381 18173 14415 18207
rect 14415 18173 14424 18207
rect 14372 18164 14424 18173
rect 16028 18164 16080 18216
rect 17224 18232 17276 18284
rect 17960 18164 18012 18216
rect 22560 18368 22612 18420
rect 22652 18368 22704 18420
rect 24492 18368 24544 18420
rect 20352 18300 20404 18352
rect 22836 18300 22888 18352
rect 26792 18368 26844 18420
rect 18604 18232 18656 18284
rect 18696 18207 18748 18216
rect 18696 18173 18705 18207
rect 18705 18173 18739 18207
rect 18739 18173 18748 18207
rect 18696 18164 18748 18173
rect 20352 18164 20404 18216
rect 20904 18207 20956 18216
rect 20904 18173 20906 18207
rect 20906 18173 20956 18207
rect 20904 18164 20956 18173
rect 21272 18275 21324 18284
rect 21272 18241 21281 18275
rect 21281 18241 21315 18275
rect 21315 18241 21324 18275
rect 21272 18232 21324 18241
rect 26608 18343 26660 18352
rect 26608 18309 26617 18343
rect 26617 18309 26651 18343
rect 26651 18309 26660 18343
rect 26608 18300 26660 18309
rect 25964 18232 26016 18284
rect 12624 18096 12676 18148
rect 13636 18096 13688 18148
rect 23664 18164 23716 18216
rect 23848 18164 23900 18216
rect 24124 18164 24176 18216
rect 24308 18164 24360 18216
rect 24676 18164 24728 18216
rect 30380 18232 30432 18284
rect 13912 18028 13964 18080
rect 14648 18028 14700 18080
rect 14832 18071 14884 18080
rect 14832 18037 14847 18071
rect 14847 18037 14881 18071
rect 14881 18037 14884 18071
rect 14832 18028 14884 18037
rect 16212 18071 16264 18080
rect 16212 18037 16221 18071
rect 16221 18037 16255 18071
rect 16255 18037 16264 18071
rect 16212 18028 16264 18037
rect 16672 18028 16724 18080
rect 18328 18071 18380 18080
rect 18328 18037 18337 18071
rect 18337 18037 18371 18071
rect 18371 18037 18380 18071
rect 18328 18028 18380 18037
rect 22192 18028 22244 18080
rect 22376 18071 22428 18080
rect 22376 18037 22385 18071
rect 22385 18037 22419 18071
rect 22419 18037 22428 18071
rect 22376 18028 22428 18037
rect 24492 18028 24544 18080
rect 25136 18028 25188 18080
rect 26148 18028 26200 18080
rect 27436 18096 27488 18148
rect 27804 18096 27856 18148
rect 29184 18164 29236 18216
rect 29368 18164 29420 18216
rect 28908 18096 28960 18148
rect 28816 18071 28868 18080
rect 28816 18037 28825 18071
rect 28825 18037 28859 18071
rect 28859 18037 28868 18071
rect 28816 18028 28868 18037
rect 29092 18028 29144 18080
rect 29736 18028 29788 18080
rect 30196 18028 30248 18080
rect 7988 17926 8040 17978
rect 8052 17926 8104 17978
rect 8116 17926 8168 17978
rect 8180 17926 8232 17978
rect 8244 17926 8296 17978
rect 15578 17926 15630 17978
rect 15642 17926 15694 17978
rect 15706 17926 15758 17978
rect 15770 17926 15822 17978
rect 15834 17926 15886 17978
rect 23168 17926 23220 17978
rect 23232 17926 23284 17978
rect 23296 17926 23348 17978
rect 23360 17926 23412 17978
rect 23424 17926 23476 17978
rect 30758 17926 30810 17978
rect 30822 17926 30874 17978
rect 30886 17926 30938 17978
rect 30950 17926 31002 17978
rect 31014 17926 31066 17978
rect 1124 17756 1176 17808
rect 848 17688 900 17740
rect 1676 17663 1728 17672
rect 1676 17629 1678 17663
rect 1678 17629 1728 17663
rect 1676 17620 1728 17629
rect 3148 17688 3200 17740
rect 2412 17620 2464 17672
rect 1216 17484 1268 17536
rect 1952 17484 2004 17536
rect 4528 17824 4580 17876
rect 4620 17824 4672 17876
rect 3516 17756 3568 17808
rect 6368 17824 6420 17876
rect 6736 17824 6788 17876
rect 7840 17824 7892 17876
rect 8484 17867 8536 17876
rect 8484 17833 8493 17867
rect 8493 17833 8527 17867
rect 8527 17833 8536 17867
rect 8484 17824 8536 17833
rect 10140 17824 10192 17876
rect 11060 17824 11112 17876
rect 12164 17824 12216 17876
rect 3884 17663 3936 17672
rect 3884 17629 3886 17663
rect 3886 17629 3936 17663
rect 3884 17620 3936 17629
rect 5816 17688 5868 17740
rect 5264 17620 5316 17672
rect 5540 17620 5592 17672
rect 8576 17688 8628 17740
rect 6092 17620 6144 17672
rect 7012 17620 7064 17672
rect 8668 17663 8720 17672
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 9036 17663 9088 17672
rect 9036 17629 9038 17663
rect 9038 17629 9088 17663
rect 9036 17620 9088 17629
rect 9220 17688 9272 17740
rect 9864 17688 9916 17740
rect 11428 17756 11480 17808
rect 11244 17620 11296 17672
rect 11520 17663 11572 17672
rect 11520 17629 11529 17663
rect 11529 17629 11563 17663
rect 11563 17629 11572 17663
rect 11520 17620 11572 17629
rect 16212 17824 16264 17876
rect 16488 17824 16540 17876
rect 16120 17756 16172 17808
rect 16672 17731 16724 17740
rect 16672 17697 16681 17731
rect 16681 17697 16715 17731
rect 16715 17697 16724 17731
rect 16672 17688 16724 17697
rect 23296 17824 23348 17876
rect 20536 17756 20588 17808
rect 21088 17756 21140 17808
rect 15016 17620 15068 17672
rect 15476 17620 15528 17672
rect 18328 17688 18380 17740
rect 19800 17688 19852 17740
rect 20904 17688 20956 17740
rect 26148 17824 26200 17876
rect 27068 17824 27120 17876
rect 23480 17731 23532 17740
rect 23480 17697 23489 17731
rect 23489 17697 23523 17731
rect 23523 17697 23532 17731
rect 23480 17688 23532 17697
rect 28908 17824 28960 17876
rect 29736 17756 29788 17808
rect 16948 17663 17000 17672
rect 16948 17629 16957 17663
rect 16957 17629 16991 17663
rect 16991 17629 17000 17663
rect 16948 17620 17000 17629
rect 17500 17663 17552 17672
rect 17500 17629 17502 17663
rect 17502 17629 17552 17663
rect 3792 17484 3844 17536
rect 4068 17484 4120 17536
rect 5908 17484 5960 17536
rect 9496 17484 9548 17536
rect 10692 17484 10744 17536
rect 10968 17484 11020 17536
rect 16396 17552 16448 17604
rect 17500 17620 17552 17629
rect 15936 17484 15988 17536
rect 17684 17484 17736 17536
rect 17960 17484 18012 17536
rect 20444 17620 20496 17672
rect 21088 17620 21140 17672
rect 21272 17663 21324 17672
rect 21272 17629 21281 17663
rect 21281 17629 21315 17663
rect 21315 17629 21324 17663
rect 21272 17620 21324 17629
rect 22928 17620 22980 17672
rect 24492 17663 24544 17672
rect 24492 17629 24494 17663
rect 24494 17629 24544 17663
rect 20812 17527 20864 17536
rect 20812 17493 20821 17527
rect 20821 17493 20855 17527
rect 20855 17493 20864 17527
rect 20812 17484 20864 17493
rect 23572 17595 23624 17604
rect 23572 17561 23581 17595
rect 23581 17561 23615 17595
rect 23615 17561 23624 17595
rect 23572 17552 23624 17561
rect 23020 17484 23072 17536
rect 23112 17527 23164 17536
rect 23112 17493 23121 17527
rect 23121 17493 23155 17527
rect 23155 17493 23164 17527
rect 23112 17484 23164 17493
rect 23756 17484 23808 17536
rect 24492 17620 24544 17629
rect 24768 17620 24820 17672
rect 28908 17731 28960 17740
rect 28908 17697 28917 17731
rect 28917 17697 28951 17731
rect 28951 17697 28960 17731
rect 28908 17688 28960 17697
rect 29184 17688 29236 17740
rect 25780 17620 25832 17672
rect 26884 17663 26936 17672
rect 26884 17629 26896 17663
rect 26896 17629 26930 17663
rect 26930 17629 26936 17663
rect 26884 17620 26936 17629
rect 24768 17484 24820 17536
rect 25780 17484 25832 17536
rect 25872 17484 25924 17536
rect 27804 17484 27856 17536
rect 30472 17663 30524 17672
rect 30472 17629 30481 17663
rect 30481 17629 30515 17663
rect 30515 17629 30524 17663
rect 30472 17620 30524 17629
rect 30104 17552 30156 17604
rect 4193 17382 4245 17434
rect 4257 17382 4309 17434
rect 4321 17382 4373 17434
rect 4385 17382 4437 17434
rect 4449 17382 4501 17434
rect 11783 17382 11835 17434
rect 11847 17382 11899 17434
rect 11911 17382 11963 17434
rect 11975 17382 12027 17434
rect 12039 17382 12091 17434
rect 19373 17382 19425 17434
rect 19437 17382 19489 17434
rect 19501 17382 19553 17434
rect 19565 17382 19617 17434
rect 19629 17382 19681 17434
rect 26963 17382 27015 17434
rect 27027 17382 27079 17434
rect 27091 17382 27143 17434
rect 27155 17382 27207 17434
rect 27219 17382 27271 17434
rect 2872 17280 2924 17332
rect 4528 17280 4580 17332
rect 9772 17280 9824 17332
rect 10508 17323 10560 17332
rect 10508 17289 10517 17323
rect 10517 17289 10551 17323
rect 10551 17289 10560 17323
rect 10508 17280 10560 17289
rect 11060 17323 11112 17332
rect 11060 17289 11069 17323
rect 11069 17289 11103 17323
rect 11103 17289 11112 17323
rect 11060 17280 11112 17289
rect 2780 17144 2832 17196
rect 3516 17144 3568 17196
rect 4068 17144 4120 17196
rect 4436 17144 4488 17196
rect 5356 17144 5408 17196
rect 6644 17144 6696 17196
rect 1216 17076 1268 17128
rect 1768 17076 1820 17128
rect 3424 17076 3476 17128
rect 3792 17076 3844 17128
rect 5908 17076 5960 17128
rect 6092 17119 6144 17128
rect 6092 17085 6101 17119
rect 6101 17085 6135 17119
rect 6135 17085 6144 17119
rect 6092 17076 6144 17085
rect 1676 16940 1728 16992
rect 8668 17119 8720 17128
rect 8668 17085 8677 17119
rect 8677 17085 8711 17119
rect 8711 17085 8720 17119
rect 8668 17076 8720 17085
rect 9496 17144 9548 17196
rect 12808 17212 12860 17264
rect 9404 17119 9456 17128
rect 9404 17085 9413 17119
rect 9413 17085 9447 17119
rect 9447 17085 9456 17119
rect 9404 17076 9456 17085
rect 12716 17144 12768 17196
rect 14188 17187 14240 17196
rect 14188 17153 14197 17187
rect 14197 17153 14231 17187
rect 14231 17153 14240 17187
rect 14188 17144 14240 17153
rect 14372 17144 14424 17196
rect 18052 17212 18104 17264
rect 16580 17144 16632 17196
rect 16764 17187 16816 17196
rect 16764 17153 16766 17187
rect 16766 17153 16816 17187
rect 16764 17144 16816 17153
rect 23112 17280 23164 17332
rect 28816 17280 28868 17332
rect 29736 17280 29788 17332
rect 30564 17280 30616 17332
rect 20536 17212 20588 17264
rect 10876 17119 10928 17128
rect 10876 17085 10885 17119
rect 10885 17085 10919 17119
rect 10919 17085 10928 17119
rect 10876 17076 10928 17085
rect 11244 17119 11296 17128
rect 11244 17085 11253 17119
rect 11253 17085 11287 17119
rect 11287 17085 11296 17119
rect 11244 17076 11296 17085
rect 11336 17076 11388 17128
rect 13636 17119 13688 17128
rect 13636 17085 13645 17119
rect 13645 17085 13679 17119
rect 13679 17085 13688 17119
rect 13636 17076 13688 17085
rect 14832 17076 14884 17128
rect 14924 17119 14976 17128
rect 14924 17085 14933 17119
rect 14933 17085 14967 17119
rect 14967 17085 14976 17119
rect 14924 17076 14976 17085
rect 16396 17119 16448 17128
rect 16396 17085 16405 17119
rect 16405 17085 16439 17119
rect 16439 17085 16448 17119
rect 16396 17076 16448 17085
rect 20720 17144 20772 17196
rect 21180 17144 21232 17196
rect 23388 17212 23440 17264
rect 23572 17212 23624 17264
rect 23848 17212 23900 17264
rect 28448 17212 28500 17264
rect 28632 17212 28684 17264
rect 28908 17212 28960 17264
rect 29368 17212 29420 17264
rect 22744 17144 22796 17196
rect 25136 17187 25188 17196
rect 3884 16940 3936 16992
rect 4252 16940 4304 16992
rect 4988 16940 5040 16992
rect 5816 16940 5868 16992
rect 6736 16940 6788 16992
rect 8484 16940 8536 16992
rect 9036 16940 9088 16992
rect 10416 16940 10468 16992
rect 11980 16940 12032 16992
rect 12072 16940 12124 16992
rect 14924 16940 14976 16992
rect 16120 16940 16172 16992
rect 20352 17008 20404 17060
rect 21364 17076 21416 17128
rect 23204 17076 23256 17128
rect 22560 17008 22612 17060
rect 24124 17076 24176 17128
rect 24216 17119 24268 17128
rect 24216 17085 24225 17119
rect 24225 17085 24259 17119
rect 24259 17085 24268 17119
rect 24216 17076 24268 17085
rect 24676 17076 24728 17128
rect 24768 17119 24820 17128
rect 24768 17085 24777 17119
rect 24777 17085 24811 17119
rect 24811 17085 24820 17119
rect 24768 17076 24820 17085
rect 25136 17153 25138 17187
rect 25138 17153 25188 17187
rect 25136 17144 25188 17153
rect 25320 17144 25372 17196
rect 26424 17144 26476 17196
rect 26792 17076 26844 17128
rect 27436 17144 27488 17196
rect 29184 17144 29236 17196
rect 27712 17076 27764 17128
rect 29092 17119 29144 17128
rect 29092 17085 29101 17119
rect 29101 17085 29135 17119
rect 29135 17085 29144 17119
rect 29092 17076 29144 17085
rect 30472 17076 30524 17128
rect 24492 17051 24544 17060
rect 24492 17017 24501 17051
rect 24501 17017 24535 17051
rect 24535 17017 24544 17051
rect 24492 17008 24544 17017
rect 30288 17008 30340 17060
rect 31116 17008 31168 17060
rect 19432 16940 19484 16992
rect 21180 16940 21232 16992
rect 22100 16940 22152 16992
rect 23756 16940 23808 16992
rect 23848 16983 23900 16992
rect 23848 16949 23857 16983
rect 23857 16949 23891 16983
rect 23891 16949 23900 16983
rect 23848 16940 23900 16949
rect 25136 16940 25188 16992
rect 25872 16940 25924 16992
rect 26240 16940 26292 16992
rect 26608 16983 26660 16992
rect 26608 16949 26617 16983
rect 26617 16949 26651 16983
rect 26651 16949 26660 16983
rect 26608 16940 26660 16949
rect 26700 16940 26752 16992
rect 29368 16940 29420 16992
rect 7988 16838 8040 16890
rect 8052 16838 8104 16890
rect 8116 16838 8168 16890
rect 8180 16838 8232 16890
rect 8244 16838 8296 16890
rect 15578 16838 15630 16890
rect 15642 16838 15694 16890
rect 15706 16838 15758 16890
rect 15770 16838 15822 16890
rect 15834 16838 15886 16890
rect 23168 16838 23220 16890
rect 23232 16838 23284 16890
rect 23296 16838 23348 16890
rect 23360 16838 23412 16890
rect 23424 16838 23476 16890
rect 30758 16838 30810 16890
rect 30822 16838 30874 16890
rect 30886 16838 30938 16890
rect 30950 16838 31002 16890
rect 31014 16838 31066 16890
rect 1216 16736 1268 16788
rect 664 16668 716 16720
rect 3240 16736 3292 16788
rect 4252 16736 4304 16788
rect 7012 16736 7064 16788
rect 9312 16736 9364 16788
rect 9588 16736 9640 16788
rect 3332 16668 3384 16720
rect 1676 16643 1728 16652
rect 1676 16609 1678 16643
rect 1678 16609 1728 16643
rect 1676 16600 1728 16609
rect 3056 16600 3108 16652
rect 3240 16600 3292 16652
rect 3424 16600 3476 16652
rect 5632 16711 5684 16720
rect 5632 16677 5641 16711
rect 5641 16677 5675 16711
rect 5675 16677 5684 16711
rect 5632 16668 5684 16677
rect 5908 16668 5960 16720
rect 10416 16779 10468 16788
rect 10416 16745 10425 16779
rect 10425 16745 10459 16779
rect 10459 16745 10468 16779
rect 10416 16736 10468 16745
rect 10876 16736 10928 16788
rect 12624 16736 12676 16788
rect 12808 16736 12860 16788
rect 14464 16736 14516 16788
rect 14832 16736 14884 16788
rect 15292 16736 15344 16788
rect 16120 16736 16172 16788
rect 16764 16736 16816 16788
rect 17500 16779 17552 16788
rect 17500 16745 17515 16779
rect 17515 16745 17549 16779
rect 17549 16745 17552 16779
rect 17500 16736 17552 16745
rect 18052 16736 18104 16788
rect 3792 16600 3844 16652
rect 5356 16600 5408 16652
rect 8116 16600 8168 16652
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 4068 16532 4120 16584
rect 4436 16532 4488 16584
rect 6368 16532 6420 16584
rect 4988 16464 5040 16516
rect 8208 16464 8260 16516
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 8944 16575 8996 16584
rect 8944 16541 8946 16575
rect 8946 16541 8996 16575
rect 8944 16532 8996 16541
rect 10784 16600 10836 16652
rect 9496 16532 9548 16584
rect 11336 16600 11388 16652
rect 11704 16600 11756 16652
rect 11980 16643 12032 16652
rect 11980 16609 11982 16643
rect 11982 16609 12032 16643
rect 11980 16600 12032 16609
rect 8484 16464 8536 16516
rect 12256 16532 12308 16584
rect 14188 16600 14240 16652
rect 20812 16736 20864 16788
rect 22744 16736 22796 16788
rect 20720 16668 20772 16720
rect 16580 16600 16632 16652
rect 19524 16600 19576 16652
rect 1032 16439 1084 16448
rect 1032 16405 1041 16439
rect 1041 16405 1075 16439
rect 1075 16405 1084 16439
rect 1032 16396 1084 16405
rect 3976 16396 4028 16448
rect 11060 16396 11112 16448
rect 12164 16396 12216 16448
rect 14648 16532 14700 16584
rect 17224 16532 17276 16584
rect 23848 16736 23900 16788
rect 24308 16736 24360 16788
rect 24492 16736 24544 16788
rect 26056 16779 26108 16788
rect 26056 16745 26065 16779
rect 26065 16745 26099 16779
rect 26099 16745 26108 16779
rect 26056 16736 26108 16745
rect 26884 16736 26936 16788
rect 27804 16736 27856 16788
rect 28540 16736 28592 16788
rect 29644 16779 29696 16788
rect 29644 16745 29653 16779
rect 29653 16745 29687 16779
rect 29687 16745 29696 16779
rect 29644 16736 29696 16745
rect 30380 16779 30432 16788
rect 30380 16745 30389 16779
rect 30389 16745 30423 16779
rect 30423 16745 30432 16779
rect 30380 16736 30432 16745
rect 23020 16668 23072 16720
rect 23756 16600 23808 16652
rect 23848 16600 23900 16652
rect 17684 16532 17736 16584
rect 19432 16575 19484 16584
rect 19432 16541 19441 16575
rect 19441 16541 19475 16575
rect 19475 16541 19484 16575
rect 19432 16532 19484 16541
rect 20628 16532 20680 16584
rect 21180 16532 21232 16584
rect 21272 16575 21324 16584
rect 21272 16541 21281 16575
rect 21281 16541 21315 16575
rect 21315 16541 21324 16575
rect 21272 16532 21324 16541
rect 24124 16532 24176 16584
rect 24492 16600 24544 16652
rect 30196 16668 30248 16720
rect 25780 16643 25832 16652
rect 25780 16609 25789 16643
rect 25789 16609 25823 16643
rect 25823 16609 25832 16643
rect 25780 16600 25832 16609
rect 26240 16600 26292 16652
rect 26792 16600 26844 16652
rect 27436 16600 27488 16652
rect 27620 16600 27672 16652
rect 28172 16600 28224 16652
rect 29000 16600 29052 16652
rect 27528 16532 27580 16584
rect 28448 16532 28500 16584
rect 15476 16464 15528 16516
rect 16304 16464 16356 16516
rect 16856 16464 16908 16516
rect 18512 16464 18564 16516
rect 15936 16396 15988 16448
rect 18788 16396 18840 16448
rect 18880 16439 18932 16448
rect 18880 16405 18889 16439
rect 18889 16405 18923 16439
rect 18923 16405 18932 16439
rect 18880 16396 18932 16405
rect 23480 16396 23532 16448
rect 23940 16396 23992 16448
rect 25136 16396 25188 16448
rect 25320 16439 25372 16448
rect 25320 16405 25329 16439
rect 25329 16405 25363 16439
rect 25363 16405 25372 16439
rect 25320 16396 25372 16405
rect 26424 16396 26476 16448
rect 28908 16396 28960 16448
rect 4193 16294 4245 16346
rect 4257 16294 4309 16346
rect 4321 16294 4373 16346
rect 4385 16294 4437 16346
rect 4449 16294 4501 16346
rect 11783 16294 11835 16346
rect 11847 16294 11899 16346
rect 11911 16294 11963 16346
rect 11975 16294 12027 16346
rect 12039 16294 12091 16346
rect 19373 16294 19425 16346
rect 19437 16294 19489 16346
rect 19501 16294 19553 16346
rect 19565 16294 19617 16346
rect 19629 16294 19681 16346
rect 26963 16294 27015 16346
rect 27027 16294 27079 16346
rect 27091 16294 27143 16346
rect 27155 16294 27207 16346
rect 27219 16294 27271 16346
rect 2964 16235 3016 16244
rect 2964 16201 2973 16235
rect 2973 16201 3007 16235
rect 3007 16201 3016 16235
rect 2964 16192 3016 16201
rect 1124 16056 1176 16108
rect 3516 16056 3568 16108
rect 3976 16192 4028 16244
rect 4068 16192 4120 16244
rect 8576 16192 8628 16244
rect 6644 16056 6696 16108
rect 11060 16124 11112 16176
rect 13728 16124 13780 16176
rect 8760 16056 8812 16108
rect 11520 16056 11572 16108
rect 3332 15963 3384 15972
rect 3332 15929 3341 15963
rect 3341 15929 3375 15963
rect 3375 15929 3384 15963
rect 3332 15920 3384 15929
rect 3884 15988 3936 16040
rect 4528 16031 4580 16040
rect 4528 15997 4537 16031
rect 4537 15997 4571 16031
rect 4571 15997 4580 16031
rect 4528 15988 4580 15997
rect 6092 16031 6144 16040
rect 6092 15997 6101 16031
rect 6101 15997 6135 16031
rect 6135 15997 6144 16031
rect 6092 15988 6144 15997
rect 6460 16031 6512 16040
rect 6460 15997 6462 16031
rect 6462 15997 6512 16031
rect 6460 15988 6512 15997
rect 7656 15988 7708 16040
rect 8208 15988 8260 16040
rect 9220 15988 9272 16040
rect 1400 15895 1452 15904
rect 1400 15861 1415 15895
rect 1415 15861 1449 15895
rect 1449 15861 1452 15895
rect 1400 15852 1452 15861
rect 3516 15852 3568 15904
rect 11336 15988 11388 16040
rect 11612 15988 11664 16040
rect 12348 15988 12400 16040
rect 14188 15988 14240 16040
rect 14832 16056 14884 16108
rect 14924 16056 14976 16108
rect 4160 15852 4212 15904
rect 7840 15852 7892 15904
rect 8944 15852 8996 15904
rect 10416 15895 10468 15904
rect 10416 15861 10425 15895
rect 10425 15861 10459 15895
rect 10459 15861 10468 15895
rect 10416 15852 10468 15861
rect 11152 15852 11204 15904
rect 11704 15895 11756 15904
rect 11704 15861 11719 15895
rect 11719 15861 11753 15895
rect 11753 15861 11756 15895
rect 11704 15852 11756 15861
rect 13084 15895 13136 15904
rect 13084 15861 13093 15895
rect 13093 15861 13127 15895
rect 13127 15861 13136 15895
rect 13084 15852 13136 15861
rect 13912 15920 13964 15972
rect 14280 15920 14332 15972
rect 14648 16031 14700 16040
rect 14648 15997 14657 16031
rect 14657 15997 14691 16031
rect 14691 15997 14700 16031
rect 14648 15988 14700 15997
rect 15200 16056 15252 16108
rect 20536 16192 20588 16244
rect 18512 16124 18564 16176
rect 17500 16056 17552 16108
rect 22376 16192 22428 16244
rect 24584 16192 24636 16244
rect 25964 16192 26016 16244
rect 20720 16167 20772 16176
rect 20720 16133 20729 16167
rect 20729 16133 20763 16167
rect 20763 16133 20772 16167
rect 20720 16124 20772 16133
rect 21916 16099 21968 16108
rect 21916 16065 21918 16099
rect 21918 16065 21968 16099
rect 21916 16056 21968 16065
rect 22008 16081 22060 16108
rect 22008 16056 22053 16081
rect 22053 16056 22060 16081
rect 23756 16056 23808 16108
rect 24216 16099 24268 16108
rect 24216 16065 24218 16099
rect 24218 16065 24268 16099
rect 24216 16056 24268 16065
rect 24400 16056 24452 16108
rect 24768 16056 24820 16108
rect 26056 16099 26108 16108
rect 26056 16065 26065 16099
rect 26065 16065 26099 16099
rect 26099 16065 26108 16099
rect 26056 16056 26108 16065
rect 26332 16056 26384 16108
rect 27896 16056 27948 16108
rect 15292 15988 15344 16040
rect 15384 16031 15436 16040
rect 15384 15997 15393 16031
rect 15393 15997 15427 16031
rect 15427 15997 15436 16031
rect 15384 15988 15436 15997
rect 16672 15988 16724 16040
rect 16856 16031 16908 16040
rect 16856 15997 16865 16031
rect 16865 15997 16899 16031
rect 16899 15997 16908 16031
rect 16856 15988 16908 15997
rect 17132 16031 17184 16040
rect 17132 15997 17141 16031
rect 17141 15997 17175 16031
rect 17175 15997 17184 16031
rect 17132 15988 17184 15997
rect 17224 15988 17276 16040
rect 16856 15852 16908 15904
rect 18420 15920 18472 15972
rect 18788 15988 18840 16040
rect 18788 15852 18840 15904
rect 19156 15852 19208 15904
rect 20812 15852 20864 15904
rect 21456 15988 21508 16040
rect 23020 15988 23072 16040
rect 24676 15988 24728 16040
rect 25412 15988 25464 16040
rect 31208 16192 31260 16244
rect 29092 16124 29144 16176
rect 28724 16056 28776 16108
rect 29368 16031 29420 16040
rect 29368 15997 29377 16031
rect 29377 15997 29411 16031
rect 29411 15997 29420 16031
rect 29368 15988 29420 15997
rect 29644 15988 29696 16040
rect 30196 16124 30248 16176
rect 29828 15988 29880 16040
rect 21180 15963 21232 15972
rect 21180 15929 21189 15963
rect 21189 15929 21223 15963
rect 21223 15929 21232 15963
rect 21180 15920 21232 15929
rect 23848 15920 23900 15972
rect 25688 15895 25740 15904
rect 25688 15861 25697 15895
rect 25697 15861 25731 15895
rect 25731 15861 25740 15895
rect 25688 15852 25740 15861
rect 26516 15895 26568 15904
rect 26516 15861 26531 15895
rect 26531 15861 26565 15895
rect 26565 15861 26568 15895
rect 28724 15920 28776 15972
rect 30656 15920 30708 15972
rect 26516 15852 26568 15861
rect 27896 15895 27948 15904
rect 27896 15861 27905 15895
rect 27905 15861 27939 15895
rect 27939 15861 27948 15895
rect 27896 15852 27948 15861
rect 29368 15852 29420 15904
rect 29644 15852 29696 15904
rect 7988 15750 8040 15802
rect 8052 15750 8104 15802
rect 8116 15750 8168 15802
rect 8180 15750 8232 15802
rect 8244 15750 8296 15802
rect 15578 15750 15630 15802
rect 15642 15750 15694 15802
rect 15706 15750 15758 15802
rect 15770 15750 15822 15802
rect 15834 15750 15886 15802
rect 23168 15750 23220 15802
rect 23232 15750 23284 15802
rect 23296 15750 23348 15802
rect 23360 15750 23412 15802
rect 23424 15750 23476 15802
rect 30758 15750 30810 15802
rect 30822 15750 30874 15802
rect 30886 15750 30938 15802
rect 30950 15750 31002 15802
rect 31014 15750 31066 15802
rect 1400 15580 1452 15632
rect 3148 15691 3200 15700
rect 3148 15657 3157 15691
rect 3157 15657 3191 15691
rect 3191 15657 3200 15691
rect 3148 15648 3200 15657
rect 4712 15648 4764 15700
rect 4988 15648 5040 15700
rect 10416 15648 10468 15700
rect 1124 15376 1176 15428
rect 2872 15444 2924 15496
rect 3516 15487 3568 15496
rect 3516 15453 3525 15487
rect 3525 15453 3559 15487
rect 3559 15453 3568 15487
rect 3516 15444 3568 15453
rect 3884 15487 3936 15496
rect 3884 15453 3886 15487
rect 3886 15453 3936 15487
rect 3884 15444 3936 15453
rect 4160 15444 4212 15496
rect 5448 15444 5500 15496
rect 1216 15308 1268 15360
rect 3792 15308 3844 15360
rect 6460 15512 6512 15564
rect 6092 15444 6144 15496
rect 7012 15444 7064 15496
rect 6276 15308 6328 15360
rect 8576 15555 8628 15564
rect 8576 15521 8585 15555
rect 8585 15521 8619 15555
rect 8619 15521 8628 15555
rect 8576 15512 8628 15521
rect 8944 15487 8996 15496
rect 8944 15453 8946 15487
rect 8946 15453 8996 15487
rect 8944 15444 8996 15453
rect 10784 15512 10836 15564
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 13084 15648 13136 15700
rect 14464 15648 14516 15700
rect 14648 15648 14700 15700
rect 11060 15623 11112 15632
rect 11060 15589 11069 15623
rect 11069 15589 11103 15623
rect 11103 15589 11112 15623
rect 11060 15580 11112 15589
rect 11336 15580 11388 15632
rect 11704 15580 11756 15632
rect 16396 15580 16448 15632
rect 17224 15648 17276 15700
rect 17776 15648 17828 15700
rect 12532 15444 12584 15496
rect 10600 15376 10652 15428
rect 11520 15376 11572 15428
rect 10416 15351 10468 15360
rect 10416 15317 10425 15351
rect 10425 15317 10459 15351
rect 10459 15317 10468 15351
rect 10416 15308 10468 15317
rect 11060 15308 11112 15360
rect 14188 15512 14240 15564
rect 14556 15555 14608 15564
rect 14556 15521 14565 15555
rect 14565 15521 14599 15555
rect 14599 15521 14608 15555
rect 14556 15512 14608 15521
rect 15936 15555 15988 15564
rect 15936 15521 15945 15555
rect 15945 15521 15979 15555
rect 15979 15521 15988 15555
rect 15936 15512 15988 15521
rect 18144 15512 18196 15564
rect 21824 15648 21876 15700
rect 24216 15648 24268 15700
rect 27436 15648 27488 15700
rect 29276 15648 29328 15700
rect 25964 15580 26016 15632
rect 26516 15580 26568 15632
rect 19432 15555 19484 15564
rect 19432 15521 19441 15555
rect 19441 15521 19475 15555
rect 19475 15521 19484 15555
rect 19432 15512 19484 15521
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 21364 15512 21416 15564
rect 16856 15419 16908 15428
rect 16856 15385 16865 15419
rect 16865 15385 16899 15419
rect 16899 15385 16908 15419
rect 16856 15376 16908 15385
rect 16028 15308 16080 15360
rect 17316 15444 17368 15496
rect 17500 15487 17552 15496
rect 17500 15453 17502 15487
rect 17502 15453 17552 15487
rect 17500 15444 17552 15453
rect 17684 15444 17736 15496
rect 17868 15487 17920 15496
rect 17868 15453 17877 15487
rect 17877 15453 17911 15487
rect 17911 15453 17920 15487
rect 17868 15444 17920 15453
rect 19064 15444 19116 15496
rect 20168 15444 20220 15496
rect 21640 15487 21692 15496
rect 21640 15453 21642 15487
rect 21642 15453 21692 15487
rect 21640 15444 21692 15453
rect 23756 15444 23808 15496
rect 24032 15444 24084 15496
rect 24308 15444 24360 15496
rect 25320 15444 25372 15496
rect 25964 15444 26016 15496
rect 26148 15444 26200 15496
rect 27436 15512 27488 15564
rect 27988 15512 28040 15564
rect 29644 15512 29696 15564
rect 18880 15376 18932 15428
rect 18972 15308 19024 15360
rect 20720 15308 20772 15360
rect 22192 15308 22244 15360
rect 22376 15308 22428 15360
rect 23848 15308 23900 15360
rect 24032 15308 24084 15360
rect 25504 15376 25556 15428
rect 25320 15351 25372 15360
rect 25320 15317 25329 15351
rect 25329 15317 25363 15351
rect 25363 15317 25372 15351
rect 25320 15308 25372 15317
rect 26148 15351 26200 15360
rect 26148 15317 26157 15351
rect 26157 15317 26191 15351
rect 26191 15317 26200 15351
rect 26148 15308 26200 15317
rect 28540 15444 28592 15496
rect 27988 15376 28040 15428
rect 26700 15308 26752 15360
rect 29276 15308 29328 15360
rect 4193 15206 4245 15258
rect 4257 15206 4309 15258
rect 4321 15206 4373 15258
rect 4385 15206 4437 15258
rect 4449 15206 4501 15258
rect 11783 15206 11835 15258
rect 11847 15206 11899 15258
rect 11911 15206 11963 15258
rect 11975 15206 12027 15258
rect 12039 15206 12091 15258
rect 19373 15206 19425 15258
rect 19437 15206 19489 15258
rect 19501 15206 19553 15258
rect 19565 15206 19617 15258
rect 19629 15206 19681 15258
rect 26963 15206 27015 15258
rect 27027 15206 27079 15258
rect 27091 15206 27143 15258
rect 27155 15206 27207 15258
rect 27219 15206 27271 15258
rect 2780 15147 2832 15156
rect 2780 15113 2789 15147
rect 2789 15113 2823 15147
rect 2823 15113 2832 15147
rect 2780 15104 2832 15113
rect 1124 14968 1176 15020
rect 2964 14968 3016 15020
rect 4988 15104 5040 15156
rect 6368 15104 6420 15156
rect 6460 15104 6512 15156
rect 6276 14968 6328 15020
rect 6552 14968 6604 15020
rect 3240 14943 3292 14952
rect 3240 14909 3249 14943
rect 3249 14909 3283 14943
rect 3283 14909 3292 14943
rect 3240 14900 3292 14909
rect 3792 14943 3844 14952
rect 3792 14909 3801 14943
rect 3801 14909 3835 14943
rect 3835 14909 3844 14943
rect 3792 14900 3844 14909
rect 3884 14900 3936 14952
rect 4528 14943 4580 14952
rect 4528 14909 4537 14943
rect 4537 14909 4571 14943
rect 4571 14909 4580 14943
rect 4528 14900 4580 14909
rect 6092 14943 6144 14952
rect 6092 14909 6101 14943
rect 6101 14909 6135 14943
rect 6135 14909 6144 14943
rect 6092 14900 6144 14909
rect 7012 14968 7064 15020
rect 9496 15104 9548 15156
rect 10324 15104 10376 15156
rect 12900 15104 12952 15156
rect 14188 15104 14240 15156
rect 15292 15104 15344 15156
rect 8944 15011 8996 15020
rect 8944 14977 8946 15011
rect 8946 14977 8996 15011
rect 8944 14968 8996 14977
rect 10692 14968 10744 15020
rect 1400 14807 1452 14816
rect 1400 14773 1415 14807
rect 1415 14773 1449 14807
rect 1449 14773 1452 14807
rect 5908 14832 5960 14884
rect 6920 14900 6972 14952
rect 7288 14900 7340 14952
rect 1400 14764 1452 14773
rect 6460 14764 6512 14816
rect 6736 14764 6788 14816
rect 8576 14943 8628 14952
rect 8576 14909 8585 14943
rect 8585 14909 8619 14943
rect 8619 14909 8628 14943
rect 8576 14900 8628 14909
rect 9680 14900 9732 14952
rect 11244 15036 11296 15088
rect 13084 15079 13136 15088
rect 13084 15045 13093 15079
rect 13093 15045 13127 15079
rect 13127 15045 13136 15079
rect 13084 15036 13136 15045
rect 16028 15147 16080 15156
rect 16028 15113 16037 15147
rect 16037 15113 16071 15147
rect 16071 15113 16080 15147
rect 16028 15104 16080 15113
rect 20720 15104 20772 15156
rect 11612 14968 11664 15020
rect 10416 14807 10468 14816
rect 10416 14773 10425 14807
rect 10425 14773 10459 14807
rect 10459 14773 10468 14807
rect 10416 14764 10468 14773
rect 10876 14764 10928 14816
rect 11336 14900 11388 14952
rect 11888 14900 11940 14952
rect 11980 14943 12032 14952
rect 11980 14909 11989 14943
rect 11989 14909 12023 14943
rect 12023 14909 12032 14943
rect 11980 14900 12032 14909
rect 14188 14943 14240 14952
rect 14188 14909 14197 14943
rect 14197 14909 14231 14943
rect 14231 14909 14240 14943
rect 14188 14900 14240 14909
rect 11612 14764 11664 14816
rect 11704 14807 11756 14816
rect 11704 14773 11719 14807
rect 11719 14773 11753 14807
rect 11753 14773 11756 14807
rect 11704 14764 11756 14773
rect 11888 14764 11940 14816
rect 15200 14900 15252 14952
rect 14280 14764 14332 14816
rect 14464 14764 14516 14816
rect 16396 15011 16448 15020
rect 16396 14977 16405 15011
rect 16405 14977 16439 15011
rect 16439 14977 16448 15011
rect 16396 14968 16448 14977
rect 19156 15036 19208 15088
rect 21364 15036 21416 15088
rect 18788 14968 18840 15020
rect 17960 14900 18012 14952
rect 19248 14900 19300 14952
rect 19800 14943 19852 14952
rect 19800 14909 19809 14943
rect 19809 14909 19843 14943
rect 19843 14909 19852 14943
rect 19800 14900 19852 14909
rect 20628 14900 20680 14952
rect 16396 14764 16448 14816
rect 16764 14764 16816 14816
rect 17500 14764 17552 14816
rect 20260 14807 20312 14816
rect 20260 14773 20275 14807
rect 20275 14773 20309 14807
rect 20309 14773 20312 14807
rect 20260 14764 20312 14773
rect 21180 14764 21232 14816
rect 22928 14968 22980 15020
rect 23480 15104 23532 15156
rect 23664 15036 23716 15088
rect 25320 15036 25372 15088
rect 23572 14900 23624 14952
rect 23756 14968 23808 15020
rect 24216 15011 24268 15020
rect 24216 14977 24218 15011
rect 24218 14977 24268 15011
rect 24216 14968 24268 14977
rect 27896 15104 27948 15156
rect 28172 15104 28224 15156
rect 28540 15104 28592 15156
rect 30380 15147 30432 15156
rect 30380 15113 30389 15147
rect 30389 15113 30423 15147
rect 30423 15113 30432 15147
rect 30380 15104 30432 15113
rect 27528 15036 27580 15088
rect 25964 14900 26016 14952
rect 26608 14968 26660 15020
rect 28908 15036 28960 15088
rect 29644 14968 29696 15020
rect 29368 14900 29420 14952
rect 29736 14900 29788 14952
rect 30012 14900 30064 14952
rect 31392 14900 31444 14952
rect 26148 14764 26200 14816
rect 26516 14807 26568 14816
rect 26516 14773 26531 14807
rect 26531 14773 26565 14807
rect 26565 14773 26568 14807
rect 26516 14764 26568 14773
rect 26700 14764 26752 14816
rect 29092 14875 29144 14884
rect 29092 14841 29101 14875
rect 29101 14841 29135 14875
rect 29135 14841 29144 14875
rect 29092 14832 29144 14841
rect 30380 14764 30432 14816
rect 7988 14662 8040 14714
rect 8052 14662 8104 14714
rect 8116 14662 8168 14714
rect 8180 14662 8232 14714
rect 8244 14662 8296 14714
rect 15578 14662 15630 14714
rect 15642 14662 15694 14714
rect 15706 14662 15758 14714
rect 15770 14662 15822 14714
rect 15834 14662 15886 14714
rect 23168 14662 23220 14714
rect 23232 14662 23284 14714
rect 23296 14662 23348 14714
rect 23360 14662 23412 14714
rect 23424 14662 23476 14714
rect 30758 14662 30810 14714
rect 30822 14662 30874 14714
rect 30886 14662 30938 14714
rect 30950 14662 31002 14714
rect 31014 14662 31066 14714
rect 1124 14560 1176 14612
rect 3056 14603 3108 14612
rect 3056 14569 3065 14603
rect 3065 14569 3099 14603
rect 3099 14569 3108 14603
rect 3056 14560 3108 14569
rect 3884 14560 3936 14612
rect 4712 14560 4764 14612
rect 3608 14492 3660 14544
rect 5540 14603 5592 14612
rect 5540 14569 5549 14603
rect 5549 14569 5583 14603
rect 5583 14569 5592 14603
rect 5540 14560 5592 14569
rect 5908 14560 5960 14612
rect 6920 14560 6972 14612
rect 7380 14560 7432 14612
rect 1400 14356 1452 14408
rect 3792 14424 3844 14476
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 5908 14424 5960 14476
rect 6276 14467 6328 14476
rect 6276 14433 6285 14467
rect 6285 14433 6319 14467
rect 6319 14433 6328 14467
rect 6276 14424 6328 14433
rect 940 14263 992 14272
rect 940 14229 949 14263
rect 949 14229 983 14263
rect 983 14229 992 14263
rect 940 14220 992 14229
rect 4160 14356 4212 14408
rect 3240 14220 3292 14272
rect 5632 14220 5684 14272
rect 5816 14263 5868 14272
rect 5816 14229 5825 14263
rect 5825 14229 5859 14263
rect 5859 14229 5868 14263
rect 5816 14220 5868 14229
rect 8944 14492 8996 14544
rect 9312 14560 9364 14612
rect 9680 14603 9732 14612
rect 9680 14569 9689 14603
rect 9689 14569 9723 14603
rect 9723 14569 9732 14603
rect 9680 14560 9732 14569
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 11244 14560 11296 14612
rect 11980 14560 12032 14612
rect 13452 14603 13504 14612
rect 13452 14569 13461 14603
rect 13461 14569 13495 14603
rect 13495 14569 13504 14603
rect 13452 14560 13504 14569
rect 14464 14560 14516 14612
rect 6552 14467 6604 14476
rect 6552 14433 6561 14467
rect 6561 14433 6595 14467
rect 6595 14433 6604 14467
rect 6552 14424 6604 14433
rect 8760 14424 8812 14476
rect 9036 14424 9088 14476
rect 9496 14424 9548 14476
rect 9680 14424 9732 14476
rect 10048 14424 10100 14476
rect 6552 14288 6604 14340
rect 6828 14356 6880 14408
rect 7104 14399 7156 14408
rect 7104 14365 7116 14399
rect 7116 14365 7150 14399
rect 7150 14365 7156 14399
rect 7104 14356 7156 14365
rect 7380 14399 7432 14408
rect 7380 14365 7389 14399
rect 7389 14365 7423 14399
rect 7423 14365 7432 14399
rect 7380 14356 7432 14365
rect 10324 14424 10376 14476
rect 11428 14492 11480 14544
rect 11704 14492 11756 14544
rect 9864 14220 9916 14272
rect 11152 14356 11204 14408
rect 11336 14424 11388 14476
rect 16488 14560 16540 14612
rect 11796 14356 11848 14408
rect 15936 14424 15988 14476
rect 16948 14492 17000 14544
rect 16304 14424 16356 14476
rect 19892 14560 19944 14612
rect 20168 14560 20220 14612
rect 19616 14492 19668 14544
rect 20628 14492 20680 14544
rect 21180 14560 21232 14612
rect 21640 14560 21692 14612
rect 23112 14603 23164 14612
rect 23112 14569 23121 14603
rect 23121 14569 23155 14603
rect 23155 14569 23164 14603
rect 23112 14560 23164 14569
rect 24584 14603 24636 14612
rect 24584 14569 24599 14603
rect 24599 14569 24633 14603
rect 24633 14569 24636 14603
rect 24584 14560 24636 14569
rect 25596 14560 25648 14612
rect 26148 14603 26200 14612
rect 26148 14569 26157 14603
rect 26157 14569 26191 14603
rect 26191 14569 26200 14603
rect 26148 14560 26200 14569
rect 27804 14560 27856 14612
rect 29276 14560 29328 14612
rect 30564 14560 30616 14612
rect 12348 14399 12400 14408
rect 12348 14365 12357 14399
rect 12357 14365 12391 14399
rect 12391 14365 12400 14399
rect 12348 14356 12400 14365
rect 14188 14356 14240 14408
rect 14464 14356 14516 14408
rect 16764 14356 16816 14408
rect 17500 14383 17545 14408
rect 17545 14383 17552 14408
rect 17500 14356 17552 14383
rect 19892 14467 19944 14476
rect 19892 14433 19901 14467
rect 19901 14433 19935 14467
rect 19935 14433 19944 14467
rect 19892 14424 19944 14433
rect 20168 14467 20220 14476
rect 20168 14433 20177 14467
rect 20177 14433 20211 14467
rect 20211 14433 20220 14467
rect 20168 14424 20220 14433
rect 20536 14424 20588 14476
rect 20812 14356 20864 14408
rect 23572 14424 23624 14476
rect 23756 14467 23808 14476
rect 23756 14433 23765 14467
rect 23765 14433 23799 14467
rect 23799 14433 23808 14467
rect 23756 14424 23808 14433
rect 23940 14424 23992 14476
rect 24032 14467 24084 14476
rect 24032 14433 24041 14467
rect 24041 14433 24075 14467
rect 24075 14433 24084 14467
rect 24032 14424 24084 14433
rect 25964 14424 26016 14476
rect 26516 14424 26568 14476
rect 27344 14424 27396 14476
rect 27712 14424 27764 14476
rect 21272 14399 21324 14408
rect 21272 14365 21281 14399
rect 21281 14365 21315 14399
rect 21315 14365 21324 14399
rect 21272 14356 21324 14365
rect 23848 14356 23900 14408
rect 25688 14356 25740 14408
rect 26884 14356 26936 14408
rect 29276 14356 29328 14408
rect 30656 14356 30708 14408
rect 10876 14220 10928 14272
rect 11244 14220 11296 14272
rect 12808 14220 12860 14272
rect 14188 14220 14240 14272
rect 14464 14220 14516 14272
rect 16304 14263 16356 14272
rect 16304 14229 16313 14263
rect 16313 14229 16347 14263
rect 16347 14229 16356 14263
rect 16304 14220 16356 14229
rect 20996 14288 21048 14340
rect 20720 14220 20772 14272
rect 20904 14220 20956 14272
rect 21456 14220 21508 14272
rect 24676 14220 24728 14272
rect 24860 14220 24912 14272
rect 27988 14263 28040 14272
rect 27988 14229 27997 14263
rect 27997 14229 28031 14263
rect 28031 14229 28040 14263
rect 27988 14220 28040 14229
rect 29920 14288 29972 14340
rect 29092 14220 29144 14272
rect 29644 14220 29696 14272
rect 31208 14220 31260 14272
rect 4193 14118 4245 14170
rect 4257 14118 4309 14170
rect 4321 14118 4373 14170
rect 4385 14118 4437 14170
rect 4449 14118 4501 14170
rect 11783 14118 11835 14170
rect 11847 14118 11899 14170
rect 11911 14118 11963 14170
rect 11975 14118 12027 14170
rect 12039 14118 12091 14170
rect 19373 14118 19425 14170
rect 19437 14118 19489 14170
rect 19501 14118 19553 14170
rect 19565 14118 19617 14170
rect 19629 14118 19681 14170
rect 26963 14118 27015 14170
rect 27027 14118 27079 14170
rect 27091 14118 27143 14170
rect 27155 14118 27207 14170
rect 27219 14118 27271 14170
rect 756 13880 808 13932
rect 1308 14016 1360 14068
rect 4068 14016 4120 14068
rect 5816 14016 5868 14068
rect 6736 14016 6788 14068
rect 7656 14016 7708 14068
rect 7840 13948 7892 14000
rect 9220 14016 9272 14068
rect 9404 14016 9456 14068
rect 3148 13880 3200 13932
rect 3884 13880 3936 13932
rect 6092 13923 6144 13932
rect 6092 13889 6101 13923
rect 6101 13889 6135 13923
rect 6135 13889 6144 13923
rect 6092 13880 6144 13889
rect 6644 13880 6696 13932
rect 6736 13880 6788 13932
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 3424 13812 3476 13864
rect 3516 13855 3568 13864
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 5172 13812 5224 13864
rect 6460 13855 6512 13864
rect 6460 13821 6462 13855
rect 6462 13821 6512 13855
rect 6460 13812 6512 13821
rect 7012 13880 7064 13932
rect 8760 13948 8812 14000
rect 8668 13880 8720 13932
rect 9864 13880 9916 13932
rect 6092 13744 6144 13796
rect 1584 13676 1636 13728
rect 2320 13676 2372 13728
rect 2780 13719 2832 13728
rect 2780 13685 2789 13719
rect 2789 13685 2823 13719
rect 2823 13685 2832 13719
rect 2780 13676 2832 13685
rect 3976 13676 4028 13728
rect 5540 13676 5592 13728
rect 10140 13812 10192 13864
rect 10324 13855 10376 13864
rect 10324 13821 10333 13855
rect 10333 13821 10367 13855
rect 10367 13821 10376 13855
rect 10324 13812 10376 13821
rect 10784 13880 10836 13932
rect 12164 13948 12216 14000
rect 12348 13991 12400 14000
rect 12348 13957 12357 13991
rect 12357 13957 12391 13991
rect 12391 13957 12400 13991
rect 12348 13948 12400 13957
rect 12532 14016 12584 14068
rect 12440 13880 12492 13932
rect 11428 13812 11480 13864
rect 11888 13812 11940 13864
rect 13084 13948 13136 14000
rect 13360 13991 13412 14000
rect 13360 13957 13369 13991
rect 13369 13957 13403 13991
rect 13403 13957 13412 13991
rect 13360 13948 13412 13957
rect 13452 13948 13504 14000
rect 16396 14016 16448 14068
rect 15660 13948 15712 14000
rect 17960 14016 18012 14068
rect 14096 13880 14148 13932
rect 14556 13923 14608 13932
rect 14556 13889 14558 13923
rect 14558 13889 14608 13923
rect 14556 13880 14608 13889
rect 14832 13880 14884 13932
rect 16028 13880 16080 13932
rect 16764 13923 16816 13932
rect 16764 13889 16766 13923
rect 16766 13889 16816 13923
rect 16764 13880 16816 13889
rect 21732 14016 21784 14068
rect 19524 13991 19576 14000
rect 19524 13957 19533 13991
rect 19533 13957 19567 13991
rect 19567 13957 19576 13991
rect 19524 13948 19576 13957
rect 23020 13948 23072 14000
rect 9404 13676 9456 13728
rect 9588 13676 9640 13728
rect 11520 13744 11572 13796
rect 11704 13744 11756 13796
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 13176 13855 13228 13864
rect 13176 13821 13185 13855
rect 13185 13821 13219 13855
rect 13219 13821 13228 13855
rect 13176 13812 13228 13821
rect 14280 13812 14332 13864
rect 16488 13812 16540 13864
rect 17500 13812 17552 13864
rect 18880 13855 18932 13864
rect 18880 13821 18889 13855
rect 18889 13821 18923 13855
rect 18923 13821 18932 13855
rect 18880 13812 18932 13821
rect 19156 13855 19208 13864
rect 19156 13821 19165 13855
rect 19165 13821 19199 13855
rect 19199 13821 19208 13855
rect 19156 13812 19208 13821
rect 20168 13880 20220 13932
rect 20444 13880 20496 13932
rect 20720 13880 20772 13932
rect 20996 13880 21048 13932
rect 21824 13880 21876 13932
rect 19800 13855 19852 13864
rect 19800 13821 19809 13855
rect 19809 13821 19843 13855
rect 19843 13821 19852 13855
rect 19800 13812 19852 13821
rect 20904 13812 20956 13864
rect 22008 13855 22060 13864
rect 22008 13821 22040 13855
rect 22040 13821 22060 13855
rect 22008 13812 22060 13821
rect 22192 13880 22244 13932
rect 23848 13880 23900 13932
rect 23940 13812 23992 13864
rect 24216 13880 24268 13932
rect 24584 13880 24636 13932
rect 24676 13880 24728 13932
rect 25504 13948 25556 14000
rect 27528 14016 27580 14068
rect 27620 14016 27672 14068
rect 29000 14016 29052 14068
rect 29552 14059 29604 14068
rect 29552 14025 29561 14059
rect 29561 14025 29595 14059
rect 29595 14025 29604 14059
rect 29552 14016 29604 14025
rect 26884 13880 26936 13932
rect 27068 13880 27120 13932
rect 24124 13812 24176 13864
rect 26424 13855 26476 13864
rect 26424 13821 26425 13855
rect 26425 13821 26459 13855
rect 26459 13821 26476 13855
rect 26424 13812 26476 13821
rect 27344 13880 27396 13932
rect 27620 13880 27672 13932
rect 30104 14059 30156 14068
rect 30104 14025 30113 14059
rect 30113 14025 30147 14059
rect 30147 14025 30156 14059
rect 30104 14016 30156 14025
rect 30288 14016 30340 14068
rect 10048 13719 10100 13728
rect 10048 13685 10063 13719
rect 10063 13685 10097 13719
rect 10097 13685 10100 13719
rect 10048 13676 10100 13685
rect 10692 13676 10744 13728
rect 12992 13744 13044 13796
rect 12624 13676 12676 13728
rect 13176 13676 13228 13728
rect 13820 13719 13872 13728
rect 13820 13685 13829 13719
rect 13829 13685 13863 13719
rect 13863 13685 13872 13719
rect 13820 13676 13872 13685
rect 14188 13676 14240 13728
rect 15016 13676 15068 13728
rect 19248 13744 19300 13796
rect 27436 13855 27488 13864
rect 27436 13821 27445 13855
rect 27445 13821 27479 13855
rect 27479 13821 27488 13855
rect 27436 13812 27488 13821
rect 27804 13812 27856 13864
rect 29092 13812 29144 13864
rect 29920 13948 29972 14000
rect 29828 13812 29880 13864
rect 30380 13812 30432 13864
rect 18144 13676 18196 13728
rect 19708 13676 19760 13728
rect 20260 13719 20312 13728
rect 20260 13685 20275 13719
rect 20275 13685 20309 13719
rect 20309 13685 20312 13719
rect 20260 13676 20312 13685
rect 21180 13676 21232 13728
rect 26240 13676 26292 13728
rect 26792 13676 26844 13728
rect 27712 13676 27764 13728
rect 29000 13719 29052 13728
rect 29000 13685 29009 13719
rect 29009 13685 29043 13719
rect 29043 13685 29052 13719
rect 29000 13676 29052 13685
rect 30104 13744 30156 13796
rect 30564 13676 30616 13728
rect 7988 13574 8040 13626
rect 8052 13574 8104 13626
rect 8116 13574 8168 13626
rect 8180 13574 8232 13626
rect 8244 13574 8296 13626
rect 15578 13574 15630 13626
rect 15642 13574 15694 13626
rect 15706 13574 15758 13626
rect 15770 13574 15822 13626
rect 15834 13574 15886 13626
rect 23168 13574 23220 13626
rect 23232 13574 23284 13626
rect 23296 13574 23348 13626
rect 23360 13574 23412 13626
rect 23424 13574 23476 13626
rect 30758 13574 30810 13626
rect 30822 13574 30874 13626
rect 30886 13574 30938 13626
rect 30950 13574 31002 13626
rect 31014 13574 31066 13626
rect 3976 13515 4028 13524
rect 3976 13481 3991 13515
rect 3991 13481 4025 13515
rect 4025 13481 4028 13515
rect 3976 13472 4028 13481
rect 5172 13472 5224 13524
rect 7288 13472 7340 13524
rect 8392 13472 8444 13524
rect 8576 13472 8628 13524
rect 8944 13515 8996 13524
rect 8944 13481 8953 13515
rect 8953 13481 8987 13515
rect 8987 13481 8996 13515
rect 8944 13472 8996 13481
rect 9128 13472 9180 13524
rect 9772 13472 9824 13524
rect 10324 13472 10376 13524
rect 11428 13472 11480 13524
rect 12808 13472 12860 13524
rect 13636 13472 13688 13524
rect 15200 13472 15252 13524
rect 940 13336 992 13388
rect 6276 13404 6328 13456
rect 848 13268 900 13320
rect 1308 13311 1360 13320
rect 1308 13277 1317 13311
rect 1317 13277 1351 13311
rect 1351 13277 1360 13311
rect 1308 13268 1360 13277
rect 1676 13311 1728 13320
rect 1676 13277 1678 13311
rect 1678 13277 1728 13311
rect 1676 13268 1728 13277
rect 2228 13268 2280 13320
rect 6736 13404 6788 13456
rect 6828 13404 6880 13456
rect 9864 13404 9916 13456
rect 5816 13268 5868 13320
rect 6184 13268 6236 13320
rect 6552 13268 6604 13320
rect 6920 13268 6972 13320
rect 7196 13311 7248 13320
rect 7196 13277 7208 13311
rect 7208 13277 7242 13311
rect 7242 13277 7248 13311
rect 7196 13268 7248 13277
rect 7472 13311 7524 13320
rect 7472 13277 7481 13311
rect 7481 13277 7515 13311
rect 7515 13277 7524 13311
rect 7472 13268 7524 13277
rect 4988 13200 5040 13252
rect 9220 13379 9272 13388
rect 9220 13345 9229 13379
rect 9229 13345 9263 13379
rect 9263 13345 9272 13379
rect 9220 13336 9272 13345
rect 9312 13336 9364 13388
rect 9404 13336 9456 13388
rect 11520 13404 11572 13456
rect 11612 13404 11664 13456
rect 10324 13379 10376 13388
rect 10324 13345 10333 13379
rect 10333 13345 10367 13379
rect 10367 13345 10376 13379
rect 10324 13336 10376 13345
rect 10508 13336 10560 13388
rect 10692 13336 10744 13388
rect 10968 13336 11020 13388
rect 15384 13404 15436 13456
rect 16028 13472 16080 13524
rect 16580 13515 16632 13524
rect 16580 13481 16589 13515
rect 16589 13481 16623 13515
rect 16623 13481 16632 13515
rect 16580 13472 16632 13481
rect 17500 13472 17552 13524
rect 20628 13515 20680 13524
rect 20628 13481 20637 13515
rect 20637 13481 20671 13515
rect 20671 13481 20680 13515
rect 20628 13472 20680 13481
rect 20812 13472 20864 13524
rect 21088 13472 21140 13524
rect 23848 13472 23900 13524
rect 24584 13515 24636 13524
rect 24584 13481 24599 13515
rect 24599 13481 24633 13515
rect 24633 13481 24636 13515
rect 24584 13472 24636 13481
rect 26424 13472 26476 13524
rect 27804 13472 27856 13524
rect 12072 13379 12124 13388
rect 12072 13345 12081 13379
rect 12081 13345 12115 13379
rect 12115 13345 12124 13379
rect 12072 13336 12124 13345
rect 12164 13336 12216 13388
rect 11428 13268 11480 13320
rect 11888 13268 11940 13320
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 15016 13336 15068 13388
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 14556 13268 14608 13320
rect 16764 13336 16816 13388
rect 17040 13336 17092 13388
rect 17684 13336 17736 13388
rect 16580 13268 16632 13320
rect 18144 13336 18196 13388
rect 20536 13336 20588 13388
rect 20904 13336 20956 13388
rect 1584 13132 1636 13184
rect 2228 13132 2280 13184
rect 2504 13132 2556 13184
rect 3424 13132 3476 13184
rect 3792 13132 3844 13184
rect 5448 13132 5500 13184
rect 6368 13132 6420 13184
rect 6644 13132 6696 13184
rect 9404 13132 9456 13184
rect 9496 13132 9548 13184
rect 10324 13200 10376 13252
rect 10416 13243 10468 13252
rect 10416 13209 10425 13243
rect 10425 13209 10459 13243
rect 10459 13209 10468 13243
rect 10416 13200 10468 13209
rect 10600 13200 10652 13252
rect 11244 13200 11296 13252
rect 9772 13132 9824 13184
rect 10048 13132 10100 13184
rect 10140 13175 10192 13184
rect 10140 13141 10149 13175
rect 10149 13141 10183 13175
rect 10183 13141 10192 13175
rect 10140 13132 10192 13141
rect 10508 13132 10560 13184
rect 11980 13175 12032 13184
rect 11980 13141 11989 13175
rect 11989 13141 12023 13175
rect 12023 13141 12032 13175
rect 11980 13132 12032 13141
rect 12808 13132 12860 13184
rect 13176 13132 13228 13184
rect 14372 13175 14424 13184
rect 14372 13141 14381 13175
rect 14381 13141 14415 13175
rect 14415 13141 14424 13175
rect 14372 13132 14424 13141
rect 18328 13311 18380 13320
rect 18328 13277 18337 13311
rect 18337 13277 18371 13311
rect 18371 13277 18380 13311
rect 18328 13268 18380 13277
rect 18696 13311 18748 13320
rect 18696 13277 18698 13311
rect 18698 13277 18748 13311
rect 18696 13268 18748 13277
rect 18788 13311 18840 13320
rect 18788 13277 18800 13311
rect 18800 13277 18834 13311
rect 18834 13277 18840 13311
rect 18788 13268 18840 13277
rect 19984 13268 20036 13320
rect 20720 13268 20772 13320
rect 20996 13268 21048 13320
rect 17868 13200 17920 13252
rect 21824 13379 21876 13388
rect 21824 13345 21833 13379
rect 21833 13345 21867 13379
rect 21867 13345 21876 13379
rect 21824 13336 21876 13345
rect 24216 13404 24268 13456
rect 26332 13404 26384 13456
rect 24124 13379 24176 13388
rect 24124 13345 24133 13379
rect 24133 13345 24167 13379
rect 24167 13345 24176 13379
rect 24124 13336 24176 13345
rect 25504 13336 25556 13388
rect 26056 13336 26108 13388
rect 22284 13268 22336 13320
rect 22560 13268 22612 13320
rect 17684 13132 17736 13184
rect 20352 13175 20404 13184
rect 20352 13141 20361 13175
rect 20361 13141 20395 13175
rect 20395 13141 20404 13175
rect 20352 13132 20404 13141
rect 21548 13200 21600 13252
rect 21732 13200 21784 13252
rect 21272 13132 21324 13184
rect 21916 13132 21968 13184
rect 22284 13132 22336 13184
rect 23664 13132 23716 13184
rect 25320 13268 25372 13320
rect 26608 13268 26660 13320
rect 29000 13472 29052 13524
rect 29368 13472 29420 13524
rect 27988 13336 28040 13388
rect 29368 13336 29420 13388
rect 29552 13336 29604 13388
rect 28264 13243 28316 13252
rect 28264 13209 28273 13243
rect 28273 13209 28307 13243
rect 28307 13209 28316 13243
rect 28264 13200 28316 13209
rect 25964 13132 26016 13184
rect 29092 13268 29144 13320
rect 28908 13132 28960 13184
rect 4193 13030 4245 13082
rect 4257 13030 4309 13082
rect 4321 13030 4373 13082
rect 4385 13030 4437 13082
rect 4449 13030 4501 13082
rect 11783 13030 11835 13082
rect 11847 13030 11899 13082
rect 11911 13030 11963 13082
rect 11975 13030 12027 13082
rect 12039 13030 12091 13082
rect 19373 13030 19425 13082
rect 19437 13030 19489 13082
rect 19501 13030 19553 13082
rect 19565 13030 19617 13082
rect 19629 13030 19681 13082
rect 26963 13030 27015 13082
rect 27027 13030 27079 13082
rect 27091 13030 27143 13082
rect 27155 13030 27207 13082
rect 27219 13030 27271 13082
rect 848 12928 900 12980
rect 4252 12928 4304 12980
rect 7196 12928 7248 12980
rect 7472 12928 7524 12980
rect 8852 12928 8904 12980
rect 3056 12792 3108 12844
rect 1308 12724 1360 12776
rect 1584 12724 1636 12776
rect 3792 12767 3844 12776
rect 3792 12733 3801 12767
rect 3801 12733 3835 12767
rect 3835 12733 3844 12767
rect 3792 12724 3844 12733
rect 4252 12792 4304 12844
rect 5632 12792 5684 12844
rect 6736 12792 6788 12844
rect 3424 12656 3476 12708
rect 6184 12724 6236 12776
rect 6644 12724 6696 12776
rect 1676 12588 1728 12640
rect 3976 12588 4028 12640
rect 6460 12588 6512 12640
rect 6736 12588 6788 12640
rect 9036 12860 9088 12912
rect 9312 12903 9364 12912
rect 9312 12869 9321 12903
rect 9321 12869 9355 12903
rect 9355 12869 9364 12903
rect 9312 12860 9364 12869
rect 8760 12792 8812 12844
rect 7840 12656 7892 12708
rect 9404 12724 9456 12776
rect 11244 12860 11296 12912
rect 9588 12835 9640 12844
rect 9588 12801 9597 12835
rect 9597 12801 9631 12835
rect 9631 12801 9640 12835
rect 9588 12792 9640 12801
rect 9772 12792 9824 12844
rect 10140 12792 10192 12844
rect 10416 12792 10468 12844
rect 10692 12792 10744 12844
rect 8668 12588 8720 12640
rect 9220 12656 9272 12708
rect 11244 12724 11296 12776
rect 12624 12792 12676 12844
rect 13268 12928 13320 12980
rect 15108 12928 15160 12980
rect 16488 12928 16540 12980
rect 17592 12971 17644 12980
rect 17592 12937 17601 12971
rect 17601 12937 17635 12971
rect 17635 12937 17644 12971
rect 17592 12928 17644 12937
rect 12992 12860 13044 12912
rect 19800 12928 19852 12980
rect 23388 12860 23440 12912
rect 11428 12724 11480 12776
rect 12256 12767 12308 12776
rect 12256 12733 12265 12767
rect 12265 12733 12299 12767
rect 12299 12733 12308 12767
rect 12256 12724 12308 12733
rect 12808 12767 12860 12776
rect 12808 12733 12817 12767
rect 12817 12733 12851 12767
rect 12851 12733 12860 12767
rect 12808 12724 12860 12733
rect 12992 12724 13044 12776
rect 13728 12792 13780 12844
rect 13820 12792 13872 12844
rect 16212 12833 16264 12844
rect 16212 12799 16240 12833
rect 16240 12799 16264 12833
rect 16212 12792 16264 12799
rect 18328 12792 18380 12844
rect 19064 12792 19116 12844
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 14556 12724 14608 12776
rect 10692 12588 10744 12640
rect 11244 12588 11296 12640
rect 15476 12656 15528 12708
rect 16488 12767 16540 12776
rect 16488 12733 16497 12767
rect 16497 12733 16531 12767
rect 16531 12733 16540 12767
rect 16488 12724 16540 12733
rect 16580 12724 16632 12776
rect 19432 12767 19484 12776
rect 19432 12733 19441 12767
rect 19441 12733 19475 12767
rect 19475 12733 19484 12767
rect 19432 12724 19484 12733
rect 20352 12792 20404 12844
rect 21548 12792 21600 12844
rect 20720 12724 20772 12776
rect 20904 12767 20956 12776
rect 20904 12733 20913 12767
rect 20913 12733 20947 12767
rect 20947 12733 20956 12767
rect 20904 12724 20956 12733
rect 18696 12656 18748 12708
rect 20628 12656 20680 12708
rect 23296 12767 23348 12776
rect 23296 12733 23305 12767
rect 23305 12733 23339 12767
rect 23339 12733 23348 12767
rect 23296 12724 23348 12733
rect 23756 12860 23808 12912
rect 23664 12792 23716 12844
rect 25688 12971 25740 12980
rect 25688 12937 25697 12971
rect 25697 12937 25731 12971
rect 25731 12937 25740 12971
rect 25688 12928 25740 12937
rect 24032 12792 24084 12844
rect 24216 12792 24268 12844
rect 26424 12792 26476 12844
rect 26884 12928 26936 12980
rect 27712 12928 27764 12980
rect 28448 12971 28500 12980
rect 28448 12937 28457 12971
rect 28457 12937 28491 12971
rect 28491 12937 28500 12971
rect 28448 12928 28500 12937
rect 28816 12928 28868 12980
rect 31300 12928 31352 12980
rect 26792 12792 26844 12844
rect 25412 12724 25464 12776
rect 26148 12724 26200 12776
rect 26608 12767 26660 12776
rect 26608 12733 26617 12767
rect 26617 12733 26651 12767
rect 26651 12733 26660 12767
rect 26608 12724 26660 12733
rect 13176 12631 13228 12640
rect 13176 12597 13185 12631
rect 13185 12597 13219 12631
rect 13219 12597 13228 12631
rect 13176 12588 13228 12597
rect 13636 12588 13688 12640
rect 14188 12588 14240 12640
rect 19156 12631 19208 12640
rect 19156 12597 19171 12631
rect 19171 12597 19205 12631
rect 19205 12597 19208 12631
rect 19156 12588 19208 12597
rect 20720 12631 20772 12640
rect 20720 12597 20729 12631
rect 20729 12597 20763 12631
rect 20763 12597 20772 12631
rect 20720 12588 20772 12597
rect 21640 12588 21692 12640
rect 29000 12724 29052 12776
rect 30104 12860 30156 12912
rect 29828 12767 29880 12776
rect 29828 12733 29837 12767
rect 29837 12733 29871 12767
rect 29871 12733 29880 12767
rect 29828 12724 29880 12733
rect 29920 12724 29972 12776
rect 28172 12656 28224 12708
rect 29552 12656 29604 12708
rect 24124 12588 24176 12640
rect 26332 12588 26384 12640
rect 26700 12588 26752 12640
rect 27988 12588 28040 12640
rect 28080 12588 28132 12640
rect 30012 12631 30064 12640
rect 30012 12597 30021 12631
rect 30021 12597 30055 12631
rect 30055 12597 30064 12631
rect 30012 12588 30064 12597
rect 7988 12486 8040 12538
rect 8052 12486 8104 12538
rect 8116 12486 8168 12538
rect 8180 12486 8232 12538
rect 8244 12486 8296 12538
rect 15578 12486 15630 12538
rect 15642 12486 15694 12538
rect 15706 12486 15758 12538
rect 15770 12486 15822 12538
rect 15834 12486 15886 12538
rect 23168 12486 23220 12538
rect 23232 12486 23284 12538
rect 23296 12486 23348 12538
rect 23360 12486 23412 12538
rect 23424 12486 23476 12538
rect 30758 12486 30810 12538
rect 30822 12486 30874 12538
rect 30886 12486 30938 12538
rect 30950 12486 31002 12538
rect 31014 12486 31066 12538
rect 1676 12384 1728 12436
rect 2688 12384 2740 12436
rect 3516 12316 3568 12368
rect 5632 12384 5684 12436
rect 5816 12427 5868 12436
rect 5816 12393 5825 12427
rect 5825 12393 5859 12427
rect 5859 12393 5868 12427
rect 5816 12384 5868 12393
rect 7932 12384 7984 12436
rect 10232 12384 10284 12436
rect 1308 12223 1360 12232
rect 1308 12189 1317 12223
rect 1317 12189 1351 12223
rect 1351 12189 1360 12223
rect 1308 12180 1360 12189
rect 1952 12180 2004 12232
rect 2044 12223 2096 12232
rect 2044 12189 2053 12223
rect 2053 12189 2087 12223
rect 2087 12189 2096 12223
rect 2044 12180 2096 12189
rect 4160 12248 4212 12300
rect 5908 12248 5960 12300
rect 6552 12316 6604 12368
rect 8668 12316 8720 12368
rect 10692 12316 10744 12368
rect 11704 12384 11756 12436
rect 12624 12384 12676 12436
rect 14004 12384 14056 12436
rect 15016 12384 15068 12436
rect 6828 12291 6880 12300
rect 4068 12180 4120 12232
rect 6828 12257 6830 12291
rect 6830 12257 6880 12291
rect 6828 12248 6880 12257
rect 9036 12291 9088 12300
rect 7104 12180 7156 12232
rect 7196 12223 7248 12232
rect 7196 12189 7205 12223
rect 7205 12189 7239 12223
rect 7239 12189 7248 12223
rect 7196 12180 7248 12189
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 9036 12257 9038 12291
rect 9038 12257 9088 12291
rect 9036 12248 9088 12257
rect 9312 12248 9364 12300
rect 10416 12180 10468 12232
rect 11336 12316 11388 12368
rect 11152 12291 11204 12300
rect 11152 12257 11161 12291
rect 11161 12257 11195 12291
rect 11195 12257 11204 12291
rect 11152 12248 11204 12257
rect 11520 12248 11572 12300
rect 11796 12316 11848 12368
rect 12440 12316 12492 12368
rect 12072 12248 12124 12300
rect 12256 12291 12308 12300
rect 12256 12257 12265 12291
rect 12265 12257 12299 12291
rect 12299 12257 12308 12291
rect 12256 12248 12308 12257
rect 16764 12316 16816 12368
rect 3424 12112 3476 12164
rect 6460 12112 6512 12164
rect 10784 12112 10836 12164
rect 10968 12112 11020 12164
rect 11980 12112 12032 12164
rect 2044 12044 2096 12096
rect 7196 12044 7248 12096
rect 7564 12044 7616 12096
rect 11704 12044 11756 12096
rect 12348 12087 12400 12096
rect 12348 12053 12357 12087
rect 12357 12053 12391 12087
rect 12391 12053 12400 12087
rect 12348 12044 12400 12053
rect 12532 12044 12584 12096
rect 12808 12180 12860 12232
rect 13268 12248 13320 12300
rect 13636 12248 13688 12300
rect 14004 12248 14056 12300
rect 19064 12384 19116 12436
rect 19156 12384 19208 12436
rect 19432 12384 19484 12436
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 20536 12384 20588 12436
rect 20628 12427 20680 12436
rect 20628 12393 20637 12427
rect 20637 12393 20671 12427
rect 20671 12393 20680 12427
rect 20628 12384 20680 12393
rect 16304 12223 16356 12232
rect 16304 12189 16313 12223
rect 16313 12189 16347 12223
rect 16347 12189 16356 12223
rect 16304 12180 16356 12189
rect 13544 12044 13596 12096
rect 14464 12087 14516 12096
rect 14464 12053 14473 12087
rect 14473 12053 14507 12087
rect 14507 12053 14516 12087
rect 14464 12044 14516 12053
rect 19156 12291 19208 12300
rect 19156 12257 19165 12291
rect 19165 12257 19199 12291
rect 19199 12257 19208 12291
rect 19156 12248 19208 12257
rect 16948 12223 17000 12232
rect 16948 12189 16957 12223
rect 16957 12189 16991 12223
rect 16991 12189 17000 12223
rect 16948 12180 17000 12189
rect 17316 12223 17368 12232
rect 17316 12189 17318 12223
rect 17318 12189 17368 12223
rect 17316 12180 17368 12189
rect 18052 12180 18104 12232
rect 19708 12248 19760 12300
rect 19892 12291 19944 12300
rect 19892 12257 19901 12291
rect 19901 12257 19935 12291
rect 19935 12257 19944 12291
rect 19892 12248 19944 12257
rect 19156 12112 19208 12164
rect 21272 12384 21324 12436
rect 22652 12384 22704 12436
rect 24032 12384 24084 12436
rect 24124 12384 24176 12436
rect 21180 12316 21232 12368
rect 23572 12316 23624 12368
rect 25320 12427 25372 12436
rect 25320 12393 25329 12427
rect 25329 12393 25363 12427
rect 25363 12393 25372 12427
rect 25320 12384 25372 12393
rect 26148 12384 26200 12436
rect 26792 12316 26844 12368
rect 26884 12359 26936 12368
rect 26884 12325 26893 12359
rect 26893 12325 26927 12359
rect 26927 12325 26936 12359
rect 26884 12316 26936 12325
rect 21272 12291 21324 12300
rect 21272 12257 21281 12291
rect 21281 12257 21315 12291
rect 21315 12257 21324 12291
rect 21272 12248 21324 12257
rect 24124 12248 24176 12300
rect 24308 12248 24360 12300
rect 21640 12223 21692 12232
rect 21640 12189 21642 12223
rect 21642 12189 21692 12223
rect 21640 12180 21692 12189
rect 21824 12180 21876 12232
rect 23664 12180 23716 12232
rect 23848 12223 23900 12232
rect 23848 12189 23850 12223
rect 23850 12189 23900 12223
rect 23848 12180 23900 12189
rect 23940 12223 23992 12232
rect 23940 12189 23952 12223
rect 23952 12189 23986 12223
rect 23986 12189 23992 12223
rect 25780 12248 25832 12300
rect 26148 12248 26200 12300
rect 26608 12248 26660 12300
rect 26700 12248 26752 12300
rect 27160 12384 27212 12436
rect 29184 12384 29236 12436
rect 27712 12248 27764 12300
rect 28080 12291 28132 12300
rect 28080 12257 28089 12291
rect 28089 12257 28123 12291
rect 28123 12257 28132 12291
rect 28080 12248 28132 12257
rect 30380 12291 30432 12300
rect 30380 12257 30389 12291
rect 30389 12257 30423 12291
rect 30423 12257 30432 12291
rect 30380 12248 30432 12257
rect 23940 12180 23992 12189
rect 28724 12180 28776 12232
rect 28816 12223 28868 12232
rect 28816 12189 28825 12223
rect 28825 12189 28859 12223
rect 28859 12189 28868 12223
rect 28816 12180 28868 12189
rect 29000 12180 29052 12232
rect 21548 12044 21600 12096
rect 21732 12044 21784 12096
rect 23020 12044 23072 12096
rect 23388 12044 23440 12096
rect 25872 12044 25924 12096
rect 28356 12044 28408 12096
rect 4193 11942 4245 11994
rect 4257 11942 4309 11994
rect 4321 11942 4373 11994
rect 4385 11942 4437 11994
rect 4449 11942 4501 11994
rect 11783 11942 11835 11994
rect 11847 11942 11899 11994
rect 11911 11942 11963 11994
rect 11975 11942 12027 11994
rect 12039 11942 12091 11994
rect 19373 11942 19425 11994
rect 19437 11942 19489 11994
rect 19501 11942 19553 11994
rect 19565 11942 19617 11994
rect 19629 11942 19681 11994
rect 26963 11942 27015 11994
rect 27027 11942 27079 11994
rect 27091 11942 27143 11994
rect 27155 11942 27207 11994
rect 27219 11942 27271 11994
rect 1124 11840 1176 11892
rect 1308 11840 1360 11892
rect 3884 11840 3936 11892
rect 7012 11840 7064 11892
rect 7472 11840 7524 11892
rect 7932 11840 7984 11892
rect 9036 11840 9088 11892
rect 9680 11840 9732 11892
rect 11980 11840 12032 11892
rect 12992 11840 13044 11892
rect 13360 11840 13412 11892
rect 14924 11840 14976 11892
rect 18880 11840 18932 11892
rect 19064 11840 19116 11892
rect 7656 11772 7708 11824
rect 24216 11840 24268 11892
rect 26056 11840 26108 11892
rect 1308 11747 1360 11756
rect 1308 11713 1310 11747
rect 1310 11713 1360 11747
rect 1308 11704 1360 11713
rect 2504 11704 2556 11756
rect 1216 11500 1268 11552
rect 1584 11500 1636 11552
rect 3424 11636 3476 11688
rect 3608 11636 3660 11688
rect 4068 11679 4120 11688
rect 4068 11645 4077 11679
rect 4077 11645 4111 11679
rect 4111 11645 4120 11679
rect 4068 11636 4120 11645
rect 4344 11636 4396 11688
rect 5632 11636 5684 11688
rect 5816 11704 5868 11756
rect 6184 11636 6236 11688
rect 7840 11704 7892 11756
rect 8944 11704 8996 11756
rect 9588 11704 9640 11756
rect 9864 11704 9916 11756
rect 10324 11704 10376 11756
rect 10876 11704 10928 11756
rect 12440 11704 12492 11756
rect 9128 11636 9180 11688
rect 9312 11636 9364 11688
rect 7196 11568 7248 11620
rect 3976 11500 4028 11552
rect 6552 11500 6604 11552
rect 6920 11500 6972 11552
rect 7840 11500 7892 11552
rect 8484 11568 8536 11620
rect 11428 11636 11480 11688
rect 11520 11636 11572 11688
rect 12256 11636 12308 11688
rect 13084 11704 13136 11756
rect 14096 11704 14148 11756
rect 9772 11568 9824 11620
rect 8760 11500 8812 11552
rect 9128 11500 9180 11552
rect 9588 11500 9640 11552
rect 10048 11500 10100 11552
rect 10508 11500 10560 11552
rect 11428 11500 11480 11552
rect 12624 11543 12676 11552
rect 12624 11509 12633 11543
rect 12633 11509 12667 11543
rect 12667 11509 12676 11543
rect 12624 11500 12676 11509
rect 13176 11611 13228 11620
rect 13176 11577 13185 11611
rect 13185 11577 13219 11611
rect 13219 11577 13228 11611
rect 13176 11568 13228 11577
rect 13544 11679 13596 11688
rect 13544 11645 13553 11679
rect 13553 11645 13587 11679
rect 13587 11645 13596 11679
rect 13544 11636 13596 11645
rect 16488 11636 16540 11688
rect 16856 11747 16908 11756
rect 16856 11713 16868 11747
rect 16868 11713 16902 11747
rect 16902 11713 16908 11747
rect 16856 11704 16908 11713
rect 19064 11704 19116 11756
rect 17592 11636 17644 11688
rect 18328 11636 18380 11688
rect 18972 11636 19024 11688
rect 19800 11704 19852 11756
rect 20720 11704 20772 11756
rect 21548 11704 21600 11756
rect 21824 11704 21876 11756
rect 20904 11679 20956 11688
rect 20904 11645 20913 11679
rect 20913 11645 20947 11679
rect 20947 11645 20956 11679
rect 20904 11636 20956 11645
rect 23388 11772 23440 11824
rect 15016 11568 15068 11620
rect 12900 11500 12952 11552
rect 13636 11500 13688 11552
rect 14924 11500 14976 11552
rect 23296 11636 23348 11688
rect 23664 11772 23716 11824
rect 23940 11772 23992 11824
rect 23940 11679 23992 11688
rect 23940 11645 23949 11679
rect 23949 11645 23983 11679
rect 23983 11645 23992 11679
rect 23940 11636 23992 11645
rect 23756 11568 23808 11620
rect 23848 11568 23900 11620
rect 24492 11704 24544 11756
rect 25320 11636 25372 11688
rect 26792 11840 26844 11892
rect 27528 11840 27580 11892
rect 27988 11883 28040 11892
rect 27988 11849 27997 11883
rect 27997 11849 28031 11883
rect 28031 11849 28040 11883
rect 27988 11840 28040 11849
rect 28816 11840 28868 11892
rect 29276 11840 29328 11892
rect 29736 11772 29788 11824
rect 26700 11704 26752 11756
rect 16672 11500 16724 11552
rect 17040 11500 17092 11552
rect 18420 11543 18472 11552
rect 18420 11509 18429 11543
rect 18429 11509 18463 11543
rect 18463 11509 18472 11543
rect 18420 11500 18472 11509
rect 19156 11543 19208 11552
rect 19156 11509 19171 11543
rect 19171 11509 19205 11543
rect 19205 11509 19208 11543
rect 19156 11500 19208 11509
rect 21180 11500 21232 11552
rect 21640 11500 21692 11552
rect 22100 11500 22152 11552
rect 22284 11500 22336 11552
rect 27160 11636 27212 11688
rect 29276 11704 29328 11756
rect 26608 11543 26660 11552
rect 26608 11509 26623 11543
rect 26623 11509 26657 11543
rect 26657 11509 26660 11543
rect 29644 11568 29696 11620
rect 29920 11568 29972 11620
rect 29184 11543 29236 11552
rect 26608 11500 26660 11509
rect 29184 11509 29193 11543
rect 29193 11509 29227 11543
rect 29227 11509 29236 11543
rect 29184 11500 29236 11509
rect 30104 11500 30156 11552
rect 7988 11398 8040 11450
rect 8052 11398 8104 11450
rect 8116 11398 8168 11450
rect 8180 11398 8232 11450
rect 8244 11398 8296 11450
rect 15578 11398 15630 11450
rect 15642 11398 15694 11450
rect 15706 11398 15758 11450
rect 15770 11398 15822 11450
rect 15834 11398 15886 11450
rect 23168 11398 23220 11450
rect 23232 11398 23284 11450
rect 23296 11398 23348 11450
rect 23360 11398 23412 11450
rect 23424 11398 23476 11450
rect 30758 11398 30810 11450
rect 30822 11398 30874 11450
rect 30886 11398 30938 11450
rect 30950 11398 31002 11450
rect 31014 11398 31066 11450
rect 1124 11339 1176 11348
rect 1124 11305 1133 11339
rect 1133 11305 1167 11339
rect 1167 11305 1176 11339
rect 1124 11296 1176 11305
rect 3608 11296 3660 11348
rect 4068 11296 4120 11348
rect 4528 11296 4580 11348
rect 5356 11339 5408 11348
rect 5356 11305 5365 11339
rect 5365 11305 5399 11339
rect 5399 11305 5408 11339
rect 5356 11296 5408 11305
rect 6000 11339 6052 11348
rect 6000 11305 6009 11339
rect 6009 11305 6043 11339
rect 6043 11305 6052 11339
rect 6000 11296 6052 11305
rect 6276 11296 6328 11348
rect 1584 11228 1636 11280
rect 1032 11092 1084 11144
rect 1124 11092 1176 11144
rect 1676 11092 1728 11144
rect 2964 11092 3016 11144
rect 664 11024 716 11076
rect 4344 11228 4396 11280
rect 3792 11160 3844 11212
rect 3976 11203 4028 11212
rect 3976 11169 3985 11203
rect 3985 11169 4019 11203
rect 4019 11169 4028 11203
rect 3976 11160 4028 11169
rect 3424 11092 3476 11144
rect 5540 11203 5592 11212
rect 5540 11169 5549 11203
rect 5549 11169 5583 11203
rect 5583 11169 5592 11203
rect 5540 11160 5592 11169
rect 8760 11296 8812 11348
rect 9220 11296 9272 11348
rect 9404 11339 9456 11348
rect 9404 11305 9413 11339
rect 9413 11305 9447 11339
rect 9447 11305 9456 11339
rect 9404 11296 9456 11305
rect 9496 11296 9548 11348
rect 9956 11296 10008 11348
rect 10324 11296 10376 11348
rect 11336 11296 11388 11348
rect 12164 11296 12216 11348
rect 13176 11296 13228 11348
rect 15476 11296 15528 11348
rect 16304 11296 16356 11348
rect 6552 11228 6604 11280
rect 6644 11203 6696 11212
rect 6644 11169 6653 11203
rect 6653 11169 6687 11203
rect 6687 11169 6696 11203
rect 6644 11160 6696 11169
rect 8576 11228 8628 11280
rect 7288 11160 7340 11212
rect 5632 11092 5684 11144
rect 5724 11092 5776 11144
rect 6092 11092 6144 11144
rect 8944 11160 8996 11212
rect 10784 11228 10836 11280
rect 10232 11160 10284 11212
rect 10508 11160 10560 11212
rect 8576 11024 8628 11076
rect 9864 11092 9916 11144
rect 11704 11203 11756 11212
rect 11704 11169 11713 11203
rect 11713 11169 11747 11203
rect 11747 11169 11756 11203
rect 11704 11160 11756 11169
rect 12256 11271 12308 11280
rect 12256 11237 12265 11271
rect 12265 11237 12299 11271
rect 12299 11237 12308 11271
rect 12256 11228 12308 11237
rect 14832 11271 14884 11280
rect 14832 11237 14841 11271
rect 14841 11237 14875 11271
rect 14875 11237 14884 11271
rect 14832 11228 14884 11237
rect 12808 11160 12860 11212
rect 13912 11160 13964 11212
rect 16580 11203 16632 11212
rect 16580 11169 16589 11203
rect 16589 11169 16623 11203
rect 16623 11169 16632 11203
rect 16580 11160 16632 11169
rect 12440 11135 12492 11144
rect 10416 11067 10468 11076
rect 10416 11033 10425 11067
rect 10425 11033 10459 11067
rect 10459 11033 10468 11067
rect 10416 11024 10468 11033
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 12440 11092 12492 11101
rect 12532 11135 12584 11144
rect 12532 11101 12541 11135
rect 12541 11101 12575 11135
rect 12575 11101 12584 11135
rect 12532 11092 12584 11101
rect 12992 11135 13044 11144
rect 12992 11101 13004 11135
rect 13004 11101 13038 11135
rect 13038 11101 13044 11135
rect 12992 11092 13044 11101
rect 13268 11135 13320 11144
rect 13268 11101 13277 11135
rect 13277 11101 13311 11135
rect 13311 11101 13320 11135
rect 13268 11092 13320 11101
rect 13452 11092 13504 11144
rect 14648 11092 14700 11144
rect 16948 11203 17000 11212
rect 16948 11169 16957 11203
rect 16957 11169 16991 11203
rect 16991 11169 17000 11203
rect 16948 11160 17000 11169
rect 17224 11296 17276 11348
rect 18788 11339 18840 11348
rect 18788 11305 18797 11339
rect 18797 11305 18831 11339
rect 18831 11305 18840 11339
rect 18788 11296 18840 11305
rect 19248 11296 19300 11348
rect 21088 11296 21140 11348
rect 21272 11296 21324 11348
rect 21364 11228 21416 11280
rect 18328 11160 18380 11212
rect 19248 11203 19300 11212
rect 19248 11169 19257 11203
rect 19257 11169 19291 11203
rect 19291 11169 19300 11203
rect 19248 11160 19300 11169
rect 19984 11203 20036 11212
rect 19984 11169 19993 11203
rect 19993 11169 20027 11203
rect 20027 11169 20036 11203
rect 19984 11160 20036 11169
rect 20628 11160 20680 11212
rect 22284 11228 22336 11280
rect 22836 11339 22888 11348
rect 22836 11305 22851 11339
rect 22851 11305 22885 11339
rect 22885 11305 22888 11339
rect 22836 11296 22888 11305
rect 24400 11339 24452 11348
rect 24400 11305 24409 11339
rect 24409 11305 24443 11339
rect 24443 11305 24452 11339
rect 24400 11296 24452 11305
rect 24492 11296 24544 11348
rect 29368 11296 29420 11348
rect 25320 11228 25372 11280
rect 26240 11228 26292 11280
rect 22468 11160 22520 11212
rect 22928 11160 22980 11212
rect 23204 11160 23256 11212
rect 24860 11160 24912 11212
rect 9956 10999 10008 11008
rect 9956 10965 9965 10999
rect 9965 10965 9999 10999
rect 9999 10965 10008 10999
rect 9956 10956 10008 10965
rect 10140 10999 10192 11008
rect 10140 10965 10149 10999
rect 10149 10965 10183 10999
rect 10183 10965 10192 10999
rect 10140 10956 10192 10965
rect 11060 11024 11112 11076
rect 17132 11092 17184 11144
rect 17316 11135 17368 11144
rect 17316 11101 17318 11135
rect 17318 11101 17368 11135
rect 17316 11092 17368 11101
rect 20536 11092 20588 11144
rect 23296 11092 23348 11144
rect 23756 11092 23808 11144
rect 24952 11092 25004 11144
rect 25504 11092 25556 11144
rect 25872 11160 25924 11212
rect 26148 11160 26200 11212
rect 12164 10956 12216 11008
rect 12256 10956 12308 11008
rect 14832 11024 14884 11076
rect 15476 11024 15528 11076
rect 15752 11067 15804 11076
rect 15752 11033 15761 11067
rect 15761 11033 15795 11067
rect 15795 11033 15804 11067
rect 15752 11024 15804 11033
rect 16856 11024 16908 11076
rect 18420 11024 18472 11076
rect 22376 11024 22428 11076
rect 26608 11092 26660 11144
rect 27896 11160 27948 11212
rect 28448 11160 28500 11212
rect 28908 11203 28960 11212
rect 28908 11169 28917 11203
rect 28917 11169 28951 11203
rect 28951 11169 28960 11203
rect 28908 11160 28960 11169
rect 27344 11092 27396 11144
rect 27528 11092 27580 11144
rect 14372 10999 14424 11008
rect 14372 10965 14381 10999
rect 14381 10965 14415 10999
rect 14415 10965 14424 10999
rect 14372 10956 14424 10965
rect 16948 10956 17000 11008
rect 19984 10956 20036 11008
rect 22008 10956 22060 11008
rect 22100 10956 22152 11008
rect 22744 10956 22796 11008
rect 28080 11024 28132 11076
rect 30012 11067 30064 11076
rect 30012 11033 30021 11067
rect 30021 11033 30055 11067
rect 30055 11033 30064 11067
rect 30012 11024 30064 11033
rect 24952 10956 25004 11008
rect 25320 10999 25372 11008
rect 25320 10965 25329 10999
rect 25329 10965 25363 10999
rect 25363 10965 25372 10999
rect 25320 10956 25372 10965
rect 4193 10854 4245 10906
rect 4257 10854 4309 10906
rect 4321 10854 4373 10906
rect 4385 10854 4437 10906
rect 4449 10854 4501 10906
rect 11783 10854 11835 10906
rect 11847 10854 11899 10906
rect 11911 10854 11963 10906
rect 11975 10854 12027 10906
rect 12039 10854 12091 10906
rect 19373 10854 19425 10906
rect 19437 10854 19489 10906
rect 19501 10854 19553 10906
rect 19565 10854 19617 10906
rect 19629 10854 19681 10906
rect 26963 10854 27015 10906
rect 27027 10854 27079 10906
rect 27091 10854 27143 10906
rect 27155 10854 27207 10906
rect 27219 10854 27271 10906
rect 5816 10752 5868 10804
rect 6092 10752 6144 10804
rect 6644 10752 6696 10804
rect 1124 10616 1176 10668
rect 2136 10616 2188 10668
rect 5448 10616 5500 10668
rect 1584 10548 1636 10600
rect 3332 10548 3384 10600
rect 4896 10548 4948 10600
rect 1400 10455 1452 10464
rect 1400 10421 1415 10455
rect 1415 10421 1449 10455
rect 1449 10421 1452 10455
rect 1400 10412 1452 10421
rect 1676 10412 1728 10464
rect 3976 10412 4028 10464
rect 5632 10548 5684 10600
rect 5908 10591 5960 10600
rect 5908 10557 5910 10591
rect 5910 10557 5960 10591
rect 5908 10548 5960 10557
rect 6276 10591 6328 10600
rect 6276 10557 6285 10591
rect 6285 10557 6319 10591
rect 6319 10557 6328 10591
rect 6276 10548 6328 10557
rect 6552 10548 6604 10600
rect 8944 10684 8996 10736
rect 12992 10752 13044 10804
rect 14556 10752 14608 10804
rect 14648 10752 14700 10804
rect 12900 10684 12952 10736
rect 13360 10684 13412 10736
rect 9036 10616 9088 10668
rect 9312 10616 9364 10668
rect 8760 10548 8812 10600
rect 9128 10548 9180 10600
rect 9404 10548 9456 10600
rect 9864 10616 9916 10668
rect 10692 10616 10744 10668
rect 13820 10659 13872 10668
rect 13820 10625 13829 10659
rect 13829 10625 13863 10659
rect 13863 10625 13872 10659
rect 13820 10616 13872 10625
rect 14372 10616 14424 10668
rect 7656 10523 7708 10532
rect 7656 10489 7665 10523
rect 7665 10489 7699 10523
rect 7699 10489 7708 10523
rect 7656 10480 7708 10489
rect 7748 10480 7800 10532
rect 11980 10548 12032 10600
rect 12256 10523 12308 10532
rect 12256 10489 12265 10523
rect 12265 10489 12299 10523
rect 12299 10489 12308 10523
rect 12256 10480 12308 10489
rect 12900 10591 12952 10600
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 13728 10591 13780 10600
rect 13728 10557 13737 10591
rect 13737 10557 13771 10591
rect 13771 10557 13780 10591
rect 13728 10548 13780 10557
rect 14096 10548 14148 10600
rect 16120 10548 16172 10600
rect 22744 10795 22796 10804
rect 22744 10761 22753 10795
rect 22753 10761 22787 10795
rect 22787 10761 22796 10795
rect 22744 10752 22796 10761
rect 24492 10752 24544 10804
rect 25964 10752 26016 10804
rect 19800 10684 19852 10736
rect 23572 10684 23624 10736
rect 16580 10616 16632 10668
rect 17500 10616 17552 10668
rect 22744 10616 22796 10668
rect 16488 10548 16540 10600
rect 17776 10548 17828 10600
rect 6092 10412 6144 10464
rect 6552 10412 6604 10464
rect 7564 10412 7616 10464
rect 9956 10412 10008 10464
rect 10048 10455 10100 10464
rect 10048 10421 10063 10455
rect 10063 10421 10097 10455
rect 10097 10421 10100 10455
rect 10048 10412 10100 10421
rect 11612 10412 11664 10464
rect 13912 10412 13964 10464
rect 16028 10455 16080 10464
rect 16028 10421 16037 10455
rect 16037 10421 16071 10455
rect 16071 10421 16080 10455
rect 16028 10412 16080 10421
rect 18512 10523 18564 10532
rect 18512 10489 18521 10523
rect 18521 10489 18555 10523
rect 18555 10489 18564 10523
rect 18512 10480 18564 10489
rect 19984 10591 20036 10600
rect 19984 10557 19993 10591
rect 19993 10557 20027 10591
rect 20027 10557 20036 10591
rect 19984 10548 20036 10557
rect 20352 10591 20404 10600
rect 20352 10557 20354 10591
rect 20354 10557 20404 10591
rect 20352 10548 20404 10557
rect 20720 10591 20772 10600
rect 20720 10557 20729 10591
rect 20729 10557 20763 10591
rect 20763 10557 20772 10591
rect 20720 10548 20772 10557
rect 21364 10548 21416 10600
rect 22652 10548 22704 10600
rect 23204 10548 23256 10600
rect 24308 10659 24360 10668
rect 24308 10625 24320 10659
rect 24320 10625 24354 10659
rect 24354 10625 24360 10659
rect 24308 10616 24360 10625
rect 23848 10591 23900 10600
rect 23848 10557 23857 10591
rect 23857 10557 23891 10591
rect 23891 10557 23900 10591
rect 23848 10548 23900 10557
rect 24216 10591 24268 10600
rect 24216 10557 24218 10591
rect 24218 10557 24268 10591
rect 24216 10548 24268 10557
rect 24584 10591 24636 10600
rect 24584 10557 24593 10591
rect 24593 10557 24627 10591
rect 24627 10557 24636 10591
rect 24584 10548 24636 10557
rect 25044 10548 25096 10600
rect 25320 10548 25372 10600
rect 26148 10591 26200 10600
rect 26148 10557 26157 10591
rect 26157 10557 26191 10591
rect 26191 10557 26200 10591
rect 26148 10548 26200 10557
rect 26240 10548 26292 10600
rect 29276 10616 29328 10668
rect 16672 10412 16724 10464
rect 17040 10412 17092 10464
rect 18328 10412 18380 10464
rect 19064 10412 19116 10464
rect 19156 10455 19208 10464
rect 19156 10421 19165 10455
rect 19165 10421 19199 10455
rect 19199 10421 19208 10455
rect 19156 10412 19208 10421
rect 20444 10412 20496 10464
rect 21732 10412 21784 10464
rect 24584 10412 24636 10464
rect 25688 10455 25740 10464
rect 25688 10421 25697 10455
rect 25697 10421 25731 10455
rect 25731 10421 25740 10455
rect 25688 10412 25740 10421
rect 27712 10412 27764 10464
rect 28172 10455 28224 10464
rect 28172 10421 28181 10455
rect 28181 10421 28215 10455
rect 28215 10421 28224 10455
rect 28172 10412 28224 10421
rect 28540 10455 28592 10464
rect 28540 10421 28549 10455
rect 28549 10421 28583 10455
rect 28583 10421 28592 10455
rect 28540 10412 28592 10421
rect 28724 10480 28776 10532
rect 28908 10412 28960 10464
rect 29276 10455 29328 10464
rect 29276 10421 29285 10455
rect 29285 10421 29319 10455
rect 29319 10421 29328 10455
rect 29276 10412 29328 10421
rect 29920 10480 29972 10532
rect 29644 10412 29696 10464
rect 30104 10412 30156 10464
rect 7988 10310 8040 10362
rect 8052 10310 8104 10362
rect 8116 10310 8168 10362
rect 8180 10310 8232 10362
rect 8244 10310 8296 10362
rect 15578 10310 15630 10362
rect 15642 10310 15694 10362
rect 15706 10310 15758 10362
rect 15770 10310 15822 10362
rect 15834 10310 15886 10362
rect 23168 10310 23220 10362
rect 23232 10310 23284 10362
rect 23296 10310 23348 10362
rect 23360 10310 23412 10362
rect 23424 10310 23476 10362
rect 30758 10310 30810 10362
rect 30822 10310 30874 10362
rect 30886 10310 30938 10362
rect 30950 10310 31002 10362
rect 31014 10310 31066 10362
rect 664 10208 716 10260
rect 1400 10208 1452 10260
rect 2964 10208 3016 10260
rect 3700 10208 3752 10260
rect 3976 10208 4028 10260
rect 6460 10208 6512 10260
rect 7472 10208 7524 10260
rect 8944 10208 8996 10260
rect 9312 10208 9364 10260
rect 9496 10208 9548 10260
rect 11612 10251 11664 10260
rect 11612 10217 11627 10251
rect 11627 10217 11661 10251
rect 11661 10217 11664 10251
rect 11612 10208 11664 10217
rect 11980 10208 12032 10260
rect 14096 10208 14148 10260
rect 5448 10183 5500 10192
rect 5448 10149 5457 10183
rect 5457 10149 5491 10183
rect 5491 10149 5500 10183
rect 5448 10140 5500 10149
rect 1124 10115 1176 10124
rect 1124 10081 1133 10115
rect 1133 10081 1167 10115
rect 1167 10081 1176 10115
rect 1124 10072 1176 10081
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 3056 9868 3108 9920
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 3884 10072 3936 10124
rect 6092 10140 6144 10192
rect 17500 10208 17552 10260
rect 20720 10208 20772 10260
rect 21180 10208 21232 10260
rect 18972 10140 19024 10192
rect 5724 10004 5776 10056
rect 6460 10047 6512 10056
rect 6460 10013 6469 10047
rect 6469 10013 6503 10047
rect 6503 10013 6512 10047
rect 6460 10004 6512 10013
rect 7012 10004 7064 10056
rect 7564 10004 7616 10056
rect 9036 10004 9088 10056
rect 10140 10072 10192 10124
rect 10968 10072 11020 10124
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 12256 10072 12308 10124
rect 13820 10115 13872 10124
rect 13820 10081 13829 10115
rect 13829 10081 13863 10115
rect 13863 10081 13872 10115
rect 13820 10072 13872 10081
rect 14464 10072 14516 10124
rect 14556 10115 14608 10124
rect 14556 10081 14565 10115
rect 14565 10081 14599 10115
rect 14599 10081 14608 10115
rect 14556 10072 14608 10081
rect 12532 10004 12584 10056
rect 16856 10072 16908 10124
rect 18604 10072 18656 10124
rect 19156 10072 19208 10124
rect 21364 10140 21416 10192
rect 20628 10072 20680 10124
rect 16948 10004 17000 10056
rect 18788 10004 18840 10056
rect 20444 10004 20496 10056
rect 21088 10072 21140 10124
rect 21732 10047 21784 10056
rect 21732 10013 21744 10047
rect 21744 10013 21778 10047
rect 21778 10013 21784 10047
rect 21732 10004 21784 10013
rect 22008 10115 22060 10124
rect 22008 10081 22017 10115
rect 22017 10081 22051 10115
rect 22051 10081 22060 10115
rect 22008 10072 22060 10081
rect 23020 10208 23072 10260
rect 25044 10208 25096 10260
rect 25688 10208 25740 10260
rect 25872 10208 25924 10260
rect 28264 10140 28316 10192
rect 11060 9868 11112 9920
rect 12256 9868 12308 9920
rect 12348 9868 12400 9920
rect 15016 9868 15068 9920
rect 16764 9868 16816 9920
rect 18144 9868 18196 9920
rect 20720 9868 20772 9920
rect 20812 9911 20864 9920
rect 20812 9877 20821 9911
rect 20821 9877 20855 9911
rect 20855 9877 20864 9911
rect 20812 9868 20864 9877
rect 21916 9868 21968 9920
rect 24492 10004 24544 10056
rect 25136 10004 25188 10056
rect 26148 10072 26200 10124
rect 28356 10072 28408 10124
rect 28448 10072 28500 10124
rect 26056 10004 26108 10056
rect 26240 10004 26292 10056
rect 26884 10047 26936 10056
rect 26884 10013 26896 10047
rect 26896 10013 26930 10047
rect 26930 10013 26936 10047
rect 26884 10004 26936 10013
rect 25320 9936 25372 9988
rect 25044 9868 25096 9920
rect 25964 9868 26016 9920
rect 26700 9868 26752 9920
rect 28264 9911 28316 9920
rect 28264 9877 28273 9911
rect 28273 9877 28307 9911
rect 28307 9877 28316 9911
rect 28264 9868 28316 9877
rect 28908 9868 28960 9920
rect 30104 9868 30156 9920
rect 4193 9766 4245 9818
rect 4257 9766 4309 9818
rect 4321 9766 4373 9818
rect 4385 9766 4437 9818
rect 4449 9766 4501 9818
rect 11783 9766 11835 9818
rect 11847 9766 11899 9818
rect 11911 9766 11963 9818
rect 11975 9766 12027 9818
rect 12039 9766 12091 9818
rect 19373 9766 19425 9818
rect 19437 9766 19489 9818
rect 19501 9766 19553 9818
rect 19565 9766 19617 9818
rect 19629 9766 19681 9818
rect 26963 9766 27015 9818
rect 27027 9766 27079 9818
rect 27091 9766 27143 9818
rect 27155 9766 27207 9818
rect 27219 9766 27271 9818
rect 848 9664 900 9716
rect 1860 9664 1912 9716
rect 2688 9664 2740 9716
rect 3056 9664 3108 9716
rect 5264 9664 5316 9716
rect 6276 9664 6328 9716
rect 6644 9664 6696 9716
rect 2780 9596 2832 9648
rect 1124 9528 1176 9580
rect 3240 9596 3292 9648
rect 9128 9664 9180 9716
rect 8392 9596 8444 9648
rect 10968 9707 11020 9716
rect 10968 9673 10977 9707
rect 10977 9673 11011 9707
rect 11011 9673 11020 9707
rect 10968 9664 11020 9673
rect 13912 9664 13964 9716
rect 16120 9707 16172 9716
rect 16120 9673 16129 9707
rect 16129 9673 16163 9707
rect 16163 9673 16172 9707
rect 16120 9664 16172 9673
rect 16764 9664 16816 9716
rect 17040 9664 17092 9716
rect 6368 9528 6420 9580
rect 6920 9528 6972 9580
rect 9312 9571 9364 9580
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 3332 9460 3384 9512
rect 3976 9503 4028 9512
rect 3976 9469 3978 9503
rect 3978 9469 4028 9503
rect 3976 9460 4028 9469
rect 4344 9503 4396 9512
rect 4344 9469 4353 9503
rect 4353 9469 4387 9503
rect 4387 9469 4396 9503
rect 4344 9460 4396 9469
rect 6460 9460 6512 9512
rect 7104 9460 7156 9512
rect 8484 9460 8536 9512
rect 9036 9460 9088 9512
rect 9312 9537 9314 9571
rect 9314 9537 9364 9571
rect 9312 9528 9364 9537
rect 9496 9528 9548 9580
rect 10416 9528 10468 9580
rect 11060 9528 11112 9580
rect 14096 9571 14148 9580
rect 5448 9392 5500 9444
rect 8760 9392 8812 9444
rect 1400 9367 1452 9376
rect 1400 9333 1415 9367
rect 1415 9333 1449 9367
rect 1449 9333 1452 9367
rect 1400 9324 1452 9333
rect 2044 9324 2096 9376
rect 2964 9324 3016 9376
rect 4252 9324 4304 9376
rect 5264 9324 5316 9376
rect 7472 9324 7524 9376
rect 9588 9324 9640 9376
rect 11152 9503 11204 9512
rect 11152 9469 11161 9503
rect 11161 9469 11195 9503
rect 11195 9469 11204 9503
rect 11152 9460 11204 9469
rect 10508 9392 10560 9444
rect 11888 9503 11940 9512
rect 11888 9469 11897 9503
rect 11897 9469 11931 9503
rect 11931 9469 11940 9503
rect 11888 9460 11940 9469
rect 11244 9324 11296 9376
rect 11612 9367 11664 9376
rect 11612 9333 11627 9367
rect 11627 9333 11661 9367
rect 11661 9333 11664 9367
rect 11612 9324 11664 9333
rect 12624 9324 12676 9376
rect 14096 9537 14098 9571
rect 14098 9537 14148 9571
rect 14096 9528 14148 9537
rect 14924 9528 14976 9580
rect 19892 9664 19944 9716
rect 20444 9664 20496 9716
rect 18052 9596 18104 9648
rect 20536 9639 20588 9648
rect 20536 9605 20545 9639
rect 20545 9605 20579 9639
rect 20579 9605 20588 9639
rect 20536 9596 20588 9605
rect 22744 9707 22796 9716
rect 22744 9673 22753 9707
rect 22753 9673 22787 9707
rect 22787 9673 22796 9707
rect 22744 9664 22796 9673
rect 23848 9664 23900 9716
rect 26884 9664 26936 9716
rect 27712 9664 27764 9716
rect 19156 9571 19208 9580
rect 19156 9537 19168 9571
rect 19168 9537 19202 9571
rect 19202 9537 19208 9571
rect 19156 9528 19208 9537
rect 20720 9528 20772 9580
rect 13820 9460 13872 9512
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 15476 9460 15528 9512
rect 16396 9503 16448 9512
rect 16396 9469 16405 9503
rect 16405 9469 16439 9503
rect 16439 9469 16448 9503
rect 16396 9460 16448 9469
rect 18328 9460 18380 9512
rect 18052 9392 18104 9444
rect 19800 9460 19852 9512
rect 20812 9460 20864 9512
rect 21088 9528 21140 9580
rect 21456 9528 21508 9580
rect 22560 9528 22612 9580
rect 22008 9460 22060 9512
rect 28356 9596 28408 9648
rect 24768 9528 24820 9580
rect 24860 9571 24912 9580
rect 24860 9537 24872 9571
rect 24872 9537 24906 9571
rect 24906 9537 24912 9571
rect 24860 9528 24912 9537
rect 24124 9460 24176 9512
rect 25412 9460 25464 9512
rect 15108 9324 15160 9376
rect 15384 9324 15436 9376
rect 17040 9324 17092 9376
rect 23664 9392 23716 9444
rect 28540 9528 28592 9580
rect 26056 9460 26108 9512
rect 26700 9460 26752 9512
rect 29184 9503 29236 9512
rect 29184 9469 29193 9503
rect 29193 9469 29227 9503
rect 29227 9469 29236 9503
rect 29184 9460 29236 9469
rect 25872 9392 25924 9444
rect 29000 9392 29052 9444
rect 21548 9324 21600 9376
rect 23756 9324 23808 9376
rect 23940 9324 23992 9376
rect 24124 9367 24176 9376
rect 24124 9333 24133 9367
rect 24133 9333 24167 9367
rect 24167 9333 24176 9367
rect 24124 9324 24176 9333
rect 24308 9324 24360 9376
rect 24400 9324 24452 9376
rect 26884 9324 26936 9376
rect 27344 9324 27396 9376
rect 29460 9324 29512 9376
rect 7988 9222 8040 9274
rect 8052 9222 8104 9274
rect 8116 9222 8168 9274
rect 8180 9222 8232 9274
rect 8244 9222 8296 9274
rect 15578 9222 15630 9274
rect 15642 9222 15694 9274
rect 15706 9222 15758 9274
rect 15770 9222 15822 9274
rect 15834 9222 15886 9274
rect 23168 9222 23220 9274
rect 23232 9222 23284 9274
rect 23296 9222 23348 9274
rect 23360 9222 23412 9274
rect 23424 9222 23476 9274
rect 30758 9222 30810 9274
rect 30822 9222 30874 9274
rect 30886 9222 30938 9274
rect 30950 9222 31002 9274
rect 31014 9222 31066 9274
rect 848 9163 900 9172
rect 848 9129 857 9163
rect 857 9129 891 9163
rect 891 9129 900 9163
rect 848 9120 900 9129
rect 756 8984 808 9036
rect 4252 9120 4304 9172
rect 4344 9120 4396 9172
rect 4896 9163 4948 9172
rect 4896 9129 4905 9163
rect 4905 9129 4939 9163
rect 4939 9129 4948 9163
rect 4896 9120 4948 9129
rect 5172 9163 5224 9172
rect 5172 9129 5181 9163
rect 5181 9129 5215 9163
rect 5215 9129 5224 9163
rect 5172 9120 5224 9129
rect 6184 9120 6236 9172
rect 7104 9120 7156 9172
rect 7472 9120 7524 9172
rect 7656 9120 7708 9172
rect 8116 9120 8168 9172
rect 9496 9163 9548 9172
rect 9496 9129 9505 9163
rect 9505 9129 9539 9163
rect 9539 9129 9548 9163
rect 9496 9120 9548 9129
rect 10508 9120 10560 9172
rect 11888 9120 11940 9172
rect 14096 9120 14148 9172
rect 14464 9120 14516 9172
rect 16396 9120 16448 9172
rect 17040 9120 17092 9172
rect 1400 9052 1452 9104
rect 2044 8984 2096 9036
rect 2320 8984 2372 9036
rect 3608 8984 3660 9036
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 2872 8916 2924 8968
rect 2964 8959 3016 8968
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 2964 8916 3016 8925
rect 3056 8916 3108 8968
rect 4068 8916 4120 8968
rect 5356 9027 5408 9036
rect 5356 8993 5365 9027
rect 5365 8993 5399 9027
rect 5399 8993 5408 9027
rect 5356 8984 5408 8993
rect 6092 8916 6144 8968
rect 6644 9027 6696 9036
rect 6644 8993 6653 9027
rect 6653 8993 6687 9027
rect 6687 8993 6696 9027
rect 6644 8984 6696 8993
rect 6920 9027 6972 9036
rect 6920 8993 6929 9027
rect 6929 8993 6963 9027
rect 6963 8993 6972 9027
rect 6920 8984 6972 8993
rect 7288 8984 7340 9036
rect 7472 8984 7524 9036
rect 7656 9027 7708 9036
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 9404 9052 9456 9104
rect 8208 8984 8260 9036
rect 6460 8916 6512 8968
rect 8116 8959 8168 8968
rect 8116 8925 8128 8959
rect 8128 8925 8162 8959
rect 8162 8925 8168 8959
rect 8116 8916 8168 8925
rect 8760 8916 8812 8968
rect 9496 8916 9548 8968
rect 10232 8984 10284 9036
rect 11244 9052 11296 9104
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 2780 8780 2832 8832
rect 3332 8780 3384 8832
rect 5356 8780 5408 8832
rect 5632 8780 5684 8832
rect 5816 8823 5868 8832
rect 5816 8789 5825 8823
rect 5825 8789 5859 8823
rect 5859 8789 5868 8823
rect 5816 8780 5868 8789
rect 6000 8780 6052 8832
rect 6460 8823 6512 8832
rect 6460 8789 6469 8823
rect 6469 8789 6503 8823
rect 6503 8789 6512 8823
rect 6460 8780 6512 8789
rect 6828 8780 6880 8832
rect 6920 8780 6972 8832
rect 7104 8780 7156 8832
rect 9772 8848 9824 8900
rect 13820 9027 13872 9036
rect 13820 8993 13829 9027
rect 13829 8993 13863 9027
rect 13863 8993 13872 9027
rect 13820 8984 13872 8993
rect 15936 9052 15988 9104
rect 18052 9120 18104 9172
rect 16028 8984 16080 9036
rect 11152 8959 11204 8968
rect 11152 8925 11161 8959
rect 11161 8925 11195 8959
rect 11195 8925 11204 8959
rect 11152 8916 11204 8925
rect 11520 8959 11572 8968
rect 11520 8925 11522 8959
rect 11522 8925 11572 8959
rect 11520 8916 11572 8925
rect 11704 8916 11756 8968
rect 14004 8916 14056 8968
rect 14372 8916 14424 8968
rect 15476 8916 15528 8968
rect 16856 9027 16908 9036
rect 16856 8993 16865 9027
rect 16865 8993 16899 9027
rect 16899 8993 16908 9027
rect 16856 8984 16908 8993
rect 21548 9120 21600 9172
rect 20812 9052 20864 9104
rect 18052 8984 18104 9036
rect 18144 9027 18196 9036
rect 18144 8993 18153 9027
rect 18153 8993 18187 9027
rect 18187 8993 18196 9027
rect 18144 8984 18196 8993
rect 22928 9120 22980 9172
rect 23756 9120 23808 9172
rect 24216 9120 24268 9172
rect 24860 9120 24912 9172
rect 25412 9120 25464 9172
rect 26700 9120 26752 9172
rect 26884 9163 26936 9172
rect 26884 9129 26899 9163
rect 26899 9129 26933 9163
rect 26933 9129 26936 9163
rect 26884 9120 26936 9129
rect 27528 9120 27580 9172
rect 30472 9120 30524 9172
rect 26056 9052 26108 9104
rect 20168 8916 20220 8968
rect 11060 8780 11112 8832
rect 18972 8848 19024 8900
rect 12256 8780 12308 8832
rect 12992 8823 13044 8832
rect 12992 8789 13001 8823
rect 13001 8789 13035 8823
rect 13035 8789 13044 8823
rect 12992 8780 13044 8789
rect 13360 8780 13412 8832
rect 14372 8780 14424 8832
rect 16028 8780 16080 8832
rect 18788 8780 18840 8832
rect 20628 8780 20680 8832
rect 20720 8780 20772 8832
rect 21824 8916 21876 8968
rect 21916 8916 21968 8968
rect 24216 9027 24268 9036
rect 24216 8993 24225 9027
rect 24225 8993 24259 9027
rect 24259 8993 24268 9027
rect 24216 8984 24268 8993
rect 23664 8916 23716 8968
rect 24032 8916 24084 8968
rect 23480 8780 23532 8832
rect 23756 8780 23808 8832
rect 25964 8984 26016 9036
rect 26516 8984 26568 9036
rect 28632 9027 28684 9036
rect 28632 8993 28641 9027
rect 28641 8993 28675 9027
rect 28675 8993 28684 9027
rect 28632 8984 28684 8993
rect 30012 8984 30064 9036
rect 26700 8916 26752 8968
rect 26884 8959 26936 8968
rect 26884 8925 26896 8959
rect 26896 8925 26930 8959
rect 26930 8925 26936 8959
rect 26884 8916 26936 8925
rect 27344 8916 27396 8968
rect 28540 8916 28592 8968
rect 29000 8780 29052 8832
rect 4193 8678 4245 8730
rect 4257 8678 4309 8730
rect 4321 8678 4373 8730
rect 4385 8678 4437 8730
rect 4449 8678 4501 8730
rect 11783 8678 11835 8730
rect 11847 8678 11899 8730
rect 11911 8678 11963 8730
rect 11975 8678 12027 8730
rect 12039 8678 12091 8730
rect 19373 8678 19425 8730
rect 19437 8678 19489 8730
rect 19501 8678 19553 8730
rect 19565 8678 19617 8730
rect 19629 8678 19681 8730
rect 26963 8678 27015 8730
rect 27027 8678 27079 8730
rect 27091 8678 27143 8730
rect 27155 8678 27207 8730
rect 27219 8678 27271 8730
rect 1124 8576 1176 8628
rect 2872 8576 2924 8628
rect 3056 8508 3108 8560
rect 1216 8372 1268 8424
rect 1768 8372 1820 8424
rect 2136 8372 2188 8424
rect 2688 8372 2740 8424
rect 2780 8372 2832 8424
rect 3424 8440 3476 8492
rect 6644 8576 6696 8628
rect 7012 8576 7064 8628
rect 7564 8576 7616 8628
rect 7196 8508 7248 8560
rect 5356 8372 5408 8424
rect 5448 8372 5500 8424
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 3056 8347 3108 8356
rect 3056 8313 3065 8347
rect 3065 8313 3099 8347
rect 3099 8313 3108 8347
rect 3056 8304 3108 8313
rect 1400 8279 1452 8288
rect 1400 8245 1415 8279
rect 1415 8245 1449 8279
rect 1449 8245 1452 8279
rect 1400 8236 1452 8245
rect 2320 8236 2372 8288
rect 3332 8304 3384 8356
rect 6092 8440 6144 8492
rect 5908 8415 5960 8424
rect 5908 8381 5910 8415
rect 5910 8381 5960 8415
rect 5908 8372 5960 8381
rect 6184 8372 6236 8424
rect 8392 8372 8444 8424
rect 8852 8551 8904 8560
rect 8852 8517 8861 8551
rect 8861 8517 8895 8551
rect 8895 8517 8904 8551
rect 8852 8508 8904 8517
rect 9036 8508 9088 8560
rect 10048 8576 10100 8628
rect 10784 8576 10836 8628
rect 11704 8619 11756 8628
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 19248 8576 19300 8628
rect 9312 8508 9364 8560
rect 9496 8508 9548 8560
rect 12164 8440 12216 8492
rect 12716 8440 12768 8492
rect 9404 8372 9456 8424
rect 9496 8372 9548 8424
rect 9680 8415 9732 8424
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 9680 8372 9732 8381
rect 9956 8372 10008 8424
rect 13636 8440 13688 8492
rect 14096 8483 14148 8492
rect 3240 8236 3292 8288
rect 5816 8236 5868 8288
rect 6184 8236 6236 8288
rect 7748 8279 7800 8288
rect 7748 8245 7757 8279
rect 7757 8245 7791 8279
rect 7791 8245 7800 8279
rect 7748 8236 7800 8245
rect 8852 8236 8904 8288
rect 9404 8236 9456 8288
rect 11980 8236 12032 8288
rect 12256 8304 12308 8356
rect 13268 8372 13320 8424
rect 13820 8372 13872 8424
rect 14096 8449 14098 8483
rect 14098 8449 14148 8483
rect 14096 8440 14148 8449
rect 14188 8483 14240 8492
rect 14188 8449 14200 8483
rect 14200 8449 14234 8483
rect 14234 8449 14240 8483
rect 14188 8440 14240 8449
rect 14832 8440 14884 8492
rect 18604 8440 18656 8492
rect 15200 8372 15252 8424
rect 19248 8440 19300 8492
rect 18972 8372 19024 8424
rect 20812 8372 20864 8424
rect 21456 8415 21508 8424
rect 21456 8381 21465 8415
rect 21465 8381 21499 8415
rect 21499 8381 21508 8415
rect 21456 8372 21508 8381
rect 25872 8619 25924 8628
rect 25872 8585 25881 8619
rect 25881 8585 25915 8619
rect 25915 8585 25924 8619
rect 25872 8576 25924 8585
rect 26516 8576 26568 8628
rect 23480 8508 23532 8560
rect 25412 8508 25464 8560
rect 27344 8576 27396 8628
rect 27436 8576 27488 8628
rect 24400 8440 24452 8492
rect 23848 8415 23900 8424
rect 18052 8347 18104 8356
rect 18052 8313 18061 8347
rect 18061 8313 18095 8347
rect 18095 8313 18104 8347
rect 18052 8304 18104 8313
rect 20720 8304 20772 8356
rect 23848 8381 23857 8415
rect 23857 8381 23891 8415
rect 23891 8381 23900 8415
rect 23848 8372 23900 8381
rect 23940 8372 23992 8424
rect 25320 8372 25372 8424
rect 26608 8440 26660 8492
rect 27068 8483 27120 8492
rect 27068 8449 27070 8483
rect 27070 8449 27120 8483
rect 27068 8440 27120 8449
rect 28264 8440 28316 8492
rect 28724 8440 28776 8492
rect 23664 8304 23716 8356
rect 12440 8236 12492 8288
rect 12532 8236 12584 8288
rect 12716 8236 12768 8288
rect 13176 8279 13228 8288
rect 13176 8245 13185 8279
rect 13185 8245 13219 8279
rect 13219 8245 13228 8279
rect 13176 8236 13228 8245
rect 16396 8279 16448 8288
rect 16396 8245 16411 8279
rect 16411 8245 16445 8279
rect 16445 8245 16448 8279
rect 16396 8236 16448 8245
rect 18144 8279 18196 8288
rect 18144 8245 18153 8279
rect 18153 8245 18187 8279
rect 18187 8245 18196 8279
rect 18144 8236 18196 8245
rect 18788 8236 18840 8288
rect 20996 8236 21048 8288
rect 21456 8236 21508 8288
rect 21640 8236 21692 8288
rect 23756 8236 23808 8288
rect 24308 8279 24360 8288
rect 24308 8245 24323 8279
rect 24323 8245 24357 8279
rect 24357 8245 24360 8279
rect 24308 8236 24360 8245
rect 26792 8372 26844 8424
rect 29092 8415 29144 8424
rect 29092 8381 29101 8415
rect 29101 8381 29135 8415
rect 29135 8381 29144 8415
rect 29092 8372 29144 8381
rect 29552 8304 29604 8356
rect 29736 8304 29788 8356
rect 27804 8236 27856 8288
rect 29184 8279 29236 8288
rect 29184 8245 29193 8279
rect 29193 8245 29227 8279
rect 29227 8245 29236 8279
rect 29184 8236 29236 8245
rect 30012 8236 30064 8288
rect 7988 8134 8040 8186
rect 8052 8134 8104 8186
rect 8116 8134 8168 8186
rect 8180 8134 8232 8186
rect 8244 8134 8296 8186
rect 15578 8134 15630 8186
rect 15642 8134 15694 8186
rect 15706 8134 15758 8186
rect 15770 8134 15822 8186
rect 15834 8134 15886 8186
rect 23168 8134 23220 8186
rect 23232 8134 23284 8186
rect 23296 8134 23348 8186
rect 23360 8134 23412 8186
rect 23424 8134 23476 8186
rect 30758 8134 30810 8186
rect 30822 8134 30874 8186
rect 30886 8134 30938 8186
rect 30950 8134 31002 8186
rect 31014 8134 31066 8186
rect 1676 8032 1728 8084
rect 1032 7939 1084 7948
rect 1032 7905 1041 7939
rect 1041 7905 1075 7939
rect 1075 7905 1084 7939
rect 1032 7896 1084 7905
rect 6460 7964 6512 8016
rect 1400 7828 1452 7880
rect 3332 7939 3384 7948
rect 3332 7905 3341 7939
rect 3341 7905 3375 7939
rect 3375 7905 3384 7939
rect 3332 7896 3384 7905
rect 3516 7939 3568 7948
rect 3516 7905 3525 7939
rect 3525 7905 3559 7939
rect 3559 7905 3568 7939
rect 3516 7896 3568 7905
rect 7104 7896 7156 7948
rect 7656 7896 7708 7948
rect 1952 7871 2004 7880
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 3700 7828 3752 7880
rect 4160 7828 4212 7880
rect 5816 7828 5868 7880
rect 6368 7828 6420 7880
rect 8208 7828 8260 7880
rect 1216 7692 1268 7744
rect 3332 7692 3384 7744
rect 4068 7692 4120 7744
rect 4160 7692 4212 7744
rect 5908 7692 5960 7744
rect 6736 7692 6788 7744
rect 6920 7692 6972 7744
rect 8760 7896 8812 7948
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 11980 7896 12032 7948
rect 12716 7896 12768 7948
rect 18788 8075 18840 8084
rect 18788 8041 18803 8075
rect 18803 8041 18837 8075
rect 18837 8041 18840 8075
rect 18788 8032 18840 8041
rect 20168 8075 20220 8084
rect 20168 8041 20177 8075
rect 20177 8041 20211 8075
rect 20211 8041 20220 8075
rect 20168 8032 20220 8041
rect 20812 8075 20864 8084
rect 20812 8041 20821 8075
rect 20821 8041 20855 8075
rect 20855 8041 20864 8075
rect 20812 8032 20864 8041
rect 21824 8032 21876 8084
rect 23756 8032 23808 8084
rect 27068 8032 27120 8084
rect 27988 8032 28040 8084
rect 28816 8032 28868 8084
rect 13912 7896 13964 7948
rect 8944 7828 8996 7880
rect 9128 7828 9180 7880
rect 9404 7871 9456 7880
rect 9404 7837 9413 7871
rect 9413 7837 9447 7871
rect 9447 7837 9456 7871
rect 9404 7828 9456 7837
rect 9588 7828 9640 7880
rect 11152 7692 11204 7744
rect 12992 7828 13044 7880
rect 13084 7828 13136 7880
rect 14464 7896 14516 7948
rect 18144 7896 18196 7948
rect 15016 7828 15068 7880
rect 15200 7828 15252 7880
rect 16304 7828 16356 7880
rect 16580 7871 16632 7880
rect 16580 7837 16592 7871
rect 16592 7837 16626 7871
rect 16626 7837 16632 7871
rect 16580 7828 16632 7837
rect 17500 7828 17552 7880
rect 20628 7896 20680 7948
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 19064 7871 19116 7880
rect 19064 7837 19073 7871
rect 19073 7837 19107 7871
rect 19107 7837 19116 7871
rect 19064 7828 19116 7837
rect 19156 7828 19208 7880
rect 22744 7964 22796 8016
rect 21640 7939 21692 7948
rect 21640 7905 21642 7939
rect 21642 7905 21692 7939
rect 21640 7896 21692 7905
rect 20904 7828 20956 7880
rect 21456 7828 21508 7880
rect 21916 7828 21968 7880
rect 21180 7760 21232 7812
rect 22744 7828 22796 7880
rect 23572 7896 23624 7948
rect 22836 7760 22888 7812
rect 23756 7828 23808 7880
rect 23940 7871 23992 7880
rect 23940 7837 23952 7871
rect 23952 7837 23986 7871
rect 23986 7837 23992 7871
rect 23940 7828 23992 7837
rect 24216 7871 24268 7880
rect 24216 7837 24225 7871
rect 24225 7837 24259 7871
rect 24259 7837 24268 7871
rect 24216 7828 24268 7837
rect 25688 7939 25740 7948
rect 25688 7905 25697 7939
rect 25697 7905 25731 7939
rect 25731 7905 25740 7939
rect 25688 7896 25740 7905
rect 26700 7896 26752 7948
rect 29276 7896 29328 7948
rect 30012 7939 30064 7948
rect 30012 7905 30021 7939
rect 30021 7905 30055 7939
rect 30055 7905 30064 7939
rect 30012 7896 30064 7905
rect 25872 7871 25924 7880
rect 25872 7837 25881 7871
rect 25881 7837 25915 7871
rect 25915 7837 25924 7871
rect 25872 7828 25924 7837
rect 25964 7828 26016 7880
rect 18972 7692 19024 7744
rect 20536 7735 20588 7744
rect 20536 7701 20545 7735
rect 20545 7701 20579 7735
rect 20579 7701 20588 7735
rect 20536 7692 20588 7701
rect 20628 7692 20680 7744
rect 23388 7692 23440 7744
rect 27436 7760 27488 7812
rect 25320 7735 25372 7744
rect 25320 7701 25329 7735
rect 25329 7701 25363 7735
rect 25363 7701 25372 7735
rect 25320 7692 25372 7701
rect 25504 7692 25556 7744
rect 25596 7692 25648 7744
rect 27344 7735 27396 7744
rect 27344 7701 27353 7735
rect 27353 7701 27387 7735
rect 27387 7701 27396 7735
rect 27344 7692 27396 7701
rect 27804 7828 27856 7880
rect 27896 7828 27948 7880
rect 28172 7828 28224 7880
rect 29368 7692 29420 7744
rect 29828 7735 29880 7744
rect 29828 7701 29837 7735
rect 29837 7701 29871 7735
rect 29871 7701 29880 7735
rect 29828 7692 29880 7701
rect 4193 7590 4245 7642
rect 4257 7590 4309 7642
rect 4321 7590 4373 7642
rect 4385 7590 4437 7642
rect 4449 7590 4501 7642
rect 11783 7590 11835 7642
rect 11847 7590 11899 7642
rect 11911 7590 11963 7642
rect 11975 7590 12027 7642
rect 12039 7590 12091 7642
rect 19373 7590 19425 7642
rect 19437 7590 19489 7642
rect 19501 7590 19553 7642
rect 19565 7590 19617 7642
rect 19629 7590 19681 7642
rect 26963 7590 27015 7642
rect 27027 7590 27079 7642
rect 27091 7590 27143 7642
rect 27155 7590 27207 7642
rect 27219 7590 27271 7642
rect 2412 7420 2464 7472
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 2964 7352 3016 7404
rect 10508 7420 10560 7472
rect 6552 7352 6604 7404
rect 7748 7352 7800 7404
rect 1216 7284 1268 7336
rect 2688 7284 2740 7336
rect 3516 7327 3568 7336
rect 3516 7293 3525 7327
rect 3525 7293 3559 7327
rect 3559 7293 3568 7327
rect 3516 7284 3568 7293
rect 5264 7284 5316 7336
rect 5724 7216 5776 7268
rect 1400 7191 1452 7200
rect 1400 7157 1415 7191
rect 1415 7157 1449 7191
rect 1449 7157 1452 7191
rect 1400 7148 1452 7157
rect 2780 7191 2832 7200
rect 2780 7157 2789 7191
rect 2789 7157 2823 7191
rect 2823 7157 2832 7191
rect 2780 7148 2832 7157
rect 3332 7148 3384 7200
rect 3976 7191 4028 7200
rect 3976 7157 3991 7191
rect 3991 7157 4025 7191
rect 4025 7157 4028 7191
rect 6184 7284 6236 7336
rect 8668 7352 8720 7404
rect 8760 7352 8812 7404
rect 13452 7488 13504 7540
rect 13728 7488 13780 7540
rect 11428 7352 11480 7404
rect 12348 7352 12400 7404
rect 12440 7352 12492 7404
rect 14372 7395 14424 7404
rect 14372 7361 14384 7395
rect 14384 7361 14418 7395
rect 14418 7361 14424 7395
rect 14372 7352 14424 7361
rect 14648 7395 14700 7404
rect 14648 7361 14657 7395
rect 14657 7361 14691 7395
rect 14691 7361 14700 7395
rect 14648 7352 14700 7361
rect 19800 7488 19852 7540
rect 20536 7488 20588 7540
rect 17960 7463 18012 7472
rect 17960 7429 17969 7463
rect 17969 7429 18003 7463
rect 18003 7429 18012 7463
rect 17960 7420 18012 7429
rect 9404 7327 9456 7336
rect 7564 7216 7616 7268
rect 8944 7216 8996 7268
rect 9404 7293 9406 7327
rect 9406 7293 9456 7327
rect 9404 7284 9456 7293
rect 10600 7284 10652 7336
rect 12716 7284 12768 7336
rect 13084 7284 13136 7336
rect 13912 7327 13964 7336
rect 13912 7293 13921 7327
rect 13921 7293 13955 7327
rect 13955 7293 13964 7327
rect 13912 7284 13964 7293
rect 14740 7284 14792 7336
rect 15108 7284 15160 7336
rect 16672 7352 16724 7404
rect 17040 7352 17092 7404
rect 18972 7352 19024 7404
rect 18604 7284 18656 7336
rect 20996 7284 21048 7336
rect 23388 7488 23440 7540
rect 24032 7488 24084 7540
rect 25320 7488 25372 7540
rect 26884 7488 26936 7540
rect 27896 7488 27948 7540
rect 28264 7488 28316 7540
rect 21640 7352 21692 7404
rect 21456 7327 21508 7336
rect 21456 7293 21465 7327
rect 21465 7293 21499 7327
rect 21499 7293 21508 7327
rect 21456 7284 21508 7293
rect 22192 7327 22244 7336
rect 22192 7293 22201 7327
rect 22201 7293 22235 7327
rect 22235 7293 22244 7327
rect 22192 7284 22244 7293
rect 3976 7148 4028 7157
rect 6368 7148 6420 7200
rect 6460 7148 6512 7200
rect 6736 7148 6788 7200
rect 9864 7148 9916 7200
rect 10876 7191 10928 7200
rect 10876 7157 10885 7191
rect 10885 7157 10919 7191
rect 10919 7157 10928 7191
rect 10876 7148 10928 7157
rect 12440 7148 12492 7200
rect 14004 7216 14056 7268
rect 13084 7191 13136 7200
rect 13084 7157 13093 7191
rect 13093 7157 13127 7191
rect 13127 7157 13136 7191
rect 13084 7148 13136 7157
rect 14280 7148 14332 7200
rect 14556 7148 14608 7200
rect 15292 7148 15344 7200
rect 16396 7148 16448 7200
rect 18788 7148 18840 7200
rect 19892 7148 19944 7200
rect 22652 7148 22704 7200
rect 23848 7395 23900 7404
rect 23848 7361 23857 7395
rect 23857 7361 23891 7395
rect 23891 7361 23900 7395
rect 23848 7352 23900 7361
rect 24124 7352 24176 7404
rect 28908 7420 28960 7472
rect 29460 7420 29512 7472
rect 28356 7352 28408 7404
rect 29000 7352 29052 7404
rect 25320 7284 25372 7336
rect 26056 7327 26108 7336
rect 26056 7293 26065 7327
rect 26065 7293 26099 7327
rect 26099 7293 26108 7327
rect 26056 7284 26108 7293
rect 26792 7327 26844 7336
rect 26792 7293 26801 7327
rect 26801 7293 26835 7327
rect 26835 7293 26844 7327
rect 26792 7284 26844 7293
rect 24124 7148 24176 7200
rect 24308 7191 24360 7200
rect 24308 7157 24323 7191
rect 24323 7157 24357 7191
rect 24357 7157 24360 7191
rect 24308 7148 24360 7157
rect 24492 7148 24544 7200
rect 25872 7148 25924 7200
rect 26884 7148 26936 7200
rect 27252 7148 27304 7200
rect 27896 7191 27948 7200
rect 27896 7157 27905 7191
rect 27905 7157 27939 7191
rect 27939 7157 27948 7191
rect 27896 7148 27948 7157
rect 28264 7148 28316 7200
rect 28540 7148 28592 7200
rect 29184 7148 29236 7200
rect 29276 7148 29328 7200
rect 7988 7046 8040 7098
rect 8052 7046 8104 7098
rect 8116 7046 8168 7098
rect 8180 7046 8232 7098
rect 8244 7046 8296 7098
rect 15578 7046 15630 7098
rect 15642 7046 15694 7098
rect 15706 7046 15758 7098
rect 15770 7046 15822 7098
rect 15834 7046 15886 7098
rect 23168 7046 23220 7098
rect 23232 7046 23284 7098
rect 23296 7046 23348 7098
rect 23360 7046 23412 7098
rect 23424 7046 23476 7098
rect 30758 7046 30810 7098
rect 30822 7046 30874 7098
rect 30886 7046 30938 7098
rect 30950 7046 31002 7098
rect 31014 7046 31066 7098
rect 1400 6944 1452 6996
rect 2688 6944 2740 6996
rect 1216 6808 1268 6860
rect 3424 6876 3476 6928
rect 5816 6987 5868 6996
rect 5816 6953 5825 6987
rect 5825 6953 5859 6987
rect 5859 6953 5868 6987
rect 5816 6944 5868 6953
rect 6460 6944 6512 6996
rect 9404 6944 9456 6996
rect 10508 6987 10560 6996
rect 10508 6953 10517 6987
rect 10517 6953 10551 6987
rect 10551 6953 10560 6987
rect 10508 6944 10560 6953
rect 10784 6876 10836 6928
rect 11980 6944 12032 6996
rect 3700 6851 3752 6860
rect 3700 6817 3702 6851
rect 3702 6817 3752 6851
rect 3700 6808 3752 6817
rect 5172 6808 5224 6860
rect 5448 6851 5500 6860
rect 5448 6817 5457 6851
rect 5457 6817 5491 6851
rect 5491 6817 5500 6851
rect 5448 6808 5500 6817
rect 5724 6808 5776 6860
rect 6184 6808 6236 6860
rect 1768 6740 1820 6792
rect 1124 6672 1176 6724
rect 1492 6604 1544 6656
rect 3516 6740 3568 6792
rect 6368 6808 6420 6860
rect 6000 6604 6052 6656
rect 6736 6740 6788 6792
rect 7012 6740 7064 6792
rect 7196 6851 7248 6860
rect 7196 6817 7205 6851
rect 7205 6817 7239 6851
rect 7239 6817 7248 6851
rect 7196 6808 7248 6817
rect 8760 6808 8812 6860
rect 9496 6808 9548 6860
rect 11152 6851 11204 6860
rect 11152 6817 11161 6851
rect 11161 6817 11195 6851
rect 11195 6817 11204 6851
rect 11152 6808 11204 6817
rect 11520 6851 11572 6860
rect 11520 6817 11529 6851
rect 11529 6817 11563 6851
rect 11563 6817 11572 6851
rect 11520 6808 11572 6817
rect 11612 6808 11664 6860
rect 12072 6851 12124 6860
rect 12072 6817 12081 6851
rect 12081 6817 12115 6851
rect 12115 6817 12124 6851
rect 12072 6808 12124 6817
rect 12900 6944 12952 6996
rect 14648 6944 14700 6996
rect 15108 6944 15160 6996
rect 16304 6944 16356 6996
rect 16396 6944 16448 6996
rect 14556 6919 14608 6928
rect 14556 6885 14565 6919
rect 14565 6885 14599 6919
rect 14599 6885 14608 6919
rect 14556 6876 14608 6885
rect 14924 6876 14976 6928
rect 12440 6851 12492 6860
rect 12440 6817 12442 6851
rect 12442 6817 12492 6851
rect 12440 6808 12492 6817
rect 13176 6808 13228 6860
rect 13268 6808 13320 6860
rect 8300 6715 8352 6724
rect 8300 6681 8309 6715
rect 8309 6681 8343 6715
rect 8343 6681 8352 6715
rect 8300 6672 8352 6681
rect 10600 6672 10652 6724
rect 11060 6672 11112 6724
rect 7932 6604 7984 6656
rect 8392 6604 8444 6656
rect 11612 6604 11664 6656
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 12624 6740 12676 6792
rect 13452 6740 13504 6792
rect 15752 6851 15804 6860
rect 15752 6817 15761 6851
rect 15761 6817 15795 6851
rect 15795 6817 15804 6851
rect 15752 6808 15804 6817
rect 15936 6808 15988 6860
rect 16304 6851 16356 6860
rect 16304 6817 16313 6851
rect 16313 6817 16347 6851
rect 16347 6817 16356 6851
rect 16304 6808 16356 6817
rect 16488 6808 16540 6860
rect 18972 6944 19024 6996
rect 21088 6944 21140 6996
rect 21548 6944 21600 6996
rect 23940 6987 23992 6996
rect 23940 6953 23949 6987
rect 23949 6953 23983 6987
rect 23983 6953 23992 6987
rect 23940 6944 23992 6953
rect 24124 6944 24176 6996
rect 22008 6876 22060 6928
rect 16764 6783 16816 6792
rect 16764 6749 16766 6783
rect 16766 6749 16816 6783
rect 14004 6672 14056 6724
rect 16764 6740 16816 6749
rect 17132 6783 17184 6792
rect 17132 6749 17141 6783
rect 17141 6749 17175 6783
rect 17175 6749 17184 6783
rect 17132 6740 17184 6749
rect 18236 6740 18288 6792
rect 18788 6740 18840 6792
rect 20720 6808 20772 6860
rect 20536 6740 20588 6792
rect 21364 6740 21416 6792
rect 21732 6851 21784 6860
rect 21732 6817 21741 6851
rect 21741 6817 21775 6851
rect 21775 6817 21784 6851
rect 21732 6808 21784 6817
rect 21824 6740 21876 6792
rect 21916 6783 21968 6792
rect 21916 6749 21925 6783
rect 21925 6749 21959 6783
rect 21959 6749 21968 6783
rect 21916 6740 21968 6749
rect 22376 6783 22428 6792
rect 22376 6749 22388 6783
rect 22388 6749 22422 6783
rect 22422 6749 22428 6783
rect 22652 6851 22704 6860
rect 22652 6817 22661 6851
rect 22661 6817 22695 6851
rect 22695 6817 22704 6851
rect 22652 6808 22704 6817
rect 23020 6808 23072 6860
rect 24032 6876 24084 6928
rect 26792 6944 26844 6996
rect 27988 6944 28040 6996
rect 27620 6876 27672 6928
rect 24492 6851 24544 6860
rect 24492 6817 24494 6851
rect 24494 6817 24544 6851
rect 24492 6808 24544 6817
rect 25596 6808 25648 6860
rect 25964 6808 26016 6860
rect 26516 6808 26568 6860
rect 22376 6740 22428 6749
rect 14556 6604 14608 6656
rect 15936 6647 15988 6656
rect 15936 6613 15945 6647
rect 15945 6613 15979 6647
rect 15979 6613 15988 6647
rect 15936 6604 15988 6613
rect 16120 6647 16172 6656
rect 16120 6613 16129 6647
rect 16129 6613 16163 6647
rect 16163 6613 16172 6647
rect 16120 6604 16172 6613
rect 21640 6672 21692 6724
rect 24676 6740 24728 6792
rect 26056 6740 26108 6792
rect 29644 6808 29696 6860
rect 30656 6808 30708 6860
rect 27528 6740 27580 6792
rect 27804 6740 27856 6792
rect 28080 6783 28132 6792
rect 28080 6749 28092 6783
rect 28092 6749 28126 6783
rect 28126 6749 28132 6783
rect 28080 6740 28132 6749
rect 29276 6740 29328 6792
rect 25872 6672 25924 6724
rect 21088 6604 21140 6656
rect 22192 6604 22244 6656
rect 22836 6604 22888 6656
rect 26240 6604 26292 6656
rect 26516 6604 26568 6656
rect 4193 6502 4245 6554
rect 4257 6502 4309 6554
rect 4321 6502 4373 6554
rect 4385 6502 4437 6554
rect 4449 6502 4501 6554
rect 11783 6502 11835 6554
rect 11847 6502 11899 6554
rect 11911 6502 11963 6554
rect 11975 6502 12027 6554
rect 12039 6502 12091 6554
rect 19373 6502 19425 6554
rect 19437 6502 19489 6554
rect 19501 6502 19553 6554
rect 19565 6502 19617 6554
rect 19629 6502 19681 6554
rect 26963 6502 27015 6554
rect 27027 6502 27079 6554
rect 27091 6502 27143 6554
rect 27155 6502 27207 6554
rect 27219 6502 27271 6554
rect 5448 6400 5500 6452
rect 940 6239 992 6248
rect 940 6205 949 6239
rect 949 6205 983 6239
rect 983 6205 992 6239
rect 940 6196 992 6205
rect 1676 6239 1728 6248
rect 1676 6205 1685 6239
rect 1685 6205 1719 6239
rect 1719 6205 1728 6239
rect 1676 6196 1728 6205
rect 3424 6196 3476 6248
rect 3976 6264 4028 6316
rect 6368 6400 6420 6452
rect 6644 6400 6696 6452
rect 7932 6443 7984 6452
rect 7932 6409 7941 6443
rect 7941 6409 7975 6443
rect 7975 6409 7984 6443
rect 7932 6400 7984 6409
rect 8300 6400 8352 6452
rect 9680 6400 9732 6452
rect 9864 6400 9916 6452
rect 11244 6400 11296 6452
rect 12072 6400 12124 6452
rect 12716 6400 12768 6452
rect 12992 6400 13044 6452
rect 13636 6400 13688 6452
rect 13728 6443 13780 6452
rect 13728 6409 13737 6443
rect 13737 6409 13771 6443
rect 13771 6409 13780 6443
rect 13728 6400 13780 6409
rect 14464 6400 14516 6452
rect 19064 6400 19116 6452
rect 10784 6332 10836 6384
rect 14372 6332 14424 6384
rect 6460 6307 6512 6316
rect 6460 6273 6462 6307
rect 6462 6273 6512 6307
rect 6460 6264 6512 6273
rect 6644 6264 6696 6316
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 7472 6264 7524 6316
rect 8760 6264 8812 6316
rect 9404 6264 9456 6316
rect 4804 6196 4856 6248
rect 5540 6196 5592 6248
rect 7104 6196 7156 6248
rect 8392 6239 8444 6248
rect 8392 6205 8401 6239
rect 8401 6205 8435 6239
rect 8435 6205 8444 6239
rect 8392 6196 8444 6205
rect 8852 6239 8904 6248
rect 8852 6205 8861 6239
rect 8861 6205 8895 6239
rect 8895 6205 8904 6239
rect 8852 6196 8904 6205
rect 9128 6239 9180 6248
rect 9128 6205 9137 6239
rect 9137 6205 9171 6239
rect 9171 6205 9180 6239
rect 9128 6196 9180 6205
rect 10232 6196 10284 6248
rect 11428 6196 11480 6248
rect 12072 6196 12124 6248
rect 12164 6196 12216 6248
rect 13452 6264 13504 6316
rect 14280 6264 14332 6316
rect 12808 6239 12860 6248
rect 1400 6103 1452 6112
rect 1400 6069 1415 6103
rect 1415 6069 1449 6103
rect 1449 6069 1452 6103
rect 1400 6060 1452 6069
rect 3240 6060 3292 6112
rect 3424 6060 3476 6112
rect 3700 6060 3752 6112
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 5632 6060 5684 6112
rect 5816 6060 5868 6112
rect 6368 6060 6420 6112
rect 6736 6060 6788 6112
rect 8576 6103 8628 6112
rect 8576 6069 8585 6103
rect 8585 6069 8619 6103
rect 8619 6069 8628 6103
rect 8576 6060 8628 6069
rect 9220 6060 9272 6112
rect 11060 6128 11112 6180
rect 12808 6205 12809 6239
rect 12809 6205 12843 6239
rect 12843 6205 12860 6239
rect 12808 6196 12860 6205
rect 12900 6239 12952 6248
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 13360 6239 13412 6248
rect 13360 6205 13369 6239
rect 13369 6205 13403 6239
rect 13403 6205 13412 6239
rect 13360 6196 13412 6205
rect 13636 6128 13688 6180
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 14740 6264 14792 6316
rect 14924 6307 14976 6316
rect 14924 6273 14926 6307
rect 14926 6273 14976 6307
rect 14924 6264 14976 6273
rect 15384 6264 15436 6316
rect 16856 6196 16908 6248
rect 9496 6060 9548 6112
rect 11520 6103 11572 6112
rect 11520 6069 11529 6103
rect 11529 6069 11563 6103
rect 11563 6069 11572 6103
rect 11520 6060 11572 6069
rect 11796 6060 11848 6112
rect 11980 6060 12032 6112
rect 12256 6060 12308 6112
rect 13360 6060 13412 6112
rect 16672 6128 16724 6180
rect 18788 6264 18840 6316
rect 20812 6400 20864 6452
rect 21088 6400 21140 6452
rect 21640 6400 21692 6452
rect 18512 6239 18564 6248
rect 18512 6205 18521 6239
rect 18521 6205 18555 6239
rect 18555 6205 18564 6239
rect 18512 6196 18564 6205
rect 21916 6264 21968 6316
rect 23020 6307 23072 6316
rect 23020 6273 23029 6307
rect 23029 6273 23063 6307
rect 23063 6273 23072 6307
rect 23020 6264 23072 6273
rect 23388 6307 23440 6316
rect 23388 6273 23397 6307
rect 23397 6273 23431 6307
rect 23431 6273 23440 6307
rect 23388 6264 23440 6273
rect 24216 6264 24268 6316
rect 27620 6400 27672 6452
rect 28172 6332 28224 6384
rect 20260 6239 20312 6248
rect 17868 6128 17920 6180
rect 18144 6128 18196 6180
rect 20260 6205 20262 6239
rect 20262 6205 20312 6239
rect 20260 6196 20312 6205
rect 20628 6239 20680 6248
rect 20628 6205 20637 6239
rect 20637 6205 20671 6239
rect 20671 6205 20680 6239
rect 20628 6196 20680 6205
rect 20720 6196 20772 6248
rect 15384 6060 15436 6112
rect 17316 6103 17368 6112
rect 17316 6069 17325 6103
rect 17325 6069 17359 6103
rect 17359 6069 17368 6103
rect 17316 6060 17368 6069
rect 18420 6060 18472 6112
rect 18972 6103 19024 6112
rect 18972 6069 18981 6103
rect 18981 6069 19015 6103
rect 19015 6069 19024 6103
rect 18972 6060 19024 6069
rect 19064 6060 19116 6112
rect 19524 6103 19576 6112
rect 19524 6069 19533 6103
rect 19533 6069 19567 6103
rect 19567 6069 19576 6103
rect 19524 6060 19576 6069
rect 19984 6128 20036 6180
rect 21640 6128 21692 6180
rect 21824 6128 21876 6180
rect 22560 6239 22612 6248
rect 22560 6205 22569 6239
rect 22569 6205 22603 6239
rect 22603 6205 22612 6239
rect 22560 6196 22612 6205
rect 22744 6239 22796 6248
rect 22744 6205 22753 6239
rect 22753 6205 22787 6239
rect 22787 6205 22796 6239
rect 22744 6196 22796 6205
rect 23572 6196 23624 6248
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 28540 6264 28592 6316
rect 26056 6196 26108 6248
rect 26608 6196 26660 6248
rect 25596 6128 25648 6180
rect 26424 6128 26476 6180
rect 21916 6103 21968 6112
rect 21916 6069 21925 6103
rect 21925 6069 21959 6103
rect 21959 6069 21968 6103
rect 21916 6060 21968 6069
rect 22100 6103 22152 6112
rect 22100 6069 22109 6103
rect 22109 6069 22143 6103
rect 22143 6069 22152 6103
rect 22100 6060 22152 6069
rect 22560 6060 22612 6112
rect 23848 6060 23900 6112
rect 24492 6103 24544 6112
rect 24492 6069 24507 6103
rect 24507 6069 24541 6103
rect 24541 6069 24544 6103
rect 24492 6060 24544 6069
rect 24676 6060 24728 6112
rect 28632 6196 28684 6248
rect 26976 6060 27028 6112
rect 27160 6103 27212 6112
rect 27160 6069 27175 6103
rect 27175 6069 27209 6103
rect 27209 6069 27212 6103
rect 27160 6060 27212 6069
rect 27344 6060 27396 6112
rect 27804 6060 27856 6112
rect 29276 6060 29328 6112
rect 7988 5958 8040 6010
rect 8052 5958 8104 6010
rect 8116 5958 8168 6010
rect 8180 5958 8232 6010
rect 8244 5958 8296 6010
rect 15578 5958 15630 6010
rect 15642 5958 15694 6010
rect 15706 5958 15758 6010
rect 15770 5958 15822 6010
rect 15834 5958 15886 6010
rect 23168 5958 23220 6010
rect 23232 5958 23284 6010
rect 23296 5958 23348 6010
rect 23360 5958 23412 6010
rect 23424 5958 23476 6010
rect 30758 5958 30810 6010
rect 30822 5958 30874 6010
rect 30886 5958 30938 6010
rect 30950 5958 31002 6010
rect 31014 5958 31066 6010
rect 1952 5856 2004 5908
rect 1032 5763 1084 5772
rect 1032 5729 1041 5763
rect 1041 5729 1075 5763
rect 1075 5729 1084 5763
rect 1032 5720 1084 5729
rect 1400 5720 1452 5772
rect 5172 5856 5224 5908
rect 5356 5856 5408 5908
rect 8484 5856 8536 5908
rect 8668 5856 8720 5908
rect 10784 5899 10836 5908
rect 10784 5865 10793 5899
rect 10793 5865 10827 5899
rect 10827 5865 10836 5899
rect 10784 5856 10836 5865
rect 6092 5831 6144 5840
rect 6092 5797 6101 5831
rect 6101 5797 6135 5831
rect 6135 5797 6144 5831
rect 6092 5788 6144 5797
rect 9772 5788 9824 5840
rect 940 5652 992 5704
rect 3608 5720 3660 5772
rect 4528 5720 4580 5772
rect 5540 5720 5592 5772
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 6184 5720 6236 5772
rect 6644 5720 6696 5772
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 2872 5652 2924 5704
rect 3700 5652 3752 5704
rect 4068 5652 4120 5704
rect 4712 5652 4764 5704
rect 7104 5763 7156 5772
rect 7104 5729 7113 5763
rect 7113 5729 7147 5763
rect 7147 5729 7156 5763
rect 7104 5720 7156 5729
rect 7656 5763 7708 5772
rect 7656 5729 7665 5763
rect 7665 5729 7699 5763
rect 7699 5729 7708 5763
rect 7656 5720 7708 5729
rect 7748 5720 7800 5772
rect 5448 5584 5500 5636
rect 7196 5652 7248 5704
rect 7840 5695 7892 5704
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 8392 5652 8444 5704
rect 10140 5652 10192 5704
rect 10508 5763 10560 5772
rect 10508 5729 10517 5763
rect 10517 5729 10551 5763
rect 10551 5729 10560 5763
rect 10508 5720 10560 5729
rect 10692 5788 10744 5840
rect 10784 5720 10836 5772
rect 11060 5720 11112 5772
rect 11244 5763 11296 5772
rect 11244 5729 11253 5763
rect 11253 5729 11287 5763
rect 11287 5729 11296 5763
rect 11244 5720 11296 5729
rect 11612 5763 11664 5772
rect 11612 5729 11621 5763
rect 11621 5729 11655 5763
rect 11655 5729 11664 5763
rect 11612 5720 11664 5729
rect 11980 5856 12032 5908
rect 12256 5856 12308 5908
rect 13912 5856 13964 5908
rect 20536 5899 20588 5908
rect 20536 5865 20545 5899
rect 20545 5865 20579 5899
rect 20579 5865 20588 5899
rect 20536 5856 20588 5865
rect 20628 5856 20680 5908
rect 21916 5856 21968 5908
rect 24492 5856 24544 5908
rect 26700 5856 26752 5908
rect 19984 5788 20036 5840
rect 1492 5516 1544 5568
rect 2044 5516 2096 5568
rect 3976 5516 4028 5568
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 6552 5516 6604 5568
rect 6736 5516 6788 5568
rect 7472 5559 7524 5568
rect 7472 5525 7481 5559
rect 7481 5525 7515 5559
rect 7515 5525 7524 5559
rect 7472 5516 7524 5525
rect 9496 5584 9548 5636
rect 10508 5584 10560 5636
rect 11244 5584 11296 5636
rect 13820 5695 13872 5704
rect 13820 5661 13829 5695
rect 13829 5661 13863 5695
rect 13863 5661 13872 5695
rect 13820 5652 13872 5661
rect 14188 5695 14240 5704
rect 14188 5661 14190 5695
rect 14190 5661 14240 5695
rect 14188 5652 14240 5661
rect 14372 5720 14424 5772
rect 16672 5720 16724 5772
rect 17316 5720 17368 5772
rect 18144 5720 18196 5772
rect 15936 5652 15988 5704
rect 16580 5695 16632 5704
rect 16580 5661 16592 5695
rect 16592 5661 16626 5695
rect 16626 5661 16632 5695
rect 16580 5652 16632 5661
rect 8668 5516 8720 5568
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 10968 5516 11020 5568
rect 12256 5516 12308 5568
rect 16764 5516 16816 5568
rect 18144 5559 18196 5568
rect 18144 5525 18153 5559
rect 18153 5525 18187 5559
rect 18187 5525 18196 5559
rect 18144 5516 18196 5525
rect 18512 5652 18564 5704
rect 18696 5695 18748 5704
rect 18696 5661 18698 5695
rect 18698 5661 18748 5695
rect 18696 5652 18748 5661
rect 18788 5695 18840 5704
rect 18788 5661 18800 5695
rect 18800 5661 18834 5695
rect 18834 5661 18840 5695
rect 18788 5652 18840 5661
rect 19524 5720 19576 5772
rect 21640 5720 21692 5772
rect 21824 5720 21876 5772
rect 26056 5788 26108 5840
rect 26332 5788 26384 5840
rect 21640 5584 21692 5636
rect 18604 5516 18656 5568
rect 20352 5559 20404 5568
rect 20352 5525 20361 5559
rect 20361 5525 20395 5559
rect 20395 5525 20404 5559
rect 20352 5516 20404 5525
rect 21088 5516 21140 5568
rect 21916 5695 21968 5704
rect 21916 5661 21925 5695
rect 21925 5661 21959 5695
rect 21959 5661 21968 5695
rect 21916 5652 21968 5661
rect 22284 5695 22336 5704
rect 22284 5661 22286 5695
rect 22286 5661 22336 5695
rect 22284 5652 22336 5661
rect 22560 5720 22612 5772
rect 27068 5788 27120 5840
rect 23848 5652 23900 5704
rect 24860 5695 24912 5704
rect 24860 5661 24869 5695
rect 24869 5661 24903 5695
rect 24903 5661 24912 5695
rect 24860 5652 24912 5661
rect 25872 5652 25924 5704
rect 26148 5652 26200 5704
rect 26976 5720 27028 5772
rect 27528 5856 27580 5908
rect 27344 5652 27396 5704
rect 29368 5899 29420 5908
rect 29368 5865 29377 5899
rect 29377 5865 29411 5899
rect 29411 5865 29420 5899
rect 29368 5856 29420 5865
rect 27804 5720 27856 5772
rect 28172 5652 28224 5704
rect 26792 5584 26844 5636
rect 22468 5516 22520 5568
rect 26148 5559 26200 5568
rect 26148 5525 26157 5559
rect 26157 5525 26191 5559
rect 26191 5525 26200 5559
rect 26148 5516 26200 5525
rect 26700 5559 26752 5568
rect 26700 5525 26709 5559
rect 26709 5525 26743 5559
rect 26743 5525 26752 5559
rect 26700 5516 26752 5525
rect 26884 5516 26936 5568
rect 28172 5516 28224 5568
rect 4193 5414 4245 5466
rect 4257 5414 4309 5466
rect 4321 5414 4373 5466
rect 4385 5414 4437 5466
rect 4449 5414 4501 5466
rect 11783 5414 11835 5466
rect 11847 5414 11899 5466
rect 11911 5414 11963 5466
rect 11975 5414 12027 5466
rect 12039 5414 12091 5466
rect 19373 5414 19425 5466
rect 19437 5414 19489 5466
rect 19501 5414 19553 5466
rect 19565 5414 19617 5466
rect 19629 5414 19681 5466
rect 26963 5414 27015 5466
rect 27027 5414 27079 5466
rect 27091 5414 27143 5466
rect 27155 5414 27207 5466
rect 27219 5414 27271 5466
rect 4068 5312 4120 5364
rect 4160 5312 4212 5364
rect 7472 5312 7524 5364
rect 3516 5287 3568 5296
rect 3516 5253 3525 5287
rect 3525 5253 3559 5287
rect 3559 5253 3568 5287
rect 3516 5244 3568 5253
rect 940 5151 992 5160
rect 940 5117 949 5151
rect 949 5117 983 5151
rect 983 5117 992 5151
rect 940 5108 992 5117
rect 4068 5176 4120 5228
rect 5724 5176 5776 5228
rect 9496 5312 9548 5364
rect 10692 5312 10744 5364
rect 13912 5312 13964 5364
rect 16580 5312 16632 5364
rect 17132 5312 17184 5364
rect 13636 5244 13688 5296
rect 20720 5355 20772 5364
rect 20720 5321 20729 5355
rect 20729 5321 20763 5355
rect 20763 5321 20772 5355
rect 20720 5312 20772 5321
rect 23480 5244 23532 5296
rect 25596 5312 25648 5364
rect 25964 5244 26016 5296
rect 26608 5244 26660 5296
rect 2964 5040 3016 5092
rect 3240 5040 3292 5092
rect 1400 5015 1452 5024
rect 1400 4981 1415 5015
rect 1415 4981 1449 5015
rect 1449 4981 1452 5015
rect 1400 4972 1452 4981
rect 2044 4972 2096 5024
rect 2320 4972 2372 5024
rect 3884 5151 3936 5160
rect 3884 5117 3893 5151
rect 3893 5117 3927 5151
rect 3927 5117 3936 5151
rect 3884 5108 3936 5117
rect 4160 5108 4212 5160
rect 5448 5108 5500 5160
rect 5908 5108 5960 5160
rect 8484 5108 8536 5160
rect 8668 5108 8720 5160
rect 8944 5108 8996 5160
rect 9680 5176 9732 5228
rect 13360 5176 13412 5228
rect 9588 5108 9640 5160
rect 11336 5108 11388 5160
rect 11520 5108 11572 5160
rect 13912 5176 13964 5228
rect 16120 5176 16172 5228
rect 18144 5176 18196 5228
rect 20260 5176 20312 5228
rect 21640 5219 21692 5228
rect 21640 5185 21649 5219
rect 21649 5185 21683 5219
rect 21683 5185 21692 5219
rect 21640 5176 21692 5185
rect 15936 5151 15988 5160
rect 15936 5117 15945 5151
rect 15945 5117 15979 5151
rect 15979 5117 15988 5151
rect 15936 5108 15988 5117
rect 18420 5108 18472 5160
rect 18512 5151 18564 5160
rect 18512 5117 18521 5151
rect 18521 5117 18555 5151
rect 18555 5117 18564 5151
rect 18512 5108 18564 5117
rect 18604 5108 18656 5160
rect 13820 5040 13872 5092
rect 18052 5083 18104 5092
rect 18052 5049 18061 5083
rect 18061 5049 18095 5083
rect 18095 5049 18104 5083
rect 18052 5040 18104 5049
rect 20812 5108 20864 5160
rect 21916 5108 21968 5160
rect 22008 5108 22060 5160
rect 23296 5151 23348 5160
rect 23296 5117 23305 5151
rect 23305 5117 23339 5151
rect 23339 5117 23348 5151
rect 23296 5108 23348 5117
rect 23572 5176 23624 5228
rect 25044 5176 25096 5228
rect 29000 5244 29052 5296
rect 27896 5176 27948 5228
rect 23664 5108 23716 5160
rect 6368 4972 6420 5024
rect 6828 4972 6880 5024
rect 9036 4972 9088 5024
rect 11520 4972 11572 5024
rect 11704 5015 11756 5024
rect 11704 4981 11719 5015
rect 11719 4981 11753 5015
rect 11753 4981 11756 5015
rect 11704 4972 11756 4981
rect 14188 5015 14240 5024
rect 14188 4981 14203 5015
rect 14203 4981 14237 5015
rect 14237 4981 14240 5015
rect 14188 4972 14240 4981
rect 16672 4972 16724 5024
rect 18696 4972 18748 5024
rect 20812 4972 20864 5024
rect 20904 4972 20956 5024
rect 21640 4972 21692 5024
rect 22284 4972 22336 5024
rect 22652 4972 22704 5024
rect 23112 5040 23164 5092
rect 23480 5040 23532 5092
rect 25320 5108 25372 5160
rect 25872 5108 25924 5160
rect 27436 5151 27488 5160
rect 27436 5117 27445 5151
rect 27445 5117 27479 5151
rect 27479 5117 27488 5151
rect 27436 5108 27488 5117
rect 31208 5244 31260 5296
rect 29092 5040 29144 5092
rect 29920 5108 29972 5160
rect 27344 4972 27396 5024
rect 27436 4972 27488 5024
rect 29000 5015 29052 5024
rect 29000 4981 29009 5015
rect 29009 4981 29043 5015
rect 29043 4981 29052 5015
rect 29000 4972 29052 4981
rect 7988 4870 8040 4922
rect 8052 4870 8104 4922
rect 8116 4870 8168 4922
rect 8180 4870 8232 4922
rect 8244 4870 8296 4922
rect 15578 4870 15630 4922
rect 15642 4870 15694 4922
rect 15706 4870 15758 4922
rect 15770 4870 15822 4922
rect 15834 4870 15886 4922
rect 23168 4870 23220 4922
rect 23232 4870 23284 4922
rect 23296 4870 23348 4922
rect 23360 4870 23412 4922
rect 23424 4870 23476 4922
rect 30758 4870 30810 4922
rect 30822 4870 30874 4922
rect 30886 4870 30938 4922
rect 30950 4870 31002 4922
rect 31014 4870 31066 4922
rect 1860 4768 1912 4820
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 4528 4768 4580 4820
rect 7656 4768 7708 4820
rect 8392 4768 8444 4820
rect 9496 4768 9548 4820
rect 11244 4768 11296 4820
rect 11428 4768 11480 4820
rect 11704 4768 11756 4820
rect 14188 4768 14240 4820
rect 18052 4768 18104 4820
rect 18788 4768 18840 4820
rect 20812 4768 20864 4820
rect 20904 4768 20956 4820
rect 21732 4768 21784 4820
rect 22100 4768 22152 4820
rect 22284 4768 22336 4820
rect 24676 4768 24728 4820
rect 24768 4811 24820 4820
rect 24768 4777 24777 4811
rect 24777 4777 24811 4811
rect 24811 4777 24820 4811
rect 24768 4768 24820 4777
rect 1400 4632 1452 4684
rect 940 4564 992 4616
rect 2780 4564 2832 4616
rect 3240 4428 3292 4480
rect 4160 4632 4212 4684
rect 6000 4632 6052 4684
rect 6184 4632 6236 4684
rect 6552 4632 6604 4684
rect 6920 4632 6972 4684
rect 3792 4564 3844 4616
rect 3976 4607 4028 4616
rect 3976 4573 3988 4607
rect 3988 4573 4022 4607
rect 4022 4573 4028 4607
rect 3976 4564 4028 4573
rect 5816 4564 5868 4616
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 7748 4564 7800 4616
rect 8208 4564 8260 4616
rect 9036 4632 9088 4684
rect 8944 4564 8996 4616
rect 9680 4632 9732 4684
rect 16120 4700 16172 4752
rect 5540 4471 5592 4480
rect 5540 4437 5549 4471
rect 5549 4437 5583 4471
rect 5583 4437 5592 4471
rect 5540 4428 5592 4437
rect 6828 4428 6880 4480
rect 7104 4428 7156 4480
rect 8392 4471 8444 4480
rect 8392 4437 8401 4471
rect 8401 4437 8435 4471
rect 8435 4437 8444 4471
rect 8392 4428 8444 4437
rect 11520 4675 11572 4684
rect 11520 4641 11529 4675
rect 11529 4641 11563 4675
rect 11563 4641 11572 4675
rect 11520 4632 11572 4641
rect 12256 4632 12308 4684
rect 12440 4632 12492 4684
rect 11336 4564 11388 4616
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 12164 4564 12216 4616
rect 11520 4496 11572 4548
rect 11336 4471 11388 4480
rect 11336 4437 11345 4471
rect 11345 4437 11379 4471
rect 11379 4437 11388 4471
rect 11336 4428 11388 4437
rect 12808 4428 12860 4480
rect 13820 4607 13872 4616
rect 13820 4573 13829 4607
rect 13829 4573 13863 4607
rect 13863 4573 13872 4607
rect 13820 4564 13872 4573
rect 16764 4632 16816 4684
rect 14372 4564 14424 4616
rect 16120 4607 16172 4616
rect 16120 4573 16129 4607
rect 16129 4573 16163 4607
rect 16163 4573 16172 4607
rect 16120 4564 16172 4573
rect 16488 4607 16540 4616
rect 16488 4573 16490 4607
rect 16490 4573 16540 4607
rect 16488 4564 16540 4573
rect 19064 4675 19116 4684
rect 19064 4641 19073 4675
rect 19073 4641 19107 4675
rect 19107 4641 19116 4675
rect 19064 4632 19116 4641
rect 20444 4632 20496 4684
rect 20996 4675 21048 4684
rect 20996 4641 21005 4675
rect 21005 4641 21039 4675
rect 21039 4641 21048 4675
rect 20996 4632 21048 4641
rect 21640 4632 21692 4684
rect 21916 4632 21968 4684
rect 26056 4768 26108 4820
rect 25044 4700 25096 4752
rect 25596 4700 25648 4752
rect 27252 4811 27304 4820
rect 27252 4777 27261 4811
rect 27261 4777 27295 4811
rect 27295 4777 27304 4811
rect 27252 4768 27304 4777
rect 27344 4768 27396 4820
rect 28264 4811 28316 4820
rect 28264 4777 28279 4811
rect 28279 4777 28313 4811
rect 28313 4777 28316 4811
rect 28264 4768 28316 4777
rect 14372 4428 14424 4480
rect 18512 4564 18564 4616
rect 18696 4607 18748 4616
rect 18696 4573 18698 4607
rect 18698 4573 18748 4607
rect 18696 4564 18748 4573
rect 19156 4564 19208 4616
rect 22376 4564 22428 4616
rect 22652 4564 22704 4616
rect 25136 4632 25188 4684
rect 26608 4632 26660 4684
rect 27436 4700 27488 4752
rect 27712 4700 27764 4752
rect 27344 4632 27396 4684
rect 25320 4564 25372 4616
rect 25412 4564 25464 4616
rect 27528 4632 27580 4684
rect 28908 4632 28960 4684
rect 18972 4428 19024 4480
rect 19064 4428 19116 4480
rect 21824 4496 21876 4548
rect 20076 4428 20128 4480
rect 21548 4471 21600 4480
rect 21548 4437 21557 4471
rect 21557 4437 21591 4471
rect 21591 4437 21600 4471
rect 21548 4428 21600 4437
rect 21640 4428 21692 4480
rect 27252 4496 27304 4548
rect 24308 4428 24360 4480
rect 24676 4428 24728 4480
rect 25044 4471 25096 4480
rect 25044 4437 25053 4471
rect 25053 4437 25087 4471
rect 25087 4437 25096 4471
rect 25044 4428 25096 4437
rect 25320 4471 25372 4480
rect 25320 4437 25329 4471
rect 25329 4437 25363 4471
rect 25363 4437 25372 4471
rect 25320 4428 25372 4437
rect 25504 4428 25556 4480
rect 4193 4326 4245 4378
rect 4257 4326 4309 4378
rect 4321 4326 4373 4378
rect 4385 4326 4437 4378
rect 4449 4326 4501 4378
rect 11783 4326 11835 4378
rect 11847 4326 11899 4378
rect 11911 4326 11963 4378
rect 11975 4326 12027 4378
rect 12039 4326 12091 4378
rect 19373 4326 19425 4378
rect 19437 4326 19489 4378
rect 19501 4326 19553 4378
rect 19565 4326 19617 4378
rect 19629 4326 19681 4378
rect 26963 4326 27015 4378
rect 27027 4326 27079 4378
rect 27091 4326 27143 4378
rect 27155 4326 27207 4378
rect 27219 4326 27271 4378
rect 2412 4156 2464 4208
rect 5724 4267 5776 4276
rect 5724 4233 5733 4267
rect 5733 4233 5767 4267
rect 5767 4233 5776 4267
rect 5724 4224 5776 4233
rect 8392 4224 8444 4276
rect 7656 4156 7708 4208
rect 8576 4156 8628 4208
rect 3056 4088 3108 4140
rect 940 4063 992 4072
rect 940 4029 949 4063
rect 949 4029 983 4063
rect 983 4029 992 4063
rect 940 4020 992 4029
rect 1952 4020 2004 4072
rect 2504 4020 2556 4072
rect 3332 4020 3384 4072
rect 3608 4063 3660 4072
rect 3608 4029 3617 4063
rect 3617 4029 3651 4063
rect 3651 4029 3660 4063
rect 3608 4020 3660 4029
rect 3792 4020 3844 4072
rect 4804 4088 4856 4140
rect 5540 4088 5592 4140
rect 6736 4088 6788 4140
rect 4344 4020 4396 4072
rect 5632 4020 5684 4072
rect 5908 4063 5960 4072
rect 5908 4029 5917 4063
rect 5917 4029 5951 4063
rect 5951 4029 5960 4063
rect 5908 4020 5960 4029
rect 6000 4020 6052 4072
rect 9036 4088 9088 4140
rect 9864 4156 9916 4208
rect 12164 4224 12216 4276
rect 13820 4224 13872 4276
rect 15108 4224 15160 4276
rect 16304 4224 16356 4276
rect 18144 4224 18196 4276
rect 21640 4224 21692 4276
rect 21732 4224 21784 4276
rect 23112 4224 23164 4276
rect 25136 4224 25188 4276
rect 27344 4224 27396 4276
rect 29092 4224 29144 4276
rect 14188 4156 14240 4208
rect 18236 4199 18288 4208
rect 18236 4165 18245 4199
rect 18245 4165 18279 4199
rect 18279 4165 18288 4199
rect 18236 4156 18288 4165
rect 6920 4020 6972 4072
rect 8668 4020 8720 4072
rect 10048 4088 10100 4140
rect 10140 4088 10192 4140
rect 10508 4088 10560 4140
rect 11520 4088 11572 4140
rect 11704 4088 11756 4140
rect 5264 3952 5316 4004
rect 5448 3952 5500 4004
rect 1400 3927 1452 3936
rect 1400 3893 1415 3927
rect 1415 3893 1449 3927
rect 1449 3893 1452 3927
rect 1400 3884 1452 3893
rect 1584 3884 1636 3936
rect 2688 3884 2740 3936
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 2780 3884 2832 3893
rect 6184 3884 6236 3936
rect 7748 3927 7800 3936
rect 7748 3893 7757 3927
rect 7757 3893 7791 3927
rect 7791 3893 7800 3927
rect 7748 3884 7800 3893
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 8576 3884 8628 3893
rect 9036 3927 9088 3936
rect 9036 3893 9045 3927
rect 9045 3893 9079 3927
rect 9079 3893 9088 3927
rect 9036 3884 9088 3893
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 9496 3884 9548 3936
rect 9588 3927 9640 3936
rect 9588 3893 9597 3927
rect 9597 3893 9631 3927
rect 9631 3893 9640 3927
rect 9588 3884 9640 3893
rect 9956 3952 10008 4004
rect 10692 3884 10744 3936
rect 13268 4088 13320 4140
rect 16764 4088 16816 4140
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 13636 4063 13688 4072
rect 13636 4029 13645 4063
rect 13645 4029 13679 4063
rect 13679 4029 13688 4063
rect 13636 4020 13688 4029
rect 14004 4020 14056 4072
rect 14556 4020 14608 4072
rect 14924 4063 14976 4072
rect 14924 4029 14933 4063
rect 14933 4029 14967 4063
rect 14967 4029 14976 4063
rect 14924 4020 14976 4029
rect 16212 4020 16264 4072
rect 18052 4088 18104 4140
rect 18696 4088 18748 4140
rect 20352 4088 20404 4140
rect 20536 4088 20588 4140
rect 21088 4088 21140 4140
rect 14280 3952 14332 4004
rect 18512 3952 18564 4004
rect 18788 3995 18840 4004
rect 18788 3961 18797 3995
rect 18797 3961 18831 3995
rect 18831 3961 18840 3995
rect 18788 3952 18840 3961
rect 19248 4063 19300 4072
rect 19248 4029 19257 4063
rect 19257 4029 19291 4063
rect 19291 4029 19300 4063
rect 19248 4020 19300 4029
rect 22376 4063 22428 4072
rect 22376 4029 22385 4063
rect 22385 4029 22419 4063
rect 22419 4029 22428 4063
rect 22376 4020 22428 4029
rect 23112 4063 23164 4072
rect 23112 4029 23121 4063
rect 23121 4029 23155 4063
rect 23155 4029 23164 4063
rect 23112 4020 23164 4029
rect 23848 4088 23900 4140
rect 24308 4088 24360 4140
rect 24676 4088 24728 4140
rect 26148 4088 26200 4140
rect 26792 4088 26844 4140
rect 26240 4063 26292 4072
rect 26240 4029 26249 4063
rect 26249 4029 26283 4063
rect 26283 4029 26292 4063
rect 26240 4020 26292 4029
rect 27344 4020 27396 4072
rect 19708 3952 19760 4004
rect 22100 3995 22152 4004
rect 22100 3961 22109 3995
rect 22109 3961 22143 3995
rect 22143 3961 22152 3995
rect 22100 3952 22152 3961
rect 22284 3952 22336 4004
rect 22652 3995 22704 4004
rect 22652 3961 22661 3995
rect 22661 3961 22695 3995
rect 22695 3961 22704 3995
rect 22652 3952 22704 3961
rect 11428 3884 11480 3936
rect 12440 3884 12492 3936
rect 14464 3884 14516 3936
rect 14832 3884 14884 3936
rect 16672 3884 16724 3936
rect 17868 3884 17920 3936
rect 20260 3884 20312 3936
rect 24124 3952 24176 4004
rect 24400 3884 24452 3936
rect 24492 3927 24544 3936
rect 24492 3893 24507 3927
rect 24507 3893 24541 3927
rect 24541 3893 24544 3927
rect 24492 3884 24544 3893
rect 26056 3927 26108 3936
rect 26056 3893 26065 3927
rect 26065 3893 26099 3927
rect 26099 3893 26108 3927
rect 26056 3884 26108 3893
rect 26700 3927 26752 3936
rect 26700 3893 26715 3927
rect 26715 3893 26749 3927
rect 26749 3893 26752 3927
rect 26700 3884 26752 3893
rect 28080 3927 28132 3936
rect 28080 3893 28089 3927
rect 28089 3893 28123 3927
rect 28123 3893 28132 3927
rect 28080 3884 28132 3893
rect 7988 3782 8040 3834
rect 8052 3782 8104 3834
rect 8116 3782 8168 3834
rect 8180 3782 8232 3834
rect 8244 3782 8296 3834
rect 15578 3782 15630 3834
rect 15642 3782 15694 3834
rect 15706 3782 15758 3834
rect 15770 3782 15822 3834
rect 15834 3782 15886 3834
rect 23168 3782 23220 3834
rect 23232 3782 23284 3834
rect 23296 3782 23348 3834
rect 23360 3782 23412 3834
rect 23424 3782 23476 3834
rect 30758 3782 30810 3834
rect 30822 3782 30874 3834
rect 30886 3782 30938 3834
rect 30950 3782 31002 3834
rect 31014 3782 31066 3834
rect 1584 3680 1636 3732
rect 1768 3723 1820 3732
rect 1768 3689 1783 3723
rect 1783 3689 1817 3723
rect 1817 3689 1820 3723
rect 1768 3680 1820 3689
rect 2504 3680 2556 3732
rect 2780 3680 2832 3732
rect 3792 3680 3844 3732
rect 4344 3680 4396 3732
rect 5080 3680 5132 3732
rect 5816 3723 5868 3732
rect 5816 3689 5825 3723
rect 5825 3689 5859 3723
rect 5859 3689 5868 3723
rect 5816 3680 5868 3689
rect 5908 3680 5960 3732
rect 6276 3680 6328 3732
rect 6920 3680 6972 3732
rect 8484 3680 8536 3732
rect 9680 3723 9732 3732
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 9680 3680 9732 3689
rect 9864 3680 9916 3732
rect 9956 3680 10008 3732
rect 11704 3680 11756 3732
rect 12440 3680 12492 3732
rect 14096 3680 14148 3732
rect 14188 3680 14240 3732
rect 16580 3723 16632 3732
rect 16580 3689 16595 3723
rect 16595 3689 16629 3723
rect 16629 3689 16632 3723
rect 16580 3680 16632 3689
rect 16764 3680 16816 3732
rect 20168 3680 20220 3732
rect 20260 3680 20312 3732
rect 21272 3680 21324 3732
rect 22100 3680 22152 3732
rect 23572 3680 23624 3732
rect 23756 3680 23808 3732
rect 4988 3612 5040 3664
rect 1492 3476 1544 3528
rect 2872 3544 2924 3596
rect 3516 3587 3568 3596
rect 3516 3553 3525 3587
rect 3525 3553 3559 3587
rect 3559 3553 3568 3587
rect 3516 3544 3568 3553
rect 5356 3544 5408 3596
rect 6460 3612 6512 3664
rect 6368 3587 6420 3596
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 2412 3476 2464 3528
rect 6736 3476 6788 3528
rect 7104 3544 7156 3596
rect 7564 3655 7616 3664
rect 7564 3621 7573 3655
rect 7573 3621 7607 3655
rect 7607 3621 7616 3655
rect 7564 3612 7616 3621
rect 7748 3612 7800 3664
rect 7840 3519 7892 3528
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 9036 3544 9088 3596
rect 9956 3544 10008 3596
rect 10692 3544 10744 3596
rect 8392 3476 8444 3528
rect 9496 3476 9548 3528
rect 11428 3612 11480 3664
rect 11336 3544 11388 3596
rect 11612 3519 11664 3528
rect 3700 3340 3752 3392
rect 3792 3340 3844 3392
rect 7196 3408 7248 3460
rect 8392 3340 8444 3392
rect 8484 3340 8536 3392
rect 11612 3485 11621 3519
rect 11621 3485 11655 3519
rect 11655 3485 11664 3519
rect 11612 3476 11664 3485
rect 12164 3476 12216 3528
rect 13820 3519 13872 3528
rect 13820 3485 13829 3519
rect 13829 3485 13863 3519
rect 13863 3485 13872 3519
rect 13820 3476 13872 3485
rect 14464 3544 14516 3596
rect 14372 3476 14424 3528
rect 16120 3519 16172 3528
rect 16120 3485 16129 3519
rect 16129 3485 16163 3519
rect 16163 3485 16172 3519
rect 16120 3476 16172 3485
rect 16856 3519 16908 3528
rect 16856 3485 16865 3519
rect 16865 3485 16899 3519
rect 16899 3485 16908 3519
rect 16856 3476 16908 3485
rect 18696 3519 18748 3528
rect 18696 3485 18698 3519
rect 18698 3485 18748 3519
rect 14280 3340 14332 3392
rect 17868 3408 17920 3460
rect 18696 3476 18748 3485
rect 19064 3587 19116 3596
rect 19064 3553 19073 3587
rect 19073 3553 19107 3587
rect 19107 3553 19116 3587
rect 19064 3544 19116 3553
rect 20720 3544 20772 3596
rect 20904 3544 20956 3596
rect 21824 3544 21876 3596
rect 23664 3476 23716 3528
rect 23848 3519 23900 3528
rect 23848 3485 23850 3519
rect 23850 3485 23900 3519
rect 23848 3476 23900 3485
rect 24124 3544 24176 3596
rect 24492 3544 24544 3596
rect 25412 3544 25464 3596
rect 25780 3544 25832 3596
rect 18604 3340 18656 3392
rect 18788 3340 18840 3392
rect 24676 3340 24728 3392
rect 26516 3612 26568 3664
rect 26700 3612 26752 3664
rect 27344 3723 27396 3732
rect 27344 3689 27353 3723
rect 27353 3689 27387 3723
rect 27387 3689 27396 3723
rect 27344 3680 27396 3689
rect 27528 3680 27580 3732
rect 28264 3680 28316 3732
rect 27436 3612 27488 3664
rect 26148 3544 26200 3596
rect 29828 3544 29880 3596
rect 28356 3519 28408 3528
rect 28356 3485 28368 3519
rect 28368 3485 28402 3519
rect 28402 3485 28408 3519
rect 28356 3476 28408 3485
rect 4193 3238 4245 3290
rect 4257 3238 4309 3290
rect 4321 3238 4373 3290
rect 4385 3238 4437 3290
rect 4449 3238 4501 3290
rect 11783 3238 11835 3290
rect 11847 3238 11899 3290
rect 11911 3238 11963 3290
rect 11975 3238 12027 3290
rect 12039 3238 12091 3290
rect 19373 3238 19425 3290
rect 19437 3238 19489 3290
rect 19501 3238 19553 3290
rect 19565 3238 19617 3290
rect 19629 3238 19681 3290
rect 26963 3238 27015 3290
rect 27027 3238 27079 3290
rect 27091 3238 27143 3290
rect 27155 3238 27207 3290
rect 27219 3238 27271 3290
rect 2688 3136 2740 3188
rect 3792 3136 3844 3188
rect 5632 3136 5684 3188
rect 8484 3136 8536 3188
rect 9588 3136 9640 3188
rect 11796 3136 11848 3188
rect 16856 3136 16908 3188
rect 3148 3000 3200 3052
rect 3240 3000 3292 3052
rect 1584 2932 1636 2984
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 4436 3000 4488 3052
rect 4528 3000 4580 3052
rect 3516 2864 3568 2916
rect 5264 2932 5316 2984
rect 1768 2796 1820 2848
rect 7840 3068 7892 3120
rect 17960 3068 18012 3120
rect 19248 3136 19300 3188
rect 20720 3136 20772 3188
rect 6092 3043 6144 3052
rect 6092 3009 6101 3043
rect 6101 3009 6135 3043
rect 6135 3009 6144 3043
rect 6092 3000 6144 3009
rect 6368 3000 6420 3052
rect 6644 3000 6696 3052
rect 11796 3000 11848 3052
rect 14280 3000 14332 3052
rect 20076 3000 20128 3052
rect 21548 3000 21600 3052
rect 5448 2932 5500 2984
rect 9036 2975 9088 2984
rect 9036 2941 9045 2975
rect 9045 2941 9079 2975
rect 9079 2941 9088 2975
rect 9036 2932 9088 2941
rect 9312 2932 9364 2984
rect 11244 2975 11296 2984
rect 11244 2941 11253 2975
rect 11253 2941 11287 2975
rect 11287 2941 11296 2975
rect 11244 2932 11296 2941
rect 11612 2932 11664 2984
rect 13820 2932 13872 2984
rect 16028 2932 16080 2984
rect 17960 2932 18012 2984
rect 6000 2907 6052 2916
rect 6000 2873 6009 2907
rect 6009 2873 6043 2907
rect 6043 2873 6052 2907
rect 6000 2864 6052 2873
rect 18604 2932 18656 2984
rect 20444 2932 20496 2984
rect 20904 2975 20956 2984
rect 20904 2941 20913 2975
rect 20913 2941 20947 2975
rect 20947 2941 20956 2975
rect 20904 2932 20956 2941
rect 21732 2932 21784 2984
rect 22376 3136 22428 3188
rect 25412 3136 25464 3188
rect 26056 3136 26108 3188
rect 22652 3068 22704 3120
rect 23848 3068 23900 3120
rect 24400 3000 24452 3052
rect 24768 3000 24820 3052
rect 26148 3068 26200 3120
rect 28632 3179 28684 3188
rect 28632 3145 28641 3179
rect 28641 3145 28675 3179
rect 28675 3145 28684 3179
rect 28632 3136 28684 3145
rect 29460 3136 29512 3188
rect 29736 3136 29788 3188
rect 26792 3000 26844 3052
rect 27620 3000 27672 3052
rect 23664 2932 23716 2984
rect 25688 2932 25740 2984
rect 26148 2932 26200 2984
rect 26240 2975 26292 2984
rect 26240 2941 26249 2975
rect 26249 2941 26283 2975
rect 26283 2941 26292 2975
rect 26240 2932 26292 2941
rect 26608 2932 26660 2984
rect 28264 2932 28316 2984
rect 6828 2796 6880 2848
rect 7564 2796 7616 2848
rect 9128 2796 9180 2848
rect 9496 2839 9548 2848
rect 9496 2805 9511 2839
rect 9511 2805 9545 2839
rect 9545 2805 9548 2839
rect 9496 2796 9548 2805
rect 11704 2839 11756 2848
rect 11704 2805 11719 2839
rect 11719 2805 11753 2839
rect 11753 2805 11756 2839
rect 11704 2796 11756 2805
rect 14188 2839 14240 2848
rect 14188 2805 14203 2839
rect 14203 2805 14237 2839
rect 14237 2805 14240 2839
rect 14188 2796 14240 2805
rect 15384 2796 15436 2848
rect 16304 2796 16356 2848
rect 16580 2796 16632 2848
rect 18696 2796 18748 2848
rect 21272 2796 21324 2848
rect 21732 2796 21784 2848
rect 23848 2796 23900 2848
rect 24124 2796 24176 2848
rect 26700 2839 26752 2848
rect 26700 2805 26715 2839
rect 26715 2805 26749 2839
rect 26749 2805 26752 2839
rect 26700 2796 26752 2805
rect 27344 2796 27396 2848
rect 7988 2694 8040 2746
rect 8052 2694 8104 2746
rect 8116 2694 8168 2746
rect 8180 2694 8232 2746
rect 8244 2694 8296 2746
rect 15578 2694 15630 2746
rect 15642 2694 15694 2746
rect 15706 2694 15758 2746
rect 15770 2694 15822 2746
rect 15834 2694 15886 2746
rect 23168 2694 23220 2746
rect 23232 2694 23284 2746
rect 23296 2694 23348 2746
rect 23360 2694 23412 2746
rect 23424 2694 23476 2746
rect 30758 2694 30810 2746
rect 30822 2694 30874 2746
rect 30886 2694 30938 2746
rect 30950 2694 31002 2746
rect 31014 2694 31066 2746
rect 940 2524 992 2576
rect 1124 2456 1176 2508
rect 1768 2635 1820 2644
rect 1768 2601 1783 2635
rect 1783 2601 1817 2635
rect 1817 2601 1820 2635
rect 1768 2592 1820 2601
rect 3148 2635 3200 2644
rect 3148 2601 3157 2635
rect 3157 2601 3191 2635
rect 3191 2601 3200 2635
rect 3148 2592 3200 2601
rect 1676 2456 1728 2508
rect 2320 2456 2372 2508
rect 4712 2592 4764 2644
rect 6000 2592 6052 2644
rect 3332 2456 3384 2508
rect 4528 2456 4580 2508
rect 4712 2456 4764 2508
rect 5908 2524 5960 2576
rect 5816 2499 5868 2508
rect 5816 2465 5825 2499
rect 5825 2465 5859 2499
rect 5859 2465 5868 2499
rect 5816 2456 5868 2465
rect 6368 2456 6420 2508
rect 6460 2499 6512 2508
rect 6460 2465 6469 2499
rect 6469 2465 6503 2499
rect 6503 2465 6512 2499
rect 6460 2456 6512 2465
rect 3976 2431 4028 2440
rect 3976 2397 3988 2431
rect 3988 2397 4022 2431
rect 4022 2397 4028 2431
rect 3976 2388 4028 2397
rect 6828 2592 6880 2644
rect 9128 2635 9180 2644
rect 9128 2601 9143 2635
rect 9143 2601 9177 2635
rect 9177 2601 9180 2635
rect 9128 2592 9180 2601
rect 11244 2635 11296 2644
rect 11244 2601 11253 2635
rect 11253 2601 11287 2635
rect 11287 2601 11296 2635
rect 11244 2592 11296 2601
rect 11704 2592 11756 2644
rect 12440 2592 12492 2644
rect 13728 2592 13780 2644
rect 14188 2592 14240 2644
rect 16580 2635 16632 2644
rect 16580 2601 16595 2635
rect 16595 2601 16629 2635
rect 16629 2601 16632 2635
rect 16580 2592 16632 2601
rect 18236 2592 18288 2644
rect 20996 2592 21048 2644
rect 21272 2592 21324 2644
rect 6736 2456 6788 2508
rect 7196 2499 7248 2508
rect 7196 2465 7205 2499
rect 7205 2465 7239 2499
rect 7239 2465 7248 2499
rect 7196 2456 7248 2465
rect 9312 2456 9364 2508
rect 11888 2456 11940 2508
rect 5632 2320 5684 2372
rect 6368 2320 6420 2372
rect 7288 2252 7340 2304
rect 11244 2388 11296 2440
rect 11612 2431 11664 2440
rect 11612 2397 11621 2431
rect 11621 2397 11655 2431
rect 11655 2397 11664 2431
rect 11612 2388 11664 2397
rect 11796 2388 11848 2440
rect 12164 2388 12216 2440
rect 9036 2252 9088 2304
rect 11980 2252 12032 2304
rect 12348 2252 12400 2304
rect 13728 2388 13780 2440
rect 14096 2388 14148 2440
rect 16028 2388 16080 2440
rect 17776 2388 17828 2440
rect 18512 2388 18564 2440
rect 18696 2431 18748 2440
rect 18696 2397 18698 2431
rect 18698 2397 18748 2431
rect 18696 2388 18748 2397
rect 19156 2456 19208 2508
rect 20536 2499 20588 2508
rect 20536 2465 20545 2499
rect 20545 2465 20579 2499
rect 20579 2465 20588 2499
rect 20536 2456 20588 2465
rect 20812 2456 20864 2508
rect 26700 2592 26752 2644
rect 28816 2635 28868 2644
rect 28816 2601 28825 2635
rect 28825 2601 28859 2635
rect 28859 2601 28868 2635
rect 28816 2592 28868 2601
rect 29368 2635 29420 2644
rect 29368 2601 29377 2635
rect 29377 2601 29411 2635
rect 29411 2601 29420 2635
rect 29368 2592 29420 2601
rect 23664 2524 23716 2576
rect 26424 2524 26476 2576
rect 13176 2320 13228 2372
rect 21180 2388 21232 2440
rect 23756 2456 23808 2508
rect 24032 2456 24084 2508
rect 21916 2388 21968 2440
rect 22008 2431 22060 2440
rect 22008 2397 22017 2431
rect 22017 2397 22051 2431
rect 22051 2397 22060 2431
rect 22008 2388 22060 2397
rect 24860 2499 24912 2508
rect 24860 2465 24869 2499
rect 24869 2465 24903 2499
rect 24903 2465 24912 2499
rect 24860 2456 24912 2465
rect 24308 2388 24360 2440
rect 24492 2431 24544 2440
rect 24492 2397 24494 2431
rect 24494 2397 24544 2431
rect 24492 2388 24544 2397
rect 24676 2388 24728 2440
rect 25688 2388 25740 2440
rect 26240 2388 26292 2440
rect 27068 2456 27120 2508
rect 29092 2524 29144 2576
rect 29460 2524 29512 2576
rect 26976 2388 27028 2440
rect 28816 2456 28868 2508
rect 29736 2456 29788 2508
rect 13728 2252 13780 2304
rect 21272 2320 21324 2372
rect 16672 2252 16724 2304
rect 19248 2252 19300 2304
rect 20628 2252 20680 2304
rect 20996 2252 21048 2304
rect 23480 2320 23532 2372
rect 23020 2252 23072 2304
rect 24308 2252 24360 2304
rect 26608 2252 26660 2304
rect 29552 2388 29604 2440
rect 29092 2363 29144 2372
rect 29092 2329 29101 2363
rect 29101 2329 29135 2363
rect 29135 2329 29144 2363
rect 29092 2320 29144 2329
rect 28264 2295 28316 2304
rect 28264 2261 28273 2295
rect 28273 2261 28307 2295
rect 28307 2261 28316 2295
rect 28264 2252 28316 2261
rect 4193 2150 4245 2202
rect 4257 2150 4309 2202
rect 4321 2150 4373 2202
rect 4385 2150 4437 2202
rect 4449 2150 4501 2202
rect 11783 2150 11835 2202
rect 11847 2150 11899 2202
rect 11911 2150 11963 2202
rect 11975 2150 12027 2202
rect 12039 2150 12091 2202
rect 19373 2150 19425 2202
rect 19437 2150 19489 2202
rect 19501 2150 19553 2202
rect 19565 2150 19617 2202
rect 19629 2150 19681 2202
rect 26963 2150 27015 2202
rect 27027 2150 27079 2202
rect 27091 2150 27143 2202
rect 27155 2150 27207 2202
rect 27219 2150 27271 2202
rect 1308 2048 1360 2100
rect 2872 2048 2924 2100
rect 3976 2048 4028 2100
rect 4620 2048 4672 2100
rect 6644 2048 6696 2100
rect 8852 2048 8904 2100
rect 10968 2048 11020 2100
rect 11980 2048 12032 2100
rect 12072 2048 12124 2100
rect 13176 2048 13228 2100
rect 14096 2048 14148 2100
rect 14556 2048 14608 2100
rect 3424 1980 3476 2032
rect 17960 2048 18012 2100
rect 21456 2048 21508 2100
rect 22008 2048 22060 2100
rect 2596 1912 2648 1964
rect 2136 1844 2188 1896
rect 3332 1844 3384 1896
rect 3700 1912 3752 1964
rect 4068 1912 4120 1964
rect 4252 1955 4304 1964
rect 4252 1921 4261 1955
rect 4261 1921 4295 1955
rect 4295 1921 4304 1955
rect 4252 1912 4304 1921
rect 6276 1912 6328 1964
rect 6368 1955 6420 1964
rect 6368 1921 6380 1955
rect 6380 1921 6414 1955
rect 6414 1921 6420 1955
rect 6368 1912 6420 1921
rect 9036 1955 9088 1964
rect 9036 1921 9045 1955
rect 9045 1921 9079 1955
rect 9079 1921 9088 1955
rect 9036 1912 9088 1921
rect 9220 1912 9272 1964
rect 9496 1955 9548 1964
rect 9496 1921 9508 1955
rect 9508 1921 9542 1955
rect 9542 1921 9548 1955
rect 9496 1912 9548 1921
rect 11796 1912 11848 1964
rect 11980 1955 12032 1964
rect 11980 1921 11989 1955
rect 11989 1921 12023 1955
rect 12023 1921 12032 1955
rect 11980 1912 12032 1921
rect 13636 1955 13688 1964
rect 13636 1921 13645 1955
rect 13645 1921 13679 1955
rect 13679 1921 13688 1955
rect 13636 1912 13688 1921
rect 14004 1955 14056 1964
rect 14004 1921 14006 1955
rect 14006 1921 14056 1955
rect 14004 1912 14056 1921
rect 3792 1844 3844 1896
rect 6184 1844 6236 1896
rect 8484 1887 8536 1896
rect 8484 1853 8493 1887
rect 8493 1853 8527 1887
rect 8527 1853 8536 1887
rect 8484 1844 8536 1853
rect 9772 1887 9824 1896
rect 9772 1853 9781 1887
rect 9781 1853 9815 1887
rect 9815 1853 9824 1887
rect 9772 1844 9824 1853
rect 11244 1887 11296 1896
rect 11244 1853 11253 1887
rect 11253 1853 11287 1887
rect 11287 1853 11296 1887
rect 11244 1844 11296 1853
rect 18512 1980 18564 2032
rect 19156 1955 19208 1964
rect 19156 1921 19168 1955
rect 19168 1921 19202 1955
rect 19202 1921 19208 1955
rect 19156 1912 19208 1921
rect 21456 1912 21508 1964
rect 23480 1980 23532 2032
rect 14372 1887 14424 1896
rect 14372 1853 14381 1887
rect 14381 1853 14415 1887
rect 14415 1853 14424 1887
rect 14372 1844 14424 1853
rect 15936 1844 15988 1896
rect 18236 1887 18288 1896
rect 18236 1853 18245 1887
rect 18245 1853 18279 1887
rect 18279 1853 18288 1887
rect 18236 1844 18288 1853
rect 18328 1844 18380 1896
rect 17960 1819 18012 1828
rect 17960 1785 17969 1819
rect 17969 1785 18003 1819
rect 18003 1785 18012 1819
rect 17960 1776 18012 1785
rect 1768 1708 1820 1760
rect 4712 1708 4764 1760
rect 6552 1708 6604 1760
rect 12072 1708 12124 1760
rect 13636 1708 13688 1760
rect 16580 1708 16632 1760
rect 18972 1844 19024 1896
rect 19432 1887 19484 1896
rect 19432 1853 19441 1887
rect 19441 1853 19475 1887
rect 19475 1853 19484 1887
rect 19432 1844 19484 1853
rect 20720 1776 20772 1828
rect 20812 1776 20864 1828
rect 22744 1844 22796 1896
rect 22928 1844 22980 1896
rect 23296 1887 23348 1896
rect 23296 1853 23305 1887
rect 23305 1853 23339 1887
rect 23339 1853 23348 1887
rect 23296 1844 23348 1853
rect 23480 1844 23532 1896
rect 23940 1776 23992 1828
rect 19064 1708 19116 1760
rect 19248 1708 19300 1760
rect 21180 1708 21232 1760
rect 22836 1708 22888 1760
rect 23664 1708 23716 1760
rect 24400 1844 24452 1896
rect 24768 1955 24820 1964
rect 24768 1921 24780 1955
rect 24780 1921 24814 1955
rect 24814 1921 24820 1955
rect 24768 1912 24820 1921
rect 25044 1955 25096 1964
rect 25044 1921 25053 1955
rect 25053 1921 25087 1955
rect 25087 1921 25096 1955
rect 25044 1912 25096 1921
rect 26332 2091 26384 2100
rect 26332 2057 26341 2091
rect 26341 2057 26375 2091
rect 26375 2057 26384 2091
rect 26332 2048 26384 2057
rect 27436 2048 27488 2100
rect 27896 2048 27948 2100
rect 28632 2048 28684 2100
rect 28724 2091 28776 2100
rect 28724 2057 28733 2091
rect 28733 2057 28767 2091
rect 28767 2057 28776 2091
rect 28724 2048 28776 2057
rect 29184 2023 29236 2032
rect 29184 1989 29193 2023
rect 29193 1989 29227 2023
rect 29227 1989 29236 2023
rect 29184 1980 29236 1989
rect 27344 1912 27396 1964
rect 29276 1912 29328 1964
rect 24216 1708 24268 1760
rect 24584 1708 24636 1760
rect 26976 1844 27028 1896
rect 27804 1844 27856 1896
rect 28908 1844 28960 1896
rect 27068 1708 27120 1760
rect 27528 1708 27580 1760
rect 27712 1708 27764 1760
rect 28816 1708 28868 1760
rect 30012 1844 30064 1896
rect 7988 1606 8040 1658
rect 8052 1606 8104 1658
rect 8116 1606 8168 1658
rect 8180 1606 8232 1658
rect 8244 1606 8296 1658
rect 15578 1606 15630 1658
rect 15642 1606 15694 1658
rect 15706 1606 15758 1658
rect 15770 1606 15822 1658
rect 15834 1606 15886 1658
rect 23168 1606 23220 1658
rect 23232 1606 23284 1658
rect 23296 1606 23348 1658
rect 23360 1606 23412 1658
rect 23424 1606 23476 1658
rect 30758 1606 30810 1658
rect 30822 1606 30874 1658
rect 30886 1606 30938 1658
rect 30950 1606 31002 1658
rect 31014 1606 31066 1658
rect 1768 1547 1820 1556
rect 1768 1513 1783 1547
rect 1783 1513 1817 1547
rect 1817 1513 1820 1547
rect 1768 1504 1820 1513
rect 3792 1504 3844 1556
rect 4620 1504 4672 1556
rect 5540 1547 5592 1556
rect 5540 1513 5549 1547
rect 5549 1513 5583 1547
rect 5583 1513 5592 1547
rect 5540 1504 5592 1513
rect 6828 1504 6880 1556
rect 5080 1436 5132 1488
rect 9036 1504 9088 1556
rect 11704 1504 11756 1556
rect 12256 1504 12308 1556
rect 13636 1547 13688 1556
rect 13636 1513 13645 1547
rect 13645 1513 13679 1547
rect 13679 1513 13688 1547
rect 13636 1504 13688 1513
rect 14096 1504 14148 1556
rect 16580 1547 16632 1556
rect 16580 1513 16595 1547
rect 16595 1513 16629 1547
rect 16629 1513 16632 1547
rect 16580 1504 16632 1513
rect 18696 1504 18748 1556
rect 19432 1504 19484 1556
rect 21180 1504 21232 1556
rect 22744 1504 22796 1556
rect 24492 1504 24544 1556
rect 1216 1411 1268 1420
rect 1216 1377 1225 1411
rect 1225 1377 1259 1411
rect 1259 1377 1268 1411
rect 1216 1368 1268 1377
rect 1308 1411 1360 1420
rect 1308 1377 1317 1411
rect 1317 1377 1351 1411
rect 1351 1377 1360 1411
rect 1308 1368 1360 1377
rect 1952 1368 2004 1420
rect 2044 1343 2096 1352
rect 2044 1309 2053 1343
rect 2053 1309 2087 1343
rect 2087 1309 2096 1343
rect 2044 1300 2096 1309
rect 3332 1300 3384 1352
rect 3884 1300 3936 1352
rect 4068 1300 4120 1352
rect 5356 1300 5408 1352
rect 5816 1411 5868 1420
rect 5816 1377 5825 1411
rect 5825 1377 5859 1411
rect 5859 1377 5868 1411
rect 5816 1368 5868 1377
rect 6460 1411 6512 1420
rect 6460 1377 6469 1411
rect 6469 1377 6503 1411
rect 6503 1377 6512 1411
rect 6460 1368 6512 1377
rect 8668 1411 8720 1420
rect 8668 1377 8677 1411
rect 8677 1377 8711 1411
rect 8711 1377 8720 1411
rect 8668 1368 8720 1377
rect 9496 1368 9548 1420
rect 11152 1368 11204 1420
rect 11520 1411 11572 1420
rect 11520 1377 11529 1411
rect 11529 1377 11563 1411
rect 11563 1377 11572 1411
rect 11520 1368 11572 1377
rect 11612 1411 11664 1420
rect 11612 1377 11621 1411
rect 11621 1377 11655 1411
rect 11655 1377 11664 1411
rect 11612 1368 11664 1377
rect 12256 1368 12308 1420
rect 13544 1368 13596 1420
rect 9036 1343 9088 1352
rect 9036 1309 9038 1343
rect 9038 1309 9088 1343
rect 9036 1300 9088 1309
rect 9220 1300 9272 1352
rect 9312 1300 9364 1352
rect 12164 1300 12216 1352
rect 14004 1300 14056 1352
rect 16028 1300 16080 1352
rect 16856 1343 16908 1352
rect 16856 1309 16865 1343
rect 16865 1309 16899 1343
rect 16899 1309 16908 1343
rect 16856 1300 16908 1309
rect 18512 1300 18564 1352
rect 20720 1411 20772 1420
rect 20720 1377 20729 1411
rect 20729 1377 20763 1411
rect 20763 1377 20772 1411
rect 20720 1368 20772 1377
rect 20812 1368 20864 1420
rect 20996 1411 21048 1420
rect 20996 1377 21005 1411
rect 21005 1377 21039 1411
rect 21039 1377 21048 1411
rect 20996 1368 21048 1377
rect 23572 1368 23624 1420
rect 24032 1368 24084 1420
rect 27252 1504 27304 1556
rect 27528 1504 27580 1556
rect 28632 1504 28684 1556
rect 22836 1300 22888 1352
rect 23480 1343 23532 1352
rect 23480 1309 23489 1343
rect 23489 1309 23523 1343
rect 23523 1309 23532 1343
rect 23480 1300 23532 1309
rect 23940 1343 23992 1352
rect 23940 1309 23952 1343
rect 23952 1309 23986 1343
rect 23986 1309 23992 1343
rect 23940 1300 23992 1309
rect 24584 1300 24636 1352
rect 25596 1411 25648 1420
rect 25596 1377 25605 1411
rect 25605 1377 25639 1411
rect 25639 1377 25648 1411
rect 25596 1368 25648 1377
rect 25688 1368 25740 1420
rect 26608 1411 26660 1420
rect 26608 1377 26617 1411
rect 26617 1377 26651 1411
rect 26651 1377 26660 1411
rect 26608 1368 26660 1377
rect 26976 1411 27028 1420
rect 26976 1377 26985 1411
rect 26985 1377 27019 1411
rect 27019 1377 27028 1411
rect 26976 1368 27028 1377
rect 27436 1368 27488 1420
rect 27804 1368 27856 1420
rect 29736 1411 29788 1420
rect 29736 1377 29745 1411
rect 29745 1377 29779 1411
rect 29779 1377 29788 1411
rect 29736 1368 29788 1377
rect 8024 1164 8076 1216
rect 9772 1164 9824 1216
rect 12348 1164 12400 1216
rect 14280 1164 14332 1216
rect 19432 1164 19484 1216
rect 21916 1164 21968 1216
rect 26332 1232 26384 1284
rect 27712 1300 27764 1352
rect 28080 1300 28132 1352
rect 28172 1300 28224 1352
rect 23848 1164 23900 1216
rect 24400 1164 24452 1216
rect 26700 1207 26752 1216
rect 26700 1173 26709 1207
rect 26709 1173 26743 1207
rect 26743 1173 26752 1207
rect 26700 1164 26752 1173
rect 26884 1164 26936 1216
rect 29828 1164 29880 1216
rect 29920 1207 29972 1216
rect 29920 1173 29929 1207
rect 29929 1173 29963 1207
rect 29963 1173 29972 1207
rect 29920 1164 29972 1173
rect 4193 1062 4245 1114
rect 4257 1062 4309 1114
rect 4321 1062 4373 1114
rect 4385 1062 4437 1114
rect 4449 1062 4501 1114
rect 11783 1062 11835 1114
rect 11847 1062 11899 1114
rect 11911 1062 11963 1114
rect 11975 1062 12027 1114
rect 12039 1062 12091 1114
rect 19373 1062 19425 1114
rect 19437 1062 19489 1114
rect 19501 1062 19553 1114
rect 19565 1062 19617 1114
rect 19629 1062 19681 1114
rect 26963 1062 27015 1114
rect 27027 1062 27079 1114
rect 27091 1062 27143 1114
rect 27155 1062 27207 1114
rect 27219 1062 27271 1114
rect 3332 960 3384 1012
rect 3516 1003 3568 1012
rect 3516 969 3525 1003
rect 3525 969 3559 1003
rect 3559 969 3568 1003
rect 3516 960 3568 969
rect 4804 960 4856 1012
rect 4988 960 5040 1012
rect 5264 960 5316 1012
rect 1492 824 1544 876
rect 9220 960 9272 1012
rect 10968 1003 11020 1012
rect 10968 969 10977 1003
rect 10977 969 11011 1003
rect 11011 969 11020 1003
rect 10968 960 11020 969
rect 8300 892 8352 944
rect 5172 824 5224 876
rect 6460 824 6512 876
rect 6644 824 6696 876
rect 6736 824 6788 876
rect 7288 824 7340 876
rect 3608 756 3660 808
rect 5632 799 5684 808
rect 5632 765 5641 799
rect 5641 765 5675 799
rect 5675 765 5684 799
rect 5632 756 5684 765
rect 6000 799 6052 808
rect 6000 765 6009 799
rect 6009 765 6043 799
rect 6043 765 6052 799
rect 6000 756 6052 765
rect 3792 620 3844 672
rect 4252 663 4304 672
rect 4252 629 4261 663
rect 4261 629 4295 663
rect 4295 629 4304 663
rect 4252 620 4304 629
rect 8024 756 8076 808
rect 8668 867 8720 876
rect 8668 833 8677 867
rect 8677 833 8711 867
rect 8711 833 8720 867
rect 8668 824 8720 833
rect 9036 867 9088 876
rect 9036 833 9038 867
rect 9038 833 9088 867
rect 9036 824 9088 833
rect 8576 799 8628 808
rect 8576 765 8585 799
rect 8585 765 8619 799
rect 8619 765 8628 799
rect 8576 756 8628 765
rect 9404 867 9456 876
rect 9404 833 9413 867
rect 9413 833 9447 867
rect 9447 833 9456 867
rect 9404 824 9456 833
rect 14372 960 14424 1012
rect 16856 960 16908 1012
rect 17776 960 17828 1012
rect 11796 824 11848 876
rect 13636 824 13688 876
rect 11152 799 11204 808
rect 11152 765 11161 799
rect 11161 765 11195 799
rect 11195 765 11204 799
rect 11152 756 11204 765
rect 10232 688 10284 740
rect 11888 756 11940 808
rect 18236 935 18288 944
rect 18236 901 18245 935
rect 18245 901 18279 935
rect 18279 901 18288 935
rect 18236 892 18288 901
rect 14280 824 14332 876
rect 12992 756 13044 808
rect 13820 799 13872 808
rect 13820 765 13829 799
rect 13829 765 13863 799
rect 13863 765 13872 799
rect 13820 756 13872 765
rect 14556 799 14608 808
rect 14556 765 14565 799
rect 14565 765 14599 799
rect 14599 765 14608 799
rect 14556 756 14608 765
rect 15384 756 15436 808
rect 20720 960 20772 1012
rect 18880 892 18932 944
rect 19156 824 19208 876
rect 19340 867 19392 876
rect 19340 833 19342 867
rect 19342 833 19392 867
rect 19340 824 19392 833
rect 19524 824 19576 876
rect 20720 824 20772 876
rect 17040 756 17092 808
rect 17132 799 17184 808
rect 17132 765 17141 799
rect 17141 765 17175 799
rect 17175 765 17184 799
rect 17132 756 17184 765
rect 21272 935 21324 944
rect 21272 901 21281 935
rect 21281 901 21315 935
rect 21315 901 21324 935
rect 21272 892 21324 901
rect 23480 960 23532 1012
rect 24584 960 24636 1012
rect 25688 1003 25740 1012
rect 25688 969 25697 1003
rect 25697 969 25731 1003
rect 25731 969 25740 1003
rect 25688 960 25740 969
rect 21916 824 21968 876
rect 23020 824 23072 876
rect 23572 824 23624 876
rect 6828 620 6880 672
rect 11612 620 11664 672
rect 13084 663 13136 672
rect 13084 629 13093 663
rect 13093 629 13127 663
rect 13127 629 13136 663
rect 13084 620 13136 629
rect 14464 620 14516 672
rect 16488 620 16540 672
rect 21364 688 21416 740
rect 22192 756 22244 808
rect 23848 799 23900 808
rect 23848 765 23857 799
rect 23857 765 23891 799
rect 23891 765 23900 799
rect 23848 756 23900 765
rect 26700 960 26752 1012
rect 28540 1003 28592 1012
rect 28540 969 28549 1003
rect 28549 969 28583 1003
rect 28583 969 28592 1003
rect 28540 960 28592 969
rect 29460 1003 29512 1012
rect 29460 969 29469 1003
rect 29469 969 29503 1003
rect 29503 969 29512 1003
rect 29460 960 29512 969
rect 29000 892 29052 944
rect 26884 824 26936 876
rect 28264 824 28316 876
rect 26332 756 26384 808
rect 27344 756 27396 808
rect 29092 824 29144 876
rect 29368 756 29420 808
rect 20444 620 20496 672
rect 22008 663 22060 672
rect 22008 629 22023 663
rect 22023 629 22057 663
rect 22057 629 22060 663
rect 22008 620 22060 629
rect 22192 620 22244 672
rect 23664 620 23716 672
rect 23940 620 23992 672
rect 24492 620 24544 672
rect 27528 620 27580 672
rect 7988 518 8040 570
rect 8052 518 8104 570
rect 8116 518 8168 570
rect 8180 518 8232 570
rect 8244 518 8296 570
rect 15578 518 15630 570
rect 15642 518 15694 570
rect 15706 518 15758 570
rect 15770 518 15822 570
rect 15834 518 15886 570
rect 23168 518 23220 570
rect 23232 518 23284 570
rect 23296 518 23348 570
rect 23360 518 23412 570
rect 23424 518 23476 570
rect 30758 518 30810 570
rect 30822 518 30874 570
rect 30886 518 30938 570
rect 30950 518 31002 570
rect 31014 518 31066 570
rect 1492 416 1544 468
rect 2044 416 2096 468
rect 5632 416 5684 468
rect 6000 416 6052 468
rect 10232 416 10284 468
rect 8576 348 8628 400
rect 10784 348 10836 400
rect 3976 280 4028 332
rect 14464 416 14516 468
rect 17132 416 17184 468
rect 19156 416 19208 468
rect 19524 416 19576 468
rect 22100 416 22152 468
rect 24308 416 24360 468
rect 13636 348 13688 400
rect 22928 348 22980 400
rect 7656 212 7708 264
rect 10784 212 10836 264
rect 12992 280 13044 332
rect 13084 280 13136 332
rect 17040 280 17092 332
rect 22100 280 22152 332
rect 22192 280 22244 332
rect 13820 144 13872 196
rect 16488 144 16540 196
rect 23756 144 23808 196
rect 22100 76 22152 128
rect 24216 76 24268 128
rect 3884 8 3936 60
rect 16212 8 16264 60
rect 18880 8 18932 60
<< metal2 >>
rect 8208 22296 8260 22302
rect 5078 22264 5134 22273
rect 5000 22222 5078 22250
rect 2502 21992 2558 22001
rect 2502 21927 2558 21936
rect 2136 21888 2188 21894
rect 2136 21830 2188 21836
rect 846 21584 902 21593
rect 846 21519 902 21528
rect 860 21146 888 21519
rect 2148 21486 2176 21830
rect 2516 21690 2544 21927
rect 4193 21788 4501 21797
rect 4193 21786 4199 21788
rect 4255 21786 4279 21788
rect 4335 21786 4359 21788
rect 4415 21786 4439 21788
rect 4495 21786 4501 21788
rect 4255 21734 4257 21786
rect 4437 21734 4439 21786
rect 4193 21732 4199 21734
rect 4255 21732 4279 21734
rect 4335 21732 4359 21734
rect 4415 21732 4439 21734
rect 4495 21732 4501 21734
rect 4193 21723 4501 21732
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 2872 21684 2924 21690
rect 2924 21644 3004 21672
rect 2872 21626 2924 21632
rect 2136 21480 2188 21486
rect 2136 21422 2188 21428
rect 1400 21412 1452 21418
rect 1400 21354 1452 21360
rect 2780 21412 2832 21418
rect 2780 21354 2832 21360
rect 848 21140 900 21146
rect 848 21082 900 21088
rect 1216 20392 1268 20398
rect 1216 20334 1268 20340
rect 1228 19922 1256 20334
rect 1412 20262 1440 21354
rect 1492 21344 1544 21350
rect 1492 21286 1544 21292
rect 1504 20942 1532 21286
rect 1858 21040 1914 21049
rect 1858 20975 1914 20984
rect 1872 20942 1900 20975
rect 1492 20936 1544 20942
rect 1492 20878 1544 20884
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1780 20602 1808 20878
rect 1768 20596 1820 20602
rect 1768 20538 1820 20544
rect 2792 20398 2820 21354
rect 1676 20392 1728 20398
rect 1676 20334 1728 20340
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 1400 20256 1452 20262
rect 1400 20198 1452 20204
rect 664 19916 716 19922
rect 664 19858 716 19864
rect 1216 19916 1268 19922
rect 1216 19858 1268 19864
rect 676 19825 704 19858
rect 662 19816 718 19825
rect 662 19751 718 19760
rect 676 16726 704 19751
rect 848 19712 900 19718
rect 848 19654 900 19660
rect 860 19514 888 19654
rect 848 19508 900 19514
rect 848 19450 900 19456
rect 1228 19310 1256 19858
rect 1688 19417 1716 20334
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1780 20058 1808 20198
rect 1768 20052 1820 20058
rect 1768 19994 1820 20000
rect 1674 19408 1730 19417
rect 1674 19343 1730 19352
rect 1216 19304 1268 19310
rect 1216 19246 1268 19252
rect 1032 18624 1084 18630
rect 1032 18566 1084 18572
rect 1044 17785 1072 18566
rect 1228 18426 1256 19246
rect 1780 19174 1808 19994
rect 2872 19916 2924 19922
rect 2872 19858 2924 19864
rect 1860 19848 1912 19854
rect 1912 19808 2176 19836
rect 1860 19790 1912 19796
rect 1768 19168 1820 19174
rect 1768 19110 1820 19116
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1308 18760 1360 18766
rect 1308 18702 1360 18708
rect 1216 18420 1268 18426
rect 1216 18362 1268 18368
rect 1216 18216 1268 18222
rect 1216 18158 1268 18164
rect 1122 17912 1178 17921
rect 1122 17847 1178 17856
rect 1136 17814 1164 17847
rect 1124 17808 1176 17814
rect 1030 17776 1086 17785
rect 848 17740 900 17746
rect 1124 17750 1176 17756
rect 1030 17711 1086 17720
rect 848 17682 900 17688
rect 664 16720 716 16726
rect 664 16662 716 16668
rect 676 14521 704 16662
rect 662 14512 718 14521
rect 662 14447 718 14456
rect 676 11082 704 14447
rect 756 13932 808 13938
rect 756 13874 808 13880
rect 664 11076 716 11082
rect 664 11018 716 11024
rect 676 10266 704 11018
rect 664 10260 716 10266
rect 664 10202 716 10208
rect 768 9042 796 13874
rect 860 13326 888 17682
rect 1228 17542 1256 18158
rect 1216 17536 1268 17542
rect 1216 17478 1268 17484
rect 1228 17134 1256 17478
rect 1216 17128 1268 17134
rect 1216 17070 1268 17076
rect 1228 16794 1256 17070
rect 1216 16788 1268 16794
rect 1216 16730 1268 16736
rect 1032 16448 1084 16454
rect 1032 16390 1084 16396
rect 940 14272 992 14278
rect 940 14214 992 14220
rect 952 13394 980 14214
rect 940 13388 992 13394
rect 940 13330 992 13336
rect 848 13320 900 13326
rect 848 13262 900 13268
rect 860 12986 888 13262
rect 848 12980 900 12986
rect 848 12922 900 12928
rect 1044 11150 1072 16390
rect 1124 16108 1176 16114
rect 1124 16050 1176 16056
rect 1136 15434 1164 16050
rect 1124 15428 1176 15434
rect 1124 15370 1176 15376
rect 1136 15026 1164 15370
rect 1216 15360 1268 15366
rect 1216 15302 1268 15308
rect 1124 15020 1176 15026
rect 1124 14962 1176 14968
rect 1136 14618 1164 14962
rect 1124 14612 1176 14618
rect 1124 14554 1176 14560
rect 1124 11892 1176 11898
rect 1124 11834 1176 11840
rect 1136 11354 1164 11834
rect 1228 11558 1256 15302
rect 1320 14074 1348 18702
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1412 15638 1440 15846
rect 1400 15632 1452 15638
rect 1400 15574 1452 15580
rect 1412 14822 1440 15574
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 1412 14414 1440 14758
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1308 14068 1360 14074
rect 1308 14010 1360 14016
rect 1596 13734 1624 18906
rect 1780 18086 1808 19110
rect 1952 18760 2004 18766
rect 1952 18702 2004 18708
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1768 18080 1820 18086
rect 1768 18022 1820 18028
rect 1688 17678 1716 18022
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1688 16998 1716 17614
rect 1964 17542 1992 18702
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1768 17128 1820 17134
rect 1768 17070 1820 17076
rect 2042 17096 2098 17105
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1688 16658 1716 16934
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1676 13864 1728 13870
rect 1674 13832 1676 13841
rect 1728 13832 1730 13841
rect 1674 13767 1730 13776
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1308 13320 1360 13326
rect 1308 13262 1360 13268
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1320 12782 1348 13262
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1596 12782 1624 13126
rect 1308 12776 1360 12782
rect 1308 12718 1360 12724
rect 1584 12776 1636 12782
rect 1584 12718 1636 12724
rect 1320 12238 1348 12718
rect 1688 12646 1716 13262
rect 1676 12640 1728 12646
rect 1780 12617 1808 17070
rect 2042 17031 2098 17040
rect 2056 16590 2084 17031
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1964 13569 1992 14350
rect 1950 13560 2006 13569
rect 1950 13495 2006 13504
rect 1676 12582 1728 12588
rect 1766 12608 1822 12617
rect 1688 12442 1716 12582
rect 1766 12543 1822 12552
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1308 12232 1360 12238
rect 1308 12174 1360 12180
rect 1320 11898 1348 12174
rect 1308 11892 1360 11898
rect 1308 11834 1360 11840
rect 1688 11778 1716 12378
rect 1950 12336 2006 12345
rect 1950 12271 2006 12280
rect 1964 12238 1992 12271
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2056 12102 2084 12174
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2148 11801 2176 19808
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2504 19304 2556 19310
rect 2504 19246 2556 19252
rect 2412 17672 2464 17678
rect 2412 17614 2464 17620
rect 2424 16697 2452 17614
rect 2410 16688 2466 16697
rect 2410 16623 2466 16632
rect 2226 16008 2282 16017
rect 2226 15943 2282 15952
rect 2240 13326 2268 15943
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12753 2268 13126
rect 2226 12744 2282 12753
rect 2226 12679 2282 12688
rect 1320 11762 1716 11778
rect 1308 11756 1716 11762
rect 1360 11750 1716 11756
rect 1308 11698 1360 11704
rect 1216 11552 1268 11558
rect 1216 11494 1268 11500
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1124 11348 1176 11354
rect 1124 11290 1176 11296
rect 1136 11150 1164 11290
rect 1596 11286 1624 11494
rect 1584 11280 1636 11286
rect 1584 11222 1636 11228
rect 1688 11150 1716 11750
rect 2134 11792 2190 11801
rect 2134 11727 2190 11736
rect 1032 11144 1084 11150
rect 1032 11086 1084 11092
rect 1124 11144 1176 11150
rect 1124 11086 1176 11092
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1136 10674 1164 11086
rect 1124 10668 1176 10674
rect 1124 10610 1176 10616
rect 1136 10130 1164 10610
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1412 10266 1440 10406
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 1124 10124 1176 10130
rect 1124 10066 1176 10072
rect 848 9716 900 9722
rect 848 9658 900 9664
rect 860 9178 888 9658
rect 1136 9586 1164 10066
rect 1124 9580 1176 9586
rect 1124 9522 1176 9528
rect 1412 9382 1440 10202
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 848 9172 900 9178
rect 848 9114 900 9120
rect 1412 9110 1440 9318
rect 1400 9104 1452 9110
rect 1596 9058 1624 10542
rect 1688 10470 1716 11086
rect 2134 10704 2190 10713
rect 2134 10639 2136 10648
rect 2188 10639 2190 10648
rect 2136 10610 2188 10616
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1872 9722 1900 9998
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1400 9046 1452 9052
rect 756 9036 808 9042
rect 756 8978 808 8984
rect 1504 9030 1624 9058
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1124 8628 1176 8634
rect 1124 8570 1176 8576
rect 1032 7948 1084 7954
rect 1032 7890 1084 7896
rect 1044 7857 1072 7890
rect 1030 7848 1086 7857
rect 1030 7783 1086 7792
rect 1136 6730 1164 8570
rect 1216 8424 1268 8430
rect 1216 8366 1268 8372
rect 1228 7750 1256 8366
rect 1412 8294 1440 8910
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 7886 1440 8230
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1216 7744 1268 7750
rect 1216 7686 1268 7692
rect 1228 7342 1256 7686
rect 1216 7336 1268 7342
rect 1216 7278 1268 7284
rect 1228 6866 1256 7278
rect 1412 7206 1440 7822
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1412 7002 1440 7142
rect 1400 6996 1452 7002
rect 1400 6938 1452 6944
rect 1216 6860 1268 6866
rect 1216 6802 1268 6808
rect 1124 6724 1176 6730
rect 1176 6684 1256 6712
rect 1124 6666 1176 6672
rect 940 6248 992 6254
rect 940 6190 992 6196
rect 952 5710 980 6190
rect 1122 6080 1178 6089
rect 1122 6015 1178 6024
rect 1032 5772 1084 5778
rect 1032 5714 1084 5720
rect 940 5704 992 5710
rect 940 5646 992 5652
rect 952 5166 980 5646
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 952 4729 980 5102
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 952 4622 980 4655
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 952 4078 980 4558
rect 940 4072 992 4078
rect 940 4014 992 4020
rect 952 2582 980 4014
rect 940 2576 992 2582
rect 940 2518 992 2524
rect 1044 2258 1072 5714
rect 1136 2514 1164 6015
rect 1124 2508 1176 2514
rect 1124 2450 1176 2456
rect 1044 2230 1164 2258
rect 1136 1465 1164 2230
rect 1122 1456 1178 1465
rect 1228 1426 1256 6684
rect 1504 6662 1532 9030
rect 1688 8090 1716 9454
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2056 9042 2084 9318
rect 2044 9036 2096 9042
rect 2044 8978 2096 8984
rect 1768 8424 1820 8430
rect 2136 8424 2188 8430
rect 1820 8384 1900 8412
rect 1768 8366 1820 8372
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1768 6792 1820 6798
rect 1766 6760 1768 6769
rect 1820 6760 1822 6769
rect 1766 6695 1822 6704
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1676 6248 1728 6254
rect 1676 6190 1728 6196
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1412 5778 1440 6054
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1412 5030 1440 5714
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1412 4690 1440 4966
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1412 3942 1440 4626
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 1412 2774 1440 3878
rect 1504 3534 1532 5510
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1596 3738 1624 3878
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1492 3528 1544 3534
rect 1492 3470 1544 3476
rect 1596 2990 1624 3674
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 1688 2774 1716 6190
rect 1872 4826 1900 8384
rect 2136 8366 2188 8372
rect 2042 8120 2098 8129
rect 2042 8055 2098 8064
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1964 5914 1992 7822
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2056 5794 2084 8055
rect 1964 5766 2084 5794
rect 1860 4820 1912 4826
rect 1860 4762 1912 4768
rect 1964 4078 1992 5766
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2056 5574 2084 5646
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 1780 2854 1808 3674
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 1412 2746 1532 2774
rect 1504 2394 1532 2746
rect 1596 2746 1716 2774
rect 1596 2666 1624 2746
rect 1596 2638 1716 2666
rect 1688 2514 1716 2638
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 1780 2394 1808 2586
rect 1504 2366 1808 2394
rect 1308 2100 1360 2106
rect 1308 2042 1360 2048
rect 1320 1426 1348 2042
rect 1768 1760 1820 1766
rect 1768 1702 1820 1708
rect 1780 1562 1808 1702
rect 1768 1556 1820 1562
rect 1768 1498 1820 1504
rect 2056 1442 2084 4966
rect 2148 1902 2176 8366
rect 2240 3777 2268 12679
rect 2332 9042 2360 13670
rect 2516 13190 2544 19246
rect 2792 18426 2820 19314
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 2594 16144 2650 16153
rect 2594 16079 2650 16088
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2608 12050 2636 16079
rect 2700 12442 2728 18158
rect 2884 17338 2912 19858
rect 2976 19242 3004 21644
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 3068 19310 3096 21490
rect 3240 21480 3292 21486
rect 3976 21480 4028 21486
rect 3240 21422 3292 21428
rect 3620 21428 3976 21434
rect 3620 21422 4028 21428
rect 3252 20942 3280 21422
rect 3620 21406 4016 21422
rect 3240 20936 3292 20942
rect 3240 20878 3292 20884
rect 3516 20936 3568 20942
rect 3516 20878 3568 20884
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 2964 19236 3016 19242
rect 2964 19178 3016 19184
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2792 15162 2820 17138
rect 2976 16250 3004 18226
rect 3160 17921 3188 19246
rect 3146 17912 3202 17921
rect 3146 17847 3202 17856
rect 3148 17740 3200 17746
rect 3148 17682 3200 17688
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2962 15464 3018 15473
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2516 12022 2636 12050
rect 2516 11762 2544 12022
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2594 8528 2650 8537
rect 2594 8463 2650 8472
rect 2320 8288 2372 8294
rect 2320 8230 2372 8236
rect 2332 5030 2360 8230
rect 2412 7472 2464 7478
rect 2412 7414 2464 7420
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2424 4298 2452 7414
rect 2332 4270 2452 4298
rect 2226 3768 2282 3777
rect 2226 3703 2282 3712
rect 2332 2514 2360 4270
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 2424 3534 2452 4150
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2516 3738 2544 4014
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 2608 1970 2636 8463
rect 2700 8430 2728 9658
rect 2792 9654 2820 13670
rect 2884 11665 2912 15438
rect 2962 15399 3018 15408
rect 2976 15026 3004 15399
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 3068 14618 3096 16594
rect 3160 15706 3188 17682
rect 3252 16794 3280 20402
rect 3528 19854 3556 20878
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3344 18057 3372 18566
rect 3436 18426 3464 18702
rect 3516 18692 3568 18698
rect 3516 18634 3568 18640
rect 3528 18465 3556 18634
rect 3514 18456 3570 18465
rect 3424 18420 3476 18426
rect 3514 18391 3570 18400
rect 3424 18362 3476 18368
rect 3514 18320 3570 18329
rect 3436 18278 3514 18306
rect 3330 18048 3386 18057
rect 3330 17983 3386 17992
rect 3436 17134 3464 18278
rect 3514 18255 3570 18264
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3528 17814 3556 18158
rect 3516 17808 3568 17814
rect 3516 17750 3568 17756
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 3332 16720 3384 16726
rect 3332 16662 3384 16668
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3148 15700 3200 15706
rect 3148 15642 3200 15648
rect 3252 14958 3280 16594
rect 3344 15978 3372 16662
rect 3436 16658 3464 17070
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3528 16114 3556 17138
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3332 15972 3384 15978
rect 3332 15914 3384 15920
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3528 15502 3556 15846
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 3240 14952 3292 14958
rect 3620 14929 3648 21406
rect 3700 21344 3752 21350
rect 3700 21286 3752 21292
rect 3712 21146 3740 21286
rect 3700 21140 3752 21146
rect 3700 21082 3752 21088
rect 3712 20942 3740 21082
rect 3700 20936 3752 20942
rect 3700 20878 3752 20884
rect 3792 20936 3844 20942
rect 4068 20936 4120 20942
rect 3792 20878 3844 20884
rect 4066 20904 4068 20913
rect 4120 20904 4122 20913
rect 3712 19938 3740 20878
rect 3804 20058 3832 20878
rect 4066 20839 4122 20848
rect 4193 20700 4501 20709
rect 4193 20698 4199 20700
rect 4255 20698 4279 20700
rect 4335 20698 4359 20700
rect 4415 20698 4439 20700
rect 4495 20698 4501 20700
rect 4255 20646 4257 20698
rect 4437 20646 4439 20698
rect 4193 20644 4199 20646
rect 4255 20644 4279 20646
rect 4335 20644 4359 20646
rect 4415 20644 4439 20646
rect 4495 20644 4501 20646
rect 4193 20635 4501 20644
rect 4712 20392 4764 20398
rect 4710 20360 4712 20369
rect 4896 20392 4948 20398
rect 4764 20360 4766 20369
rect 3976 20324 4028 20330
rect 4710 20295 4766 20304
rect 4816 20340 4896 20346
rect 4816 20334 4948 20340
rect 4816 20318 4936 20334
rect 3976 20266 4028 20272
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3712 19910 3924 19938
rect 3896 19854 3924 19910
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3712 19446 3740 19790
rect 3700 19440 3752 19446
rect 3700 19382 3752 19388
rect 3896 19310 3924 19790
rect 3988 19514 4016 20266
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 4620 20256 4672 20262
rect 4620 20198 4672 20204
rect 4264 20058 4292 20198
rect 4252 20052 4304 20058
rect 4252 19994 4304 20000
rect 4193 19612 4501 19621
rect 4193 19610 4199 19612
rect 4255 19610 4279 19612
rect 4335 19610 4359 19612
rect 4415 19610 4439 19612
rect 4495 19610 4501 19612
rect 4255 19558 4257 19610
rect 4437 19558 4439 19610
rect 4193 19556 4199 19558
rect 4255 19556 4279 19558
rect 4335 19556 4359 19558
rect 4415 19556 4439 19558
rect 4495 19556 4501 19558
rect 4193 19547 4501 19556
rect 4632 19514 4660 20198
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 4252 19440 4304 19446
rect 4252 19382 4304 19388
rect 3792 19304 3844 19310
rect 3792 19246 3844 19252
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3700 18828 3752 18834
rect 3700 18770 3752 18776
rect 3712 18630 3740 18770
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3240 14894 3292 14900
rect 3606 14920 3662 14929
rect 3606 14855 3662 14864
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 3608 14544 3660 14550
rect 3608 14486 3660 14492
rect 2962 14376 3018 14385
rect 2962 14311 3018 14320
rect 2870 11656 2926 11665
rect 2870 11591 2926 11600
rect 2976 11150 3004 14311
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3054 12880 3110 12889
rect 3054 12815 3056 12824
rect 3108 12815 3110 12824
rect 3056 12786 3108 12792
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2976 9382 3004 10202
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 3068 9722 3096 9862
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2792 8514 2820 8774
rect 2884 8634 2912 8910
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2792 8486 2912 8514
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2688 7336 2740 7342
rect 2792 7313 2820 8366
rect 2688 7278 2740 7284
rect 2778 7304 2834 7313
rect 2700 7002 2728 7278
rect 2778 7239 2834 7248
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2792 4622 2820 7142
rect 2884 5710 2912 8486
rect 2976 8265 3004 8910
rect 3068 8566 3096 8910
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 2962 8256 3018 8265
rect 2962 8191 3018 8200
rect 2962 7440 3018 7449
rect 2962 7375 2964 7384
rect 3016 7375 3018 7384
rect 2964 7346 3016 7352
rect 2962 6896 3018 6905
rect 2962 6831 3018 6840
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2976 5098 3004 6831
rect 2964 5092 3016 5098
rect 2964 5034 3016 5040
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 3068 4146 3096 8298
rect 3160 4826 3188 13874
rect 3252 9654 3280 14214
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3436 13190 3464 13806
rect 3528 13274 3556 13806
rect 3620 13433 3648 14486
rect 3606 13424 3662 13433
rect 3606 13359 3662 13368
rect 3606 13288 3662 13297
rect 3528 13246 3606 13274
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3436 12714 3464 13126
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3436 12170 3464 12650
rect 3528 12374 3556 13246
rect 3606 13223 3662 13232
rect 3516 12368 3568 12374
rect 3516 12310 3568 12316
rect 3424 12164 3476 12170
rect 3424 12106 3476 12112
rect 3436 11694 3464 12106
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3436 11150 3464 11630
rect 3620 11354 3648 11630
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3712 11257 3740 18566
rect 3804 18329 3832 19246
rect 3790 18320 3846 18329
rect 3896 18290 3924 19246
rect 4264 19242 4292 19382
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4434 19272 4490 19281
rect 4252 19236 4304 19242
rect 4252 19178 4304 19184
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 3976 18828 4028 18834
rect 3976 18770 4028 18776
rect 3988 18426 4016 18770
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 3790 18255 3846 18264
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 4080 18222 4108 19110
rect 4172 18884 4200 19110
rect 4356 19009 4384 19246
rect 4724 19242 4752 19790
rect 4816 19242 4844 20318
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4434 19207 4490 19216
rect 4620 19236 4672 19242
rect 4342 19000 4398 19009
rect 4342 18935 4398 18944
rect 4448 18952 4476 19207
rect 4620 19178 4672 19184
rect 4712 19236 4764 19242
rect 4712 19178 4764 19184
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 4632 19145 4660 19178
rect 4618 19136 4674 19145
rect 4908 19122 4936 20198
rect 5000 19242 5028 22222
rect 11152 22296 11204 22302
rect 8208 22238 8260 22244
rect 11150 22264 11152 22273
rect 12256 22296 12308 22302
rect 11204 22264 11206 22273
rect 5078 22199 5134 22208
rect 6460 22228 6512 22234
rect 6460 22170 6512 22176
rect 6092 22160 6144 22166
rect 6092 22102 6144 22108
rect 6104 21622 6132 22102
rect 6472 21690 6500 22170
rect 6644 21956 6696 21962
rect 6644 21898 6696 21904
rect 6460 21684 6512 21690
rect 6460 21626 6512 21632
rect 6092 21616 6144 21622
rect 6092 21558 6144 21564
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 5092 20466 5120 21286
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5080 19848 5132 19854
rect 5080 19790 5132 19796
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 5092 19378 5120 19790
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 4988 19236 5040 19242
rect 4988 19178 5040 19184
rect 4618 19071 4674 19080
rect 4724 19094 4936 19122
rect 4448 18924 4568 18952
rect 4172 18856 4476 18884
rect 4172 18766 4200 18856
rect 4160 18760 4212 18766
rect 4448 18737 4476 18856
rect 4160 18702 4212 18708
rect 4250 18728 4306 18737
rect 4434 18728 4490 18737
rect 4344 18692 4396 18698
rect 4306 18672 4344 18680
rect 4250 18663 4344 18672
rect 4264 18652 4344 18663
rect 4540 18698 4568 18924
rect 4724 18884 4752 19094
rect 4632 18856 4752 18884
rect 4802 18864 4858 18873
rect 4632 18698 4660 18856
rect 4724 18808 4802 18816
rect 4724 18799 4858 18808
rect 4896 18828 4948 18834
rect 4724 18788 4844 18799
rect 4724 18698 4752 18788
rect 4896 18770 4948 18776
rect 4434 18663 4490 18672
rect 4528 18692 4580 18698
rect 4344 18634 4396 18640
rect 4528 18634 4580 18640
rect 4620 18692 4672 18698
rect 4620 18634 4672 18640
rect 4712 18692 4764 18698
rect 4712 18634 4764 18640
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4193 18524 4501 18533
rect 4193 18522 4199 18524
rect 4255 18522 4279 18524
rect 4335 18522 4359 18524
rect 4415 18522 4439 18524
rect 4495 18522 4501 18524
rect 4255 18470 4257 18522
rect 4437 18470 4439 18522
rect 4193 18468 4199 18470
rect 4255 18468 4279 18470
rect 4335 18468 4359 18470
rect 4415 18468 4439 18470
rect 4495 18468 4501 18470
rect 4193 18459 4501 18468
rect 4816 18426 4844 18566
rect 4804 18420 4856 18426
rect 4908 18408 4936 18770
rect 5184 18426 5212 19790
rect 5460 19718 5488 20334
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 5446 19408 5502 19417
rect 5552 19378 5580 20742
rect 5446 19343 5502 19352
rect 5540 19372 5592 19378
rect 5356 19236 5408 19242
rect 5356 19178 5408 19184
rect 5172 18420 5224 18426
rect 4908 18380 5028 18408
rect 4804 18362 4856 18368
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 4526 18184 4582 18193
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3804 17134 3832 17478
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3804 16658 3832 17070
rect 3896 16998 3924 17614
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 3988 16697 4016 18158
rect 4582 18142 4660 18170
rect 4526 18119 4582 18128
rect 4632 17882 4660 18142
rect 4816 17954 4844 18362
rect 4894 18184 4950 18193
rect 4894 18119 4950 18128
rect 4724 17926 4844 17954
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4540 17649 4568 17818
rect 4526 17640 4582 17649
rect 4526 17575 4582 17584
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 4080 17202 4108 17478
rect 4193 17436 4501 17445
rect 4193 17434 4199 17436
rect 4255 17434 4279 17436
rect 4335 17434 4359 17436
rect 4415 17434 4439 17436
rect 4495 17434 4501 17436
rect 4255 17382 4257 17434
rect 4437 17382 4439 17434
rect 4193 17380 4199 17382
rect 4255 17380 4279 17382
rect 4335 17380 4359 17382
rect 4415 17380 4439 17382
rect 4495 17380 4501 17382
rect 4193 17371 4501 17380
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 4436 17196 4488 17202
rect 4436 17138 4488 17144
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4264 16794 4292 16934
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 3974 16688 4030 16697
rect 3792 16652 3844 16658
rect 3974 16623 4030 16632
rect 3792 16594 3844 16600
rect 4448 16590 4476 17138
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 3976 16448 4028 16454
rect 3976 16390 4028 16396
rect 3988 16250 4016 16390
rect 4080 16250 4108 16526
rect 4193 16348 4501 16357
rect 4193 16346 4199 16348
rect 4255 16346 4279 16348
rect 4335 16346 4359 16348
rect 4415 16346 4439 16348
rect 4495 16346 4501 16348
rect 4255 16294 4257 16346
rect 4437 16294 4439 16346
rect 4193 16292 4199 16294
rect 4255 16292 4279 16294
rect 4335 16292 4359 16294
rect 4415 16292 4439 16294
rect 4495 16292 4501 16294
rect 4193 16283 4501 16292
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 4540 16046 4568 17274
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 4528 16040 4580 16046
rect 4528 15982 4580 15988
rect 3896 15502 3924 15982
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4172 15502 4200 15846
rect 4724 15706 4752 17926
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 14958 3832 15302
rect 3896 14958 3924 15438
rect 4193 15260 4501 15269
rect 4193 15258 4199 15260
rect 4255 15258 4279 15260
rect 4335 15258 4359 15260
rect 4415 15258 4439 15260
rect 4495 15258 4501 15260
rect 4255 15206 4257 15258
rect 4437 15206 4439 15258
rect 4193 15204 4199 15206
rect 4255 15204 4279 15206
rect 4335 15204 4359 15206
rect 4415 15204 4439 15206
rect 4495 15204 4501 15206
rect 4193 15195 4501 15204
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 3804 14482 3832 14894
rect 3896 14618 3924 14894
rect 4158 14648 4214 14657
rect 3884 14612 3936 14618
rect 4158 14583 4214 14592
rect 3884 14554 3936 14560
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 4172 14414 4200 14583
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4193 14172 4501 14181
rect 4193 14170 4199 14172
rect 4255 14170 4279 14172
rect 4335 14170 4359 14172
rect 4415 14170 4439 14172
rect 4495 14170 4501 14172
rect 4255 14118 4257 14170
rect 4437 14118 4439 14170
rect 4193 14116 4199 14118
rect 4255 14116 4279 14118
rect 4335 14116 4359 14118
rect 4415 14116 4439 14118
rect 4495 14116 4501 14118
rect 4193 14107 4501 14116
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3804 12782 3832 13126
rect 3792 12776 3844 12782
rect 3792 12718 3844 12724
rect 3896 11898 3924 13874
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3988 13530 4016 13670
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 3988 12646 4016 13466
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3988 12220 4016 12582
rect 4080 12322 4108 14010
rect 4193 13084 4501 13093
rect 4193 13082 4199 13084
rect 4255 13082 4279 13084
rect 4335 13082 4359 13084
rect 4415 13082 4439 13084
rect 4495 13082 4501 13084
rect 4255 13030 4257 13082
rect 4437 13030 4439 13082
rect 4193 13028 4199 13030
rect 4255 13028 4279 13030
rect 4335 13028 4359 13030
rect 4415 13028 4439 13030
rect 4495 13028 4501 13030
rect 4193 13019 4501 13028
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4264 12850 4292 12922
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4080 12306 4200 12322
rect 4080 12300 4212 12306
rect 4080 12294 4160 12300
rect 4160 12242 4212 12248
rect 4068 12232 4120 12238
rect 3988 12192 4068 12220
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3988 11558 4016 12192
rect 4068 12174 4120 12180
rect 4193 11996 4501 12005
rect 4193 11994 4199 11996
rect 4255 11994 4279 11996
rect 4335 11994 4359 11996
rect 4415 11994 4439 11996
rect 4495 11994 4501 11996
rect 4255 11942 4257 11994
rect 4437 11942 4439 11994
rect 4193 11940 4199 11942
rect 4255 11940 4279 11942
rect 4335 11940 4359 11942
rect 4415 11940 4439 11942
rect 4495 11940 4501 11942
rect 4193 11931 4501 11940
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3698 11248 3754 11257
rect 3988 11218 4016 11494
rect 4080 11354 4108 11630
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4356 11286 4384 11630
rect 4540 11354 4568 14894
rect 4724 14618 4752 15642
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4908 13025 4936 18119
rect 5000 16998 5028 18380
rect 5172 18362 5224 18368
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 5276 18193 5304 18362
rect 5262 18184 5318 18193
rect 5262 18119 5318 18128
rect 5262 18048 5318 18057
rect 5092 18006 5262 18034
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 4988 16516 5040 16522
rect 4988 16458 5040 16464
rect 5000 15706 5028 16458
rect 4988 15700 5040 15706
rect 4988 15642 5040 15648
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 5000 13258 5028 15098
rect 4988 13252 5040 13258
rect 4988 13194 5040 13200
rect 5092 13161 5120 18006
rect 5262 17983 5318 17992
rect 5170 17912 5226 17921
rect 5170 17847 5226 17856
rect 5184 13977 5212 17847
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 5170 13968 5226 13977
rect 5170 13903 5226 13912
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5184 13530 5212 13806
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5078 13152 5134 13161
rect 5078 13087 5134 13096
rect 4894 13016 4950 13025
rect 4894 12951 4950 12960
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 3698 11183 3754 11192
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3436 10690 3464 11086
rect 3344 10662 3464 10690
rect 3344 10606 3372 10662
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3344 10062 3372 10542
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3712 10146 3740 10202
rect 3804 10146 3832 11154
rect 3988 10470 4016 11154
rect 4193 10908 4501 10917
rect 4193 10906 4199 10908
rect 4255 10906 4279 10908
rect 4335 10906 4359 10908
rect 4415 10906 4439 10908
rect 4495 10906 4501 10908
rect 4255 10854 4257 10906
rect 4437 10854 4439 10906
rect 4193 10852 4199 10854
rect 4255 10852 4279 10854
rect 4335 10852 4359 10854
rect 4415 10852 4439 10854
rect 4495 10852 4501 10854
rect 4193 10843 4501 10852
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3988 10266 4016 10406
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3712 10130 3924 10146
rect 3712 10124 3936 10130
rect 3712 10118 3884 10124
rect 3884 10066 3936 10072
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 3344 9518 3372 9998
rect 3988 9518 4016 10202
rect 4193 9820 4501 9829
rect 4193 9818 4199 9820
rect 4255 9818 4279 9820
rect 4335 9818 4359 9820
rect 4415 9818 4439 9820
rect 4495 9818 4501 9820
rect 4255 9766 4257 9818
rect 4437 9766 4439 9818
rect 4193 9764 4199 9766
rect 4255 9764 4279 9766
rect 4335 9764 4359 9766
rect 4415 9764 4439 9766
rect 4495 9764 4501 9766
rect 4193 9755 4501 9764
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4264 9178 4292 9318
rect 4356 9178 4384 9454
rect 4908 9178 4936 10542
rect 4986 10024 5042 10033
rect 5042 9982 5120 10010
rect 4986 9959 5042 9968
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3344 8362 3372 8774
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3252 6118 3280 8230
rect 3330 7984 3386 7993
rect 3330 7919 3332 7928
rect 3384 7919 3386 7928
rect 3332 7890 3384 7896
rect 3330 7848 3386 7857
rect 3330 7783 3386 7792
rect 3344 7750 3372 7783
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3344 7206 3372 7686
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3240 5092 3292 5098
rect 3240 5034 3292 5040
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3252 4729 3280 5034
rect 3238 4720 3294 4729
rect 3238 4655 3294 4664
rect 3238 4584 3294 4593
rect 3238 4519 3294 4528
rect 3252 4486 3280 4519
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2686 4040 2742 4049
rect 2686 3975 2742 3984
rect 2700 3942 2728 3975
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2686 3768 2742 3777
rect 2792 3738 2820 3878
rect 2686 3703 2742 3712
rect 2780 3732 2832 3738
rect 2700 3194 2728 3703
rect 2780 3674 2832 3680
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2884 2106 2912 3538
rect 3252 3058 3280 4422
rect 3344 4078 3372 7142
rect 3436 6934 3464 8434
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3528 7342 3556 7890
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3424 6928 3476 6934
rect 3424 6870 3476 6876
rect 3528 6798 3556 7278
rect 3516 6792 3568 6798
rect 3436 6752 3516 6780
rect 3436 6254 3464 6752
rect 3516 6734 3568 6740
rect 3424 6248 3476 6254
rect 3476 6208 3556 6236
rect 3424 6190 3476 6196
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 5817 3464 6054
rect 3422 5808 3478 5817
rect 3422 5743 3478 5752
rect 3528 5302 3556 6208
rect 3620 5778 3648 8978
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3712 7188 3740 7822
rect 4080 7750 4108 8910
rect 4193 8732 4501 8741
rect 4193 8730 4199 8732
rect 4255 8730 4279 8732
rect 4335 8730 4359 8732
rect 4415 8730 4439 8732
rect 4495 8730 4501 8732
rect 4255 8678 4257 8730
rect 4437 8678 4439 8730
rect 4193 8676 4199 8678
rect 4255 8676 4279 8678
rect 4335 8676 4359 8678
rect 4415 8676 4439 8678
rect 4495 8676 4501 8678
rect 4193 8667 4501 8676
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4172 7750 4200 7822
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 4193 7644 4501 7653
rect 4193 7642 4199 7644
rect 4255 7642 4279 7644
rect 4335 7642 4359 7644
rect 4415 7642 4439 7644
rect 4495 7642 4501 7644
rect 4255 7590 4257 7642
rect 4437 7590 4439 7642
rect 4193 7588 4199 7590
rect 4255 7588 4279 7590
rect 4335 7588 4359 7590
rect 4415 7588 4439 7590
rect 4495 7588 4501 7590
rect 4193 7579 4501 7588
rect 3976 7200 4028 7206
rect 3712 7160 3976 7188
rect 3712 6866 3740 7160
rect 3976 7142 4028 7148
rect 4066 6896 4122 6905
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3988 6854 4066 6882
rect 3712 6118 3740 6802
rect 3988 6322 4016 6854
rect 4066 6831 4122 6840
rect 4193 6556 4501 6565
rect 4193 6554 4199 6556
rect 4255 6554 4279 6556
rect 4335 6554 4359 6556
rect 4415 6554 4439 6556
rect 4495 6554 4501 6556
rect 4255 6502 4257 6554
rect 4437 6502 4439 6554
rect 4193 6500 4199 6502
rect 4255 6500 4279 6502
rect 4335 6500 4359 6502
rect 4415 6500 4439 6502
rect 4495 6500 4501 6502
rect 4193 6491 4501 6500
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 4804 6248 4856 6254
rect 4986 6216 5042 6225
rect 4804 6190 4856 6196
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 3700 5704 3752 5710
rect 4068 5704 4120 5710
rect 3752 5652 3832 5658
rect 3700 5646 3832 5652
rect 4068 5646 4120 5652
rect 3712 5630 3832 5646
rect 3516 5296 3568 5302
rect 3516 5238 3568 5244
rect 3804 4622 3832 5630
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3804 4078 3832 4558
rect 3896 4128 3924 5102
rect 3988 4622 4016 5510
rect 4080 5370 4108 5646
rect 4193 5468 4501 5477
rect 4193 5466 4199 5468
rect 4255 5466 4279 5468
rect 4335 5466 4359 5468
rect 4415 5466 4439 5468
rect 4495 5466 4501 5468
rect 4255 5414 4257 5466
rect 4437 5414 4439 5466
rect 4193 5412 4199 5414
rect 4255 5412 4279 5414
rect 4335 5412 4359 5414
rect 4415 5412 4439 5414
rect 4495 5412 4501 5414
rect 4193 5403 4501 5412
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4172 5250 4200 5306
rect 4080 5234 4200 5250
rect 4068 5228 4200 5234
rect 4120 5222 4200 5228
rect 4068 5170 4120 5176
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4172 4690 4200 5102
rect 4540 4826 4568 5714
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4160 4684 4212 4690
rect 4080 4644 4160 4672
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3896 4100 4016 4128
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 3792 4072 3844 4078
rect 3844 4049 3924 4060
rect 3844 4040 3938 4049
rect 3844 4032 3882 4040
rect 3792 4014 3844 4020
rect 3514 3904 3570 3913
rect 3436 3862 3514 3890
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3160 2650 3188 2994
rect 3330 2680 3386 2689
rect 3148 2644 3200 2650
rect 3330 2615 3386 2624
rect 3148 2586 3200 2592
rect 3344 2514 3372 2615
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 3436 2038 3464 3862
rect 3514 3839 3570 3848
rect 3514 3768 3570 3777
rect 3514 3703 3570 3712
rect 3528 3602 3556 3703
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3424 2032 3476 2038
rect 3424 1974 3476 1980
rect 2596 1964 2648 1970
rect 2596 1906 2648 1912
rect 2136 1896 2188 1902
rect 2136 1838 2188 1844
rect 3332 1896 3384 1902
rect 3332 1838 3384 1844
rect 1964 1426 2084 1442
rect 1122 1391 1178 1400
rect 1216 1420 1268 1426
rect 1216 1362 1268 1368
rect 1308 1420 1360 1426
rect 1308 1362 1360 1368
rect 1952 1420 2084 1426
rect 2004 1414 2084 1420
rect 1952 1362 2004 1368
rect 3344 1358 3372 1838
rect 2044 1352 2096 1358
rect 2044 1294 2096 1300
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 1492 876 1544 882
rect 1492 818 1544 824
rect 1504 474 1532 818
rect 2056 474 2084 1294
rect 3344 1018 3372 1294
rect 3528 1018 3556 2858
rect 3332 1012 3384 1018
rect 3332 954 3384 960
rect 3516 1012 3568 1018
rect 3516 954 3568 960
rect 3620 814 3648 4014
rect 3882 3975 3938 3984
rect 3988 3777 4016 4100
rect 3974 3768 4030 3777
rect 3792 3732 3844 3738
rect 3844 3692 3924 3720
rect 3974 3703 4030 3712
rect 3792 3674 3844 3680
rect 3896 3652 3924 3692
rect 4080 3652 4108 4644
rect 4160 4626 4212 4632
rect 4193 4380 4501 4389
rect 4193 4378 4199 4380
rect 4255 4378 4279 4380
rect 4335 4378 4359 4380
rect 4415 4378 4439 4380
rect 4495 4378 4501 4380
rect 4255 4326 4257 4378
rect 4437 4326 4439 4378
rect 4193 4324 4199 4326
rect 4255 4324 4279 4326
rect 4335 4324 4359 4326
rect 4415 4324 4439 4326
rect 4495 4324 4501 4326
rect 4193 4315 4501 4324
rect 4344 4072 4396 4078
rect 4540 4060 4568 4762
rect 4396 4032 4568 4060
rect 4344 4014 4396 4020
rect 4356 3738 4384 4014
rect 4724 3913 4752 5646
rect 4816 4146 4844 6190
rect 4908 6174 4986 6202
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4710 3904 4766 3913
rect 4908 3890 4936 6174
rect 4986 6151 5042 6160
rect 5092 5930 5120 9982
rect 5276 9722 5304 17614
rect 5368 17202 5396 19178
rect 5460 19122 5488 19343
rect 5540 19314 5592 19320
rect 5644 19224 5672 21422
rect 6656 21418 6684 21898
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 6932 21690 6960 21830
rect 6920 21684 6972 21690
rect 6920 21626 6972 21632
rect 8220 21622 8248 22238
rect 10048 22228 10100 22234
rect 10048 22170 10100 22176
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 11060 22228 11112 22234
rect 12256 22238 12308 22244
rect 24124 22296 24176 22302
rect 24124 22238 24176 22244
rect 11150 22199 11206 22208
rect 11060 22170 11112 22176
rect 9404 22160 9456 22166
rect 10060 22137 10088 22170
rect 10980 22137 11008 22170
rect 9404 22102 9456 22108
rect 10046 22128 10102 22137
rect 8574 21856 8630 21865
rect 8312 21814 8574 21842
rect 8208 21616 8260 21622
rect 8208 21558 8260 21564
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 6644 21412 6696 21418
rect 6644 21354 6696 21360
rect 6092 21140 6144 21146
rect 6092 21082 6144 21088
rect 6644 21140 6696 21146
rect 6644 21082 6696 21088
rect 5908 21072 5960 21078
rect 5908 21014 5960 21020
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5828 19961 5856 20878
rect 5814 19952 5870 19961
rect 5814 19887 5870 19896
rect 5828 19854 5856 19887
rect 5816 19848 5868 19854
rect 5816 19790 5868 19796
rect 5920 19394 5948 21014
rect 5998 20632 6054 20641
rect 5998 20567 6054 20576
rect 6012 20534 6040 20567
rect 6000 20528 6052 20534
rect 6000 20470 6052 20476
rect 6104 19836 6132 21082
rect 6552 20936 6604 20942
rect 6552 20878 6604 20884
rect 6460 20800 6512 20806
rect 6564 20777 6592 20878
rect 6460 20742 6512 20748
rect 6550 20768 6606 20777
rect 6472 20466 6500 20742
rect 6550 20703 6606 20712
rect 6656 20602 6684 21082
rect 6932 20602 6960 21490
rect 7288 21480 7340 21486
rect 7288 21422 7340 21428
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 6184 19848 6236 19854
rect 6104 19808 6184 19836
rect 6184 19790 6236 19796
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6196 19514 6224 19790
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 5920 19366 6132 19394
rect 5644 19196 5856 19224
rect 5460 19094 5672 19122
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5460 17241 5488 18770
rect 5552 18465 5580 18906
rect 5538 18456 5594 18465
rect 5644 18426 5672 19094
rect 5828 18850 5856 19196
rect 5908 19168 5960 19174
rect 6000 19168 6052 19174
rect 5908 19110 5960 19116
rect 5998 19136 6000 19145
rect 6052 19136 6054 19145
rect 5920 18970 5948 19110
rect 5998 19071 6054 19080
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 5736 18822 5856 18850
rect 5908 18828 5960 18834
rect 5538 18391 5594 18400
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5538 18320 5594 18329
rect 5538 18255 5540 18264
rect 5592 18255 5594 18264
rect 5632 18284 5684 18290
rect 5540 18226 5592 18232
rect 5632 18226 5684 18232
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5446 17232 5502 17241
rect 5356 17196 5408 17202
rect 5446 17167 5502 17176
rect 5356 17138 5408 17144
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5368 11354 5396 16594
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5460 13841 5488 15438
rect 5552 14618 5580 17614
rect 5644 16726 5672 18226
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5736 16425 5764 18822
rect 5908 18770 5960 18776
rect 5814 18728 5870 18737
rect 5920 18714 5948 18770
rect 6104 18737 6132 19366
rect 6196 18970 6224 19450
rect 6564 19417 6592 19790
rect 6734 19544 6790 19553
rect 6734 19479 6790 19488
rect 6550 19408 6606 19417
rect 6460 19372 6512 19378
rect 6550 19343 6606 19352
rect 6460 19314 6512 19320
rect 6276 19304 6328 19310
rect 6276 19246 6328 19252
rect 6184 18964 6236 18970
rect 6184 18906 6236 18912
rect 6184 18760 6236 18766
rect 5870 18686 5948 18714
rect 6090 18728 6146 18737
rect 5814 18663 5870 18672
rect 6184 18702 6236 18708
rect 6090 18663 6146 18672
rect 5828 17746 5856 18663
rect 5908 18352 5960 18358
rect 6104 18306 6132 18663
rect 5908 18294 5960 18300
rect 5920 17785 5948 18294
rect 6012 18278 6132 18306
rect 6012 18222 6040 18278
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 5998 18048 6054 18057
rect 5998 17983 6054 17992
rect 5906 17776 5962 17785
rect 5816 17740 5868 17746
rect 5906 17711 5962 17720
rect 5816 17682 5868 17688
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5920 17134 5948 17478
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 5722 16416 5778 16425
rect 5722 16351 5778 16360
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 5632 14272 5684 14278
rect 5736 14260 5764 16351
rect 5828 14464 5856 16934
rect 5920 16726 5948 17070
rect 5908 16720 5960 16726
rect 5908 16662 5960 16668
rect 5908 14884 5960 14890
rect 5908 14826 5960 14832
rect 5920 14618 5948 14826
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 5908 14476 5960 14482
rect 5828 14436 5908 14464
rect 5908 14418 5960 14424
rect 5684 14232 5764 14260
rect 5816 14272 5868 14278
rect 5632 14214 5684 14220
rect 5816 14214 5868 14220
rect 5828 14074 5856 14214
rect 5920 14113 5948 14418
rect 5906 14104 5962 14113
rect 5816 14068 5868 14074
rect 5906 14039 5962 14048
rect 5816 14010 5868 14016
rect 5446 13832 5502 13841
rect 5446 13767 5502 13776
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5448 13184 5500 13190
rect 5552 13138 5580 13670
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5500 13132 5580 13138
rect 5448 13126 5580 13132
rect 5460 13110 5580 13126
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5552 11218 5580 13110
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5644 12442 5672 12786
rect 5722 12472 5778 12481
rect 5632 12436 5684 12442
rect 5828 12442 5856 13262
rect 5722 12407 5778 12416
rect 5816 12436 5868 12442
rect 5632 12378 5684 12384
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5644 11150 5672 11630
rect 5736 11150 5764 12407
rect 5816 12378 5868 12384
rect 5920 12306 5948 14039
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5460 10198 5488 10610
rect 5644 10606 5672 11086
rect 5828 10810 5856 11698
rect 6012 11354 6040 17983
rect 6104 17678 6132 18158
rect 6196 18086 6224 18702
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 6104 17134 6132 17614
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 6092 16040 6144 16046
rect 6092 15982 6144 15988
rect 6104 15502 6132 15982
rect 6092 15496 6144 15502
rect 6288 15484 6316 19246
rect 6472 18834 6500 19314
rect 6642 18864 6698 18873
rect 6460 18828 6512 18834
rect 6642 18799 6698 18808
rect 6460 18770 6512 18776
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6380 17882 6408 18702
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 6656 17202 6684 18799
rect 6748 18426 6776 19479
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6736 18080 6788 18086
rect 6840 18057 6868 20334
rect 6918 19952 6974 19961
rect 6918 19887 6920 19896
rect 6972 19887 6974 19896
rect 6920 19858 6972 19864
rect 7116 19514 7144 20334
rect 7300 19825 7328 21422
rect 8312 21350 8340 21814
rect 8574 21791 8630 21800
rect 9416 21690 9444 22102
rect 9956 22092 10008 22098
rect 10966 22128 11022 22137
rect 10046 22063 10102 22072
rect 10416 22092 10468 22098
rect 9956 22034 10008 22040
rect 10966 22063 11022 22072
rect 10416 22034 10468 22040
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 8576 21616 8628 21622
rect 8628 21576 8892 21604
rect 8576 21558 8628 21564
rect 8864 21486 8892 21576
rect 8576 21480 8628 21486
rect 8576 21422 8628 21428
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8484 21412 8536 21418
rect 8484 21354 8536 21360
rect 8300 21344 8352 21350
rect 8496 21321 8524 21354
rect 8300 21286 8352 21292
rect 8482 21312 8538 21321
rect 7988 21244 8296 21253
rect 8482 21247 8538 21256
rect 7988 21242 7994 21244
rect 8050 21242 8074 21244
rect 8130 21242 8154 21244
rect 8210 21242 8234 21244
rect 8290 21242 8296 21244
rect 8050 21190 8052 21242
rect 8232 21190 8234 21242
rect 7988 21188 7994 21190
rect 8050 21188 8074 21190
rect 8130 21188 8154 21190
rect 8210 21188 8234 21190
rect 8290 21188 8296 21190
rect 7988 21179 8296 21188
rect 7840 21072 7892 21078
rect 7840 21014 7892 21020
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7668 19854 7696 20742
rect 7760 20534 7788 20946
rect 7748 20528 7800 20534
rect 7748 20470 7800 20476
rect 7656 19848 7708 19854
rect 7286 19816 7342 19825
rect 7656 19790 7708 19796
rect 7286 19751 7342 19760
rect 7760 19718 7788 20470
rect 7852 20058 7880 21014
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8404 20233 8432 20334
rect 8390 20224 8446 20233
rect 7988 20156 8296 20165
rect 8390 20159 8446 20168
rect 7988 20154 7994 20156
rect 8050 20154 8074 20156
rect 8130 20154 8154 20156
rect 8210 20154 8234 20156
rect 8290 20154 8296 20156
rect 8050 20102 8052 20154
rect 8232 20102 8234 20154
rect 7988 20100 7994 20102
rect 8050 20100 8074 20102
rect 8130 20100 8154 20102
rect 8210 20100 8234 20102
rect 8290 20100 8296 20102
rect 7988 20091 8296 20100
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 8404 19990 8432 20159
rect 8392 19984 8444 19990
rect 8392 19926 8444 19932
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 8220 19514 8248 19858
rect 8392 19848 8444 19854
rect 8588 19836 8616 21422
rect 9312 21412 9364 21418
rect 9312 21354 9364 21360
rect 8668 21344 8720 21350
rect 9324 21321 9352 21354
rect 8668 21286 8720 21292
rect 9310 21312 9366 21321
rect 8680 21010 8708 21286
rect 9310 21247 9366 21256
rect 8758 21040 8814 21049
rect 8668 21004 8720 21010
rect 8758 20975 8814 20984
rect 8668 20946 8720 20952
rect 8772 20942 8800 20975
rect 8760 20936 8812 20942
rect 8760 20878 8812 20884
rect 8852 20936 8904 20942
rect 8852 20878 8904 20884
rect 8864 20641 8892 20878
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8850 20632 8906 20641
rect 8850 20567 8906 20576
rect 8668 20256 8720 20262
rect 8668 20198 8720 20204
rect 8444 19808 8616 19836
rect 8392 19790 8444 19796
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 8208 19508 8260 19514
rect 8208 19450 8260 19456
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6932 18601 6960 19314
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 7484 18970 7512 19110
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7472 18760 7524 18766
rect 7472 18702 7524 18708
rect 6918 18592 6974 18601
rect 6918 18527 6974 18536
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6932 18329 6960 18362
rect 6918 18320 6974 18329
rect 6918 18255 6974 18264
rect 7378 18320 7434 18329
rect 7378 18255 7434 18264
rect 6736 18022 6788 18028
rect 6826 18048 6882 18057
rect 6748 17882 6776 18022
rect 6826 17983 6882 17992
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6748 16998 6776 17818
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 7024 16794 7052 17614
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6092 15438 6144 15444
rect 6196 15456 6316 15484
rect 6104 15201 6132 15438
rect 6090 15192 6146 15201
rect 6090 15127 6146 15136
rect 6104 14958 6132 15127
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 6104 13938 6132 14894
rect 6196 14249 6224 15456
rect 6276 15360 6328 15366
rect 6276 15302 6328 15308
rect 6288 15026 6316 15302
rect 6380 15162 6408 16526
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6472 15570 6500 15982
rect 6656 15609 6684 16050
rect 6642 15600 6698 15609
rect 6460 15564 6512 15570
rect 6642 15535 6698 15544
rect 6460 15506 6512 15512
rect 6472 15162 6500 15506
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 6642 15328 6698 15337
rect 6642 15263 6698 15272
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6472 14822 6500 15098
rect 6550 15056 6606 15065
rect 6550 14991 6552 15000
rect 6604 14991 6606 15000
rect 6552 14962 6604 14968
rect 6460 14816 6512 14822
rect 6274 14784 6330 14793
rect 6460 14758 6512 14764
rect 6274 14719 6330 14728
rect 6288 14482 6316 14719
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6182 14240 6238 14249
rect 6182 14175 6238 14184
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 6092 13796 6144 13802
rect 6092 13738 6144 13744
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6104 11150 6132 13738
rect 6288 13462 6316 14418
rect 6472 13870 6500 14758
rect 6550 14512 6606 14521
rect 6550 14447 6552 14456
rect 6604 14447 6606 14456
rect 6552 14418 6604 14424
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6276 13456 6328 13462
rect 6276 13398 6328 13404
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6196 12782 6224 13262
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 5632 10600 5684 10606
rect 5632 10542 5684 10548
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5264 9716 5316 9722
rect 5644 9674 5672 10542
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5264 9658 5316 9664
rect 5552 9646 5672 9674
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 5184 6866 5212 9114
rect 5276 7342 5304 9318
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5368 8838 5396 8978
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5354 8664 5410 8673
rect 5354 8599 5410 8608
rect 5368 8430 5396 8599
rect 5460 8430 5488 9386
rect 5552 8430 5580 9646
rect 5630 8936 5686 8945
rect 5630 8871 5686 8880
rect 5644 8838 5672 8871
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5354 6488 5410 6497
rect 5276 6446 5354 6474
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 4710 3839 4766 3848
rect 4816 3862 4936 3890
rect 5000 5902 5120 5930
rect 5184 5914 5212 6054
rect 5172 5908 5224 5914
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 3698 3632 3754 3641
rect 3896 3624 4108 3652
rect 3698 3567 3754 3576
rect 3712 3398 3740 3567
rect 3882 3496 3938 3505
rect 3882 3431 3938 3440
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3804 3194 3832 3334
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3896 3058 3924 3431
rect 4193 3292 4501 3301
rect 4193 3290 4199 3292
rect 4255 3290 4279 3292
rect 4335 3290 4359 3292
rect 4415 3290 4439 3292
rect 4495 3290 4501 3292
rect 4255 3238 4257 3290
rect 4437 3238 4439 3290
rect 4193 3236 4199 3238
rect 4255 3236 4279 3238
rect 4335 3236 4359 3238
rect 4415 3236 4439 3238
rect 4495 3236 4501 3238
rect 4193 3227 4501 3236
rect 4526 3088 4582 3097
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 4436 3052 4488 3058
rect 4526 3023 4528 3032
rect 4436 2994 4488 3000
rect 4580 3023 4582 3032
rect 4528 2994 4580 3000
rect 3698 2816 3754 2825
rect 3698 2751 3754 2760
rect 4448 2774 4476 2994
rect 3712 1970 3740 2751
rect 4448 2746 4660 2774
rect 4526 2544 4582 2553
rect 4526 2479 4528 2488
rect 4580 2479 4582 2488
rect 4528 2450 4580 2456
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 3988 2106 4016 2382
rect 4193 2204 4501 2213
rect 4193 2202 4199 2204
rect 4255 2202 4279 2204
rect 4335 2202 4359 2204
rect 4415 2202 4439 2204
rect 4495 2202 4501 2204
rect 4255 2150 4257 2202
rect 4437 2150 4439 2202
rect 4193 2148 4199 2150
rect 4255 2148 4279 2150
rect 4335 2148 4359 2150
rect 4415 2148 4439 2150
rect 4495 2148 4501 2150
rect 4193 2139 4501 2148
rect 4632 2106 4660 2746
rect 4712 2644 4764 2650
rect 4816 2632 4844 3862
rect 5000 3754 5028 5902
rect 5172 5850 5224 5856
rect 5170 5400 5226 5409
rect 5170 5335 5226 5344
rect 4908 3726 5028 3754
rect 5080 3732 5132 3738
rect 4908 3516 4936 3726
rect 5080 3674 5132 3680
rect 4988 3664 5040 3670
rect 4986 3632 4988 3641
rect 5040 3632 5042 3641
rect 4986 3567 5042 3576
rect 4908 3488 5028 3516
rect 4764 2604 4844 2632
rect 4712 2586 4764 2592
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 4620 2100 4672 2106
rect 4620 2042 4672 2048
rect 4250 2000 4306 2009
rect 3700 1964 3752 1970
rect 4068 1964 4120 1970
rect 3700 1906 3752 1912
rect 3988 1924 4068 1952
rect 3792 1896 3844 1902
rect 3792 1838 3844 1844
rect 3804 1562 3832 1838
rect 3792 1556 3844 1562
rect 3792 1498 3844 1504
rect 3608 808 3660 814
rect 3608 750 3660 756
rect 3804 678 3832 1498
rect 3884 1352 3936 1358
rect 3884 1294 3936 1300
rect 3792 672 3844 678
rect 3792 614 3844 620
rect 1492 468 1544 474
rect 1492 410 1544 416
rect 2044 468 2096 474
rect 2044 410 2096 416
rect 3896 66 3924 1294
rect 3988 338 4016 1924
rect 4250 1935 4252 1944
rect 4068 1906 4120 1912
rect 4304 1935 4306 1944
rect 4252 1906 4304 1912
rect 4724 1766 4752 2450
rect 4712 1760 4764 1766
rect 4618 1728 4674 1737
rect 4712 1702 4764 1708
rect 4618 1663 4674 1672
rect 4632 1562 4660 1663
rect 4620 1556 4672 1562
rect 4620 1498 4672 1504
rect 4068 1352 4120 1358
rect 4066 1320 4068 1329
rect 4120 1320 4122 1329
rect 4066 1255 4122 1264
rect 4193 1116 4501 1125
rect 4193 1114 4199 1116
rect 4255 1114 4279 1116
rect 4335 1114 4359 1116
rect 4415 1114 4439 1116
rect 4495 1114 4501 1116
rect 4255 1062 4257 1114
rect 4437 1062 4439 1114
rect 4193 1060 4199 1062
rect 4255 1060 4279 1062
rect 4335 1060 4359 1062
rect 4415 1060 4439 1062
rect 4495 1060 4501 1062
rect 4193 1051 4501 1060
rect 4816 1018 4844 2604
rect 5000 1018 5028 3488
rect 5092 1494 5120 3674
rect 5184 2553 5212 5335
rect 5276 4010 5304 6446
rect 5460 6458 5488 6802
rect 5354 6423 5410 6432
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5540 6248 5592 6254
rect 5644 6236 5672 8774
rect 5736 7546 5764 9998
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5828 8294 5856 8774
rect 5920 8430 5948 10542
rect 6104 10470 6132 10746
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 6104 9058 6132 10134
rect 6196 9178 6224 11630
rect 6288 11354 6316 13398
rect 6564 13326 6592 14282
rect 6656 13938 6684 15263
rect 7024 15026 7052 15438
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6748 14657 6776 14758
rect 6734 14648 6790 14657
rect 6932 14618 6960 14894
rect 7300 14793 7328 14894
rect 7286 14784 7342 14793
rect 7286 14719 7342 14728
rect 7392 14618 7420 18255
rect 7484 17921 7512 18702
rect 7576 18329 7604 19450
rect 8206 19408 8262 19417
rect 8206 19343 8208 19352
rect 8260 19343 8262 19352
rect 8208 19314 8260 19320
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7562 18320 7618 18329
rect 7562 18255 7618 18264
rect 7668 18086 7696 19246
rect 7760 18766 7788 19246
rect 7840 19236 7892 19242
rect 7840 19178 7892 19184
rect 7748 18760 7800 18766
rect 7748 18702 7800 18708
rect 7746 18592 7802 18601
rect 7746 18527 7802 18536
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7470 17912 7526 17921
rect 7470 17847 7526 17856
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 6734 14583 6790 14592
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6748 13938 6776 14010
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6840 13462 6868 14350
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7024 13841 7052 13874
rect 7010 13832 7066 13841
rect 7010 13767 7066 13776
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 6552 13320 6604 13326
rect 6748 13308 6776 13398
rect 6920 13320 6972 13326
rect 6748 13297 6868 13308
rect 6552 13262 6604 13268
rect 6734 13288 6868 13297
rect 6790 13280 6868 13288
rect 6734 13223 6790 13232
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6644 13184 6696 13190
rect 6696 13144 6776 13172
rect 6644 13126 6696 13132
rect 6380 12481 6408 13126
rect 6748 12850 6776 13144
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6644 12776 6696 12782
rect 6840 12730 6868 13280
rect 6920 13262 6972 13268
rect 6644 12718 6696 12724
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 6366 12472 6422 12481
rect 6366 12407 6422 12416
rect 6472 12170 6500 12582
rect 6552 12368 6604 12374
rect 6656 12322 6684 12718
rect 6748 12702 6868 12730
rect 6748 12646 6776 12702
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6604 12316 6684 12322
rect 6552 12310 6684 12316
rect 6564 12294 6684 12310
rect 6460 12164 6512 12170
rect 6512 12124 6592 12152
rect 6460 12106 6512 12112
rect 6564 11558 6592 12124
rect 6552 11552 6604 11558
rect 6552 11494 6604 11500
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6564 11286 6592 11494
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6564 10606 6592 11222
rect 6656 11218 6684 12294
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6656 10810 6684 11154
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6276 10600 6328 10606
rect 6552 10600 6604 10606
rect 6276 10542 6328 10548
rect 6472 10548 6552 10554
rect 6472 10542 6604 10548
rect 6288 9722 6316 10542
rect 6472 10526 6592 10542
rect 6472 10266 6500 10526
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 6460 10056 6512 10062
rect 6380 10016 6460 10044
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6380 9586 6408 10016
rect 6460 9998 6512 10004
rect 6564 9674 6592 10406
rect 6472 9646 6592 9674
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6104 9030 6316 9058
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5724 7268 5776 7274
rect 5724 7210 5776 7216
rect 5736 6866 5764 7210
rect 5828 7002 5856 7822
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5592 6208 5672 6236
rect 5540 6190 5592 6196
rect 5552 6089 5580 6190
rect 5632 6112 5684 6118
rect 5538 6080 5594 6089
rect 5632 6054 5684 6060
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5538 6015 5594 6024
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5368 3602 5396 5850
rect 5552 5778 5580 6015
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5460 5166 5488 5578
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5448 5160 5500 5166
rect 5552 5137 5580 5510
rect 5448 5102 5500 5108
rect 5538 5128 5594 5137
rect 5538 5063 5594 5072
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 4146 5580 4422
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5644 4078 5672 6054
rect 5828 5778 5856 6054
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5736 4282 5764 5170
rect 5920 5166 5948 7686
rect 6012 6662 6040 8774
rect 6104 8498 6132 8910
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6196 8294 6224 8366
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6182 7440 6238 7449
rect 6182 7375 6238 7384
rect 6196 7342 6224 7375
rect 6184 7336 6236 7342
rect 6288 7313 6316 9030
rect 6380 8956 6408 9522
rect 6472 9518 6500 9646
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6656 9042 6684 9658
rect 6644 9036 6696 9042
rect 6748 9024 6776 12582
rect 6828 12300 6880 12306
rect 6932 12288 6960 13262
rect 7116 12594 7144 14350
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7208 12986 7236 13262
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7300 12696 7328 13466
rect 7392 12764 7420 14350
rect 7668 14074 7696 15982
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7470 13560 7526 13569
rect 7526 13518 7604 13546
rect 7470 13495 7526 13504
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7484 12986 7512 13262
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7392 12736 7512 12764
rect 6880 12260 6960 12288
rect 7024 12566 7144 12594
rect 7208 12668 7328 12696
rect 7208 12594 7236 12668
rect 7208 12566 7239 12594
rect 6828 12242 6880 12248
rect 7024 11898 7052 12566
rect 7102 12472 7158 12481
rect 7211 12434 7239 12566
rect 7102 12407 7158 12416
rect 7116 12238 7144 12407
rect 7208 12406 7239 12434
rect 7208 12322 7236 12406
rect 7208 12294 7328 12322
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7208 12102 7236 12174
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7194 11656 7250 11665
rect 7194 11591 7196 11600
rect 7248 11591 7250 11600
rect 7196 11562 7248 11568
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 9586 6960 11494
rect 7300 11218 7328 12294
rect 7484 11898 7512 12736
rect 7576 12102 7604 13518
rect 7760 12696 7788 18527
rect 7852 17882 7880 19178
rect 7988 19068 8296 19077
rect 7988 19066 7994 19068
rect 8050 19066 8074 19068
rect 8130 19066 8154 19068
rect 8210 19066 8234 19068
rect 8290 19066 8296 19068
rect 8050 19014 8052 19066
rect 8232 19014 8234 19066
rect 7988 19012 7994 19014
rect 8050 19012 8074 19014
rect 8130 19012 8154 19014
rect 8210 19012 8234 19014
rect 8290 19012 8296 19014
rect 7988 19003 8296 19012
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 8208 18624 8260 18630
rect 8206 18592 8208 18601
rect 8260 18592 8262 18601
rect 8206 18527 8262 18536
rect 8312 18290 8340 18634
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 7988 17980 8296 17989
rect 7988 17978 7994 17980
rect 8050 17978 8074 17980
rect 8130 17978 8154 17980
rect 8210 17978 8234 17980
rect 8290 17978 8296 17980
rect 8050 17926 8052 17978
rect 8232 17926 8234 17978
rect 7988 17924 7994 17926
rect 8050 17924 8074 17926
rect 8130 17924 8154 17926
rect 8210 17924 8234 17926
rect 8290 17924 8296 17926
rect 7988 17915 8296 17924
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7988 16892 8296 16901
rect 7988 16890 7994 16892
rect 8050 16890 8074 16892
rect 8130 16890 8154 16892
rect 8210 16890 8234 16892
rect 8290 16890 8296 16892
rect 8050 16838 8052 16890
rect 8232 16838 8234 16890
rect 7988 16836 7994 16838
rect 8050 16836 8074 16838
rect 8130 16836 8154 16838
rect 8210 16836 8234 16838
rect 8290 16836 8296 16838
rect 7988 16827 8296 16836
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 7840 15904 7892 15910
rect 8128 15892 8156 16594
rect 8404 16561 8432 19790
rect 8484 19712 8536 19718
rect 8482 19680 8484 19689
rect 8536 19680 8538 19689
rect 8482 19615 8538 19624
rect 8496 18630 8524 19615
rect 8680 19514 8708 20198
rect 8956 19854 8984 20742
rect 9586 20496 9642 20505
rect 9586 20431 9642 20440
rect 9496 20392 9548 20398
rect 9034 20360 9090 20369
rect 9090 20318 9168 20346
rect 9496 20334 9548 20340
rect 9034 20295 9090 20304
rect 9036 19916 9088 19922
rect 9036 19858 9088 19864
rect 8852 19848 8904 19854
rect 8852 19790 8904 19796
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 8864 19514 8892 19790
rect 9048 19553 9076 19858
rect 9034 19544 9090 19553
rect 8668 19508 8720 19514
rect 8668 19450 8720 19456
rect 8852 19508 8904 19514
rect 9034 19479 9090 19488
rect 8852 19450 8904 19456
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8588 18902 8616 19314
rect 8680 18902 8708 19450
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8576 18896 8628 18902
rect 8576 18838 8628 18844
rect 8668 18896 8720 18902
rect 8668 18838 8720 18844
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8576 18624 8628 18630
rect 8772 18578 8800 19110
rect 8628 18572 8800 18578
rect 8576 18566 8800 18572
rect 8588 18550 8800 18566
rect 8484 18352 8536 18358
rect 8484 18294 8536 18300
rect 8496 17882 8524 18294
rect 8576 18148 8628 18154
rect 8576 18090 8628 18096
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8588 17746 8616 18090
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8680 17678 8708 18550
rect 8864 18426 8892 19110
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 8864 18222 8892 18362
rect 8852 18216 8904 18222
rect 8852 18158 8904 18164
rect 8864 17864 8892 18158
rect 8864 17836 9076 17864
rect 8850 17776 8906 17785
rect 8772 17734 8850 17762
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8680 17134 8708 17614
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8496 16833 8524 16934
rect 8482 16824 8538 16833
rect 8482 16759 8538 16768
rect 8390 16552 8446 16561
rect 8208 16516 8260 16522
rect 8496 16522 8524 16759
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8390 16487 8446 16496
rect 8484 16516 8536 16522
rect 8208 16458 8260 16464
rect 8484 16458 8536 16464
rect 8220 16046 8248 16458
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8128 15864 8432 15892
rect 7840 15846 7892 15852
rect 7852 14006 7880 15846
rect 7988 15804 8296 15813
rect 7988 15802 7994 15804
rect 8050 15802 8074 15804
rect 8130 15802 8154 15804
rect 8210 15802 8234 15804
rect 8290 15802 8296 15804
rect 8050 15750 8052 15802
rect 8232 15750 8234 15802
rect 7988 15748 7994 15750
rect 8050 15748 8074 15750
rect 8130 15748 8154 15750
rect 8210 15748 8234 15750
rect 8290 15748 8296 15750
rect 7988 15739 8296 15748
rect 7988 14716 8296 14725
rect 7988 14714 7994 14716
rect 8050 14714 8074 14716
rect 8130 14714 8154 14716
rect 8210 14714 8234 14716
rect 8290 14714 8296 14716
rect 8050 14662 8052 14714
rect 8232 14662 8234 14714
rect 7988 14660 7994 14662
rect 8050 14660 8074 14662
rect 8130 14660 8154 14662
rect 8210 14660 8234 14662
rect 8290 14660 8296 14662
rect 7988 14651 8296 14660
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 7988 13628 8296 13637
rect 7988 13626 7994 13628
rect 8050 13626 8074 13628
rect 8130 13626 8154 13628
rect 8210 13626 8234 13628
rect 8290 13626 8296 13628
rect 8050 13574 8052 13626
rect 8232 13574 8234 13626
rect 7988 13572 7994 13574
rect 8050 13572 8074 13574
rect 8130 13572 8154 13574
rect 8210 13572 8234 13574
rect 8290 13572 8296 13574
rect 7988 13563 8296 13572
rect 8404 13530 8432 15864
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 7840 12708 7892 12714
rect 7760 12668 7840 12696
rect 7840 12650 7892 12656
rect 7654 12608 7710 12617
rect 7654 12543 7710 12552
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7668 11830 7696 12543
rect 7988 12540 8296 12549
rect 7988 12538 7994 12540
rect 8050 12538 8074 12540
rect 8130 12538 8154 12540
rect 8210 12538 8234 12540
rect 8290 12538 8296 12540
rect 8050 12486 8052 12538
rect 8232 12486 8234 12538
rect 7988 12484 7994 12486
rect 8050 12484 8074 12486
rect 8130 12484 8154 12486
rect 8210 12484 8234 12486
rect 8290 12484 8296 12486
rect 7988 12475 8296 12484
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7944 11898 7972 12378
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7656 11824 7708 11830
rect 7656 11766 7708 11772
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7852 11642 7880 11698
rect 7760 11614 7880 11642
rect 8496 11626 8524 16458
rect 8588 16250 8616 16526
rect 8576 16244 8628 16250
rect 8576 16186 8628 16192
rect 8588 15570 8616 16186
rect 8772 16114 8800 17734
rect 8850 17711 8906 17720
rect 9048 17678 9076 17836
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 8850 17096 8906 17105
rect 8850 17031 8906 17040
rect 8760 16108 8812 16114
rect 8680 16068 8760 16096
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8588 15201 8616 15506
rect 8574 15192 8630 15201
rect 8574 15127 8630 15136
rect 8588 14958 8616 15127
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8680 14113 8708 16068
rect 8760 16050 8812 16056
rect 8758 14648 8814 14657
rect 8758 14583 8814 14592
rect 8772 14482 8800 14583
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8666 14104 8722 14113
rect 8666 14039 8722 14048
rect 8680 13938 8708 14039
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8484 11620 8536 11626
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7760 10996 7788 11614
rect 8484 11562 8536 11568
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7576 10968 7788 10996
rect 7576 10470 7604 10968
rect 7656 10532 7708 10538
rect 7656 10474 7708 10480
rect 7748 10532 7800 10538
rect 7748 10474 7800 10480
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6920 9036 6972 9042
rect 6748 8996 6920 9024
rect 6644 8978 6696 8984
rect 6920 8978 6972 8984
rect 6460 8968 6512 8974
rect 6380 8928 6460 8956
rect 6932 8945 6960 8978
rect 6460 8910 6512 8916
rect 6918 8936 6974 8945
rect 6918 8871 6974 8880
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6472 8129 6500 8774
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6458 8120 6514 8129
rect 6458 8055 6514 8064
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6184 7278 6236 7284
rect 6274 7304 6330 7313
rect 6274 7239 6330 7248
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 6092 5840 6144 5846
rect 6090 5808 6092 5817
rect 6144 5808 6146 5817
rect 6196 5778 6224 6802
rect 6288 6100 6316 7239
rect 6380 7206 6408 7822
rect 6472 7206 6500 7958
rect 6550 7440 6606 7449
rect 6550 7375 6552 7384
rect 6604 7375 6606 7384
rect 6552 7346 6604 7352
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6380 6866 6408 7142
rect 6472 7002 6500 7142
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 6380 6458 6408 6802
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6472 6322 6500 6938
rect 6656 6458 6684 8570
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6748 7206 6776 7686
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6656 6202 6684 6258
rect 6472 6174 6684 6202
rect 6368 6112 6420 6118
rect 6288 6072 6368 6100
rect 6368 6054 6420 6060
rect 6090 5743 6146 5752
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6380 5250 6408 6054
rect 6472 5681 6500 6174
rect 6748 6118 6776 6734
rect 6840 6322 6868 8774
rect 6932 8673 6960 8774
rect 6918 8664 6974 8673
rect 7024 8634 7052 9998
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7116 9178 7144 9454
rect 7484 9382 7512 10202
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7484 9178 7512 9318
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7470 9072 7526 9081
rect 7288 9036 7340 9042
rect 7470 9007 7472 9016
rect 7288 8978 7340 8984
rect 7524 9007 7526 9016
rect 7472 8978 7524 8984
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 6918 8599 6974 8608
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7010 8392 7066 8401
rect 7010 8327 7066 8336
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 6905 6960 7686
rect 6918 6896 6974 6905
rect 6918 6831 6974 6840
rect 7024 6798 7052 8327
rect 7116 7954 7144 8774
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7208 6866 7236 8502
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 7104 6248 7156 6254
rect 7300 6236 7328 8978
rect 7484 6322 7512 8978
rect 7576 8634 7604 9998
rect 7668 9178 7696 10474
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7656 9036 7708 9042
rect 7760 9024 7788 10474
rect 7708 8996 7788 9024
rect 7656 8978 7708 8984
rect 7852 8820 7880 11494
rect 7988 11452 8296 11461
rect 7988 11450 7994 11452
rect 8050 11450 8074 11452
rect 8130 11450 8154 11452
rect 8210 11450 8234 11452
rect 8290 11450 8296 11452
rect 8050 11398 8052 11450
rect 8232 11398 8234 11450
rect 7988 11396 7994 11398
rect 8050 11396 8074 11398
rect 8130 11396 8154 11398
rect 8210 11396 8234 11398
rect 8290 11396 8296 11398
rect 7988 11387 8296 11396
rect 7988 10364 8296 10373
rect 7988 10362 7994 10364
rect 8050 10362 8074 10364
rect 8130 10362 8154 10364
rect 8210 10362 8234 10364
rect 8290 10362 8296 10364
rect 8050 10310 8052 10362
rect 8232 10310 8234 10362
rect 7988 10308 7994 10310
rect 8050 10308 8074 10310
rect 8130 10308 8154 10310
rect 8210 10308 8234 10310
rect 8290 10308 8296 10310
rect 7988 10299 8296 10308
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 7988 9276 8296 9285
rect 7988 9274 7994 9276
rect 8050 9274 8074 9276
rect 8130 9274 8154 9276
rect 8210 9274 8234 9276
rect 8290 9274 8296 9276
rect 8050 9222 8052 9274
rect 8232 9222 8234 9274
rect 7988 9220 7994 9222
rect 8050 9220 8074 9222
rect 8130 9220 8154 9222
rect 8210 9220 8234 9222
rect 8290 9220 8296 9222
rect 7988 9211 8296 9220
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8128 8974 8156 9114
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8220 8820 8248 8978
rect 7852 8792 8248 8820
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 8404 8430 8432 9590
rect 8496 9518 8524 11562
rect 8588 11286 8616 13466
rect 8772 12850 8800 13942
rect 8864 12986 8892 17031
rect 9048 16998 9076 17614
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8956 15910 8984 16526
rect 8944 15904 8996 15910
rect 8944 15846 8996 15852
rect 8956 15502 8984 15846
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8956 15026 8984 15438
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8956 14550 8984 14962
rect 8944 14544 8996 14550
rect 8944 14486 8996 14492
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 8942 14240 8998 14249
rect 8942 14175 8998 14184
rect 8956 13530 8984 14175
rect 8944 13524 8996 13530
rect 8944 13466 8996 13472
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 9048 12918 9076 14418
rect 9140 13530 9168 20318
rect 9508 20233 9536 20334
rect 9494 20224 9550 20233
rect 9494 20159 9550 20168
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9232 19281 9260 19790
rect 9218 19272 9274 19281
rect 9218 19207 9274 19216
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9218 18184 9274 18193
rect 9218 18119 9274 18128
rect 9232 17746 9260 18119
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 9218 17640 9274 17649
rect 9218 17575 9274 17584
rect 9232 16425 9260 17575
rect 9416 17218 9444 18702
rect 9508 18630 9536 20159
rect 9600 20058 9628 20431
rect 9588 20052 9640 20058
rect 9588 19994 9640 20000
rect 9968 19786 9996 22034
rect 10230 21992 10286 22001
rect 10230 21927 10286 21936
rect 10244 21894 10272 21927
rect 10232 21888 10284 21894
rect 10232 21830 10284 21836
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 10336 21622 10364 21830
rect 10324 21616 10376 21622
rect 10324 21558 10376 21564
rect 10428 21486 10456 22034
rect 10966 21584 11022 21593
rect 10966 21519 11022 21528
rect 10416 21480 10468 21486
rect 10416 21422 10468 21428
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 10784 21480 10836 21486
rect 10784 21422 10836 21428
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 10598 21040 10654 21049
rect 10508 21004 10560 21010
rect 10598 20975 10654 20984
rect 10508 20946 10560 20952
rect 10520 20602 10548 20946
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 9956 19780 10008 19786
rect 9956 19722 10008 19728
rect 10244 19514 10272 20334
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 10336 19514 10364 19654
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9496 18624 9548 18630
rect 9600 18601 9628 18702
rect 9496 18566 9548 18572
rect 9586 18592 9642 18601
rect 9508 18408 9536 18566
rect 9586 18527 9642 18536
rect 9678 18456 9734 18465
rect 9588 18420 9640 18426
rect 9508 18380 9588 18408
rect 9678 18391 9734 18400
rect 9588 18362 9640 18368
rect 9692 18290 9720 18391
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9876 17746 9904 18906
rect 10322 18864 10378 18873
rect 10322 18799 10378 18808
rect 10232 18692 10284 18698
rect 10232 18634 10284 18640
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9678 17504 9734 17513
rect 9324 17190 9444 17218
rect 9508 17202 9536 17478
rect 9734 17462 9904 17490
rect 9678 17439 9734 17448
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9496 17196 9548 17202
rect 9324 16794 9352 17190
rect 9496 17138 9548 17144
rect 9404 17128 9456 17134
rect 9784 17105 9812 17274
rect 9404 17070 9456 17076
rect 9770 17096 9826 17105
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9218 16416 9274 16425
rect 9218 16351 9274 16360
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9232 14074 9260 15982
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9324 14618 9352 15438
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9416 14074 9444 17070
rect 9770 17031 9826 17040
rect 9494 16824 9550 16833
rect 9588 16788 9640 16794
rect 9550 16768 9588 16776
rect 9494 16759 9588 16768
rect 9508 16748 9588 16759
rect 9588 16730 9640 16736
rect 9678 16688 9734 16697
rect 9734 16646 9812 16674
rect 9678 16623 9734 16632
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9508 16425 9536 16526
rect 9494 16416 9550 16425
rect 9494 16351 9550 16360
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9508 14482 9536 15098
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9692 14618 9720 14894
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9692 13954 9720 14418
rect 9508 13926 9720 13954
rect 9218 13832 9274 13841
rect 9274 13790 9352 13818
rect 9218 13767 9274 13776
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9324 13394 9352 13790
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9416 13394 9444 13670
rect 9220 13388 9272 13394
rect 9140 13348 9220 13376
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8668 12640 8720 12646
rect 9048 12617 9076 12854
rect 9034 12608 9090 12617
rect 8668 12582 8720 12588
rect 8680 12374 8708 12582
rect 8956 12566 9034 12594
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8680 11540 8708 12174
rect 8956 11762 8984 12566
rect 9034 12543 9090 12552
rect 9036 12300 9088 12306
rect 9036 12242 9088 12248
rect 9048 11898 9076 12242
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8760 11552 8812 11558
rect 8680 11512 8760 11540
rect 8760 11494 8812 11500
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8588 9081 8616 11018
rect 8772 10606 8800 11290
rect 8956 11218 8984 11698
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 9048 10826 9076 11834
rect 9140 11694 9168 13348
rect 9220 13330 9272 13336
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9416 13274 9444 13330
rect 9232 13246 9444 13274
rect 9232 12714 9260 13246
rect 9508 13190 9536 13926
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9496 13184 9548 13190
rect 9496 13126 9548 13132
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8956 10798 9076 10826
rect 8956 10742 8984 10798
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8956 10266 8984 10678
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 9048 10062 9076 10610
rect 9140 10606 9168 11494
rect 9232 11354 9260 12650
rect 9324 12306 9352 12854
rect 9416 12782 9444 13126
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9402 11792 9458 11801
rect 9402 11727 9458 11736
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 9324 10674 9352 11630
rect 9416 11354 9444 11727
rect 9508 11354 9536 13126
rect 9600 12850 9628 13670
rect 9784 13530 9812 16646
rect 9876 14362 9904 17462
rect 9968 14618 9996 18158
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10060 14482 10088 18022
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 9876 14334 9996 14362
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 13938 9904 14214
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9784 12850 9812 13126
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9600 12696 9628 12786
rect 9600 12668 9720 12696
rect 9692 12594 9720 12668
rect 9600 12566 9720 12594
rect 9600 11762 9628 12566
rect 9680 11892 9732 11898
rect 9784 11880 9812 12786
rect 9732 11852 9812 11880
rect 9680 11834 9732 11840
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9600 11558 9628 11698
rect 9784 11626 9812 11852
rect 9876 11762 9904 13398
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9968 11354 9996 14334
rect 10152 13870 10180 17818
rect 10244 14634 10272 18634
rect 10336 15162 10364 18799
rect 10508 18760 10560 18766
rect 10508 18702 10560 18708
rect 10520 17338 10548 18702
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10428 16794 10456 16934
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10506 16552 10562 16561
rect 10506 16487 10562 16496
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10428 15706 10456 15846
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10414 15464 10470 15473
rect 10414 15399 10470 15408
rect 10428 15366 10456 15399
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10322 14648 10378 14657
rect 10244 14606 10322 14634
rect 10322 14583 10378 14592
rect 10322 14512 10378 14521
rect 10322 14447 10324 14456
rect 10376 14447 10378 14456
rect 10324 14418 10376 14424
rect 10322 14240 10378 14249
rect 10244 14198 10322 14226
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 10060 13190 10088 13670
rect 10244 13376 10272 14198
rect 10322 14175 10378 14184
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10336 13530 10364 13806
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10428 13433 10456 14758
rect 10414 13424 10470 13433
rect 10324 13388 10376 13394
rect 10244 13348 10324 13376
rect 10520 13394 10548 16487
rect 10612 15434 10640 20975
rect 10704 19417 10732 21422
rect 10796 21321 10824 21422
rect 10782 21312 10838 21321
rect 10782 21247 10838 21256
rect 10888 20874 10916 21422
rect 10980 21078 11008 21519
rect 11072 21486 11100 22170
rect 12268 21962 12296 22238
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 22468 22228 22520 22234
rect 22468 22170 22520 22176
rect 14004 22092 14056 22098
rect 14004 22034 14056 22040
rect 14280 22092 14332 22098
rect 14280 22034 14332 22040
rect 13818 21992 13874 22001
rect 12072 21956 12124 21962
rect 12256 21956 12308 21962
rect 12124 21916 12204 21944
rect 12072 21898 12124 21904
rect 11783 21788 12091 21797
rect 11783 21786 11789 21788
rect 11845 21786 11869 21788
rect 11925 21786 11949 21788
rect 12005 21786 12029 21788
rect 12085 21786 12091 21788
rect 11845 21734 11847 21786
rect 12027 21734 12029 21786
rect 11783 21732 11789 21734
rect 11845 21732 11869 21734
rect 11925 21732 11949 21734
rect 12005 21732 12029 21734
rect 12085 21732 12091 21734
rect 11783 21723 12091 21732
rect 11256 21644 11560 21672
rect 11256 21486 11284 21644
rect 11428 21548 11480 21554
rect 11428 21490 11480 21496
rect 11060 21480 11112 21486
rect 11060 21422 11112 21428
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 10968 21072 11020 21078
rect 10968 21014 11020 21020
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 10876 20868 10928 20874
rect 10876 20810 10928 20816
rect 10888 20602 10916 20810
rect 10966 20632 11022 20641
rect 10876 20596 10928 20602
rect 10966 20567 10968 20576
rect 10876 20538 10928 20544
rect 11020 20567 11022 20576
rect 10968 20538 11020 20544
rect 10888 19922 10916 20538
rect 11072 20482 11100 20878
rect 11072 20454 11192 20482
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10876 19916 10928 19922
rect 10876 19858 10928 19864
rect 10690 19408 10746 19417
rect 10690 19343 10746 19352
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10980 19334 11008 20334
rect 10692 19304 10744 19310
rect 10690 19272 10692 19281
rect 10744 19272 10746 19281
rect 10690 19207 10746 19216
rect 10704 18698 10732 19207
rect 10796 18902 10824 19314
rect 10980 19306 11100 19334
rect 11164 19310 11192 20454
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 11256 20058 11284 20334
rect 11244 20052 11296 20058
rect 11244 19994 11296 20000
rect 11244 19938 11296 19944
rect 11244 19880 11296 19886
rect 11256 19310 11284 19880
rect 10784 18896 10836 18902
rect 10784 18838 10836 18844
rect 10692 18692 10744 18698
rect 10692 18634 10744 18640
rect 10692 18080 10744 18086
rect 10690 18048 10692 18057
rect 10744 18048 10746 18057
rect 10690 17983 10746 17992
rect 11072 17882 11100 19306
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11242 18864 11298 18873
rect 11242 18799 11298 18808
rect 11256 18766 11284 18799
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11058 17776 11114 17785
rect 11058 17711 11114 17720
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10600 15428 10652 15434
rect 10600 15370 10652 15376
rect 10598 15192 10654 15201
rect 10598 15127 10654 15136
rect 10414 13359 10470 13368
rect 10508 13388 10560 13394
rect 10324 13330 10376 13336
rect 10508 13330 10560 13336
rect 10336 13258 10364 13330
rect 10612 13258 10640 15127
rect 10704 15026 10732 17478
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10782 16824 10838 16833
rect 10888 16794 10916 17070
rect 10782 16759 10838 16768
rect 10876 16788 10928 16794
rect 10796 16658 10824 16759
rect 10876 16730 10928 16736
rect 10980 16674 11008 17478
rect 11072 17338 11100 17711
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 11058 16960 11114 16969
rect 11058 16895 11114 16904
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10888 16646 11008 16674
rect 10782 15872 10838 15881
rect 10782 15807 10838 15816
rect 10796 15570 10824 15807
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10888 14822 10916 16646
rect 11072 16454 11100 16895
rect 11164 16640 11192 18566
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11256 17134 11284 17614
rect 11348 17134 11376 21286
rect 11440 20806 11468 21490
rect 11532 20942 11560 21644
rect 11704 21480 11756 21486
rect 11704 21422 11756 21428
rect 11612 21344 11664 21350
rect 11610 21312 11612 21321
rect 11664 21312 11666 21321
rect 11610 21247 11666 21256
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 11428 20800 11480 20806
rect 11428 20742 11480 20748
rect 11532 20058 11560 20878
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11440 19009 11468 19790
rect 11532 19174 11560 19994
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11426 19000 11482 19009
rect 11426 18935 11482 18944
rect 11440 17814 11468 18935
rect 11624 18902 11652 20198
rect 11612 18896 11664 18902
rect 11612 18838 11664 18844
rect 11520 18760 11572 18766
rect 11520 18702 11572 18708
rect 11428 17808 11480 17814
rect 11428 17750 11480 17756
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 11256 16776 11284 17070
rect 11256 16748 11376 16776
rect 11348 16658 11376 16748
rect 11336 16652 11388 16658
rect 11164 16612 11284 16640
rect 11150 16552 11206 16561
rect 11150 16487 11206 16496
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 11072 15638 11100 16118
rect 11164 15910 11192 16487
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11164 15745 11192 15846
rect 11150 15736 11206 15745
rect 11150 15671 11206 15680
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 11060 15360 11112 15366
rect 11058 15328 11060 15337
rect 11112 15328 11114 15337
rect 11058 15263 11114 15272
rect 11256 15178 11284 16612
rect 11336 16594 11388 16600
rect 11348 16046 11376 16594
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11348 15638 11376 15982
rect 11336 15632 11388 15638
rect 11336 15574 11388 15580
rect 11164 15150 11284 15178
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10888 14278 10916 14758
rect 11164 14498 11192 15150
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11256 14618 11284 15030
rect 11348 14958 11376 15574
rect 11336 14952 11388 14958
rect 11336 14894 11388 14900
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11440 14550 11468 17750
rect 11532 17678 11560 18702
rect 11624 18290 11652 18838
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11716 17921 11744 21422
rect 12176 21049 12204 21916
rect 12256 21898 12308 21904
rect 12716 21956 12768 21962
rect 13818 21927 13874 21936
rect 12716 21898 12768 21904
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 12254 21584 12310 21593
rect 12254 21519 12310 21528
rect 12162 21040 12218 21049
rect 12162 20975 12218 20984
rect 12268 20806 12296 21519
rect 12348 21344 12400 21350
rect 12348 21286 12400 21292
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 11783 20700 12091 20709
rect 11783 20698 11789 20700
rect 11845 20698 11869 20700
rect 11925 20698 11949 20700
rect 12005 20698 12029 20700
rect 12085 20698 12091 20700
rect 11845 20646 11847 20698
rect 12027 20646 12029 20698
rect 11783 20644 11789 20646
rect 11845 20644 11869 20646
rect 11925 20644 11949 20646
rect 12005 20644 12029 20646
rect 12085 20644 12091 20646
rect 11783 20635 12091 20644
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 11783 19612 12091 19621
rect 11783 19610 11789 19612
rect 11845 19610 11869 19612
rect 11925 19610 11949 19612
rect 12005 19610 12029 19612
rect 12085 19610 12091 19612
rect 11845 19558 11847 19610
rect 12027 19558 12029 19610
rect 11783 19556 11789 19558
rect 11845 19556 11869 19558
rect 11925 19556 11949 19558
rect 12005 19556 12029 19558
rect 12085 19556 12091 19558
rect 11783 19547 12091 19556
rect 12268 19310 12296 19790
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 11783 18524 12091 18533
rect 11783 18522 11789 18524
rect 11845 18522 11869 18524
rect 11925 18522 11949 18524
rect 12005 18522 12029 18524
rect 12085 18522 12091 18524
rect 11845 18470 11847 18522
rect 12027 18470 12029 18522
rect 11783 18468 11789 18470
rect 11845 18468 11869 18470
rect 11925 18468 11949 18470
rect 12005 18468 12029 18470
rect 12085 18468 12091 18470
rect 11783 18459 12091 18468
rect 11702 17912 11758 17921
rect 12176 17882 12204 18702
rect 11702 17847 11758 17856
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11783 17436 12091 17445
rect 11783 17434 11789 17436
rect 11845 17434 11869 17436
rect 11925 17434 11949 17436
rect 12005 17434 12029 17436
rect 12085 17434 12091 17436
rect 11845 17382 11847 17434
rect 12027 17382 12029 17434
rect 11783 17380 11789 17382
rect 11845 17380 11869 17382
rect 11925 17380 11949 17382
rect 12005 17380 12029 17382
rect 12085 17380 12091 17382
rect 11783 17371 12091 17380
rect 11532 17292 12112 17320
rect 11532 16114 11560 17292
rect 12084 16998 12112 17292
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11992 16674 12020 16934
rect 12176 16674 12204 17818
rect 12254 17096 12310 17105
rect 12254 17031 12310 17040
rect 11992 16658 12204 16674
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11980 16652 12204 16658
rect 12032 16646 12204 16652
rect 11980 16594 12032 16600
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11520 15428 11572 15434
rect 11520 15370 11572 15376
rect 11428 14544 11480 14550
rect 11072 14482 11376 14498
rect 11428 14486 11480 14492
rect 11072 14476 11388 14482
rect 11072 14470 11336 14476
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10704 13394 10732 13670
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10324 13252 10376 13258
rect 10324 13194 10376 13200
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10600 13252 10652 13258
rect 10600 13194 10652 13200
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10152 12968 10180 13126
rect 10152 12940 10364 12968
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10152 12594 10180 12786
rect 10152 12566 10272 12594
rect 10244 12442 10272 12566
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10336 11762 10364 12940
rect 10428 12850 10456 13194
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10416 12232 10468 12238
rect 10414 12200 10416 12209
rect 10468 12200 10470 12209
rect 10414 12135 10470 12144
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10520 11558 10548 13126
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10704 12646 10732 12786
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10692 12368 10744 12374
rect 10692 12310 10744 12316
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9954 11248 10010 11257
rect 9954 11183 10010 11192
rect 9864 11144 9916 11150
rect 9586 11112 9642 11121
rect 9508 11070 9586 11098
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9048 9518 9076 9998
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8574 9072 8630 9081
rect 8574 9007 8630 9016
rect 8772 8974 8800 9386
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8852 8560 8904 8566
rect 8850 8528 8852 8537
rect 9036 8560 9088 8566
rect 8904 8528 8906 8537
rect 9140 8548 9168 9658
rect 9324 9586 9352 10202
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9324 8650 9352 9522
rect 9416 9110 9444 10542
rect 9508 10266 9536 11070
rect 9864 11086 9916 11092
rect 9586 11047 9642 11056
rect 9876 10674 9904 11086
rect 9968 11014 9996 11183
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 10060 10470 10088 11494
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9508 9178 9536 9522
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9324 8622 9444 8650
rect 9088 8520 9168 8548
rect 9312 8560 9364 8566
rect 9036 8502 9088 8508
rect 9312 8502 9364 8508
rect 8850 8463 8906 8472
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 7748 8288 7800 8294
rect 7654 8256 7710 8265
rect 7748 8230 7800 8236
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 7654 8191 7710 8200
rect 7668 7954 7696 8191
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7760 7410 7788 8230
rect 7988 8188 8296 8197
rect 7988 8186 7994 8188
rect 8050 8186 8074 8188
rect 8130 8186 8154 8188
rect 8210 8186 8234 8188
rect 8290 8186 8296 8188
rect 8050 8134 8052 8186
rect 8232 8134 8234 8186
rect 7988 8132 7994 8134
rect 8050 8132 8074 8134
rect 8130 8132 8154 8134
rect 8210 8132 8234 8134
rect 8290 8132 8296 8134
rect 7988 8123 8296 8132
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8208 7880 8260 7886
rect 8206 7848 8208 7857
rect 8260 7848 8262 7857
rect 8206 7783 8262 7792
rect 8772 7410 8800 7890
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 7562 7304 7618 7313
rect 7562 7239 7564 7248
rect 7616 7239 7618 7248
rect 7564 7210 7616 7216
rect 7988 7100 8296 7109
rect 7988 7098 7994 7100
rect 8050 7098 8074 7100
rect 8130 7098 8154 7100
rect 8210 7098 8234 7100
rect 8290 7098 8296 7100
rect 8050 7046 8052 7098
rect 8232 7046 8234 7098
rect 7988 7044 7994 7046
rect 8050 7044 8074 7046
rect 8130 7044 8154 7046
rect 8210 7044 8234 7046
rect 8290 7044 8296 7046
rect 7988 7035 8296 7044
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7944 6458 7972 6598
rect 8312 6458 8340 6666
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 8404 6254 8432 6598
rect 7156 6208 7328 6236
rect 8392 6248 8444 6254
rect 7104 6190 7156 6196
rect 8392 6190 8444 6196
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 7116 5778 7144 6190
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 7988 6012 8296 6021
rect 7988 6010 7994 6012
rect 8050 6010 8074 6012
rect 8130 6010 8154 6012
rect 8210 6010 8234 6012
rect 8290 6010 8296 6012
rect 8050 5958 8052 6010
rect 8232 5958 8234 6010
rect 7988 5956 7994 5958
rect 8050 5956 8074 5958
rect 8130 5956 8154 5958
rect 8210 5956 8234 5958
rect 8290 5956 8296 5958
rect 7988 5947 8296 5956
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 7104 5772 7156 5778
rect 7104 5714 7156 5720
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 6458 5672 6514 5681
rect 6458 5607 6514 5616
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6380 5222 6500 5250
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6000 4684 6052 4690
rect 6184 4684 6236 4690
rect 6052 4644 6184 4672
rect 6000 4626 6052 4632
rect 6184 4626 6236 4632
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5460 3074 5488 3946
rect 5828 3738 5856 4558
rect 5920 4078 5948 4558
rect 6012 4078 6040 4626
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 5920 3777 5948 4014
rect 5906 3768 5962 3777
rect 5816 3732 5868 3738
rect 5906 3703 5908 3712
rect 5816 3674 5868 3680
rect 5960 3703 5962 3712
rect 5908 3674 5960 3680
rect 6012 3618 6040 4014
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 5920 3590 6040 3618
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5276 3046 5488 3074
rect 5276 2990 5304 3046
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5460 2774 5488 2926
rect 5276 2746 5488 2774
rect 5170 2544 5226 2553
rect 5170 2479 5226 2488
rect 5080 1488 5132 1494
rect 5080 1430 5132 1436
rect 5170 1456 5226 1465
rect 5170 1391 5226 1400
rect 4804 1012 4856 1018
rect 4804 954 4856 960
rect 4988 1012 5040 1018
rect 4988 954 5040 960
rect 5184 882 5212 1391
rect 5276 1018 5304 2746
rect 5354 2544 5410 2553
rect 5354 2479 5410 2488
rect 5368 1358 5396 2479
rect 5644 2378 5672 3130
rect 5920 2582 5948 3590
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 5998 2952 6054 2961
rect 5998 2887 6000 2896
rect 6052 2887 6054 2896
rect 6000 2858 6052 2864
rect 5998 2680 6054 2689
rect 6104 2632 6132 2994
rect 6054 2624 6132 2632
rect 5998 2615 6000 2624
rect 6052 2604 6132 2624
rect 6000 2586 6052 2592
rect 5908 2576 5960 2582
rect 5908 2518 5960 2524
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 5538 2000 5594 2009
rect 5538 1935 5594 1944
rect 5552 1562 5580 1935
rect 5540 1556 5592 1562
rect 5540 1498 5592 1504
rect 5828 1426 5856 2450
rect 6196 1902 6224 3878
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6288 1970 6316 3674
rect 6380 3602 6408 4966
rect 6472 3670 6500 5222
rect 6564 4690 6592 5510
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6656 4570 6684 5714
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6564 4542 6684 4570
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6380 3058 6408 3538
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6472 2632 6500 3606
rect 6564 2825 6592 4542
rect 6748 4146 6776 5510
rect 6826 5128 6882 5137
rect 6882 5086 6960 5114
rect 6826 5063 6882 5072
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6840 4486 6868 4966
rect 6932 4690 6960 5086
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 7116 4486 7144 5714
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7208 4593 7236 5646
rect 7472 5568 7524 5574
rect 7472 5510 7524 5516
rect 7484 5370 7512 5510
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7668 4826 7696 5714
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7760 4622 7788 5714
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 7748 4616 7800 4622
rect 7194 4584 7250 4593
rect 7748 4558 7800 4564
rect 7194 4519 7250 4528
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6932 3738 6960 4014
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 6918 3632 6974 3641
rect 7116 3618 7144 4422
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 6974 3602 7144 3618
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 6974 3596 7156 3602
rect 6974 3590 7104 3596
rect 6918 3567 6974 3576
rect 7104 3538 7156 3544
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6550 2816 6606 2825
rect 6550 2751 6606 2760
rect 6380 2604 6500 2632
rect 6380 2514 6408 2604
rect 6368 2508 6420 2514
rect 6368 2450 6420 2456
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 6368 2372 6420 2378
rect 6368 2314 6420 2320
rect 6380 1970 6408 2314
rect 6276 1964 6328 1970
rect 6276 1906 6328 1912
rect 6368 1964 6420 1970
rect 6368 1906 6420 1912
rect 6184 1896 6236 1902
rect 6184 1838 6236 1844
rect 6472 1426 6500 2450
rect 6656 2106 6684 2994
rect 6748 2514 6776 3470
rect 7196 3460 7248 3466
rect 7196 3402 7248 3408
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6840 2650 6868 2790
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6552 1760 6604 1766
rect 6550 1728 6552 1737
rect 6604 1728 6606 1737
rect 6550 1663 6606 1672
rect 6840 1562 6868 2586
rect 7208 2514 7236 3402
rect 7576 2854 7604 3606
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 6828 1556 6880 1562
rect 6828 1498 6880 1504
rect 5816 1420 5868 1426
rect 5816 1362 5868 1368
rect 6460 1420 6512 1426
rect 6460 1362 6512 1368
rect 5356 1352 5408 1358
rect 5356 1294 5408 1300
rect 5264 1012 5316 1018
rect 5264 954 5316 960
rect 6472 882 6500 1362
rect 6734 1320 6790 1329
rect 6734 1255 6790 1264
rect 6642 1048 6698 1057
rect 6642 983 6698 992
rect 6656 882 6684 983
rect 6748 882 6776 1255
rect 5172 876 5224 882
rect 5172 818 5224 824
rect 6460 876 6512 882
rect 6460 818 6512 824
rect 6644 876 6696 882
rect 6644 818 6696 824
rect 6736 876 6788 882
rect 6736 818 6788 824
rect 5632 808 5684 814
rect 5632 750 5684 756
rect 6000 808 6052 814
rect 6000 750 6052 756
rect 4252 672 4304 678
rect 4252 614 4304 620
rect 4264 377 4292 614
rect 5644 474 5672 750
rect 6012 474 6040 750
rect 6840 678 6868 1498
rect 7300 882 7328 2246
rect 7288 876 7340 882
rect 7288 818 7340 824
rect 6828 672 6880 678
rect 6828 614 6880 620
rect 5632 468 5684 474
rect 5632 410 5684 416
rect 6000 468 6052 474
rect 6000 410 6052 416
rect 4250 368 4306 377
rect 3976 332 4028 338
rect 4250 303 4306 312
rect 3976 274 4028 280
rect 7668 270 7696 4150
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7760 3670 7788 3878
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 7852 3534 7880 5646
rect 7988 4924 8296 4933
rect 7988 4922 7994 4924
rect 8050 4922 8074 4924
rect 8130 4922 8154 4924
rect 8210 4922 8234 4924
rect 8290 4922 8296 4924
rect 8050 4870 8052 4922
rect 8232 4870 8234 4922
rect 7988 4868 7994 4870
rect 8050 4868 8074 4870
rect 8130 4868 8154 4870
rect 8210 4868 8234 4870
rect 8290 4868 8296 4870
rect 7988 4859 8296 4868
rect 8404 4826 8432 5646
rect 8496 5166 8524 5850
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8208 4616 8260 4622
rect 8206 4584 8208 4593
rect 8260 4584 8262 4593
rect 8206 4519 8262 4528
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8404 4282 8432 4422
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 7988 3836 8296 3845
rect 7988 3834 7994 3836
rect 8050 3834 8074 3836
rect 8130 3834 8154 3836
rect 8210 3834 8234 3836
rect 8290 3834 8296 3836
rect 8050 3782 8052 3834
rect 8232 3782 8234 3834
rect 7988 3780 7994 3782
rect 8050 3780 8074 3782
rect 8130 3780 8154 3782
rect 8210 3780 8234 3782
rect 8290 3780 8296 3782
rect 7988 3771 8296 3780
rect 8496 3738 8524 5102
rect 8588 4214 8616 6054
rect 8680 5914 8708 7346
rect 8772 6866 8800 7346
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8772 6322 8800 6802
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8864 6254 8892 8230
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8956 7274 8984 7822
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8680 5166 8708 5510
rect 8850 5264 8906 5273
rect 8772 5222 8850 5250
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8772 4729 8800 5222
rect 8850 5199 8906 5208
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 8758 4720 8814 4729
rect 8758 4655 8814 4664
rect 8666 4584 8722 4593
rect 8666 4519 8722 4528
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8680 4078 8708 4519
rect 8668 4072 8720 4078
rect 8574 4040 8630 4049
rect 8668 4014 8720 4020
rect 8574 3975 8630 3984
rect 8588 3942 8616 3975
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 7852 3126 7880 3470
rect 8404 3398 8432 3470
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8496 3194 8524 3334
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 8588 2774 8616 3878
rect 7988 2748 8296 2757
rect 7988 2746 7994 2748
rect 8050 2746 8074 2748
rect 8130 2746 8154 2748
rect 8210 2746 8234 2748
rect 8290 2746 8296 2748
rect 8050 2694 8052 2746
rect 8232 2694 8234 2746
rect 7988 2692 7994 2694
rect 8050 2692 8074 2694
rect 8130 2692 8154 2694
rect 8210 2692 8234 2694
rect 8290 2692 8296 2694
rect 7988 2683 8296 2692
rect 8496 2746 8616 2774
rect 8772 2774 8800 4655
rect 8956 4622 8984 5102
rect 9048 5030 9076 8502
rect 9324 8378 9352 8502
rect 9416 8430 9444 8622
rect 9508 8566 9536 8910
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9232 8350 9352 8378
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 9496 8424 9548 8430
rect 9600 8412 9628 9318
rect 9772 8900 9824 8906
rect 9772 8842 9824 8848
rect 9680 8424 9732 8430
rect 9600 8384 9680 8412
rect 9496 8366 9548 8372
rect 9680 8366 9732 8372
rect 9232 7936 9260 8350
rect 9404 8288 9456 8294
rect 9508 8276 9536 8366
rect 9784 8276 9812 8842
rect 9968 8430 9996 10406
rect 10152 10130 10180 10950
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10244 9042 10272 11154
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9508 8248 9812 8276
rect 9404 8230 9456 8236
rect 9416 8106 9444 8230
rect 9416 8078 9536 8106
rect 9232 7908 9352 7936
rect 9128 7880 9180 7886
rect 9324 7868 9352 7908
rect 9404 7880 9456 7886
rect 9324 7840 9404 7868
rect 9128 7822 9180 7828
rect 9404 7822 9456 7828
rect 9140 7721 9168 7822
rect 9126 7712 9182 7721
rect 9126 7647 9182 7656
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9416 7002 9444 7278
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9416 6322 9444 6938
rect 9508 6866 9536 8078
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9600 7721 9628 7822
rect 9586 7712 9642 7721
rect 9586 7647 9642 7656
rect 9692 6882 9720 8248
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9496 6860 9548 6866
rect 9692 6854 9812 6882
rect 9496 6802 9548 6808
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9128 6248 9180 6254
rect 9126 6216 9128 6225
rect 9180 6216 9182 6225
rect 9126 6151 9182 6160
rect 9220 6112 9272 6118
rect 9496 6112 9548 6118
rect 9272 6072 9444 6100
rect 9220 6054 9272 6060
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 9048 4690 9076 4966
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8956 3754 8984 4558
rect 9048 4146 9076 4626
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9036 3936 9088 3942
rect 9312 3936 9364 3942
rect 9088 3896 9260 3924
rect 9036 3878 9088 3884
rect 8956 3726 9076 3754
rect 9048 3602 9076 3726
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 9048 2990 9076 3538
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 8772 2746 8892 2774
rect 8496 1902 8524 2746
rect 8864 2106 8892 2746
rect 9048 2310 9076 2926
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9140 2650 9168 2790
rect 9232 2774 9260 3896
rect 9312 3878 9364 3884
rect 9324 2990 9352 3878
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9232 2746 9352 2774
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 8852 2100 8904 2106
rect 8852 2042 8904 2048
rect 9048 1970 9076 2246
rect 9036 1964 9088 1970
rect 9036 1906 9088 1912
rect 9140 1952 9168 2586
rect 9324 2514 9352 2746
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 9220 1964 9272 1970
rect 9140 1924 9220 1952
rect 8484 1896 8536 1902
rect 8484 1838 8536 1844
rect 7988 1660 8296 1669
rect 7988 1658 7994 1660
rect 8050 1658 8074 1660
rect 8130 1658 8154 1660
rect 8210 1658 8234 1660
rect 8290 1658 8296 1660
rect 8050 1606 8052 1658
rect 8232 1606 8234 1658
rect 7988 1604 7994 1606
rect 8050 1604 8074 1606
rect 8130 1604 8154 1606
rect 8210 1604 8234 1606
rect 8290 1604 8296 1606
rect 7988 1595 8296 1604
rect 9048 1562 9076 1906
rect 9036 1556 9088 1562
rect 9036 1498 9088 1504
rect 8668 1420 8720 1426
rect 8668 1362 8720 1368
rect 8024 1216 8076 1222
rect 8024 1158 8076 1164
rect 8298 1184 8354 1193
rect 8036 814 8064 1158
rect 8298 1119 8354 1128
rect 8312 950 8340 1119
rect 8300 944 8352 950
rect 8300 886 8352 892
rect 8680 882 8708 1362
rect 9036 1352 9088 1358
rect 9140 1340 9168 1924
rect 9220 1906 9272 1912
rect 9088 1312 9168 1340
rect 9220 1352 9272 1358
rect 9036 1294 9088 1300
rect 9220 1294 9272 1300
rect 9312 1352 9364 1358
rect 9312 1294 9364 1300
rect 9048 882 9076 1294
rect 9232 1018 9260 1294
rect 9324 1193 9352 1294
rect 9310 1184 9366 1193
rect 9310 1119 9366 1128
rect 9220 1012 9272 1018
rect 9220 954 9272 960
rect 9416 882 9444 6072
rect 9496 6054 9548 6060
rect 9508 5642 9536 6054
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9508 5370 9536 5578
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9692 5234 9720 6394
rect 9784 5846 9812 6854
rect 9876 6458 9904 7142
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 10060 5658 10088 8570
rect 10230 7032 10286 7041
rect 10230 6967 10286 6976
rect 10244 6254 10272 6967
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 9876 5630 10088 5658
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9588 5160 9640 5166
rect 9508 5120 9588 5148
rect 9508 4826 9536 5120
rect 9588 5102 9640 5108
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9508 3942 9536 4762
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9508 3534 9536 3878
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9508 2854 9536 3470
rect 9600 3194 9628 3878
rect 9692 3738 9720 4626
rect 9876 4214 9904 5630
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9876 3738 9904 4150
rect 10060 4146 10088 5510
rect 10152 4146 10180 5646
rect 10336 5545 10364 11290
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 10428 9586 10456 11018
rect 10520 10418 10548 11154
rect 10704 10674 10732 12310
rect 10796 12170 10824 13874
rect 10888 13274 10916 14214
rect 11072 13784 11100 14470
rect 11336 14418 11388 14424
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 10980 13756 11100 13784
rect 10980 13394 11008 13756
rect 11058 13696 11114 13705
rect 11058 13631 11114 13640
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10888 13246 11008 13274
rect 10874 12880 10930 12889
rect 10874 12815 10930 12824
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10782 11792 10838 11801
rect 10888 11762 10916 12815
rect 10980 12170 11008 13246
rect 11072 12753 11100 13631
rect 11058 12744 11114 12753
rect 11058 12679 11114 12688
rect 11164 12306 11192 14350
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 13258 11284 14214
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11440 13530 11468 13806
rect 11532 13802 11560 15370
rect 11624 15026 11652 15982
rect 11716 15910 11744 16594
rect 12268 16590 12296 17031
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12164 16448 12216 16454
rect 12162 16416 12164 16425
rect 12216 16416 12218 16425
rect 11783 16348 12091 16357
rect 12162 16351 12218 16360
rect 11783 16346 11789 16348
rect 11845 16346 11869 16348
rect 11925 16346 11949 16348
rect 12005 16346 12029 16348
rect 12085 16346 12091 16348
rect 11845 16294 11847 16346
rect 12027 16294 12029 16346
rect 11783 16292 11789 16294
rect 11845 16292 11869 16294
rect 11925 16292 11949 16294
rect 12005 16292 12029 16294
rect 12085 16292 12091 16294
rect 11783 16283 12091 16292
rect 12360 16046 12388 21286
rect 12438 20904 12494 20913
rect 12438 20839 12494 20848
rect 12452 19174 12480 20839
rect 12636 20346 12664 21830
rect 12728 21690 12756 21898
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12820 21690 12848 21830
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 13832 21554 13860 21927
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13360 21480 13412 21486
rect 13360 21422 13412 21428
rect 12636 20318 12756 20346
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12544 18426 12572 19790
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12636 16794 12664 18090
rect 12728 17202 12756 20318
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 13280 19446 13308 20198
rect 13268 19440 13320 19446
rect 13268 19382 13320 19388
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 12806 18048 12862 18057
rect 12806 17983 12862 17992
rect 12820 17270 12848 17983
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12806 16824 12862 16833
rect 12624 16788 12676 16794
rect 12806 16759 12808 16768
rect 12624 16730 12676 16736
rect 12860 16759 12862 16768
rect 12808 16730 12860 16736
rect 12348 16040 12400 16046
rect 12268 16000 12348 16028
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11716 15638 11744 15846
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11716 14822 11744 15574
rect 11783 15260 12091 15269
rect 11783 15258 11789 15260
rect 11845 15258 11869 15260
rect 11925 15258 11949 15260
rect 12005 15258 12029 15260
rect 12085 15258 12091 15260
rect 11845 15206 11847 15258
rect 12027 15206 12029 15258
rect 11783 15204 11789 15206
rect 11845 15204 11869 15206
rect 11925 15204 11949 15206
rect 12005 15204 12029 15206
rect 12085 15204 12091 15206
rect 11783 15195 12091 15204
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 11900 14822 11928 14894
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11624 13462 11652 14758
rect 11716 14550 11744 14758
rect 11704 14544 11756 14550
rect 11900 14498 11928 14758
rect 11992 14618 12020 14894
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11704 14486 11756 14492
rect 11716 14056 11744 14486
rect 11808 14470 11928 14498
rect 11808 14414 11836 14470
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11783 14172 12091 14181
rect 11783 14170 11789 14172
rect 11845 14170 11869 14172
rect 11925 14170 11949 14172
rect 12005 14170 12029 14172
rect 12085 14170 12091 14172
rect 11845 14118 11847 14170
rect 12027 14118 12029 14170
rect 11783 14116 11789 14118
rect 11845 14116 11869 14118
rect 11925 14116 11949 14118
rect 12005 14116 12029 14118
rect 12085 14116 12091 14118
rect 11783 14107 12091 14116
rect 11716 14028 11928 14056
rect 11900 13870 11928 14028
rect 12164 14000 12216 14006
rect 11978 13968 12034 13977
rect 12034 13926 12112 13954
rect 12164 13942 12216 13948
rect 11978 13903 12034 13912
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11978 13832 12034 13841
rect 11704 13796 11756 13802
rect 11978 13767 12034 13776
rect 11704 13738 11756 13744
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 11242 13016 11298 13025
rect 11242 12951 11298 12960
rect 11256 12918 11284 12951
rect 11244 12912 11296 12918
rect 11244 12854 11296 12860
rect 11440 12782 11468 13262
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11256 12646 11284 12718
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11336 12368 11388 12374
rect 11440 12356 11468 12718
rect 11388 12328 11468 12356
rect 11336 12310 11388 12316
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 10968 12164 11020 12170
rect 10968 12106 11020 12112
rect 10782 11727 10838 11736
rect 10876 11756 10928 11762
rect 10796 11286 10824 11727
rect 10876 11698 10928 11704
rect 11058 11656 11114 11665
rect 11058 11591 11114 11600
rect 10874 11384 10930 11393
rect 10874 11319 10930 11328
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10782 10432 10838 10441
rect 10520 10390 10782 10418
rect 10782 10367 10838 10376
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10508 9444 10560 9450
rect 10508 9386 10560 9392
rect 10520 9178 10548 9386
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10796 9042 10824 10367
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10796 8634 10824 8978
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10520 7002 10548 7414
rect 10600 7336 10652 7342
rect 10888 7324 10916 11319
rect 11072 11082 11100 11591
rect 11348 11354 11376 12310
rect 11532 12306 11560 13398
rect 11610 13016 11666 13025
rect 11610 12951 11666 12960
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11532 11694 11560 12242
rect 11624 12209 11652 12951
rect 11716 12442 11744 13738
rect 11888 13320 11940 13326
rect 11794 13288 11850 13297
rect 11850 13268 11888 13274
rect 11850 13262 11940 13268
rect 11850 13246 11928 13262
rect 11794 13223 11850 13232
rect 11992 13190 12020 13767
rect 12084 13394 12112 13926
rect 12176 13394 12204 13942
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11783 13084 12091 13093
rect 11783 13082 11789 13084
rect 11845 13082 11869 13084
rect 11925 13082 11949 13084
rect 12005 13082 12029 13084
rect 12085 13082 12091 13084
rect 11845 13030 11847 13082
rect 12027 13030 12029 13082
rect 11783 13028 11789 13030
rect 11845 13028 11869 13030
rect 11925 13028 11949 13030
rect 12005 13028 12029 13030
rect 12085 13028 12091 13030
rect 11783 13019 12091 13028
rect 12268 12866 12296 16000
rect 12348 15982 12400 15988
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12360 14006 12388 14350
rect 12544 14074 12572 15438
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12452 13161 12480 13874
rect 12636 13734 12664 16730
rect 12912 15162 12940 18702
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13096 18329 13124 18362
rect 13082 18320 13138 18329
rect 13082 18255 13138 18264
rect 13372 17785 13400 21422
rect 13728 21344 13780 21350
rect 13556 21304 13728 21332
rect 13556 19310 13584 21304
rect 13728 21286 13780 21292
rect 13818 21312 13874 21321
rect 13818 21247 13874 21256
rect 13832 20942 13860 21247
rect 14016 21078 14044 22034
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14094 21448 14150 21457
rect 14094 21383 14150 21392
rect 14004 21072 14056 21078
rect 14004 21014 14056 21020
rect 13912 21004 13964 21010
rect 13912 20946 13964 20952
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 13924 20058 13952 20946
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 13648 19310 13676 19994
rect 14108 19310 14136 21383
rect 14200 21298 14228 21830
rect 14292 21486 14320 22034
rect 14280 21480 14332 21486
rect 14280 21422 14332 21428
rect 14200 21270 14320 21298
rect 14188 21072 14240 21078
rect 14188 21014 14240 21020
rect 14200 20602 14228 21014
rect 14292 20874 14320 21270
rect 14372 21004 14424 21010
rect 14372 20946 14424 20952
rect 14280 20868 14332 20874
rect 14280 20810 14332 20816
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14200 19854 14228 20538
rect 14292 20398 14320 20810
rect 14384 20602 14412 20946
rect 14372 20596 14424 20602
rect 14372 20538 14424 20544
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14476 19854 14504 22170
rect 22480 22137 22508 22170
rect 23756 22160 23808 22166
rect 19338 22128 19394 22137
rect 22466 22128 22522 22137
rect 19338 22063 19340 22072
rect 19392 22063 19394 22072
rect 19708 22092 19760 22098
rect 19340 22034 19392 22040
rect 19708 22034 19760 22040
rect 21088 22092 21140 22098
rect 23756 22102 23808 22108
rect 22466 22063 22522 22072
rect 21088 22034 21140 22040
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 18880 21888 18932 21894
rect 18880 21830 18932 21836
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 14556 21684 14608 21690
rect 14556 21626 14608 21632
rect 14568 21486 14596 21626
rect 16868 21554 16896 21830
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 14556 21480 14608 21486
rect 14556 21422 14608 21428
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14188 19848 14240 19854
rect 14464 19848 14516 19854
rect 14240 19796 14412 19802
rect 14188 19790 14412 19796
rect 14464 19790 14516 19796
rect 14554 19816 14610 19825
rect 14200 19774 14412 19790
rect 14278 19408 14334 19417
rect 14278 19343 14334 19352
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13636 19304 13688 19310
rect 13636 19246 13688 19252
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13450 18864 13506 18873
rect 13450 18799 13506 18808
rect 13464 18426 13492 18799
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13634 18184 13690 18193
rect 13634 18119 13636 18128
rect 13688 18119 13690 18128
rect 13636 18090 13688 18096
rect 13358 17776 13414 17785
rect 13358 17711 13414 17720
rect 13634 17232 13690 17241
rect 13634 17167 13690 17176
rect 13648 17134 13676 17167
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 13648 16561 13676 17070
rect 13634 16552 13690 16561
rect 13634 16487 13690 16496
rect 13174 16416 13230 16425
rect 13174 16351 13230 16360
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13096 15706 13124 15846
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 13084 15088 13136 15094
rect 13082 15056 13084 15065
rect 13136 15056 13138 15065
rect 13082 14991 13138 15000
rect 12714 14512 12770 14521
rect 12714 14447 12770 14456
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12438 13152 12494 13161
rect 12438 13087 12494 13096
rect 12268 12838 12480 12866
rect 12256 12776 12308 12782
rect 12308 12736 12388 12764
rect 12256 12718 12308 12724
rect 11794 12608 11850 12617
rect 11794 12543 11850 12552
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11808 12374 11836 12543
rect 12360 12481 12388 12736
rect 12346 12472 12402 12481
rect 12346 12407 12402 12416
rect 12452 12374 12480 12838
rect 11796 12368 11848 12374
rect 12440 12368 12492 12374
rect 11796 12310 11848 12316
rect 11978 12336 12034 12345
rect 12440 12310 12492 12316
rect 11978 12271 12034 12280
rect 12072 12300 12124 12306
rect 11610 12200 11666 12209
rect 11992 12170 12020 12271
rect 12072 12242 12124 12248
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 11610 12135 11666 12144
rect 11980 12164 12032 12170
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11440 11558 11468 11630
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11624 10470 11652 12135
rect 11980 12106 12032 12112
rect 11704 12096 11756 12102
rect 12084 12084 12112 12242
rect 12084 12056 12204 12084
rect 11704 12038 11756 12044
rect 11716 11218 11744 12038
rect 11783 11996 12091 12005
rect 11783 11994 11789 11996
rect 11845 11994 11869 11996
rect 11925 11994 11949 11996
rect 12005 11994 12029 11996
rect 12085 11994 12091 11996
rect 11845 11942 11847 11994
rect 12027 11942 12029 11994
rect 11783 11940 11789 11942
rect 11845 11940 11869 11942
rect 11925 11940 11949 11942
rect 12005 11940 12029 11942
rect 12085 11940 12091 11942
rect 11783 11931 12091 11940
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11992 11801 12020 11834
rect 11978 11792 12034 11801
rect 11978 11727 12034 11736
rect 12176 11354 12204 12056
rect 12268 11694 12296 12242
rect 12544 12102 12572 13262
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12636 12442 12664 12786
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12728 12345 12756 14447
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 13082 14240 13138 14249
rect 12820 13530 12848 14214
rect 13082 14175 13138 14184
rect 13096 14006 13124 14175
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 13188 13870 13216 16351
rect 13740 16182 13768 18226
rect 13728 16176 13780 16182
rect 13728 16118 13780 16124
rect 13832 15881 13860 18566
rect 13924 18086 13952 18906
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 14016 16969 14044 19110
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14200 18426 14228 18770
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 14002 16960 14058 16969
rect 14002 16895 14058 16904
rect 14200 16658 14228 17138
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14200 16046 14228 16594
rect 14188 16040 14240 16046
rect 14188 15982 14240 15988
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 13818 15872 13874 15881
rect 13818 15807 13874 15816
rect 13450 15600 13506 15609
rect 13450 15535 13506 15544
rect 13464 14618 13492 15535
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13924 14226 13952 15914
rect 14200 15570 14228 15982
rect 14292 15978 14320 19343
rect 14384 18834 14412 19774
rect 14554 19751 14610 19760
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14384 17202 14412 18158
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14280 15972 14332 15978
rect 14280 15914 14332 15920
rect 14476 15706 14504 16730
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14200 15162 14228 15506
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14200 14958 14228 15098
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14200 14414 14228 14894
rect 14476 14822 14504 15642
rect 14568 15570 14596 19751
rect 14660 19514 14688 21422
rect 16396 21412 16448 21418
rect 16396 21354 16448 21360
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 15578 21244 15886 21253
rect 15578 21242 15584 21244
rect 15640 21242 15664 21244
rect 15720 21242 15744 21244
rect 15800 21242 15824 21244
rect 15880 21242 15886 21244
rect 15640 21190 15642 21242
rect 15822 21190 15824 21242
rect 15578 21188 15584 21190
rect 15640 21188 15664 21190
rect 15720 21188 15744 21190
rect 15800 21188 15824 21190
rect 15880 21188 15886 21190
rect 15578 21179 15886 21188
rect 16132 21146 16160 21286
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 15568 21072 15620 21078
rect 15936 21072 15988 21078
rect 15620 21020 15936 21026
rect 15568 21014 15988 21020
rect 15580 20998 15976 21014
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 15198 20632 15254 20641
rect 15108 20596 15160 20602
rect 15198 20567 15200 20576
rect 15108 20538 15160 20544
rect 15252 20567 15254 20576
rect 15200 20538 15252 20544
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 14844 20058 14872 20266
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 15120 19700 15148 20538
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15200 19712 15252 19718
rect 15120 19672 15200 19700
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14660 16590 14688 18022
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14660 15706 14688 15982
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14188 14408 14240 14414
rect 14108 14368 14188 14396
rect 13924 14198 14044 14226
rect 13360 14000 13412 14006
rect 13452 14000 13504 14006
rect 13360 13942 13412 13948
rect 13450 13968 13452 13977
rect 13504 13968 13506 13977
rect 12900 13864 12952 13870
rect 13176 13864 13228 13870
rect 12900 13806 12952 13812
rect 13096 13824 13176 13852
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12912 13433 12940 13806
rect 12992 13796 13044 13802
rect 12992 13738 13044 13744
rect 12898 13424 12954 13433
rect 12898 13359 12954 13368
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12820 12782 12848 13126
rect 13004 12918 13032 13738
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 12714 12336 12770 12345
rect 12714 12271 12770 12280
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12360 11937 12388 12038
rect 12346 11928 12402 11937
rect 12346 11863 12402 11872
rect 12438 11792 12494 11801
rect 12438 11727 12440 11736
rect 12492 11727 12494 11736
rect 12440 11698 12492 11704
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12268 11286 12296 11630
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 12544 11150 12572 12038
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12820 11540 12848 12174
rect 13004 11898 13032 12718
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 13096 11762 13124 13824
rect 13372 13841 13400 13942
rect 13450 13903 13506 13912
rect 13176 13806 13228 13812
rect 13358 13832 13414 13841
rect 13358 13767 13414 13776
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13188 13190 13216 13670
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13280 12986 13308 13262
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 13188 12434 13216 12582
rect 13188 12406 13308 12434
rect 13280 12306 13308 12406
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13556 12102 13584 12718
rect 13648 12646 13676 13466
rect 13832 13297 13860 13670
rect 13818 13288 13874 13297
rect 13818 13223 13874 13232
rect 13818 13152 13874 13161
rect 13818 13087 13874 13096
rect 13832 12850 13860 13087
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13648 12306 13676 12582
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13174 11928 13230 11937
rect 13230 11886 13308 11914
rect 13174 11863 13230 11872
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 12900 11552 12952 11558
rect 12820 11512 12900 11540
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12346 10976 12402 10985
rect 11783 10908 12091 10917
rect 11783 10906 11789 10908
rect 11845 10906 11869 10908
rect 11925 10906 11949 10908
rect 12005 10906 12029 10908
rect 12085 10906 12091 10908
rect 11845 10854 11847 10906
rect 12027 10854 12029 10906
rect 11783 10852 11789 10854
rect 11845 10852 11869 10854
rect 11925 10852 11949 10854
rect 12005 10852 12029 10854
rect 12085 10852 12091 10854
rect 11783 10843 12091 10852
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11426 10296 11482 10305
rect 11992 10266 12020 10542
rect 11426 10231 11482 10240
rect 11612 10260 11664 10266
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10980 9722 11008 10066
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 11072 9586 11100 9862
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11164 9518 11192 9998
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11164 8974 11192 9454
rect 11244 9376 11296 9382
rect 11296 9336 11376 9364
rect 11244 9318 11296 9324
rect 11242 9208 11298 9217
rect 11242 9143 11298 9152
rect 11256 9110 11284 9143
rect 11244 9104 11296 9110
rect 11244 9046 11296 9052
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10888 7296 11008 7324
rect 10600 7278 10652 7284
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10612 6730 10640 7278
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10784 6928 10836 6934
rect 10784 6870 10836 6876
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10506 6624 10562 6633
rect 10506 6559 10562 6568
rect 10520 5778 10548 6559
rect 10796 6390 10824 6870
rect 10888 6769 10916 7142
rect 10874 6760 10930 6769
rect 10874 6695 10930 6704
rect 10784 6384 10836 6390
rect 10784 6326 10836 6332
rect 10782 6080 10838 6089
rect 10782 6015 10838 6024
rect 10796 5914 10824 6015
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10520 5642 10548 5714
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10322 5536 10378 5545
rect 10322 5471 10378 5480
rect 10520 4146 10548 5578
rect 10704 5370 10732 5782
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9968 3738 9996 3946
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9968 3602 9996 3674
rect 10704 3602 10732 3878
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9496 1964 9548 1970
rect 9496 1906 9548 1912
rect 9508 1426 9536 1906
rect 9772 1896 9824 1902
rect 9772 1838 9824 1844
rect 9496 1420 9548 1426
rect 9496 1362 9548 1368
rect 9784 1222 9812 1838
rect 9772 1216 9824 1222
rect 9772 1158 9824 1164
rect 8668 876 8720 882
rect 8668 818 8720 824
rect 9036 876 9088 882
rect 9036 818 9088 824
rect 9404 876 9456 882
rect 9404 818 9456 824
rect 8024 808 8076 814
rect 8024 750 8076 756
rect 8576 808 8628 814
rect 8576 750 8628 756
rect 7988 572 8296 581
rect 7988 570 7994 572
rect 8050 570 8074 572
rect 8130 570 8154 572
rect 8210 570 8234 572
rect 8290 570 8296 572
rect 8050 518 8052 570
rect 8232 518 8234 570
rect 7988 516 7994 518
rect 8050 516 8074 518
rect 8130 516 8154 518
rect 8210 516 8234 518
rect 8290 516 8296 518
rect 7988 507 8296 516
rect 8588 406 8616 750
rect 10232 740 10284 746
rect 10232 682 10284 688
rect 10244 474 10272 682
rect 10232 468 10284 474
rect 10232 410 10284 416
rect 10796 406 10824 5714
rect 10980 5658 11008 7296
rect 11072 6730 11100 8774
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11164 7313 11192 7686
rect 11150 7304 11206 7313
rect 11150 7239 11206 7248
rect 11152 6860 11204 6866
rect 11256 6848 11284 9046
rect 11348 6882 11376 9336
rect 11440 8786 11468 10231
rect 11612 10202 11664 10208
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11624 9382 11652 10202
rect 11783 9820 12091 9829
rect 11783 9818 11789 9820
rect 11845 9818 11869 9820
rect 11925 9818 11949 9820
rect 12005 9818 12029 9820
rect 12085 9818 12091 9820
rect 11845 9766 11847 9818
rect 12027 9766 12029 9818
rect 11783 9764 11789 9766
rect 11845 9764 11869 9766
rect 11925 9764 11949 9766
rect 12005 9764 12029 9766
rect 12085 9764 12091 9766
rect 11783 9755 12091 9764
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11520 8968 11572 8974
rect 11624 8956 11652 9318
rect 11900 9178 11928 9454
rect 12176 9217 12204 10950
rect 12268 10538 12296 10950
rect 12346 10911 12402 10920
rect 12256 10532 12308 10538
rect 12256 10474 12308 10480
rect 12254 10296 12310 10305
rect 12254 10231 12310 10240
rect 12268 10130 12296 10231
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12360 10010 12388 10911
rect 12452 10146 12480 11086
rect 12636 10441 12664 11494
rect 12820 11218 12848 11512
rect 12900 11494 12952 11500
rect 13188 11354 13216 11562
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12820 11121 12848 11154
rect 13280 11150 13308 11886
rect 13360 11892 13412 11898
rect 13412 11852 13492 11880
rect 13360 11834 13412 11840
rect 13464 11150 13492 11852
rect 13556 11694 13584 12038
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13648 11558 13676 12242
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 12992 11144 13044 11150
rect 12806 11112 12862 11121
rect 12992 11086 13044 11092
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 12806 11047 12862 11056
rect 13004 10810 13032 11086
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 12912 10606 12940 10678
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12622 10432 12678 10441
rect 12622 10367 12678 10376
rect 13266 10432 13322 10441
rect 13266 10367 13322 10376
rect 12452 10118 12756 10146
rect 12268 9982 12388 10010
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12268 9926 12296 9982
rect 12256 9920 12308 9926
rect 12256 9862 12308 9868
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12162 9208 12218 9217
rect 11888 9172 11940 9178
rect 12162 9143 12218 9152
rect 11888 9114 11940 9120
rect 11572 8928 11652 8956
rect 11704 8968 11756 8974
rect 11520 8910 11572 8916
rect 11704 8910 11756 8916
rect 11440 8758 11560 8786
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11440 7410 11468 7890
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11532 7324 11560 8758
rect 11716 8634 11744 8910
rect 11783 8732 12091 8741
rect 11783 8730 11789 8732
rect 11845 8730 11869 8732
rect 11925 8730 11949 8732
rect 12005 8730 12029 8732
rect 12085 8730 12091 8732
rect 11845 8678 11847 8730
rect 12027 8678 12029 8730
rect 11783 8676 11789 8678
rect 11845 8676 11869 8678
rect 11925 8676 11949 8678
rect 12005 8676 12029 8678
rect 12085 8676 12091 8678
rect 11783 8667 12091 8676
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 12176 8498 12204 9143
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12268 8362 12296 8774
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11992 7954 12020 8230
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11783 7644 12091 7653
rect 11783 7642 11789 7644
rect 11845 7642 11869 7644
rect 11925 7642 11949 7644
rect 12005 7642 12029 7644
rect 12085 7642 12091 7644
rect 11845 7590 11847 7642
rect 12027 7590 12029 7642
rect 11783 7588 11789 7590
rect 11845 7588 11869 7590
rect 11925 7588 11949 7590
rect 12005 7588 12029 7590
rect 12085 7588 12091 7590
rect 11783 7579 12091 7588
rect 12360 7410 12388 9862
rect 12544 8294 12572 9998
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12452 7410 12480 8230
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 11532 7296 11744 7324
rect 11518 6896 11574 6905
rect 11348 6854 11518 6882
rect 11204 6820 11284 6848
rect 11518 6831 11520 6840
rect 11152 6802 11204 6808
rect 11572 6831 11574 6840
rect 11612 6860 11664 6866
rect 11520 6802 11572 6808
rect 11612 6802 11664 6808
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 11072 5778 11100 6122
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 10888 5630 11008 5658
rect 10888 5273 10916 5630
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10874 5264 10930 5273
rect 10874 5199 10930 5208
rect 10980 2825 11008 5510
rect 10966 2816 11022 2825
rect 10966 2751 11022 2760
rect 10968 2100 11020 2106
rect 10968 2042 11020 2048
rect 10980 1018 11008 2042
rect 11164 1426 11192 6802
rect 11624 6662 11652 6802
rect 11716 6662 11744 7296
rect 12452 7290 12480 7346
rect 12084 7262 12480 7290
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11992 6746 12020 6938
rect 12084 6866 12112 7262
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 6866 12480 7142
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12636 6798 12664 9318
rect 12728 8498 12756 10118
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 12716 8492 12768 8498
rect 12768 8452 12848 8480
rect 12716 8434 12768 8440
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12728 7954 12756 8230
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12624 6792 12676 6798
rect 11992 6718 12204 6746
rect 12624 6734 12676 6740
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11610 6488 11666 6497
rect 11244 6452 11296 6458
rect 11610 6423 11666 6432
rect 11244 6394 11296 6400
rect 11256 5778 11284 6394
rect 11428 6248 11480 6254
rect 11426 6216 11428 6225
rect 11624 6225 11652 6423
rect 11480 6216 11482 6225
rect 11426 6151 11482 6160
rect 11610 6216 11666 6225
rect 11610 6151 11666 6160
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11244 5772 11296 5778
rect 11296 5732 11468 5760
rect 11244 5714 11296 5720
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11256 4826 11284 5578
rect 11336 5160 11388 5166
rect 11336 5102 11388 5108
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11348 4622 11376 5102
rect 11440 4826 11468 5732
rect 11532 5166 11560 6054
rect 11716 5953 11744 6598
rect 11783 6556 12091 6565
rect 11783 6554 11789 6556
rect 11845 6554 11869 6556
rect 11925 6554 11949 6556
rect 12005 6554 12029 6556
rect 12085 6554 12091 6556
rect 11845 6502 11847 6554
rect 12027 6502 12029 6554
rect 11783 6500 11789 6502
rect 11845 6500 11869 6502
rect 11925 6500 11949 6502
rect 12005 6500 12029 6502
rect 12085 6500 12091 6502
rect 11783 6491 12091 6500
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12084 6254 12112 6394
rect 12176 6254 12204 6718
rect 12728 6458 12756 7278
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12820 6254 12848 8452
rect 13004 7886 13032 8774
rect 13280 8430 13308 10367
rect 13372 8838 13400 10678
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 13096 7342 13124 7822
rect 13084 7336 13136 7342
rect 12898 7304 12954 7313
rect 12954 7262 13032 7290
rect 13084 7278 13136 7284
rect 12898 7239 12954 7248
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12912 6254 12940 6938
rect 13004 6458 13032 7262
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 13096 7041 13124 7142
rect 13082 7032 13138 7041
rect 13082 6967 13138 6976
rect 13188 6866 13216 8230
rect 13176 6860 13228 6866
rect 13176 6802 13228 6808
rect 13268 6860 13320 6866
rect 13372 6848 13400 8774
rect 13464 8294 13492 11086
rect 13740 10606 13768 12786
rect 14016 12442 14044 14198
rect 14108 13938 14136 14368
rect 14188 14350 14240 14356
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 14200 13734 14228 14214
rect 14292 13870 14320 14758
rect 14476 14618 14504 14758
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14476 14498 14504 14554
rect 14476 14470 14596 14498
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14476 14278 14504 14350
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14568 13938 14596 14470
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14568 13326 14596 13874
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 14188 12640 14240 12646
rect 14188 12582 14240 12588
rect 14004 12436 14056 12442
rect 13832 12396 14004 12424
rect 13832 10985 13860 12396
rect 14004 12378 14056 12384
rect 14002 12336 14058 12345
rect 14002 12271 14004 12280
rect 14056 12271 14058 12280
rect 14004 12242 14056 12248
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13818 10976 13874 10985
rect 13818 10911 13874 10920
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13832 10130 13860 10610
rect 13924 10470 13952 11154
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 13832 9518 13860 10066
rect 13924 9722 13952 10406
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13832 9042 13860 9454
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13464 8266 13584 8294
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 7546 13492 7686
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13556 7154 13584 8266
rect 13320 6820 13400 6848
rect 13464 7126 13584 7154
rect 13268 6802 13320 6808
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11702 5944 11758 5953
rect 11702 5879 11758 5888
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11532 4690 11560 4966
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11532 4554 11560 4626
rect 11624 4622 11652 5714
rect 11808 5556 11836 6054
rect 11992 5914 12020 6054
rect 11980 5908 12032 5914
rect 12084 5896 12112 6190
rect 12256 6112 12308 6118
rect 12308 6072 12480 6100
rect 12256 6054 12308 6060
rect 12256 5908 12308 5914
rect 12084 5868 12256 5896
rect 11980 5850 12032 5856
rect 12256 5850 12308 5856
rect 11716 5528 11836 5556
rect 12256 5568 12308 5574
rect 11716 5030 11744 5528
rect 12256 5510 12308 5516
rect 11783 5468 12091 5477
rect 11783 5466 11789 5468
rect 11845 5466 11869 5468
rect 11925 5466 11949 5468
rect 12005 5466 12029 5468
rect 12085 5466 12091 5468
rect 11845 5414 11847 5466
rect 12027 5414 12029 5466
rect 11783 5412 11789 5414
rect 11845 5412 11869 5414
rect 11925 5412 11949 5414
rect 12005 5412 12029 5414
rect 12085 5412 12091 5414
rect 11783 5403 12091 5412
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 4826 11744 4966
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11348 3602 11376 4422
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11440 3670 11468 3878
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 11336 3596 11388 3602
rect 11336 3538 11388 3544
rect 11244 2984 11296 2990
rect 11244 2926 11296 2932
rect 11256 2650 11284 2926
rect 11426 2680 11482 2689
rect 11244 2644 11296 2650
rect 11426 2615 11482 2624
rect 11244 2586 11296 2592
rect 11256 2446 11284 2586
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11256 1902 11284 2382
rect 11244 1896 11296 1902
rect 11244 1838 11296 1844
rect 11152 1420 11204 1426
rect 11152 1362 11204 1368
rect 10968 1012 11020 1018
rect 10968 954 11020 960
rect 11164 814 11192 1362
rect 11440 1057 11468 2615
rect 11532 1426 11560 4082
rect 11624 3534 11652 4558
rect 11716 4146 11744 4762
rect 12268 4690 12296 5510
rect 12452 4690 12480 6072
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 11783 4380 12091 4389
rect 11783 4378 11789 4380
rect 11845 4378 11869 4380
rect 11925 4378 11949 4380
rect 12005 4378 12029 4380
rect 12085 4378 12091 4380
rect 11845 4326 11847 4378
rect 12027 4326 12029 4378
rect 11783 4324 11789 4326
rect 11845 4324 11869 4326
rect 11925 4324 11949 4326
rect 12005 4324 12029 4326
rect 12085 4324 12091 4326
rect 11783 4315 12091 4324
rect 12176 4282 12204 4558
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12254 4312 12310 4321
rect 12164 4276 12216 4282
rect 12254 4247 12310 4256
rect 12164 4218 12216 4224
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11716 3738 11744 4082
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11624 2990 11652 3470
rect 11612 2984 11664 2990
rect 11612 2926 11664 2932
rect 11716 2854 11744 3674
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 11783 3292 12091 3301
rect 11783 3290 11789 3292
rect 11845 3290 11869 3292
rect 11925 3290 11949 3292
rect 12005 3290 12029 3292
rect 12085 3290 12091 3292
rect 11845 3238 11847 3290
rect 12027 3238 12029 3290
rect 11783 3236 11789 3238
rect 11845 3236 11869 3238
rect 11925 3236 11949 3238
rect 12005 3236 12029 3238
rect 12085 3236 12091 3238
rect 11783 3227 12091 3236
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11808 3058 11836 3130
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11794 2816 11850 2825
rect 11716 2650 11744 2790
rect 11794 2751 11850 2760
rect 11704 2644 11756 2650
rect 11704 2586 11756 2592
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11624 1426 11652 2382
rect 11716 1952 11744 2586
rect 11808 2446 11836 2751
rect 12176 2632 12204 3470
rect 12268 2689 12296 4247
rect 12820 4078 12848 4422
rect 13280 4146 13308 6802
rect 13464 6798 13492 7126
rect 13542 7032 13598 7041
rect 13542 6967 13598 6976
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13358 6624 13414 6633
rect 13358 6559 13414 6568
rect 13372 6254 13400 6559
rect 13464 6322 13492 6734
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13372 5234 13400 6054
rect 13556 5681 13584 6967
rect 13648 6458 13676 8434
rect 13832 8430 13860 8978
rect 14016 8974 14044 12242
rect 14094 11792 14150 11801
rect 14094 11727 14096 11736
rect 14148 11727 14150 11736
rect 14096 11698 14148 11704
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14108 10266 14136 10542
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14108 9586 14136 10202
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14108 9178 14136 9522
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 14016 8378 14044 8910
rect 14108 8498 14136 9114
rect 14200 8498 14228 12582
rect 14384 12434 14412 13126
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14292 12406 14412 12434
rect 14292 8956 14320 12406
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14384 10674 14412 10950
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14476 10130 14504 12038
rect 14568 11393 14596 12718
rect 14752 12434 14780 19654
rect 15016 18760 15068 18766
rect 15120 18748 15148 19672
rect 15200 19654 15252 19660
rect 15396 19514 15424 20198
rect 15578 20156 15886 20165
rect 15578 20154 15584 20156
rect 15640 20154 15664 20156
rect 15720 20154 15744 20156
rect 15800 20154 15824 20156
rect 15880 20154 15886 20156
rect 15640 20102 15642 20154
rect 15822 20102 15824 20154
rect 15578 20100 15584 20102
rect 15640 20100 15664 20102
rect 15720 20100 15744 20102
rect 15800 20100 15824 20102
rect 15880 20100 15886 20102
rect 15578 20091 15886 20100
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15384 19508 15436 19514
rect 15384 19450 15436 19456
rect 15856 19378 15884 19654
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15948 19310 15976 20402
rect 16224 20330 16252 20946
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16212 20324 16264 20330
rect 16212 20266 16264 20272
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 16040 19310 16068 19858
rect 16224 19854 16252 20266
rect 16316 19922 16344 20878
rect 16408 20602 16436 21354
rect 16776 20913 16804 21354
rect 16762 20904 16818 20913
rect 16762 20839 16818 20848
rect 16764 20800 16816 20806
rect 16684 20760 16764 20788
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16578 20496 16634 20505
rect 16578 20431 16634 20440
rect 16396 20392 16448 20398
rect 16396 20334 16448 20340
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16118 19272 16174 19281
rect 15578 19068 15886 19077
rect 15578 19066 15584 19068
rect 15640 19066 15664 19068
rect 15720 19066 15744 19068
rect 15800 19066 15824 19068
rect 15880 19066 15886 19068
rect 15640 19014 15642 19066
rect 15822 19014 15824 19066
rect 15578 19012 15584 19014
rect 15640 19012 15664 19014
rect 15720 19012 15744 19014
rect 15800 19012 15824 19014
rect 15880 19012 15886 19014
rect 15578 19003 15886 19012
rect 15948 18986 15976 19246
rect 16118 19207 16174 19216
rect 15948 18958 16068 18986
rect 15292 18896 15344 18902
rect 15292 18838 15344 18844
rect 15068 18720 15148 18748
rect 15016 18702 15068 18708
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 14844 17134 14872 18022
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14844 16794 14872 17070
rect 14936 16998 14964 17070
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 14832 16788 14884 16794
rect 14884 16748 14964 16776
rect 14832 16730 14884 16736
rect 14936 16114 14964 16748
rect 15028 16697 15056 17614
rect 15304 16794 15332 18838
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 15578 17980 15886 17989
rect 15578 17978 15584 17980
rect 15640 17978 15664 17980
rect 15720 17978 15744 17980
rect 15800 17978 15824 17980
rect 15880 17978 15886 17980
rect 15640 17926 15642 17978
rect 15822 17926 15824 17978
rect 15578 17924 15584 17926
rect 15640 17924 15664 17926
rect 15720 17924 15744 17926
rect 15800 17924 15824 17926
rect 15880 17924 15886 17926
rect 15578 17915 15886 17924
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15014 16688 15070 16697
rect 15014 16623 15070 16632
rect 15488 16522 15516 17614
rect 15948 17542 15976 18770
rect 16040 18222 16068 18958
rect 16132 18902 16160 19207
rect 16120 18896 16172 18902
rect 16120 18838 16172 18844
rect 16224 18714 16252 19790
rect 16316 18834 16344 19858
rect 16408 18970 16436 20334
rect 16592 20058 16620 20431
rect 16580 20052 16632 20058
rect 16580 19994 16632 20000
rect 16684 19786 16712 20760
rect 16764 20742 16816 20748
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16486 19272 16542 19281
rect 16486 19207 16542 19216
rect 16396 18964 16448 18970
rect 16396 18906 16448 18912
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 16396 18760 16448 18766
rect 16132 18708 16396 18714
rect 16132 18702 16448 18708
rect 16132 18686 16436 18702
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 16132 17814 16160 18686
rect 16396 18420 16448 18426
rect 16396 18362 16448 18368
rect 16212 18080 16264 18086
rect 16408 18057 16436 18362
rect 16212 18022 16264 18028
rect 16394 18048 16450 18057
rect 16224 17882 16252 18022
rect 16394 17983 16450 17992
rect 16500 17882 16528 19207
rect 16684 18850 16712 19722
rect 16684 18834 16804 18850
rect 16960 18834 16988 19790
rect 17040 19236 17092 19242
rect 17040 19178 17092 19184
rect 16672 18828 16804 18834
rect 16724 18822 16804 18828
rect 16672 18770 16724 18776
rect 16672 18692 16724 18698
rect 16672 18634 16724 18640
rect 16684 18086 16712 18634
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 16684 17746 16712 18022
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16776 17660 16804 18822
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16948 17672 17000 17678
rect 16776 17632 16948 17660
rect 16948 17614 17000 17620
rect 16396 17604 16448 17610
rect 16396 17546 16448 17552
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 16408 17134 16436 17546
rect 17052 17490 17080 19178
rect 16960 17462 17080 17490
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16120 16992 16172 16998
rect 16120 16934 16172 16940
rect 15578 16892 15886 16901
rect 15578 16890 15584 16892
rect 15640 16890 15664 16892
rect 15720 16890 15744 16892
rect 15800 16890 15824 16892
rect 15880 16890 15886 16892
rect 15640 16838 15642 16890
rect 15822 16838 15824 16890
rect 15578 16836 15584 16838
rect 15640 16836 15664 16838
rect 15720 16836 15744 16838
rect 15800 16836 15824 16838
rect 15880 16836 15886 16838
rect 15578 16827 15886 16836
rect 16132 16794 16160 16934
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 15476 16516 15528 16522
rect 15476 16458 15528 16464
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 14844 15892 14872 16050
rect 15212 15892 15240 16050
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 14844 15864 15240 15892
rect 15304 15162 15332 15982
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15200 14952 15252 14958
rect 14830 14920 14886 14929
rect 15200 14894 15252 14900
rect 14830 14855 14886 14864
rect 14844 13938 14872 14855
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 13394 15056 13670
rect 15212 13530 15240 14894
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15396 13462 15424 15982
rect 15578 15804 15886 15813
rect 15578 15802 15584 15804
rect 15640 15802 15664 15804
rect 15720 15802 15744 15804
rect 15800 15802 15824 15804
rect 15880 15802 15886 15804
rect 15640 15750 15642 15802
rect 15822 15750 15824 15802
rect 15578 15748 15584 15750
rect 15640 15748 15664 15750
rect 15720 15748 15744 15750
rect 15800 15748 15824 15750
rect 15880 15748 15886 15750
rect 15578 15739 15886 15748
rect 15948 15570 15976 16390
rect 15936 15564 15988 15570
rect 15936 15506 15988 15512
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 16040 15162 16068 15302
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 15578 14716 15886 14725
rect 15578 14714 15584 14716
rect 15640 14714 15664 14716
rect 15720 14714 15744 14716
rect 15800 14714 15824 14716
rect 15880 14714 15886 14716
rect 15640 14662 15642 14714
rect 15822 14662 15824 14714
rect 15578 14660 15584 14662
rect 15640 14660 15664 14662
rect 15720 14660 15744 14662
rect 15800 14660 15824 14662
rect 15880 14660 15886 14662
rect 15578 14651 15886 14660
rect 16316 14600 16344 16458
rect 16408 15638 16436 17070
rect 16592 16810 16620 17138
rect 16592 16782 16712 16810
rect 16776 16794 16804 17138
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16396 15632 16448 15638
rect 16396 15574 16448 15580
rect 16408 15026 16436 15574
rect 16396 15020 16448 15026
rect 16448 14980 16528 15008
rect 16396 14962 16448 14968
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16224 14572 16344 14600
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15672 13841 15700 13942
rect 15658 13832 15714 13841
rect 15658 13767 15714 13776
rect 15578 13628 15886 13637
rect 15578 13626 15584 13628
rect 15640 13626 15664 13628
rect 15720 13626 15744 13628
rect 15800 13626 15824 13628
rect 15880 13626 15886 13628
rect 15640 13574 15642 13626
rect 15822 13574 15824 13626
rect 15578 13572 15584 13574
rect 15640 13572 15664 13574
rect 15720 13572 15744 13574
rect 15800 13572 15824 13574
rect 15880 13572 15886 13574
rect 15578 13563 15886 13572
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15016 12436 15068 12442
rect 14752 12406 14872 12434
rect 14844 11880 14872 12406
rect 15016 12378 15068 12384
rect 14924 11892 14976 11898
rect 14844 11852 14924 11880
rect 14554 11384 14610 11393
rect 14554 11319 14610 11328
rect 14844 11286 14872 11852
rect 14924 11834 14976 11840
rect 15028 11626 15056 12378
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14660 10810 14688 11086
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14568 10130 14596 10746
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14476 9178 14504 9454
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 14372 8968 14424 8974
rect 14292 8928 14372 8956
rect 14372 8910 14424 8916
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14016 8350 14136 8378
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13740 6458 13768 7482
rect 13924 7342 13952 7890
rect 13912 7336 13964 7342
rect 13910 7304 13912 7313
rect 13964 7304 13966 7313
rect 13910 7239 13966 7248
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 14016 6730 14044 7210
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13542 5672 13598 5681
rect 13542 5607 13598 5616
rect 13648 5302 13676 6122
rect 13912 5908 13964 5914
rect 14016 5896 14044 6666
rect 14108 6254 14136 8350
rect 14384 7410 14412 8774
rect 14844 8498 14872 11018
rect 14936 9586 14964 11494
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14464 7948 14516 7954
rect 14516 7908 14596 7936
rect 14464 7890 14516 7896
rect 14462 7848 14518 7857
rect 14462 7783 14518 7792
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14292 6322 14320 7142
rect 14476 6458 14504 7783
rect 14568 7206 14596 7908
rect 15028 7886 15056 9862
rect 15120 9382 15148 12922
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15488 11354 15516 12650
rect 15578 12540 15886 12549
rect 15578 12538 15584 12540
rect 15640 12538 15664 12540
rect 15720 12538 15744 12540
rect 15800 12538 15824 12540
rect 15880 12538 15886 12540
rect 15640 12486 15642 12538
rect 15822 12486 15824 12538
rect 15578 12484 15584 12486
rect 15640 12484 15664 12486
rect 15720 12484 15744 12486
rect 15800 12484 15824 12486
rect 15880 12484 15886 12486
rect 15578 12475 15886 12484
rect 15578 11452 15886 11461
rect 15578 11450 15584 11452
rect 15640 11450 15664 11452
rect 15720 11450 15744 11452
rect 15800 11450 15824 11452
rect 15880 11450 15886 11452
rect 15640 11398 15642 11450
rect 15822 11398 15824 11450
rect 15578 11396 15584 11398
rect 15640 11396 15664 11398
rect 15720 11396 15744 11398
rect 15800 11396 15824 11398
rect 15880 11396 15886 11398
rect 15578 11387 15886 11396
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15750 11112 15806 11121
rect 15476 11076 15528 11082
rect 15750 11047 15752 11056
rect 15476 11018 15528 11024
rect 15804 11047 15806 11056
rect 15752 11018 15804 11024
rect 15488 9518 15516 11018
rect 15578 10364 15886 10373
rect 15578 10362 15584 10364
rect 15640 10362 15664 10364
rect 15720 10362 15744 10364
rect 15800 10362 15824 10364
rect 15880 10362 15886 10364
rect 15640 10310 15642 10362
rect 15822 10310 15824 10362
rect 15578 10308 15584 10310
rect 15640 10308 15664 10310
rect 15720 10308 15744 10310
rect 15800 10308 15824 10310
rect 15880 10308 15886 10310
rect 15578 10299 15886 10308
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15108 9376 15160 9382
rect 15108 9318 15160 9324
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15200 8424 15252 8430
rect 15120 8384 15200 8412
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14568 6934 14596 7142
rect 14660 7002 14688 7346
rect 15120 7342 15148 8384
rect 15200 8366 15252 8372
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 14740 7336 14792 7342
rect 15108 7336 15160 7342
rect 14740 7278 14792 7284
rect 15106 7304 15108 7313
rect 15160 7304 15162 7313
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14556 6928 14608 6934
rect 14556 6870 14608 6876
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 13964 5868 14044 5896
rect 13912 5850 13964 5856
rect 14384 5778 14412 6326
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13648 4078 13676 5238
rect 13832 5098 13860 5646
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13924 5234 13952 5306
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13832 4622 13860 5034
rect 14200 5030 14228 5646
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14200 4826 14228 4966
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13832 4282 13860 4558
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12452 3738 12480 3878
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 13832 3534 13860 4218
rect 14200 4214 14228 4762
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14384 4486 14412 4558
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14188 4208 14240 4214
rect 14188 4150 14240 4156
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13910 3496 13966 3505
rect 13832 2990 13860 3470
rect 14016 3482 14044 4014
rect 14200 3738 14228 4150
rect 14568 4078 14596 6598
rect 14752 6322 14780 7278
rect 15106 7239 15162 7248
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 14924 6928 14976 6934
rect 14924 6870 14976 6876
rect 14936 6322 14964 6870
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 15120 4282 15148 6938
rect 15212 4593 15240 7822
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15304 7041 15332 7142
rect 15290 7032 15346 7041
rect 15290 6967 15346 6976
rect 15290 6488 15346 6497
rect 15290 6423 15346 6432
rect 15304 6089 15332 6423
rect 15396 6322 15424 9318
rect 15488 8974 15516 9454
rect 15578 9276 15886 9285
rect 15578 9274 15584 9276
rect 15640 9274 15664 9276
rect 15720 9274 15744 9276
rect 15800 9274 15824 9276
rect 15880 9274 15886 9276
rect 15640 9222 15642 9274
rect 15822 9222 15824 9274
rect 15578 9220 15584 9222
rect 15640 9220 15664 9222
rect 15720 9220 15744 9222
rect 15800 9220 15824 9222
rect 15880 9220 15886 9222
rect 15578 9211 15886 9220
rect 15948 9110 15976 14418
rect 16224 13954 16252 14572
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16316 14278 16344 14418
rect 16304 14272 16356 14278
rect 16302 14240 16304 14249
rect 16356 14240 16358 14249
rect 16302 14175 16358 14184
rect 16408 14074 16436 14758
rect 16500 14618 16528 14980
rect 16592 14657 16620 16594
rect 16684 16046 16712 16782
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16854 16552 16910 16561
rect 16854 16487 16856 16496
rect 16908 16487 16910 16496
rect 16856 16458 16908 16464
rect 16868 16046 16896 16458
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16856 16040 16908 16046
rect 16856 15982 16908 15988
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16868 15434 16896 15846
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 16960 15065 16988 17462
rect 17144 16130 17172 21626
rect 17958 21584 18014 21593
rect 17958 21519 18014 21528
rect 17972 21146 18000 21519
rect 18892 21486 18920 21830
rect 19064 21616 19116 21622
rect 19064 21558 19116 21564
rect 18788 21480 18840 21486
rect 18788 21422 18840 21428
rect 18880 21480 18932 21486
rect 18880 21422 18932 21428
rect 18800 21332 18828 21422
rect 18972 21344 19024 21350
rect 18800 21304 18972 21332
rect 18972 21286 19024 21292
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 18880 20936 18932 20942
rect 18932 20896 19012 20924
rect 18880 20878 18932 20884
rect 17224 20800 17276 20806
rect 17224 20742 17276 20748
rect 17236 18290 17264 20742
rect 17960 20324 18012 20330
rect 17960 20266 18012 20272
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 17500 20256 17552 20262
rect 17500 20198 17552 20204
rect 17512 19922 17540 20198
rect 17972 19922 18000 20266
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 17960 19236 18012 19242
rect 17960 19178 18012 19184
rect 17684 18760 17736 18766
rect 17972 18737 18000 19178
rect 18248 18873 18276 19246
rect 18234 18864 18290 18873
rect 18234 18799 18290 18808
rect 17684 18702 17736 18708
rect 17958 18728 18014 18737
rect 17696 18426 17724 18702
rect 17958 18663 18014 18672
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17960 18216 18012 18222
rect 18340 18170 18368 19246
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 17960 18158 18012 18164
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17512 16794 17540 17614
rect 17972 17542 18000 18158
rect 18248 18142 18368 18170
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17052 16102 17172 16130
rect 17052 15473 17080 16102
rect 17236 16046 17264 16526
rect 17512 16114 17540 16730
rect 17696 16590 17724 17478
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 18064 16794 18092 17206
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 18248 16425 18276 18142
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 18340 17746 18368 18022
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 18234 16416 18290 16425
rect 18234 16351 18290 16360
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17038 15464 17094 15473
rect 17038 15399 17094 15408
rect 16946 15056 17002 15065
rect 16946 14991 17002 15000
rect 16764 14816 16816 14822
rect 16764 14758 16816 14764
rect 16578 14648 16634 14657
rect 16488 14612 16540 14618
rect 16578 14583 16634 14592
rect 16488 14554 16540 14560
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16028 13932 16080 13938
rect 16224 13926 16344 13954
rect 16028 13874 16080 13880
rect 16040 13530 16068 13874
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15488 6848 15516 8910
rect 15578 8188 15886 8197
rect 15578 8186 15584 8188
rect 15640 8186 15664 8188
rect 15720 8186 15744 8188
rect 15800 8186 15824 8188
rect 15880 8186 15886 8188
rect 15640 8134 15642 8186
rect 15822 8134 15824 8186
rect 15578 8132 15584 8134
rect 15640 8132 15664 8134
rect 15720 8132 15744 8134
rect 15800 8132 15824 8134
rect 15880 8132 15886 8134
rect 15578 8123 15886 8132
rect 15578 7100 15886 7109
rect 15578 7098 15584 7100
rect 15640 7098 15664 7100
rect 15720 7098 15744 7100
rect 15800 7098 15824 7100
rect 15880 7098 15886 7100
rect 15640 7046 15642 7098
rect 15822 7046 15824 7098
rect 15578 7044 15584 7046
rect 15640 7044 15664 7046
rect 15720 7044 15744 7046
rect 15800 7044 15824 7046
rect 15880 7044 15886 7046
rect 15578 7035 15886 7044
rect 15948 6866 15976 9046
rect 16040 9042 16068 10406
rect 16132 9722 16160 10542
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 15752 6860 15804 6866
rect 15488 6820 15752 6848
rect 15752 6802 15804 6808
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15764 6769 15792 6802
rect 15750 6760 15806 6769
rect 15750 6695 15806 6704
rect 15936 6656 15988 6662
rect 15936 6598 15988 6604
rect 15948 6361 15976 6598
rect 15934 6352 15990 6361
rect 15384 6316 15436 6322
rect 15934 6287 15990 6296
rect 15384 6258 15436 6264
rect 15384 6112 15436 6118
rect 15290 6080 15346 6089
rect 15384 6054 15436 6060
rect 15290 6015 15346 6024
rect 15198 4584 15254 4593
rect 15198 4519 15254 4528
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 14556 4072 14608 4078
rect 14924 4072 14976 4078
rect 14556 4014 14608 4020
rect 14922 4040 14924 4049
rect 14976 4040 14978 4049
rect 14280 4004 14332 4010
rect 14922 3975 14978 3984
rect 14280 3946 14332 3952
rect 14292 3890 14320 3946
rect 14464 3936 14516 3942
rect 14292 3862 14412 3890
rect 14464 3878 14516 3884
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14108 3505 14136 3674
rect 13966 3454 14044 3482
rect 14094 3496 14150 3505
rect 13910 3431 13966 3440
rect 14094 3431 14150 3440
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13832 2774 13860 2926
rect 14200 2854 14228 3674
rect 14384 3534 14412 3862
rect 14476 3602 14504 3878
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14372 3528 14424 3534
rect 14844 3505 14872 3878
rect 14372 3470 14424 3476
rect 14830 3496 14886 3505
rect 14830 3431 14886 3440
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14292 3058 14320 3334
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 15396 2854 15424 6054
rect 15578 6012 15886 6021
rect 15578 6010 15584 6012
rect 15640 6010 15664 6012
rect 15720 6010 15744 6012
rect 15800 6010 15824 6012
rect 15880 6010 15886 6012
rect 15640 5958 15642 6010
rect 15822 5958 15824 6010
rect 15578 5956 15584 5958
rect 15640 5956 15664 5958
rect 15720 5956 15744 5958
rect 15800 5956 15824 5958
rect 15880 5956 15886 5958
rect 15578 5947 15886 5956
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15948 5166 15976 5646
rect 16040 5409 16068 8774
rect 16224 8294 16252 12786
rect 16316 12238 16344 13926
rect 16500 13870 16528 14554
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16592 13530 16620 14583
rect 16776 14414 16804 14758
rect 16960 14550 16988 14991
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16776 13938 16804 14350
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 17052 13394 17080 15399
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16500 12782 16528 12922
rect 16592 12782 16620 13262
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16132 8266 16252 8294
rect 16132 7993 16160 8266
rect 16118 7984 16174 7993
rect 16316 7970 16344 11290
rect 16500 10606 16528 11630
rect 16592 11218 16620 12718
rect 16776 12374 16804 13330
rect 16764 12368 16816 12374
rect 16764 12310 16816 12316
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16776 11762 16896 11778
rect 16776 11756 16908 11762
rect 16776 11750 16856 11756
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16684 11121 16712 11494
rect 16670 11112 16726 11121
rect 16670 11047 16726 11056
rect 16578 10704 16634 10713
rect 16578 10639 16580 10648
rect 16632 10639 16634 10648
rect 16580 10610 16632 10616
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16408 9178 16436 9454
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16118 7919 16174 7928
rect 16224 7942 16344 7970
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16132 6361 16160 6598
rect 16118 6352 16174 6361
rect 16118 6287 16174 6296
rect 16224 5817 16252 7942
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16316 7002 16344 7822
rect 16408 7206 16436 8230
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16408 7002 16436 7142
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16302 6896 16358 6905
rect 16500 6866 16528 10542
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16578 10160 16634 10169
rect 16578 10095 16634 10104
rect 16592 7886 16620 10095
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16684 7410 16712 10406
rect 16776 10033 16804 11750
rect 16856 11698 16908 11704
rect 16960 11218 16988 12174
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16868 10130 16896 11018
rect 16960 11014 16988 11154
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16960 10062 16988 10950
rect 17052 10470 17080 11494
rect 17144 11336 17172 15982
rect 17236 15706 17264 15982
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17314 15600 17370 15609
rect 17314 15535 17370 15544
rect 17328 15502 17356 15535
rect 17512 15502 17540 16050
rect 18432 15978 18460 18906
rect 18524 18902 18552 19110
rect 18512 18896 18564 18902
rect 18512 18838 18564 18844
rect 18616 18290 18644 19654
rect 18708 19378 18736 20198
rect 18800 19922 18828 20266
rect 18788 19916 18840 19922
rect 18788 19858 18840 19864
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18800 19258 18828 19858
rect 18708 19230 18828 19258
rect 18708 18630 18736 19230
rect 18984 18873 19012 20896
rect 18970 18864 19026 18873
rect 18970 18799 19026 18808
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18604 18284 18656 18290
rect 18604 18226 18656 18232
rect 18708 18222 18736 18566
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 18512 16516 18564 16522
rect 18512 16458 18564 16464
rect 18524 16182 18552 16458
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18512 16176 18564 16182
rect 18512 16118 18564 16124
rect 18800 16046 18828 16390
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18420 15972 18472 15978
rect 18420 15914 18472 15920
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17512 14822 17540 15438
rect 17696 15337 17724 15438
rect 17682 15328 17738 15337
rect 17682 15263 17738 15272
rect 17788 14929 17816 15642
rect 18142 15600 18198 15609
rect 18142 15535 18144 15544
rect 18196 15535 18198 15544
rect 18144 15506 18196 15512
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17774 14920 17830 14929
rect 17774 14855 17830 14864
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17498 14512 17554 14521
rect 17498 14447 17554 14456
rect 17512 14414 17540 14447
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 17512 13530 17540 13806
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17590 13424 17646 13433
rect 17590 13359 17646 13368
rect 17684 13388 17736 13394
rect 17604 12986 17632 13359
rect 17684 13330 17736 13336
rect 17696 13190 17724 13330
rect 17880 13258 17908 15438
rect 18800 15026 18828 15846
rect 18892 15434 18920 16390
rect 19076 15502 19104 21558
rect 19260 21554 19288 21830
rect 19373 21788 19681 21797
rect 19373 21786 19379 21788
rect 19435 21786 19459 21788
rect 19515 21786 19539 21788
rect 19595 21786 19619 21788
rect 19675 21786 19681 21788
rect 19435 21734 19437 21786
rect 19617 21734 19619 21786
rect 19373 21732 19379 21734
rect 19435 21732 19459 21734
rect 19515 21732 19539 21734
rect 19595 21732 19619 21734
rect 19675 21732 19681 21734
rect 19373 21723 19681 21732
rect 19720 21672 19748 22034
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19628 21644 19748 21672
rect 19628 21554 19656 21644
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19616 21548 19668 21554
rect 19616 21490 19668 21496
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19260 20466 19288 20878
rect 19373 20700 19681 20709
rect 19373 20698 19379 20700
rect 19435 20698 19459 20700
rect 19515 20698 19539 20700
rect 19595 20698 19619 20700
rect 19675 20698 19681 20700
rect 19435 20646 19437 20698
rect 19617 20646 19619 20698
rect 19373 20644 19379 20646
rect 19435 20644 19459 20646
rect 19515 20644 19539 20646
rect 19595 20644 19619 20646
rect 19675 20644 19681 20646
rect 19373 20635 19681 20644
rect 19904 20641 19932 21966
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 20364 21729 20392 21898
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20350 21720 20406 21729
rect 20350 21655 20406 21664
rect 20548 21350 20576 21830
rect 21100 21690 21128 22034
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 21456 21956 21508 21962
rect 21456 21898 21508 21904
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 21468 21554 21496 21898
rect 22376 21684 22428 21690
rect 22376 21626 22428 21632
rect 22006 21584 22062 21593
rect 21456 21548 21508 21554
rect 22006 21519 22008 21528
rect 21456 21490 21508 21496
rect 22060 21519 22062 21528
rect 22008 21490 22060 21496
rect 20720 21480 20772 21486
rect 20720 21422 20772 21428
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20628 21004 20680 21010
rect 20628 20946 20680 20952
rect 19890 20632 19946 20641
rect 19890 20567 19946 20576
rect 19248 20460 19300 20466
rect 19248 20402 19300 20408
rect 20640 20398 20668 20946
rect 20628 20392 20680 20398
rect 20628 20334 20680 20340
rect 20628 19916 20680 19922
rect 20628 19858 20680 19864
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 19800 19712 19852 19718
rect 19800 19654 19852 19660
rect 19373 19612 19681 19621
rect 19373 19610 19379 19612
rect 19435 19610 19459 19612
rect 19515 19610 19539 19612
rect 19595 19610 19619 19612
rect 19675 19610 19681 19612
rect 19435 19558 19437 19610
rect 19617 19558 19619 19610
rect 19373 19556 19379 19558
rect 19435 19556 19459 19558
rect 19515 19556 19539 19558
rect 19595 19556 19619 19558
rect 19675 19556 19681 19558
rect 19373 19547 19681 19556
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 18880 15428 18932 15434
rect 18880 15370 18932 15376
rect 18972 15360 19024 15366
rect 18878 15328 18934 15337
rect 18934 15308 18972 15314
rect 18934 15302 19024 15308
rect 18934 15286 19012 15302
rect 18878 15263 18934 15272
rect 19168 15094 19196 15846
rect 19156 15088 19208 15094
rect 19156 15030 19208 15036
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 19260 14958 19288 19246
rect 19373 18524 19681 18533
rect 19373 18522 19379 18524
rect 19435 18522 19459 18524
rect 19515 18522 19539 18524
rect 19595 18522 19619 18524
rect 19675 18522 19681 18524
rect 19435 18470 19437 18522
rect 19617 18470 19619 18522
rect 19373 18468 19379 18470
rect 19435 18468 19459 18470
rect 19515 18468 19539 18470
rect 19595 18468 19619 18470
rect 19675 18468 19681 18470
rect 19373 18459 19681 18468
rect 19812 17746 19840 19654
rect 20088 19514 20116 19790
rect 20444 19712 20496 19718
rect 20444 19654 20496 19660
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 20456 19310 20484 19654
rect 20640 19514 20668 19858
rect 20732 19786 20760 21422
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21284 21146 21312 21286
rect 22204 21146 22232 21422
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 21180 20936 21232 20942
rect 21180 20878 21232 20884
rect 21192 20466 21220 20878
rect 22296 20754 22324 21422
rect 22020 20726 22324 20754
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 20720 19780 20772 19786
rect 20720 19722 20772 19728
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 20456 18834 20484 19246
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20364 18358 20392 18702
rect 20456 18698 20484 18770
rect 20444 18692 20496 18698
rect 20444 18634 20496 18640
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 19982 17776 20038 17785
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19904 17734 19982 17762
rect 19373 17436 19681 17445
rect 19373 17434 19379 17436
rect 19435 17434 19459 17436
rect 19515 17434 19539 17436
rect 19595 17434 19619 17436
rect 19675 17434 19681 17436
rect 19435 17382 19437 17434
rect 19617 17382 19619 17434
rect 19373 17380 19379 17382
rect 19435 17380 19459 17382
rect 19515 17380 19539 17382
rect 19595 17380 19619 17382
rect 19675 17380 19681 17382
rect 19373 17371 19681 17380
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19522 16960 19578 16969
rect 19444 16590 19472 16934
rect 19522 16895 19578 16904
rect 19536 16658 19564 16895
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19373 16348 19681 16357
rect 19373 16346 19379 16348
rect 19435 16346 19459 16348
rect 19515 16346 19539 16348
rect 19595 16346 19619 16348
rect 19675 16346 19681 16348
rect 19435 16294 19437 16346
rect 19617 16294 19619 16346
rect 19373 16292 19379 16294
rect 19435 16292 19459 16294
rect 19515 16292 19539 16294
rect 19595 16292 19619 16294
rect 19675 16292 19681 16294
rect 19373 16283 19681 16292
rect 19432 15564 19484 15570
rect 19484 15524 19840 15552
rect 19432 15506 19484 15512
rect 19373 15260 19681 15269
rect 19373 15258 19379 15260
rect 19435 15258 19459 15260
rect 19515 15258 19539 15260
rect 19595 15258 19619 15260
rect 19675 15258 19681 15260
rect 19435 15206 19437 15258
rect 19617 15206 19619 15258
rect 19373 15204 19379 15206
rect 19435 15204 19459 15206
rect 19515 15204 19539 15206
rect 19595 15204 19619 15206
rect 19675 15204 19681 15206
rect 19373 15195 19681 15204
rect 19812 15201 19840 15524
rect 19798 15192 19854 15201
rect 19798 15127 19854 15136
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 19800 14952 19852 14958
rect 19800 14894 19852 14900
rect 17972 14074 18000 14894
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18880 13864 18932 13870
rect 19156 13864 19208 13870
rect 18880 13806 18932 13812
rect 19154 13832 19156 13841
rect 19208 13832 19210 13841
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18156 13394 18184 13670
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17316 12232 17368 12238
rect 17696 12209 17724 13126
rect 18340 12850 18368 13262
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 18052 12232 18104 12238
rect 17316 12174 17368 12180
rect 17682 12200 17738 12209
rect 17224 11348 17276 11354
rect 17144 11308 17224 11336
rect 17224 11290 17276 11296
rect 17328 11150 17356 12174
rect 18052 12174 18104 12180
rect 17682 12135 17738 12144
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 16948 10056 17000 10062
rect 16762 10024 16818 10033
rect 16948 9998 17000 10004
rect 16762 9959 16818 9968
rect 16764 9920 16816 9926
rect 16816 9880 16896 9908
rect 16764 9862 16816 9868
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16302 6831 16304 6840
rect 16356 6831 16358 6840
rect 16488 6860 16540 6866
rect 16304 6802 16356 6808
rect 16488 6802 16540 6808
rect 16500 6769 16528 6802
rect 16776 6798 16804 9658
rect 16868 9042 16896 9880
rect 17052 9722 17080 10406
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 17052 9178 17080 9318
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 16764 6792 16816 6798
rect 16486 6760 16542 6769
rect 16764 6734 16816 6740
rect 16486 6695 16542 6704
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16210 5808 16266 5817
rect 16684 5778 16712 6122
rect 16776 6100 16804 6734
rect 16868 6254 16896 8978
rect 17040 7404 17092 7410
rect 17144 7392 17172 11086
rect 17328 10656 17356 11086
rect 17500 10668 17552 10674
rect 17328 10628 17500 10656
rect 17500 10610 17552 10616
rect 17512 10266 17540 10610
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17092 7364 17172 7392
rect 17040 7346 17092 7352
rect 17052 6633 17080 7346
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17038 6624 17094 6633
rect 17038 6559 17094 6568
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16776 6072 16896 6100
rect 16210 5743 16266 5752
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16026 5400 16082 5409
rect 16592 5370 16620 5646
rect 16026 5335 16082 5344
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 15578 4924 15886 4933
rect 15578 4922 15584 4924
rect 15640 4922 15664 4924
rect 15720 4922 15744 4924
rect 15800 4922 15824 4924
rect 15880 4922 15886 4924
rect 15640 4870 15642 4922
rect 15822 4870 15824 4922
rect 15578 4868 15584 4870
rect 15640 4868 15664 4870
rect 15720 4868 15744 4870
rect 15800 4868 15824 4870
rect 15880 4868 15886 4870
rect 15578 4859 15886 4868
rect 15948 4604 15976 5102
rect 16132 4758 16160 5170
rect 16684 5030 16712 5714
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 16120 4616 16172 4622
rect 15948 4576 16120 4604
rect 16120 4558 16172 4564
rect 16488 4616 16540 4622
rect 16684 4604 16712 4966
rect 16776 4690 16804 5510
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16540 4576 16712 4604
rect 16488 4558 16540 4564
rect 15578 3836 15886 3845
rect 15578 3834 15584 3836
rect 15640 3834 15664 3836
rect 15720 3834 15744 3836
rect 15800 3834 15824 3836
rect 15880 3834 15886 3836
rect 15640 3782 15642 3834
rect 15822 3782 15824 3834
rect 15578 3780 15584 3782
rect 15640 3780 15664 3782
rect 15720 3780 15744 3782
rect 15800 3780 15824 3782
rect 15880 3780 15886 3782
rect 15578 3771 15886 3780
rect 16132 3534 16160 4558
rect 16302 4448 16358 4457
rect 16302 4383 16358 4392
rect 16316 4282 16344 4383
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16120 3528 16172 3534
rect 16040 3488 16120 3516
rect 16040 2990 16068 3488
rect 16120 3470 16172 3476
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 13740 2746 13860 2774
rect 11992 2604 12204 2632
rect 12254 2680 12310 2689
rect 13740 2650 13768 2746
rect 14200 2650 14228 2790
rect 12254 2615 12310 2624
rect 12440 2644 12492 2650
rect 11888 2508 11940 2514
rect 11888 2450 11940 2456
rect 11796 2440 11848 2446
rect 11900 2417 11928 2450
rect 11796 2382 11848 2388
rect 11886 2408 11942 2417
rect 11886 2343 11942 2352
rect 11992 2310 12020 2604
rect 12440 2586 12492 2592
rect 13728 2644 13780 2650
rect 14188 2644 14240 2650
rect 13728 2586 13780 2592
rect 14016 2604 14188 2632
rect 12164 2440 12216 2446
rect 12452 2417 12480 2586
rect 13740 2446 13768 2586
rect 13728 2440 13780 2446
rect 12164 2382 12216 2388
rect 12438 2408 12494 2417
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11783 2204 12091 2213
rect 11783 2202 11789 2204
rect 11845 2202 11869 2204
rect 11925 2202 11949 2204
rect 12005 2202 12029 2204
rect 12085 2202 12091 2204
rect 11845 2150 11847 2202
rect 12027 2150 12029 2202
rect 11783 2148 11789 2150
rect 11845 2148 11869 2150
rect 11925 2148 11949 2150
rect 12005 2148 12029 2150
rect 12085 2148 12091 2150
rect 11783 2139 12091 2148
rect 11980 2100 12032 2106
rect 11980 2042 12032 2048
rect 12072 2100 12124 2106
rect 12072 2042 12124 2048
rect 11992 1970 12020 2042
rect 11796 1964 11848 1970
rect 11716 1924 11796 1952
rect 11716 1562 11744 1924
rect 11796 1906 11848 1912
rect 11980 1964 12032 1970
rect 11980 1906 12032 1912
rect 12084 1766 12112 2042
rect 12072 1760 12124 1766
rect 12072 1702 12124 1708
rect 11704 1556 11756 1562
rect 11704 1498 11756 1504
rect 12176 1442 12204 2382
rect 13648 2388 13728 2394
rect 13648 2382 13780 2388
rect 12438 2343 12494 2352
rect 13176 2372 13228 2378
rect 13176 2314 13228 2320
rect 13648 2366 13768 2382
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12256 1556 12308 1562
rect 12256 1498 12308 1504
rect 11520 1420 11572 1426
rect 11520 1362 11572 1368
rect 11612 1420 11664 1426
rect 11612 1362 11664 1368
rect 11716 1414 12204 1442
rect 12268 1426 12296 1498
rect 12256 1420 12308 1426
rect 11426 1048 11482 1057
rect 11426 983 11482 992
rect 11152 808 11204 814
rect 11716 762 11744 1414
rect 12256 1362 12308 1368
rect 12164 1352 12216 1358
rect 12164 1294 12216 1300
rect 11783 1116 12091 1125
rect 11783 1114 11789 1116
rect 11845 1114 11869 1116
rect 11925 1114 11949 1116
rect 12005 1114 12029 1116
rect 12085 1114 12091 1116
rect 11845 1062 11847 1114
rect 12027 1062 12029 1114
rect 11783 1060 11789 1062
rect 11845 1060 11869 1062
rect 11925 1060 11949 1062
rect 12005 1060 12029 1062
rect 12085 1060 12091 1062
rect 11783 1051 12091 1060
rect 11794 912 11850 921
rect 11794 847 11796 856
rect 11848 847 11850 856
rect 11796 818 11848 824
rect 11152 750 11204 756
rect 11624 734 11744 762
rect 11888 808 11940 814
rect 12176 762 12204 1294
rect 12360 1222 12388 2246
rect 13188 2106 13216 2314
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 13648 1970 13676 2366
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13636 1964 13688 1970
rect 13636 1906 13688 1912
rect 13648 1850 13676 1906
rect 13556 1822 13676 1850
rect 13556 1426 13584 1822
rect 13636 1760 13688 1766
rect 13636 1702 13688 1708
rect 13648 1562 13676 1702
rect 13636 1556 13688 1562
rect 13636 1498 13688 1504
rect 13544 1420 13596 1426
rect 13544 1362 13596 1368
rect 13740 1340 13768 2246
rect 14016 1970 14044 2604
rect 14188 2586 14240 2592
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14108 2106 14136 2382
rect 14096 2100 14148 2106
rect 14096 2042 14148 2048
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 14004 1964 14056 1970
rect 14004 1906 14056 1912
rect 14016 1578 14044 1906
rect 14372 1896 14424 1902
rect 14372 1838 14424 1844
rect 14016 1562 14136 1578
rect 14016 1556 14148 1562
rect 14016 1550 14096 1556
rect 14096 1498 14148 1504
rect 14004 1352 14056 1358
rect 13740 1312 14004 1340
rect 14004 1294 14056 1300
rect 12348 1216 12400 1222
rect 12348 1158 12400 1164
rect 14280 1216 14332 1222
rect 14280 1158 14332 1164
rect 14292 882 14320 1158
rect 14384 1018 14412 1838
rect 14372 1012 14424 1018
rect 14372 954 14424 960
rect 13636 876 13688 882
rect 13636 818 13688 824
rect 14280 876 14332 882
rect 14280 818 14332 824
rect 11940 756 12204 762
rect 11888 750 12204 756
rect 12992 808 13044 814
rect 12992 750 13044 756
rect 11900 734 12204 750
rect 11624 678 11652 734
rect 11612 672 11664 678
rect 11612 614 11664 620
rect 8576 400 8628 406
rect 8576 342 8628 348
rect 10784 400 10836 406
rect 10784 342 10836 348
rect 10796 270 10824 342
rect 13004 338 13032 750
rect 13084 672 13136 678
rect 13084 614 13136 620
rect 13096 338 13124 614
rect 13648 406 13676 818
rect 14568 814 14596 2042
rect 15396 814 15424 2790
rect 15578 2748 15886 2757
rect 15578 2746 15584 2748
rect 15640 2746 15664 2748
rect 15720 2746 15744 2748
rect 15800 2746 15824 2748
rect 15880 2746 15886 2748
rect 15640 2694 15642 2746
rect 15822 2694 15824 2746
rect 15578 2692 15584 2694
rect 15640 2692 15664 2694
rect 15720 2692 15744 2694
rect 15800 2692 15824 2694
rect 15880 2692 15886 2694
rect 15578 2683 15886 2692
rect 16040 2446 16068 2926
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 16040 1986 16068 2382
rect 15948 1958 16068 1986
rect 15948 1902 15976 1958
rect 15936 1896 15988 1902
rect 15936 1838 15988 1844
rect 15578 1660 15886 1669
rect 15578 1658 15584 1660
rect 15640 1658 15664 1660
rect 15720 1658 15744 1660
rect 15800 1658 15824 1660
rect 15880 1658 15886 1660
rect 15640 1606 15642 1658
rect 15822 1606 15824 1658
rect 15578 1604 15584 1606
rect 15640 1604 15664 1606
rect 15720 1604 15744 1606
rect 15800 1604 15824 1606
rect 15880 1604 15886 1606
rect 15578 1595 15886 1604
rect 16040 1358 16068 1958
rect 16028 1352 16080 1358
rect 16028 1294 16080 1300
rect 13820 808 13872 814
rect 13820 750 13872 756
rect 14556 808 14608 814
rect 14556 750 14608 756
rect 15384 808 15436 814
rect 15384 750 15436 756
rect 13636 400 13688 406
rect 13636 342 13688 348
rect 12992 332 13044 338
rect 12992 274 13044 280
rect 13084 332 13136 338
rect 13084 274 13136 280
rect 7656 264 7708 270
rect 7656 206 7708 212
rect 10784 264 10836 270
rect 10784 206 10836 212
rect 13832 202 13860 750
rect 14464 672 14516 678
rect 14464 614 14516 620
rect 14476 474 14504 614
rect 15578 572 15886 581
rect 15578 570 15584 572
rect 15640 570 15664 572
rect 15720 570 15744 572
rect 15800 570 15824 572
rect 15880 570 15886 572
rect 15640 518 15642 570
rect 15822 518 15824 570
rect 15578 516 15584 518
rect 15640 516 15664 518
rect 15720 516 15744 518
rect 15800 516 15824 518
rect 15880 516 15886 518
rect 15578 507 15886 516
rect 14464 468 14516 474
rect 14464 410 14516 416
rect 13820 196 13872 202
rect 13820 138 13872 144
rect 16224 66 16252 4014
rect 16592 3738 16620 4576
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16592 2854 16620 3674
rect 16304 2848 16356 2854
rect 16302 2816 16304 2825
rect 16580 2848 16632 2854
rect 16356 2816 16358 2825
rect 16580 2790 16632 2796
rect 16302 2751 16358 2760
rect 16592 2650 16620 2790
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16592 1766 16620 2586
rect 16684 2310 16712 3878
rect 16776 3738 16804 4082
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16868 3618 16896 6072
rect 17144 5370 17172 6734
rect 17512 6497 17540 7822
rect 17498 6488 17554 6497
rect 17498 6423 17554 6432
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17328 5778 17356 6054
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17512 4729 17540 6423
rect 17604 5137 17632 11630
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17788 5273 17816 10542
rect 18064 9654 18092 12174
rect 18340 11694 18368 12786
rect 18708 12714 18736 13262
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18328 11688 18380 11694
rect 18328 11630 18380 11636
rect 18340 11218 18368 11630
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18328 11212 18380 11218
rect 18328 11154 18380 11160
rect 18432 11082 18460 11494
rect 18800 11354 18828 13262
rect 18892 12434 18920 13806
rect 19260 13802 19288 14894
rect 19706 14784 19762 14793
rect 19706 14719 19762 14728
rect 19614 14648 19670 14657
rect 19614 14583 19670 14592
rect 19628 14550 19656 14583
rect 19616 14544 19668 14550
rect 19616 14486 19668 14492
rect 19373 14172 19681 14181
rect 19373 14170 19379 14172
rect 19435 14170 19459 14172
rect 19515 14170 19539 14172
rect 19595 14170 19619 14172
rect 19675 14170 19681 14172
rect 19435 14118 19437 14170
rect 19617 14118 19619 14170
rect 19373 14116 19379 14118
rect 19435 14116 19459 14118
rect 19515 14116 19539 14118
rect 19595 14116 19619 14118
rect 19675 14116 19681 14118
rect 19373 14107 19681 14116
rect 19524 14000 19576 14006
rect 19522 13968 19524 13977
rect 19576 13968 19578 13977
rect 19522 13903 19578 13912
rect 19154 13767 19210 13776
rect 19248 13796 19300 13802
rect 19248 13738 19300 13744
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 18970 12472 19026 12481
rect 18892 12416 18970 12434
rect 19076 12442 19104 12786
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19168 12442 19196 12582
rect 18892 12407 19026 12416
rect 19064 12436 19116 12442
rect 18892 12406 19012 12407
rect 18892 11898 18920 12406
rect 19064 12378 19116 12384
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19156 12300 19208 12306
rect 19260 12288 19288 13738
rect 19720 13734 19748 14719
rect 19812 13870 19840 14894
rect 19904 14618 19932 17734
rect 19982 17711 20038 17720
rect 20364 17066 20392 18158
rect 20456 17678 20484 18634
rect 20536 17808 20588 17814
rect 20536 17750 20588 17756
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20548 17270 20576 17750
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20640 16590 20668 19450
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 21376 19334 21404 20538
rect 21560 19922 21588 20538
rect 22020 20262 22048 20726
rect 22008 20256 22060 20262
rect 22008 20198 22060 20204
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 21548 19916 21600 19922
rect 21548 19858 21600 19864
rect 22100 19712 22152 19718
rect 22006 19680 22062 19689
rect 21928 19638 22006 19666
rect 21928 19378 21956 19638
rect 22100 19654 22152 19660
rect 22006 19615 22062 19624
rect 22112 19378 22140 19654
rect 22204 19446 22232 19994
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 21916 19372 21968 19378
rect 20732 18970 20760 19314
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20720 18624 20772 18630
rect 20720 18566 20772 18572
rect 20732 17202 20760 18566
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 20916 17746 20944 18158
rect 21100 17814 21128 19314
rect 21376 19306 21496 19334
rect 21916 19314 21968 19320
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 21178 18320 21234 18329
rect 21178 18255 21234 18264
rect 21272 18284 21324 18290
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 20812 17536 20864 17542
rect 20812 17478 20864 17484
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20824 16794 20852 17478
rect 21100 16980 21128 17614
rect 21192 17202 21220 18255
rect 21272 18226 21324 18232
rect 21284 17785 21312 18226
rect 21270 17776 21326 17785
rect 21270 17711 21326 17720
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 21284 17116 21312 17614
rect 21364 17128 21416 17134
rect 21284 17088 21364 17116
rect 21180 16992 21232 16998
rect 21100 16952 21180 16980
rect 21180 16934 21232 16940
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20534 16416 20590 16425
rect 20534 16351 20590 16360
rect 20548 16250 20576 16351
rect 20536 16244 20588 16250
rect 20536 16186 20588 16192
rect 20732 16182 20760 16662
rect 21192 16590 21220 16934
rect 21284 16590 21312 17088
rect 21364 17070 21416 17076
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 21272 16584 21324 16590
rect 21468 16572 21496 19306
rect 22388 19242 22416 21626
rect 22480 21554 22508 21966
rect 23664 21956 23716 21962
rect 23664 21898 23716 21904
rect 23572 21888 23624 21894
rect 23570 21856 23572 21865
rect 23624 21856 23626 21865
rect 23570 21791 23626 21800
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 23584 21486 23612 21791
rect 23204 21480 23256 21486
rect 23202 21448 23204 21457
rect 23572 21480 23624 21486
rect 23256 21448 23258 21457
rect 23572 21422 23624 21428
rect 23202 21383 23258 21392
rect 22744 21344 22796 21350
rect 22928 21344 22980 21350
rect 22796 21292 22876 21298
rect 22744 21286 22876 21292
rect 22928 21286 22980 21292
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 22756 21270 22876 21286
rect 22848 21078 22876 21270
rect 22836 21072 22888 21078
rect 22836 21014 22888 21020
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22558 20360 22614 20369
rect 22558 20295 22614 20304
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22480 19854 22508 20198
rect 22468 19848 22520 19854
rect 22468 19790 22520 19796
rect 22468 19712 22520 19718
rect 22466 19680 22468 19689
rect 22520 19680 22522 19689
rect 22466 19615 22522 19624
rect 22376 19236 22428 19242
rect 22376 19178 22428 19184
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 21652 18834 21680 19110
rect 22572 18902 22600 20295
rect 22560 18896 22612 18902
rect 22560 18838 22612 18844
rect 21640 18828 21692 18834
rect 21640 18770 21692 18776
rect 22190 18456 22246 18465
rect 22664 18426 22692 20742
rect 22756 19990 22784 20742
rect 22836 20052 22888 20058
rect 22836 19994 22888 20000
rect 22744 19984 22796 19990
rect 22744 19926 22796 19932
rect 22744 19236 22796 19242
rect 22744 19178 22796 19184
rect 22756 18698 22784 19178
rect 22744 18692 22796 18698
rect 22744 18634 22796 18640
rect 22190 18391 22246 18400
rect 22560 18420 22612 18426
rect 22204 18086 22232 18391
rect 22560 18362 22612 18368
rect 22652 18420 22704 18426
rect 22652 18362 22704 18368
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22100 16992 22152 16998
rect 22098 16960 22100 16969
rect 22152 16960 22154 16969
rect 22098 16895 22154 16904
rect 21546 16688 21602 16697
rect 21602 16646 21680 16674
rect 21546 16623 21602 16632
rect 21468 16544 21588 16572
rect 21272 16526 21324 16532
rect 20720 16176 20772 16182
rect 20720 16118 20772 16124
rect 21192 15978 21220 16526
rect 21180 15972 21232 15978
rect 21180 15914 21232 15920
rect 20812 15904 20864 15910
rect 20810 15872 20812 15881
rect 20864 15872 20866 15881
rect 20810 15807 20866 15816
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20180 14618 20208 15438
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20732 15162 20760 15302
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20628 14952 20680 14958
rect 20442 14920 20498 14929
rect 20628 14894 20680 14900
rect 20442 14855 20498 14864
rect 20260 14816 20312 14822
rect 20260 14758 20312 14764
rect 19892 14612 19944 14618
rect 19892 14554 19944 14560
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 19892 14476 19944 14482
rect 19892 14418 19944 14424
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 19904 14113 19932 14418
rect 20180 14249 20208 14418
rect 20166 14240 20222 14249
rect 20166 14175 20222 14184
rect 19890 14104 19946 14113
rect 19890 14039 19946 14048
rect 20180 13938 20208 14175
rect 20168 13932 20220 13938
rect 19904 13892 20168 13920
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 19708 13728 19760 13734
rect 19708 13670 19760 13676
rect 19373 13084 19681 13093
rect 19373 13082 19379 13084
rect 19435 13082 19459 13084
rect 19515 13082 19539 13084
rect 19595 13082 19619 13084
rect 19675 13082 19681 13084
rect 19435 13030 19437 13082
rect 19617 13030 19619 13082
rect 19373 13028 19379 13030
rect 19435 13028 19459 13030
rect 19515 13028 19539 13030
rect 19595 13028 19619 13030
rect 19675 13028 19681 13030
rect 19373 13019 19681 13028
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19444 12442 19472 12718
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19720 12306 19748 13670
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19208 12260 19288 12288
rect 19708 12300 19760 12306
rect 19156 12242 19208 12248
rect 19708 12242 19760 12248
rect 19156 12164 19208 12170
rect 19156 12106 19208 12112
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19076 11762 19104 11834
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18420 11076 18472 11082
rect 18420 11018 18472 11024
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 18064 9178 18092 9386
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 18064 9042 18092 9114
rect 18156 9042 18184 9862
rect 18340 9518 18368 10406
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 18052 9036 18104 9042
rect 18052 8978 18104 8984
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18524 8945 18552 10474
rect 18984 10198 19012 11630
rect 19168 11558 19196 12106
rect 19373 11996 19681 12005
rect 19373 11994 19379 11996
rect 19435 11994 19459 11996
rect 19515 11994 19539 11996
rect 19595 11994 19619 11996
rect 19675 11994 19681 11996
rect 19435 11942 19437 11994
rect 19617 11942 19619 11994
rect 19373 11940 19379 11942
rect 19435 11940 19459 11942
rect 19515 11940 19539 11942
rect 19595 11940 19619 11942
rect 19675 11940 19681 11942
rect 19373 11931 19681 11940
rect 19812 11762 19840 12922
rect 19904 12306 19932 13892
rect 20168 13874 20220 13880
rect 20272 13734 20300 14758
rect 20456 13938 20484 14855
rect 20640 14550 20668 14894
rect 21192 14822 21220 15914
rect 21284 15570 21312 16526
rect 21456 16040 21508 16046
rect 21456 15982 21508 15988
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21192 14618 21220 14758
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 20628 14544 20680 14550
rect 20628 14486 20680 14492
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 20548 13410 20576 14418
rect 21284 14414 21312 15506
rect 21376 15473 21404 15506
rect 21362 15464 21418 15473
rect 21362 15399 21418 15408
rect 21364 15088 21416 15094
rect 21364 15030 21416 15036
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20732 13938 20760 14214
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20626 13832 20682 13841
rect 20626 13767 20682 13776
rect 20640 13530 20668 13767
rect 20824 13530 20852 14350
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20916 13870 20944 14214
rect 21008 13938 21036 14282
rect 21376 14090 21404 15030
rect 21468 14278 21496 15982
rect 21560 14498 21588 16544
rect 21652 15586 21680 16646
rect 21914 16280 21970 16289
rect 22388 16250 22416 18022
rect 22572 17066 22600 18362
rect 22848 18358 22876 19994
rect 22940 19242 22968 21286
rect 22928 19236 22980 19242
rect 22928 19178 22980 19184
rect 22926 19136 22982 19145
rect 22926 19071 22982 19080
rect 22940 18850 22968 19071
rect 23032 18970 23060 21286
rect 23168 21244 23476 21253
rect 23168 21242 23174 21244
rect 23230 21242 23254 21244
rect 23310 21242 23334 21244
rect 23390 21242 23414 21244
rect 23470 21242 23476 21244
rect 23230 21190 23232 21242
rect 23412 21190 23414 21242
rect 23168 21188 23174 21190
rect 23230 21188 23254 21190
rect 23310 21188 23334 21190
rect 23390 21188 23414 21190
rect 23470 21188 23476 21190
rect 23168 21179 23476 21188
rect 23112 21004 23164 21010
rect 23112 20946 23164 20952
rect 23124 20534 23152 20946
rect 23112 20528 23164 20534
rect 23112 20470 23164 20476
rect 23124 20330 23152 20470
rect 23112 20324 23164 20330
rect 23112 20266 23164 20272
rect 23480 20324 23532 20330
rect 23532 20284 23612 20312
rect 23480 20266 23532 20272
rect 23168 20156 23476 20165
rect 23168 20154 23174 20156
rect 23230 20154 23254 20156
rect 23310 20154 23334 20156
rect 23390 20154 23414 20156
rect 23470 20154 23476 20156
rect 23230 20102 23232 20154
rect 23412 20102 23414 20154
rect 23168 20100 23174 20102
rect 23230 20100 23254 20102
rect 23310 20100 23334 20102
rect 23390 20100 23414 20102
rect 23470 20100 23476 20102
rect 23168 20091 23476 20100
rect 23110 19952 23166 19961
rect 23584 19922 23612 20284
rect 23110 19887 23166 19896
rect 23572 19916 23624 19922
rect 23124 19854 23152 19887
rect 23572 19858 23624 19864
rect 23112 19848 23164 19854
rect 23112 19790 23164 19796
rect 23676 19446 23704 21898
rect 23664 19440 23716 19446
rect 23664 19382 23716 19388
rect 23572 19304 23624 19310
rect 23572 19246 23624 19252
rect 23168 19068 23476 19077
rect 23168 19066 23174 19068
rect 23230 19066 23254 19068
rect 23310 19066 23334 19068
rect 23390 19066 23414 19068
rect 23470 19066 23476 19068
rect 23230 19014 23232 19066
rect 23412 19014 23414 19066
rect 23168 19012 23174 19014
rect 23230 19012 23254 19014
rect 23310 19012 23334 19014
rect 23390 19012 23414 19014
rect 23470 19012 23476 19014
rect 23168 19003 23476 19012
rect 23020 18964 23072 18970
rect 23020 18906 23072 18912
rect 23478 18864 23534 18873
rect 22940 18822 23060 18850
rect 22928 18624 22980 18630
rect 22928 18566 22980 18572
rect 22836 18352 22888 18358
rect 22836 18294 22888 18300
rect 22940 17678 22968 18566
rect 23032 18057 23060 18822
rect 23478 18799 23534 18808
rect 23492 18698 23520 18799
rect 23480 18692 23532 18698
rect 23480 18634 23532 18640
rect 23018 18048 23074 18057
rect 23018 17983 23074 17992
rect 22928 17672 22980 17678
rect 22928 17614 22980 17620
rect 23032 17626 23060 17983
rect 23168 17980 23476 17989
rect 23168 17978 23174 17980
rect 23230 17978 23254 17980
rect 23310 17978 23334 17980
rect 23390 17978 23414 17980
rect 23470 17978 23476 17980
rect 23230 17926 23232 17978
rect 23412 17926 23414 17978
rect 23168 17924 23174 17926
rect 23230 17924 23254 17926
rect 23310 17924 23334 17926
rect 23390 17924 23414 17926
rect 23470 17924 23476 17926
rect 23168 17915 23476 17924
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23032 17598 23244 17626
rect 23020 17536 23072 17542
rect 23020 17478 23072 17484
rect 23112 17536 23164 17542
rect 23112 17478 23164 17484
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22560 17060 22612 17066
rect 22560 17002 22612 17008
rect 22756 16794 22784 17138
rect 22926 17096 22982 17105
rect 22926 17031 22982 17040
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 21914 16215 21970 16224
rect 22376 16244 22428 16250
rect 21928 16114 21956 16215
rect 22376 16186 22428 16192
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 21822 15872 21878 15881
rect 21822 15807 21878 15816
rect 21836 15706 21864 15807
rect 21824 15700 21876 15706
rect 21824 15642 21876 15648
rect 22020 15609 22048 16050
rect 22006 15600 22062 15609
rect 21652 15558 21772 15586
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21652 14618 21680 15438
rect 21640 14612 21692 14618
rect 21640 14554 21692 14560
rect 21560 14470 21680 14498
rect 21456 14272 21508 14278
rect 21456 14214 21508 14220
rect 21100 14062 21404 14090
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 20904 13864 20956 13870
rect 20904 13806 20956 13812
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20548 13394 20944 13410
rect 20536 13388 20956 13394
rect 20588 13382 20904 13388
rect 20536 13330 20588 13336
rect 20904 13330 20956 13336
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19996 12442 20024 13262
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 20364 12850 20392 13126
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20548 12442 20576 13330
rect 21008 13326 21036 13874
rect 21100 13530 21128 14062
rect 21180 13728 21232 13734
rect 21180 13670 21232 13676
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 20732 12782 20760 13262
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20628 12708 20680 12714
rect 20628 12650 20680 12656
rect 20640 12442 20668 12650
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 19892 12300 19944 12306
rect 19892 12242 19944 12248
rect 20732 11762 20760 12582
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20916 11694 20944 12718
rect 21192 12481 21220 13670
rect 21548 13252 21600 13258
rect 21548 13194 21600 13200
rect 21272 13184 21324 13190
rect 21270 13152 21272 13161
rect 21324 13152 21326 13161
rect 21270 13087 21326 13096
rect 21178 12472 21234 12481
rect 21284 12442 21312 13087
rect 21560 12850 21588 13194
rect 21548 12844 21600 12850
rect 21548 12786 21600 12792
rect 21652 12730 21680 14470
rect 21744 14074 21772 15558
rect 22006 15535 22062 15544
rect 22192 15360 22244 15366
rect 22192 15302 22244 15308
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 21732 14068 21784 14074
rect 21732 14010 21784 14016
rect 22204 13938 22232 15302
rect 22388 14793 22416 15302
rect 22940 15026 22968 17031
rect 23032 16726 23060 17478
rect 23124 17338 23152 17478
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23216 17134 23244 17598
rect 23308 17513 23336 17818
rect 23478 17776 23534 17785
rect 23478 17711 23480 17720
rect 23532 17711 23534 17720
rect 23480 17682 23532 17688
rect 23584 17610 23612 19246
rect 23676 18222 23704 19382
rect 23664 18216 23716 18222
rect 23664 18158 23716 18164
rect 23768 18034 23796 22102
rect 23940 21956 23992 21962
rect 23940 21898 23992 21904
rect 23952 21622 23980 21898
rect 24136 21894 24164 22238
rect 25596 22228 25648 22234
rect 25596 22170 25648 22176
rect 25412 22024 25464 22030
rect 25412 21966 25464 21972
rect 24124 21888 24176 21894
rect 24124 21830 24176 21836
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 23846 20632 23902 20641
rect 23846 20567 23902 20576
rect 23860 19334 23888 20567
rect 23952 20058 23980 21422
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 23938 19952 23994 19961
rect 23938 19887 23940 19896
rect 23992 19887 23994 19896
rect 23940 19858 23992 19864
rect 23860 19306 24072 19334
rect 24044 19242 24072 19306
rect 24032 19236 24084 19242
rect 24032 19178 24084 19184
rect 24044 19145 24072 19178
rect 24136 19174 24164 21830
rect 24214 21720 24270 21729
rect 24214 21655 24270 21664
rect 24124 19168 24176 19174
rect 24030 19136 24086 19145
rect 24124 19110 24176 19116
rect 24030 19071 24086 19080
rect 23940 18828 23992 18834
rect 23940 18770 23992 18776
rect 23848 18760 23900 18766
rect 23848 18702 23900 18708
rect 23860 18601 23888 18702
rect 23846 18592 23902 18601
rect 23846 18527 23902 18536
rect 23848 18216 23900 18222
rect 23848 18158 23900 18164
rect 23676 18006 23796 18034
rect 23572 17604 23624 17610
rect 23572 17546 23624 17552
rect 23294 17504 23350 17513
rect 23294 17439 23350 17448
rect 23388 17264 23440 17270
rect 23386 17232 23388 17241
rect 23572 17264 23624 17270
rect 23440 17232 23442 17241
rect 23572 17206 23624 17212
rect 23386 17167 23442 17176
rect 23204 17128 23256 17134
rect 23204 17070 23256 17076
rect 23168 16892 23476 16901
rect 23168 16890 23174 16892
rect 23230 16890 23254 16892
rect 23310 16890 23334 16892
rect 23390 16890 23414 16892
rect 23470 16890 23476 16892
rect 23230 16838 23232 16890
rect 23412 16838 23414 16890
rect 23168 16836 23174 16838
rect 23230 16836 23254 16838
rect 23310 16836 23334 16838
rect 23390 16836 23414 16838
rect 23470 16836 23476 16838
rect 23168 16827 23476 16836
rect 23020 16720 23072 16726
rect 23020 16662 23072 16668
rect 23478 16688 23534 16697
rect 23478 16623 23534 16632
rect 23492 16454 23520 16623
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 23020 16040 23072 16046
rect 23020 15982 23072 15988
rect 22928 15020 22980 15026
rect 22928 14962 22980 14968
rect 22374 14784 22430 14793
rect 22374 14719 22430 14728
rect 23032 14006 23060 15982
rect 23168 15804 23476 15813
rect 23168 15802 23174 15804
rect 23230 15802 23254 15804
rect 23310 15802 23334 15804
rect 23390 15802 23414 15804
rect 23470 15802 23476 15804
rect 23230 15750 23232 15802
rect 23412 15750 23414 15802
rect 23168 15748 23174 15750
rect 23230 15748 23254 15750
rect 23310 15748 23334 15750
rect 23390 15748 23414 15750
rect 23470 15748 23476 15750
rect 23168 15739 23476 15748
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23492 14804 23520 15098
rect 23584 14958 23612 17206
rect 23676 15094 23704 18006
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23768 16998 23796 17478
rect 23860 17270 23888 18158
rect 23848 17264 23900 17270
rect 23848 17206 23900 17212
rect 23756 16992 23808 16998
rect 23756 16934 23808 16940
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 23768 16658 23796 16934
rect 23860 16794 23888 16934
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23846 16688 23902 16697
rect 23756 16652 23808 16658
rect 23846 16623 23848 16632
rect 23756 16594 23808 16600
rect 23900 16623 23902 16632
rect 23848 16594 23900 16600
rect 23768 16114 23796 16594
rect 23952 16454 23980 18770
rect 24136 18222 24164 19110
rect 24124 18216 24176 18222
rect 24124 18158 24176 18164
rect 24122 17232 24178 17241
rect 24122 17167 24178 17176
rect 24136 17134 24164 17167
rect 24228 17134 24256 21655
rect 24490 21584 24546 21593
rect 25424 21554 25452 21966
rect 25504 21616 25556 21622
rect 25504 21558 25556 21564
rect 24490 21519 24492 21528
rect 24544 21519 24546 21528
rect 24584 21548 24636 21554
rect 24492 21490 24544 21496
rect 24584 21490 24636 21496
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 24596 20890 24624 21490
rect 24768 21480 24820 21486
rect 24768 21422 24820 21428
rect 24412 20862 24624 20890
rect 24412 20330 24440 20862
rect 24492 20800 24544 20806
rect 24492 20742 24544 20748
rect 24400 20324 24452 20330
rect 24400 20266 24452 20272
rect 24400 19304 24452 19310
rect 24400 19246 24452 19252
rect 24308 18760 24360 18766
rect 24308 18702 24360 18708
rect 24320 18222 24348 18702
rect 24412 18630 24440 19246
rect 24504 19174 24532 20742
rect 24780 20262 24808 21422
rect 25044 21344 25096 21350
rect 25044 21286 25096 21292
rect 25056 21078 25084 21286
rect 25134 21176 25190 21185
rect 25134 21111 25190 21120
rect 25044 21072 25096 21078
rect 25044 21014 25096 21020
rect 25148 21010 25176 21111
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 25148 20398 25176 20946
rect 25424 20913 25452 21490
rect 25410 20904 25466 20913
rect 25410 20839 25466 20848
rect 25136 20392 25188 20398
rect 25516 20369 25544 21558
rect 25608 21298 25636 22170
rect 27988 22092 28040 22098
rect 27988 22034 28040 22040
rect 25688 21888 25740 21894
rect 25688 21830 25740 21836
rect 25700 21486 25728 21830
rect 26963 21788 27271 21797
rect 26963 21786 26969 21788
rect 27025 21786 27049 21788
rect 27105 21786 27129 21788
rect 27185 21786 27209 21788
rect 27265 21786 27271 21788
rect 27025 21734 27027 21786
rect 27207 21734 27209 21786
rect 26963 21732 26969 21734
rect 27025 21732 27049 21734
rect 27105 21732 27129 21734
rect 27185 21732 27209 21734
rect 27265 21732 27271 21734
rect 25870 21720 25926 21729
rect 26963 21723 27271 21732
rect 25870 21655 25926 21664
rect 25780 21548 25832 21554
rect 25780 21490 25832 21496
rect 25688 21480 25740 21486
rect 25792 21457 25820 21490
rect 25688 21422 25740 21428
rect 25778 21448 25834 21457
rect 25778 21383 25834 21392
rect 25688 21344 25740 21350
rect 25608 21292 25688 21298
rect 25608 21286 25740 21292
rect 25608 21270 25728 21286
rect 25700 20398 25728 21270
rect 25884 21078 25912 21655
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 27436 21344 27488 21350
rect 27436 21286 27488 21292
rect 27448 21162 27476 21286
rect 27356 21134 27476 21162
rect 25872 21072 25924 21078
rect 25872 21014 25924 21020
rect 26620 20998 26924 21026
rect 26620 20466 26648 20998
rect 26896 20942 26924 20998
rect 26700 20936 26752 20942
rect 26700 20878 26752 20884
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26884 20936 26936 20942
rect 26884 20878 26936 20884
rect 26424 20460 26476 20466
rect 26424 20402 26476 20408
rect 26608 20460 26660 20466
rect 26608 20402 26660 20408
rect 25688 20392 25740 20398
rect 25136 20334 25188 20340
rect 25502 20360 25558 20369
rect 24768 20256 24820 20262
rect 24768 20198 24820 20204
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24676 19848 24728 19854
rect 24676 19790 24728 19796
rect 24688 19514 24716 19790
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 24492 19168 24544 19174
rect 24492 19110 24544 19116
rect 24400 18624 24452 18630
rect 24400 18566 24452 18572
rect 24504 18426 24532 19110
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24492 18420 24544 18426
rect 24492 18362 24544 18368
rect 24308 18216 24360 18222
rect 24308 18158 24360 18164
rect 24492 18080 24544 18086
rect 24492 18022 24544 18028
rect 24504 17921 24532 18022
rect 24490 17912 24546 17921
rect 24490 17847 24546 17856
rect 24492 17672 24544 17678
rect 24492 17614 24544 17620
rect 24124 17128 24176 17134
rect 24124 17070 24176 17076
rect 24216 17128 24268 17134
rect 24216 17070 24268 17076
rect 24228 16946 24256 17070
rect 24504 17066 24532 17614
rect 24492 17060 24544 17066
rect 24492 17002 24544 17008
rect 24044 16918 24256 16946
rect 23940 16448 23992 16454
rect 23938 16416 23940 16425
rect 23992 16416 23994 16425
rect 23938 16351 23994 16360
rect 23756 16108 23808 16114
rect 23756 16050 23808 16056
rect 23768 15502 23796 16050
rect 23848 15972 23900 15978
rect 23848 15914 23900 15920
rect 23860 15858 23888 15914
rect 24044 15858 24072 16918
rect 24504 16794 24532 17002
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 24492 16788 24544 16794
rect 24492 16730 24544 16736
rect 24124 16584 24176 16590
rect 24320 16538 24348 16730
rect 24492 16652 24544 16658
rect 24124 16526 24176 16532
rect 23860 15830 24072 15858
rect 23846 15736 23902 15745
rect 23846 15671 23902 15680
rect 23756 15496 23808 15502
rect 23756 15438 23808 15444
rect 23664 15088 23716 15094
rect 23664 15030 23716 15036
rect 23768 15026 23796 15438
rect 23860 15366 23888 15671
rect 24032 15496 24084 15502
rect 24032 15438 24084 15444
rect 24044 15366 24072 15438
rect 23848 15360 23900 15366
rect 23848 15302 23900 15308
rect 24032 15360 24084 15366
rect 24032 15302 24084 15308
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23572 14952 23624 14958
rect 23572 14894 23624 14900
rect 23492 14776 23612 14804
rect 23168 14716 23476 14725
rect 23168 14714 23174 14716
rect 23230 14714 23254 14716
rect 23310 14714 23334 14716
rect 23390 14714 23414 14716
rect 23470 14714 23476 14716
rect 23230 14662 23232 14714
rect 23412 14662 23414 14714
rect 23168 14660 23174 14662
rect 23230 14660 23254 14662
rect 23310 14660 23334 14662
rect 23390 14660 23414 14662
rect 23470 14660 23476 14662
rect 23168 14651 23476 14660
rect 23112 14612 23164 14618
rect 23112 14554 23164 14560
rect 23124 14521 23152 14554
rect 23110 14512 23166 14521
rect 23584 14482 23612 14776
rect 24030 14784 24086 14793
rect 24030 14719 24086 14728
rect 23938 14512 23994 14521
rect 23110 14447 23166 14456
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23756 14476 23808 14482
rect 24044 14482 24072 14719
rect 23938 14447 23940 14456
rect 23756 14418 23808 14424
rect 23992 14447 23994 14456
rect 24032 14476 24084 14482
rect 23940 14418 23992 14424
rect 24032 14418 24084 14424
rect 23020 14000 23072 14006
rect 23020 13942 23072 13948
rect 21824 13932 21876 13938
rect 21824 13874 21876 13880
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 21836 13394 21864 13874
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 22020 13433 22048 13806
rect 23168 13628 23476 13637
rect 23168 13626 23174 13628
rect 23230 13626 23254 13628
rect 23310 13626 23334 13628
rect 23390 13626 23414 13628
rect 23470 13626 23476 13628
rect 23230 13574 23232 13626
rect 23412 13574 23414 13626
rect 23168 13572 23174 13574
rect 23230 13572 23254 13574
rect 23310 13572 23334 13574
rect 23390 13572 23414 13574
rect 23470 13572 23476 13574
rect 23168 13563 23476 13572
rect 22006 13424 22062 13433
rect 21824 13388 21876 13394
rect 22006 13359 22062 13368
rect 21824 13330 21876 13336
rect 22284 13320 22336 13326
rect 22284 13262 22336 13268
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 21732 13252 21784 13258
rect 21732 13194 21784 13200
rect 21560 12702 21680 12730
rect 21178 12407 21234 12416
rect 21272 12436 21324 12442
rect 21192 12374 21220 12407
rect 21272 12378 21324 12384
rect 21180 12368 21232 12374
rect 21180 12310 21232 12316
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 20904 11688 20956 11694
rect 21284 11676 21312 12242
rect 21560 12209 21588 12702
rect 21640 12640 21692 12646
rect 21640 12582 21692 12588
rect 21652 12238 21680 12582
rect 21640 12232 21692 12238
rect 21546 12200 21602 12209
rect 21640 12174 21692 12180
rect 21546 12135 21602 12144
rect 21548 12096 21600 12102
rect 21548 12038 21600 12044
rect 21560 11762 21588 12038
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 20956 11648 21312 11676
rect 20904 11630 20956 11636
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 19260 11218 19288 11290
rect 19798 11248 19854 11257
rect 19248 11212 19300 11218
rect 19798 11183 19854 11192
rect 19984 11212 20036 11218
rect 19248 11154 19300 11160
rect 19373 10908 19681 10917
rect 19373 10906 19379 10908
rect 19435 10906 19459 10908
rect 19515 10906 19539 10908
rect 19595 10906 19619 10908
rect 19675 10906 19681 10908
rect 19435 10854 19437 10906
rect 19617 10854 19619 10906
rect 19373 10852 19379 10854
rect 19435 10852 19459 10854
rect 19515 10852 19539 10854
rect 19595 10852 19619 10854
rect 19675 10852 19681 10854
rect 19373 10843 19681 10852
rect 19812 10742 19840 11183
rect 19984 11154 20036 11160
rect 20628 11212 20680 11218
rect 20628 11154 20680 11160
rect 19996 11121 20024 11154
rect 20536 11144 20588 11150
rect 19982 11112 20038 11121
rect 20536 11086 20588 11092
rect 19982 11047 20038 11056
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 19800 10736 19852 10742
rect 19800 10678 19852 10684
rect 19996 10606 20024 10950
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 20352 10600 20404 10606
rect 20442 10568 20498 10577
rect 20404 10548 20442 10554
rect 20352 10542 20442 10548
rect 20364 10526 20442 10542
rect 20442 10503 20498 10512
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19156 10464 19208 10470
rect 19156 10406 19208 10412
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 18972 10192 19024 10198
rect 18972 10134 19024 10140
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18510 8936 18566 8945
rect 18510 8871 18566 8880
rect 18616 8498 18644 10066
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18800 8838 18828 9998
rect 19076 9674 19104 10406
rect 19168 10130 19196 10406
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 20456 10062 20484 10406
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 19373 9820 19681 9829
rect 19373 9818 19379 9820
rect 19435 9818 19459 9820
rect 19515 9818 19539 9820
rect 19595 9818 19619 9820
rect 19675 9818 19681 9820
rect 19435 9766 19437 9818
rect 19617 9766 19619 9818
rect 19373 9764 19379 9766
rect 19435 9764 19459 9766
rect 19515 9764 19539 9766
rect 19595 9764 19619 9766
rect 19675 9764 19681 9766
rect 19373 9755 19681 9764
rect 20456 9722 20484 9998
rect 18984 9646 19104 9674
rect 19892 9716 19944 9722
rect 19892 9658 19944 9664
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 18984 9500 19012 9646
rect 19156 9580 19208 9586
rect 19208 9540 19288 9568
rect 19156 9522 19208 9528
rect 18984 9472 19104 9500
rect 18972 8900 19024 8906
rect 18972 8842 19024 8848
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18604 8492 18656 8498
rect 18524 8452 18604 8480
rect 18050 8392 18106 8401
rect 18050 8327 18052 8336
rect 18104 8327 18106 8336
rect 18052 8298 18104 8304
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18156 7954 18184 8230
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17972 7585 18000 7686
rect 17958 7576 18014 7585
rect 17958 7511 18014 7520
rect 17960 7472 18012 7478
rect 17958 7440 17960 7449
rect 18012 7440 18014 7449
rect 17958 7375 18014 7384
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 17868 6180 17920 6186
rect 17868 6122 17920 6128
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 17774 5264 17830 5273
rect 17774 5199 17830 5208
rect 17590 5128 17646 5137
rect 17590 5063 17646 5072
rect 17498 4720 17554 4729
rect 17880 4706 17908 6122
rect 18156 5778 18184 6122
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18156 5234 18184 5510
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18052 5092 18104 5098
rect 18052 5034 18104 5040
rect 18064 4826 18092 5034
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 17880 4678 18000 4706
rect 17498 4655 17554 4664
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 16776 3590 16896 3618
rect 16776 3505 16804 3590
rect 16856 3528 16908 3534
rect 16762 3496 16818 3505
rect 16856 3470 16908 3476
rect 16762 3431 16818 3440
rect 16868 3194 16896 3470
rect 17880 3466 17908 3878
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17972 3126 18000 4678
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 18052 4140 18104 4146
rect 18156 4128 18184 4218
rect 18248 4214 18276 6734
rect 18524 6254 18552 8452
rect 18604 8434 18656 8440
rect 18984 8430 19012 8842
rect 19076 8786 19104 9472
rect 19076 8758 19196 8786
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18788 8288 18840 8294
rect 18788 8230 18840 8236
rect 18800 8090 18828 8230
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18604 7336 18656 7342
rect 18602 7304 18604 7313
rect 18656 7304 18658 7313
rect 18602 7239 18658 7248
rect 18800 7206 18828 8026
rect 18984 7750 19012 8366
rect 19168 7886 19196 8758
rect 19260 8634 19288 9540
rect 19800 9512 19852 9518
rect 19800 9454 19852 9460
rect 19373 8732 19681 8741
rect 19373 8730 19379 8732
rect 19435 8730 19459 8732
rect 19515 8730 19539 8732
rect 19595 8730 19619 8732
rect 19675 8730 19681 8732
rect 19435 8678 19437 8730
rect 19617 8678 19619 8730
rect 19373 8676 19379 8678
rect 19435 8676 19459 8678
rect 19515 8676 19539 8678
rect 19595 8676 19619 8678
rect 19675 8676 19681 8678
rect 19373 8667 19681 8676
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19260 8401 19288 8434
rect 19246 8392 19302 8401
rect 19246 8327 19302 8336
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18984 7410 19012 7686
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18800 6798 18828 7142
rect 18984 7002 19012 7346
rect 18972 6996 19024 7002
rect 18972 6938 19024 6944
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18800 6322 18828 6734
rect 19076 6458 19104 7822
rect 19373 7644 19681 7653
rect 19373 7642 19379 7644
rect 19435 7642 19459 7644
rect 19515 7642 19539 7644
rect 19595 7642 19619 7644
rect 19675 7642 19681 7644
rect 19435 7590 19437 7642
rect 19617 7590 19619 7642
rect 19373 7588 19379 7590
rect 19435 7588 19459 7590
rect 19515 7588 19539 7590
rect 19595 7588 19619 7590
rect 19675 7588 19681 7590
rect 19373 7579 19681 7588
rect 19812 7546 19840 9454
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19904 7206 19932 9658
rect 20548 9654 20576 11086
rect 20640 10130 20668 11154
rect 20720 10600 20772 10606
rect 20720 10542 20772 10548
rect 20732 10266 20760 10542
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 21100 10130 21128 11290
rect 21192 10266 21220 11494
rect 21284 11354 21312 11648
rect 21652 11558 21680 12174
rect 21744 12102 21772 13194
rect 22296 13190 22324 13262
rect 21916 13184 21968 13190
rect 21916 13126 21968 13132
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 21928 13025 21956 13126
rect 21914 13016 21970 13025
rect 21914 12951 21970 12960
rect 22572 12434 22600 13262
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23388 12912 23440 12918
rect 23388 12854 23440 12860
rect 23296 12776 23348 12782
rect 23294 12744 23296 12753
rect 23348 12744 23350 12753
rect 23294 12679 23350 12688
rect 23400 12628 23428 12854
rect 23676 12850 23704 13126
rect 23768 12918 23796 14418
rect 23848 14408 23900 14414
rect 23848 14350 23900 14356
rect 23860 13938 23888 14350
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23940 13864 23992 13870
rect 24044 13852 24072 14418
rect 24136 13977 24164 16526
rect 24228 16510 24348 16538
rect 24412 16612 24492 16640
rect 24228 16114 24256 16510
rect 24412 16114 24440 16612
rect 24492 16594 24544 16600
rect 24490 16280 24546 16289
rect 24596 16250 24624 18702
rect 24676 18216 24728 18222
rect 24676 18158 24728 18164
rect 24688 17490 24716 18158
rect 24780 17678 24808 19994
rect 25148 19922 25176 20334
rect 25688 20334 25740 20340
rect 25502 20295 25558 20304
rect 25136 19916 25188 19922
rect 25136 19858 25188 19864
rect 25596 19304 25648 19310
rect 24950 19272 25006 19281
rect 25596 19246 25648 19252
rect 24950 19207 25006 19216
rect 24964 19174 24992 19207
rect 24952 19168 25004 19174
rect 24952 19110 25004 19116
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 24964 18970 24992 19110
rect 24952 18964 25004 18970
rect 24952 18906 25004 18912
rect 25136 18080 25188 18086
rect 25136 18022 25188 18028
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24768 17536 24820 17542
rect 24688 17484 24768 17490
rect 24688 17478 24820 17484
rect 24688 17462 24808 17478
rect 24780 17134 24808 17462
rect 25148 17202 25176 18022
rect 25332 17202 25360 19110
rect 25502 18048 25558 18057
rect 25502 17983 25558 17992
rect 25136 17196 25188 17202
rect 25136 17138 25188 17144
rect 25320 17196 25372 17202
rect 25320 17138 25372 17144
rect 24676 17128 24728 17134
rect 24676 17070 24728 17076
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 24490 16215 24546 16224
rect 24584 16244 24636 16250
rect 24504 16130 24532 16215
rect 24584 16186 24636 16192
rect 24216 16108 24268 16114
rect 24216 16050 24268 16056
rect 24400 16108 24452 16114
rect 24504 16102 24624 16130
rect 24400 16050 24452 16056
rect 24228 15706 24256 16050
rect 24216 15700 24268 15706
rect 24216 15642 24268 15648
rect 24228 15026 24256 15642
rect 24308 15496 24360 15502
rect 24308 15438 24360 15444
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24122 13968 24178 13977
rect 24122 13903 24178 13912
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 23992 13824 24072 13852
rect 24124 13864 24176 13870
rect 23940 13806 23992 13812
rect 24124 13806 24176 13812
rect 23848 13524 23900 13530
rect 23848 13466 23900 13472
rect 23860 13002 23888 13466
rect 24136 13394 24164 13806
rect 24228 13462 24256 13874
rect 24216 13456 24268 13462
rect 24216 13398 24268 13404
rect 24124 13388 24176 13394
rect 24124 13330 24176 13336
rect 24320 13025 24348 15438
rect 24596 14618 24624 16102
rect 24688 16046 24716 17070
rect 25148 16998 25176 17138
rect 25136 16992 25188 16998
rect 25136 16934 25188 16940
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 25320 16448 25372 16454
rect 25320 16390 25372 16396
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 24676 16040 24728 16046
rect 24676 15982 24728 15988
rect 24584 14612 24636 14618
rect 24584 14554 24636 14560
rect 24596 13938 24624 14554
rect 24676 14272 24728 14278
rect 24676 14214 24728 14220
rect 24688 13938 24716 14214
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24596 13530 24624 13874
rect 24780 13705 24808 16050
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24766 13696 24822 13705
rect 24766 13631 24822 13640
rect 24584 13524 24636 13530
rect 24584 13466 24636 13472
rect 24306 13016 24362 13025
rect 23860 12974 24164 13002
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 23400 12600 23612 12628
rect 23168 12540 23476 12549
rect 23168 12538 23174 12540
rect 23230 12538 23254 12540
rect 23310 12538 23334 12540
rect 23390 12538 23414 12540
rect 23470 12538 23476 12540
rect 23230 12486 23232 12538
rect 23412 12486 23414 12538
rect 23168 12484 23174 12486
rect 23230 12484 23254 12486
rect 23310 12484 23334 12486
rect 23390 12484 23414 12486
rect 23470 12484 23476 12486
rect 23168 12475 23476 12484
rect 22652 12436 22704 12442
rect 22572 12406 22652 12434
rect 22652 12378 22704 12384
rect 23584 12374 23612 12600
rect 23572 12368 23624 12374
rect 23572 12310 23624 12316
rect 23676 12238 23704 12786
rect 23860 12238 23888 12974
rect 24032 12844 24084 12850
rect 23952 12804 24032 12832
rect 23952 12238 23980 12804
rect 24032 12786 24084 12792
rect 24136 12646 24164 12974
rect 24306 12951 24362 12960
rect 24216 12844 24268 12850
rect 24216 12786 24268 12792
rect 24124 12640 24176 12646
rect 24124 12582 24176 12588
rect 24136 12442 24164 12582
rect 24032 12436 24084 12442
rect 24032 12378 24084 12384
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24044 12322 24072 12378
rect 24044 12306 24164 12322
rect 24044 12300 24176 12306
rect 24044 12294 24124 12300
rect 24124 12242 24176 12248
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23848 12232 23900 12238
rect 23848 12174 23900 12180
rect 23940 12232 23992 12238
rect 23940 12174 23992 12180
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21836 11762 21864 12174
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 22100 11552 22152 11558
rect 22100 11494 22152 11500
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21364 11280 21416 11286
rect 21364 11222 21416 11228
rect 21376 10849 21404 11222
rect 22112 11014 22140 11494
rect 22296 11286 22324 11494
rect 22836 11348 22888 11354
rect 22756 11308 22836 11336
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 22466 11248 22522 11257
rect 22466 11183 22468 11192
rect 22520 11183 22522 11192
rect 22468 11154 22520 11160
rect 22376 11076 22428 11082
rect 22376 11018 22428 11024
rect 22008 11008 22060 11014
rect 22008 10950 22060 10956
rect 22100 11008 22152 11014
rect 22100 10950 22152 10956
rect 21362 10840 21418 10849
rect 21362 10775 21418 10784
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 21180 10260 21232 10266
rect 21180 10202 21232 10208
rect 21376 10198 21404 10542
rect 21732 10464 21784 10470
rect 21732 10406 21784 10412
rect 21364 10192 21416 10198
rect 21364 10134 21416 10140
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 21088 10124 21140 10130
rect 21088 10066 21140 10072
rect 21744 10062 21772 10406
rect 22020 10130 22048 10950
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 21732 10056 21784 10062
rect 21732 9998 21784 10004
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 21916 9920 21968 9926
rect 21916 9862 21968 9868
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20732 9586 20760 9862
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20824 9518 20852 9862
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20824 9110 20852 9454
rect 20812 9104 20864 9110
rect 20812 9046 20864 9052
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20180 8090 20208 8910
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20640 7954 20668 8774
rect 20732 8362 20760 8774
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20824 8090 20852 8366
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20640 7750 20668 7890
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20628 7744 20680 7750
rect 20628 7686 20680 7692
rect 20548 7546 20576 7686
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20916 7313 20944 7822
rect 21008 7342 21036 8230
rect 20996 7336 21048 7342
rect 20902 7304 20958 7313
rect 20996 7278 21048 7284
rect 20902 7239 20958 7248
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 20718 6896 20774 6905
rect 20718 6831 20720 6840
rect 20772 6831 20774 6840
rect 20720 6802 20772 6808
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 19373 6556 19681 6565
rect 19373 6554 19379 6556
rect 19435 6554 19459 6556
rect 19515 6554 19539 6556
rect 19595 6554 19619 6556
rect 19675 6554 19681 6556
rect 19435 6502 19437 6554
rect 19617 6502 19619 6554
rect 19373 6500 19379 6502
rect 19435 6500 19459 6502
rect 19515 6500 19539 6502
rect 19595 6500 19619 6502
rect 19675 6500 19681 6502
rect 19373 6491 19681 6500
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 18788 6316 18840 6322
rect 18788 6258 18840 6264
rect 18512 6248 18564 6254
rect 18340 6208 18512 6236
rect 18236 4208 18288 4214
rect 18236 4150 18288 4156
rect 18104 4100 18184 4128
rect 18052 4082 18104 4088
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 16580 1760 16632 1766
rect 16580 1702 16632 1708
rect 16592 1562 16620 1702
rect 16580 1556 16632 1562
rect 16580 1498 16632 1504
rect 16856 1352 16908 1358
rect 16856 1294 16908 1300
rect 16868 1018 16896 1294
rect 17788 1018 17816 2382
rect 17972 2106 18000 2926
rect 18236 2644 18288 2650
rect 18236 2586 18288 2592
rect 17960 2100 18012 2106
rect 17960 2042 18012 2048
rect 18248 1902 18276 2586
rect 18340 1902 18368 6208
rect 18512 6190 18564 6196
rect 20260 6248 20312 6254
rect 20260 6190 20312 6196
rect 19984 6180 20036 6186
rect 19984 6122 20036 6128
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 19064 6112 19116 6118
rect 19064 6054 19116 6060
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 18432 5166 18460 6054
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18696 5704 18748 5710
rect 18696 5646 18748 5652
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18524 5166 18552 5646
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 18616 5166 18644 5510
rect 18420 5160 18472 5166
rect 18420 5102 18472 5108
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18512 4616 18564 4622
rect 18616 4604 18644 5102
rect 18708 5030 18736 5646
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18708 4622 18736 4966
rect 18800 4826 18828 5646
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18564 4576 18644 4604
rect 18696 4616 18748 4622
rect 18512 4558 18564 4564
rect 18696 4558 18748 4564
rect 18524 4010 18552 4558
rect 18708 4146 18736 4558
rect 18984 4486 19012 6054
rect 19076 4690 19104 6054
rect 19536 5778 19564 6054
rect 19996 5846 20024 6122
rect 19984 5840 20036 5846
rect 19984 5782 20036 5788
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19373 5468 19681 5477
rect 19373 5466 19379 5468
rect 19435 5466 19459 5468
rect 19515 5466 19539 5468
rect 19595 5466 19619 5468
rect 19675 5466 19681 5468
rect 19435 5414 19437 5466
rect 19617 5414 19619 5466
rect 19373 5412 19379 5414
rect 19435 5412 19459 5414
rect 19515 5412 19539 5414
rect 19595 5412 19619 5414
rect 19675 5412 19681 5414
rect 19373 5403 19681 5412
rect 20272 5234 20300 6190
rect 20548 5914 20576 6734
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20640 5914 20668 6190
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 19064 4480 19116 4486
rect 19168 4457 19196 4558
rect 20076 4480 20128 4486
rect 19064 4422 19116 4428
rect 19154 4448 19210 4457
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18512 4004 18564 4010
rect 18512 3946 18564 3952
rect 18708 3534 18736 4082
rect 18788 4004 18840 4010
rect 18788 3946 18840 3952
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 2990 18644 3334
rect 18604 2984 18656 2990
rect 18604 2926 18656 2932
rect 18616 2774 18644 2926
rect 18708 2854 18736 3470
rect 18800 3398 18828 3946
rect 19076 3602 19104 4422
rect 20076 4422 20128 4428
rect 19154 4383 19210 4392
rect 19373 4380 19681 4389
rect 19373 4378 19379 4380
rect 19435 4378 19459 4380
rect 19515 4378 19539 4380
rect 19595 4378 19619 4380
rect 19675 4378 19681 4380
rect 19435 4326 19437 4378
rect 19617 4326 19619 4378
rect 19373 4324 19379 4326
rect 19435 4324 19459 4326
rect 19515 4324 19539 4326
rect 19595 4324 19619 4326
rect 19675 4324 19681 4326
rect 19373 4315 19681 4324
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 19064 3596 19116 3602
rect 19064 3538 19116 3544
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 19260 3194 19288 4014
rect 19708 4004 19760 4010
rect 19708 3946 19760 3952
rect 19373 3292 19681 3301
rect 19373 3290 19379 3292
rect 19435 3290 19459 3292
rect 19515 3290 19539 3292
rect 19595 3290 19619 3292
rect 19675 3290 19681 3292
rect 19435 3238 19437 3290
rect 19617 3238 19619 3290
rect 19373 3236 19379 3238
rect 19435 3236 19459 3238
rect 19515 3236 19539 3238
rect 19595 3236 19619 3238
rect 19675 3236 19681 3238
rect 19373 3227 19681 3236
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18524 2746 18644 2774
rect 18524 2446 18552 2746
rect 18708 2446 18736 2790
rect 19260 2774 19288 3130
rect 19720 3097 19748 3946
rect 19706 3088 19762 3097
rect 20088 3058 20116 4422
rect 20272 3942 20300 5170
rect 20364 4146 20392 5510
rect 20732 5370 20760 6190
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20824 5166 20852 6394
rect 20812 5160 20864 5166
rect 20732 5108 20812 5114
rect 20732 5102 20864 5108
rect 20732 5086 20852 5102
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20272 3738 20300 3878
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 19706 3023 19762 3032
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19168 2746 19288 2774
rect 20180 2774 20208 3674
rect 20456 2990 20484 4626
rect 20732 4162 20760 5086
rect 20916 5030 20944 7239
rect 21100 7002 21128 9522
rect 21468 8430 21496 9522
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21560 9178 21588 9318
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21928 8974 21956 9862
rect 22008 9512 22060 9518
rect 22008 9454 22060 9460
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21468 7886 21496 8230
rect 21652 7954 21680 8230
rect 21836 8090 21864 8910
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21456 7880 21508 7886
rect 21362 7848 21418 7857
rect 21180 7812 21232 7818
rect 21456 7822 21508 7828
rect 21362 7783 21418 7792
rect 21180 7754 21232 7760
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 21088 6656 21140 6662
rect 21088 6598 21140 6604
rect 21100 6458 21128 6598
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 21088 5568 21140 5574
rect 21088 5510 21140 5516
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20824 4826 20852 4966
rect 20916 4826 20944 4966
rect 20812 4820 20864 4826
rect 20812 4762 20864 4768
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 20548 4146 20760 4162
rect 20536 4140 20760 4146
rect 20588 4134 20760 4140
rect 20536 4082 20588 4088
rect 20732 3602 20760 4134
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20720 3188 20772 3194
rect 20640 3148 20720 3176
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 20180 2746 20300 2774
rect 19168 2514 19196 2746
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 18524 2038 18552 2382
rect 18512 2032 18564 2038
rect 18512 1974 18564 1980
rect 18236 1896 18288 1902
rect 17958 1864 18014 1873
rect 18236 1838 18288 1844
rect 18328 1896 18380 1902
rect 18328 1838 18380 1844
rect 17958 1799 17960 1808
rect 18012 1799 18014 1808
rect 17960 1770 18012 1776
rect 18524 1358 18552 1974
rect 18708 1884 18736 2382
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19260 1986 19288 2246
rect 19373 2204 19681 2213
rect 19373 2202 19379 2204
rect 19435 2202 19459 2204
rect 19515 2202 19539 2204
rect 19595 2202 19619 2204
rect 19675 2202 19681 2204
rect 19435 2150 19437 2202
rect 19617 2150 19619 2202
rect 19373 2148 19379 2150
rect 19435 2148 19459 2150
rect 19515 2148 19539 2150
rect 19595 2148 19619 2150
rect 19675 2148 19681 2150
rect 19373 2139 19681 2148
rect 19156 1964 19208 1970
rect 19076 1924 19156 1952
rect 18972 1896 19024 1902
rect 18708 1856 18972 1884
rect 18708 1562 18736 1856
rect 19076 1873 19104 1924
rect 19260 1958 19380 1986
rect 19156 1906 19208 1912
rect 18972 1838 19024 1844
rect 19062 1864 19118 1873
rect 19062 1799 19118 1808
rect 19064 1760 19116 1766
rect 19248 1760 19300 1766
rect 19116 1720 19248 1748
rect 19064 1702 19116 1708
rect 19248 1702 19300 1708
rect 18696 1556 18748 1562
rect 18696 1498 18748 1504
rect 18512 1352 18564 1358
rect 18234 1320 18290 1329
rect 18512 1294 18564 1300
rect 18878 1320 18934 1329
rect 18234 1255 18290 1264
rect 18878 1255 18934 1264
rect 16856 1012 16908 1018
rect 16856 954 16908 960
rect 17776 1012 17828 1018
rect 17776 954 17828 960
rect 18248 950 18276 1255
rect 18892 950 18920 1255
rect 19352 1204 19380 1958
rect 19432 1896 19484 1902
rect 19432 1838 19484 1844
rect 19444 1562 19472 1838
rect 19432 1556 19484 1562
rect 19432 1498 19484 1504
rect 19430 1456 19486 1465
rect 19430 1391 19486 1400
rect 19444 1222 19472 1391
rect 19260 1176 19380 1204
rect 19432 1216 19484 1222
rect 18236 944 18288 950
rect 18236 886 18288 892
rect 18880 944 18932 950
rect 18880 886 18932 892
rect 19260 898 19288 1176
rect 19432 1158 19484 1164
rect 19373 1116 19681 1125
rect 19373 1114 19379 1116
rect 19435 1114 19459 1116
rect 19515 1114 19539 1116
rect 19595 1114 19619 1116
rect 19675 1114 19681 1116
rect 19435 1062 19437 1114
rect 19617 1062 19619 1114
rect 19373 1060 19379 1062
rect 19435 1060 19459 1062
rect 19515 1060 19539 1062
rect 19595 1060 19619 1062
rect 19675 1060 19681 1062
rect 19373 1051 19681 1060
rect 17040 808 17092 814
rect 17040 750 17092 756
rect 17132 808 17184 814
rect 17132 750 17184 756
rect 16488 672 16540 678
rect 16488 614 16540 620
rect 16500 202 16528 614
rect 17052 338 17080 750
rect 17144 474 17172 750
rect 17132 468 17184 474
rect 17132 410 17184 416
rect 17040 332 17092 338
rect 17040 274 17092 280
rect 16488 196 16540 202
rect 16488 138 16540 144
rect 18892 66 18920 886
rect 19260 882 19380 898
rect 19156 876 19208 882
rect 19260 876 19392 882
rect 19260 870 19340 876
rect 19156 818 19208 824
rect 19340 818 19392 824
rect 19524 876 19576 882
rect 19524 818 19576 824
rect 19168 474 19196 818
rect 19536 474 19564 818
rect 20272 762 20300 2746
rect 20536 2508 20588 2514
rect 20640 2496 20668 3148
rect 20720 3130 20772 3136
rect 20916 2990 20944 3538
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 20916 2774 20944 2926
rect 20824 2746 20944 2774
rect 20824 2514 20852 2746
rect 21008 2650 21036 4626
rect 21100 4146 21128 5510
rect 21088 4140 21140 4146
rect 21088 4082 21140 4088
rect 21086 2816 21142 2825
rect 21192 2802 21220 7754
rect 21376 6798 21404 7783
rect 21468 7342 21496 7822
rect 21652 7410 21680 7890
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21456 7336 21508 7342
rect 21456 7278 21508 7284
rect 21928 7018 21956 7822
rect 21560 7002 21956 7018
rect 21548 6996 21956 7002
rect 21600 6990 21956 6996
rect 21548 6938 21600 6944
rect 22020 6934 22048 9454
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22008 6928 22060 6934
rect 22008 6870 22060 6876
rect 21732 6860 21784 6866
rect 21732 6802 21784 6808
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 21272 3732 21324 3738
rect 21272 3674 21324 3680
rect 21284 2854 21312 3674
rect 21142 2774 21220 2802
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 21086 2751 21142 2760
rect 20996 2644 21048 2650
rect 20996 2586 21048 2592
rect 20588 2468 20668 2496
rect 20812 2508 20864 2514
rect 20536 2450 20588 2456
rect 20812 2450 20864 2456
rect 20628 2304 20680 2310
rect 20626 2272 20628 2281
rect 20680 2272 20682 2281
rect 20626 2207 20682 2216
rect 20718 1864 20774 1873
rect 20824 1834 20852 2450
rect 21100 2394 21128 2751
rect 21284 2650 21312 2790
rect 21272 2644 21324 2650
rect 21192 2604 21272 2632
rect 21192 2446 21220 2604
rect 21272 2586 21324 2592
rect 21008 2366 21128 2394
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 21008 2310 21036 2366
rect 20996 2304 21048 2310
rect 20996 2246 21048 2252
rect 20902 2136 20958 2145
rect 20902 2071 20958 2080
rect 20718 1799 20720 1808
rect 20772 1799 20774 1808
rect 20812 1828 20864 1834
rect 20720 1770 20772 1776
rect 20812 1770 20864 1776
rect 20732 1426 20760 1770
rect 20824 1426 20852 1770
rect 20720 1420 20772 1426
rect 20720 1362 20772 1368
rect 20812 1420 20864 1426
rect 20812 1362 20864 1368
rect 20916 1306 20944 2071
rect 21008 1426 21036 2246
rect 21192 1766 21220 2382
rect 21272 2372 21324 2378
rect 21272 2314 21324 2320
rect 21180 1760 21232 1766
rect 21180 1702 21232 1708
rect 21192 1562 21220 1702
rect 21180 1556 21232 1562
rect 21180 1498 21232 1504
rect 20996 1420 21048 1426
rect 20996 1362 21048 1368
rect 20824 1278 20944 1306
rect 20718 1048 20774 1057
rect 20718 983 20720 992
rect 20772 983 20774 992
rect 20720 954 20772 960
rect 20720 876 20772 882
rect 20824 864 20852 1278
rect 21284 950 21312 2314
rect 21272 944 21324 950
rect 21272 886 21324 892
rect 20772 836 20852 864
rect 20720 818 20772 824
rect 20272 734 20484 762
rect 21376 746 21404 6734
rect 21640 6724 21692 6730
rect 21640 6666 21692 6672
rect 21652 6458 21680 6666
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21640 6180 21692 6186
rect 21640 6122 21692 6128
rect 21652 5778 21680 6122
rect 21640 5772 21692 5778
rect 21640 5714 21692 5720
rect 21640 5636 21692 5642
rect 21640 5578 21692 5584
rect 21652 5234 21680 5578
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 21640 5024 21692 5030
rect 21640 4966 21692 4972
rect 21652 4690 21680 4966
rect 21744 4826 21772 6802
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 21836 6186 21864 6734
rect 21928 6322 21956 6734
rect 22204 6662 22232 7278
rect 22388 6798 22416 11018
rect 22756 11014 22784 11308
rect 22836 11290 22888 11296
rect 22928 11212 22980 11218
rect 22848 11172 22928 11200
rect 22744 11008 22796 11014
rect 22744 10950 22796 10956
rect 22744 10804 22796 10810
rect 22848 10792 22876 11172
rect 23032 11200 23060 12038
rect 23400 11830 23428 12038
rect 23676 11830 23704 12174
rect 23388 11824 23440 11830
rect 23388 11766 23440 11772
rect 23664 11824 23716 11830
rect 23664 11766 23716 11772
rect 23296 11688 23348 11694
rect 23294 11656 23296 11665
rect 23348 11656 23350 11665
rect 23294 11591 23350 11600
rect 23400 11540 23428 11766
rect 23860 11626 23888 12174
rect 24228 11898 24256 12786
rect 24308 12300 24360 12306
rect 24308 12242 24360 12248
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 23940 11824 23992 11830
rect 24320 11778 24348 12242
rect 23992 11772 24348 11778
rect 23940 11766 24348 11772
rect 23952 11750 24348 11766
rect 24492 11756 24544 11762
rect 23952 11694 23980 11750
rect 24412 11716 24492 11744
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 23756 11620 23808 11626
rect 23756 11562 23808 11568
rect 23848 11620 23900 11626
rect 23848 11562 23900 11568
rect 23400 11512 23612 11540
rect 23168 11452 23476 11461
rect 23168 11450 23174 11452
rect 23230 11450 23254 11452
rect 23310 11450 23334 11452
rect 23390 11450 23414 11452
rect 23470 11450 23476 11452
rect 23230 11398 23232 11450
rect 23412 11398 23414 11450
rect 23168 11396 23174 11398
rect 23230 11396 23254 11398
rect 23310 11396 23334 11398
rect 23390 11396 23414 11398
rect 23470 11396 23476 11398
rect 23168 11387 23476 11396
rect 23204 11212 23256 11218
rect 23032 11172 23204 11200
rect 22928 11154 22980 11160
rect 23204 11154 23256 11160
rect 22796 10764 22876 10792
rect 22744 10746 22796 10752
rect 22926 10704 22982 10713
rect 22744 10668 22796 10674
rect 22926 10639 22982 10648
rect 22744 10610 22796 10616
rect 22652 10600 22704 10606
rect 22652 10542 22704 10548
rect 22560 9580 22612 9586
rect 22560 9522 22612 9528
rect 22376 6792 22428 6798
rect 22376 6734 22428 6740
rect 22192 6656 22244 6662
rect 22192 6598 22244 6604
rect 21916 6316 21968 6322
rect 21916 6258 21968 6264
rect 22572 6254 22600 9522
rect 22664 8004 22692 10542
rect 22756 9722 22784 10610
rect 22744 9716 22796 9722
rect 22744 9658 22796 9664
rect 22940 9178 22968 10639
rect 23216 10606 23244 11154
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 23204 10600 23256 10606
rect 23204 10542 23256 10548
rect 23308 10452 23336 11086
rect 23584 10742 23612 11512
rect 23768 11150 23796 11562
rect 24412 11354 24440 11716
rect 24492 11698 24544 11704
rect 24490 11656 24546 11665
rect 24490 11591 24546 11600
rect 24504 11354 24532 11591
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24492 11348 24544 11354
rect 24492 11290 24544 11296
rect 24872 11218 24900 14214
rect 25148 11665 25176 16390
rect 25332 15502 25360 16390
rect 25412 16040 25464 16046
rect 25412 15982 25464 15988
rect 25320 15496 25372 15502
rect 25320 15438 25372 15444
rect 25320 15360 25372 15366
rect 25320 15302 25372 15308
rect 25332 15094 25360 15302
rect 25320 15088 25372 15094
rect 25320 15030 25372 15036
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25332 12442 25360 13262
rect 25424 12782 25452 15982
rect 25516 15434 25544 17983
rect 25504 15428 25556 15434
rect 25504 15370 25556 15376
rect 25608 14618 25636 19246
rect 25700 16028 25728 20334
rect 26240 20256 26292 20262
rect 26240 20198 26292 20204
rect 26252 19145 26280 20198
rect 26238 19136 26294 19145
rect 26238 19071 26294 19080
rect 26056 18692 26108 18698
rect 26056 18634 26108 18640
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 25976 18290 26004 18566
rect 25964 18284 26016 18290
rect 25964 18226 26016 18232
rect 25780 17672 25832 17678
rect 25780 17614 25832 17620
rect 25792 17542 25820 17614
rect 25780 17536 25832 17542
rect 25872 17536 25924 17542
rect 25780 17478 25832 17484
rect 25870 17504 25872 17513
rect 25924 17504 25926 17513
rect 25792 16658 25820 17478
rect 25870 17439 25926 17448
rect 25872 16992 25924 16998
rect 25872 16934 25924 16940
rect 25780 16652 25832 16658
rect 25780 16594 25832 16600
rect 25700 16000 25820 16028
rect 25688 15904 25740 15910
rect 25688 15846 25740 15852
rect 25700 14929 25728 15846
rect 25792 15201 25820 16000
rect 25778 15192 25834 15201
rect 25778 15127 25834 15136
rect 25686 14920 25742 14929
rect 25686 14855 25742 14864
rect 25596 14612 25648 14618
rect 25596 14554 25648 14560
rect 25688 14408 25740 14414
rect 25688 14350 25740 14356
rect 25792 14362 25820 15127
rect 25884 14464 25912 16934
rect 26068 16794 26096 18634
rect 26148 18080 26200 18086
rect 26148 18022 26200 18028
rect 26160 17882 26188 18022
rect 26148 17876 26200 17882
rect 26148 17818 26200 17824
rect 26252 16998 26280 19071
rect 26436 18766 26464 20402
rect 26608 20324 26660 20330
rect 26608 20266 26660 20272
rect 26516 20256 26568 20262
rect 26516 20198 26568 20204
rect 26528 20058 26556 20198
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 26620 19281 26648 20266
rect 26712 19718 26740 20878
rect 26804 19854 26832 20878
rect 26884 20800 26936 20806
rect 26884 20742 26936 20748
rect 26792 19848 26844 19854
rect 26792 19790 26844 19796
rect 26700 19712 26752 19718
rect 26700 19654 26752 19660
rect 26606 19272 26662 19281
rect 26606 19207 26662 19216
rect 26620 18952 26648 19207
rect 26528 18924 26740 18952
rect 26424 18760 26476 18766
rect 26424 18702 26476 18708
rect 26424 18624 26476 18630
rect 26424 18566 26476 18572
rect 26436 17202 26464 18566
rect 26424 17196 26476 17202
rect 26424 17138 26476 17144
rect 26240 16992 26292 16998
rect 26240 16934 26292 16940
rect 26056 16788 26108 16794
rect 26056 16730 26108 16736
rect 25964 16244 26016 16250
rect 25964 16186 26016 16192
rect 25976 15745 26004 16186
rect 26068 16114 26096 16730
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 26056 16108 26108 16114
rect 26108 16068 26188 16096
rect 26056 16050 26108 16056
rect 25962 15736 26018 15745
rect 25962 15671 26018 15680
rect 25976 15638 26004 15671
rect 25964 15632 26016 15638
rect 25964 15574 26016 15580
rect 26160 15502 26188 16068
rect 26252 15881 26280 16594
rect 26424 16448 26476 16454
rect 26424 16390 26476 16396
rect 26332 16108 26384 16114
rect 26332 16050 26384 16056
rect 26238 15872 26294 15881
rect 26238 15807 26294 15816
rect 25964 15496 26016 15502
rect 25964 15438 26016 15444
rect 26148 15496 26200 15502
rect 26148 15438 26200 15444
rect 25976 14958 26004 15438
rect 26148 15360 26200 15366
rect 26148 15302 26200 15308
rect 25964 14952 26016 14958
rect 26160 14929 26188 15302
rect 25964 14894 26016 14900
rect 26146 14920 26202 14929
rect 26146 14855 26202 14864
rect 26148 14816 26200 14822
rect 26148 14758 26200 14764
rect 26160 14618 26188 14758
rect 26148 14612 26200 14618
rect 26148 14554 26200 14560
rect 25964 14476 26016 14482
rect 25884 14436 25964 14464
rect 25964 14418 26016 14424
rect 25504 14000 25556 14006
rect 25504 13942 25556 13948
rect 25516 13394 25544 13942
rect 25504 13388 25556 13394
rect 25504 13330 25556 13336
rect 25700 12986 25728 14350
rect 25792 14334 26004 14362
rect 25976 13190 26004 14334
rect 26252 13734 26280 15807
rect 26240 13728 26292 13734
rect 26240 13670 26292 13676
rect 26344 13462 26372 16050
rect 26436 13870 26464 16390
rect 26528 15910 26556 18924
rect 26712 18834 26740 18924
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26700 18828 26752 18834
rect 26700 18770 26752 18776
rect 26620 18442 26648 18770
rect 26620 18414 26740 18442
rect 26804 18426 26832 19790
rect 26608 18352 26660 18358
rect 26606 18320 26608 18329
rect 26660 18320 26662 18329
rect 26606 18255 26662 18264
rect 26606 17232 26662 17241
rect 26712 17218 26740 18414
rect 26792 18420 26844 18426
rect 26792 18362 26844 18368
rect 26662 17190 26740 17218
rect 26606 17167 26662 17176
rect 26804 17134 26832 18362
rect 26896 17678 26924 20742
rect 26963 20700 27271 20709
rect 26963 20698 26969 20700
rect 27025 20698 27049 20700
rect 27105 20698 27129 20700
rect 27185 20698 27209 20700
rect 27265 20698 27271 20700
rect 27025 20646 27027 20698
rect 27207 20646 27209 20698
rect 26963 20644 26969 20646
rect 27025 20644 27049 20646
rect 27105 20644 27129 20646
rect 27185 20644 27209 20646
rect 27265 20644 27271 20646
rect 26963 20635 27271 20644
rect 27068 20596 27120 20602
rect 27068 20538 27120 20544
rect 27080 20398 27108 20538
rect 27068 20392 27120 20398
rect 27068 20334 27120 20340
rect 26963 19612 27271 19621
rect 26963 19610 26969 19612
rect 27025 19610 27049 19612
rect 27105 19610 27129 19612
rect 27185 19610 27209 19612
rect 27265 19610 27271 19612
rect 27025 19558 27027 19610
rect 27207 19558 27209 19610
rect 26963 19556 26969 19558
rect 27025 19556 27049 19558
rect 27105 19556 27129 19558
rect 27185 19556 27209 19558
rect 27265 19556 27271 19558
rect 26963 19547 27271 19556
rect 27356 19334 27384 21134
rect 27436 21004 27488 21010
rect 27436 20946 27488 20952
rect 27448 20602 27476 20946
rect 27436 20596 27488 20602
rect 27436 20538 27488 20544
rect 27816 20058 27844 21422
rect 27804 20052 27856 20058
rect 27804 19994 27856 20000
rect 27620 19848 27672 19854
rect 27620 19790 27672 19796
rect 26976 19304 27028 19310
rect 26974 19272 26976 19281
rect 27264 19306 27384 19334
rect 27028 19272 27030 19281
rect 26974 19207 27030 19216
rect 27264 19156 27292 19306
rect 27632 19281 27660 19790
rect 27618 19272 27674 19281
rect 27618 19207 27674 19216
rect 27264 19128 27384 19156
rect 26963 18524 27271 18533
rect 26963 18522 26969 18524
rect 27025 18522 27049 18524
rect 27105 18522 27129 18524
rect 27185 18522 27209 18524
rect 27265 18522 27271 18524
rect 27025 18470 27027 18522
rect 27207 18470 27209 18522
rect 26963 18468 26969 18470
rect 27025 18468 27049 18470
rect 27105 18468 27129 18470
rect 27185 18468 27209 18470
rect 27265 18468 27271 18470
rect 26963 18459 27271 18468
rect 27066 17912 27122 17921
rect 27066 17847 27068 17856
rect 27120 17847 27122 17856
rect 27068 17818 27120 17824
rect 26884 17672 26936 17678
rect 26884 17614 26936 17620
rect 26963 17436 27271 17445
rect 26963 17434 26969 17436
rect 27025 17434 27049 17436
rect 27105 17434 27129 17436
rect 27185 17434 27209 17436
rect 27265 17434 27271 17436
rect 27025 17382 27027 17434
rect 27207 17382 27209 17434
rect 26963 17380 26969 17382
rect 27025 17380 27049 17382
rect 27105 17380 27129 17382
rect 27185 17380 27209 17382
rect 27265 17380 27271 17382
rect 26963 17371 27271 17380
rect 26792 17128 26844 17134
rect 26698 17096 26754 17105
rect 26792 17070 26844 17076
rect 26698 17031 26754 17040
rect 26712 16998 26740 17031
rect 26608 16992 26660 16998
rect 26608 16934 26660 16940
rect 26700 16992 26752 16998
rect 26700 16934 26752 16940
rect 26620 16697 26648 16934
rect 26884 16788 26936 16794
rect 26884 16730 26936 16736
rect 26606 16688 26662 16697
rect 26606 16623 26662 16632
rect 26792 16652 26844 16658
rect 26792 16594 26844 16600
rect 26516 15904 26568 15910
rect 26516 15846 26568 15852
rect 26528 15638 26556 15846
rect 26804 15745 26832 16594
rect 26790 15736 26846 15745
rect 26790 15671 26846 15680
rect 26516 15632 26568 15638
rect 26516 15574 26568 15580
rect 26528 14822 26556 15574
rect 26700 15360 26752 15366
rect 26804 15337 26832 15671
rect 26700 15302 26752 15308
rect 26790 15328 26846 15337
rect 26608 15020 26660 15026
rect 26608 14962 26660 14968
rect 26516 14816 26568 14822
rect 26516 14758 26568 14764
rect 26516 14476 26568 14482
rect 26516 14418 26568 14424
rect 26528 14385 26556 14418
rect 26514 14376 26570 14385
rect 26514 14311 26570 14320
rect 26424 13864 26476 13870
rect 26476 13824 26556 13852
rect 26424 13806 26476 13812
rect 26424 13524 26476 13530
rect 26424 13466 26476 13472
rect 26332 13456 26384 13462
rect 26332 13398 26384 13404
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 25964 13184 26016 13190
rect 25964 13126 26016 13132
rect 25688 12980 25740 12986
rect 25688 12922 25740 12928
rect 25412 12776 25464 12782
rect 25412 12718 25464 12724
rect 25320 12436 25372 12442
rect 25320 12378 25372 12384
rect 25780 12300 25832 12306
rect 25780 12242 25832 12248
rect 25320 11688 25372 11694
rect 25134 11656 25190 11665
rect 25320 11630 25372 11636
rect 25134 11591 25190 11600
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 24964 11014 24992 11086
rect 24952 11008 25004 11014
rect 24952 10950 25004 10956
rect 24492 10804 24544 10810
rect 24492 10746 24544 10752
rect 23572 10736 23624 10742
rect 23572 10678 23624 10684
rect 24214 10704 24270 10713
rect 24270 10674 24348 10690
rect 24270 10668 24360 10674
rect 24270 10662 24308 10668
rect 24214 10639 24270 10648
rect 24308 10610 24360 10616
rect 23848 10600 23900 10606
rect 24216 10600 24268 10606
rect 23848 10542 23900 10548
rect 24214 10568 24216 10577
rect 24268 10568 24270 10577
rect 23032 10424 23336 10452
rect 23032 10266 23060 10424
rect 23168 10364 23476 10373
rect 23168 10362 23174 10364
rect 23230 10362 23254 10364
rect 23310 10362 23334 10364
rect 23390 10362 23414 10364
rect 23470 10362 23476 10364
rect 23230 10310 23232 10362
rect 23412 10310 23414 10362
rect 23168 10308 23174 10310
rect 23230 10308 23254 10310
rect 23310 10308 23334 10310
rect 23390 10308 23414 10310
rect 23470 10308 23476 10310
rect 23168 10299 23476 10308
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 23860 9722 23888 10542
rect 24270 10526 24348 10554
rect 24214 10503 24270 10512
rect 23848 9716 23900 9722
rect 23848 9658 23900 9664
rect 24320 9674 24348 10526
rect 24504 10062 24532 10746
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24596 10470 24624 10542
rect 24584 10464 24636 10470
rect 24584 10406 24636 10412
rect 24492 10056 24544 10062
rect 24492 9998 24544 10004
rect 24320 9646 24440 9674
rect 24124 9512 24176 9518
rect 24122 9480 24124 9489
rect 24176 9480 24178 9489
rect 23664 9444 23716 9450
rect 24122 9415 24178 9424
rect 23664 9386 23716 9392
rect 23168 9276 23476 9285
rect 23168 9274 23174 9276
rect 23230 9274 23254 9276
rect 23310 9274 23334 9276
rect 23390 9274 23414 9276
rect 23470 9274 23476 9276
rect 23230 9222 23232 9274
rect 23412 9222 23414 9274
rect 23168 9220 23174 9222
rect 23230 9220 23254 9222
rect 23310 9220 23334 9222
rect 23390 9220 23414 9222
rect 23470 9220 23476 9222
rect 23168 9211 23476 9220
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 23676 9058 23704 9386
rect 24412 9382 24440 9646
rect 24766 9616 24822 9625
rect 24766 9551 24768 9560
rect 24820 9551 24822 9560
rect 24860 9580 24912 9586
rect 24768 9522 24820 9528
rect 24860 9522 24912 9528
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23940 9376 23992 9382
rect 23940 9318 23992 9324
rect 24124 9376 24176 9382
rect 24124 9318 24176 9324
rect 24308 9376 24360 9382
rect 24308 9318 24360 9324
rect 24400 9376 24452 9382
rect 24400 9318 24452 9324
rect 23768 9178 23796 9318
rect 23756 9172 23808 9178
rect 23756 9114 23808 9120
rect 23676 9030 23796 9058
rect 23664 8968 23716 8974
rect 23664 8910 23716 8916
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23492 8566 23520 8774
rect 23480 8560 23532 8566
rect 23480 8502 23532 8508
rect 23676 8362 23704 8910
rect 23768 8838 23796 9030
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 23952 8430 23980 9318
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 23940 8424 23992 8430
rect 23940 8366 23992 8372
rect 23664 8356 23716 8362
rect 23664 8298 23716 8304
rect 23756 8288 23808 8294
rect 23756 8230 23808 8236
rect 23168 8188 23476 8197
rect 23168 8186 23174 8188
rect 23230 8186 23254 8188
rect 23310 8186 23334 8188
rect 23390 8186 23414 8188
rect 23470 8186 23476 8188
rect 23230 8134 23232 8186
rect 23412 8134 23414 8186
rect 23168 8132 23174 8134
rect 23230 8132 23254 8134
rect 23310 8132 23334 8134
rect 23390 8132 23414 8134
rect 23470 8132 23476 8134
rect 23168 8123 23476 8132
rect 23768 8090 23796 8230
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 22744 8016 22796 8022
rect 22664 7976 22744 8004
rect 22744 7958 22796 7964
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22652 7200 22704 7206
rect 22756 7154 22784 7822
rect 22836 7812 22888 7818
rect 22836 7754 22888 7760
rect 22704 7148 22784 7154
rect 22652 7142 22784 7148
rect 22664 7126 22784 7142
rect 22652 6860 22704 6866
rect 22652 6802 22704 6808
rect 22664 6769 22692 6802
rect 22650 6760 22706 6769
rect 22650 6695 22706 6704
rect 22756 6254 22784 7126
rect 22848 6662 22876 7754
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23400 7546 23428 7686
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23168 7100 23476 7109
rect 23168 7098 23174 7100
rect 23230 7098 23254 7100
rect 23310 7098 23334 7100
rect 23390 7098 23414 7100
rect 23470 7098 23476 7100
rect 23230 7046 23232 7098
rect 23412 7046 23414 7098
rect 23168 7044 23174 7046
rect 23230 7044 23254 7046
rect 23310 7044 23334 7046
rect 23390 7044 23414 7046
rect 23470 7044 23476 7046
rect 23168 7035 23476 7044
rect 23020 6860 23072 6866
rect 23020 6802 23072 6808
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 23032 6322 23060 6802
rect 23386 6352 23442 6361
rect 23020 6316 23072 6322
rect 23386 6287 23388 6296
rect 23020 6258 23072 6264
rect 23440 6287 23442 6296
rect 23388 6258 23440 6264
rect 23584 6254 23612 7890
rect 23756 7880 23808 7886
rect 23756 7822 23808 7828
rect 22560 6248 22612 6254
rect 22480 6208 22560 6236
rect 21824 6180 21876 6186
rect 21824 6122 21876 6128
rect 21916 6112 21968 6118
rect 21916 6054 21968 6060
rect 22100 6112 22152 6118
rect 22100 6054 22152 6060
rect 21928 5914 21956 6054
rect 21916 5908 21968 5914
rect 21916 5850 21968 5856
rect 21836 5778 22048 5794
rect 21824 5772 22048 5778
rect 21876 5766 22048 5772
rect 21824 5714 21876 5720
rect 21916 5704 21968 5710
rect 21916 5646 21968 5652
rect 21928 5166 21956 5646
rect 22020 5166 22048 5766
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 22008 5160 22060 5166
rect 22008 5102 22060 5108
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 21640 4684 21692 4690
rect 21640 4626 21692 4632
rect 21652 4593 21680 4626
rect 21638 4584 21694 4593
rect 21638 4519 21694 4528
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21640 4480 21692 4486
rect 21640 4422 21692 4428
rect 21560 3058 21588 4422
rect 21652 4282 21680 4422
rect 21744 4282 21772 4762
rect 21928 4690 21956 5102
rect 22112 4826 22140 6054
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22374 5672 22430 5681
rect 22296 5030 22324 5646
rect 22374 5607 22430 5616
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22296 4826 22324 4966
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 22284 4820 22336 4826
rect 22284 4762 22336 4768
rect 21916 4684 21968 4690
rect 21916 4626 21968 4632
rect 21824 4548 21876 4554
rect 21824 4490 21876 4496
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21732 4276 21784 4282
rect 21732 4218 21784 4224
rect 21836 3602 21864 4490
rect 22296 4010 22324 4762
rect 22388 4622 22416 5607
rect 22480 5574 22508 6208
rect 22560 6190 22612 6196
rect 22744 6248 22796 6254
rect 22744 6190 22796 6196
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22572 5778 22600 6054
rect 23168 6012 23476 6021
rect 23168 6010 23174 6012
rect 23230 6010 23254 6012
rect 23310 6010 23334 6012
rect 23390 6010 23414 6012
rect 23470 6010 23476 6012
rect 23230 5958 23232 6010
rect 23412 5958 23414 6010
rect 23168 5956 23174 5958
rect 23230 5956 23254 5958
rect 23310 5956 23334 5958
rect 23390 5956 23414 5958
rect 23470 5956 23476 5958
rect 23168 5947 23476 5956
rect 23386 5808 23442 5817
rect 22560 5772 22612 5778
rect 23386 5743 23442 5752
rect 22560 5714 22612 5720
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 23400 5250 23428 5743
rect 23308 5222 23428 5250
rect 23480 5296 23532 5302
rect 23480 5238 23532 5244
rect 23308 5166 23336 5222
rect 23296 5160 23348 5166
rect 23124 5108 23296 5114
rect 23124 5102 23348 5108
rect 23124 5098 23336 5102
rect 23492 5098 23520 5238
rect 23572 5228 23624 5234
rect 23572 5170 23624 5176
rect 23112 5092 23336 5098
rect 23164 5086 23336 5092
rect 23480 5092 23532 5098
rect 23112 5034 23164 5040
rect 23480 5034 23532 5040
rect 22652 5024 22704 5030
rect 22652 4966 22704 4972
rect 22664 4622 22692 4966
rect 23168 4924 23476 4933
rect 23168 4922 23174 4924
rect 23230 4922 23254 4924
rect 23310 4922 23334 4924
rect 23390 4922 23414 4924
rect 23470 4922 23476 4924
rect 23230 4870 23232 4922
rect 23412 4870 23414 4922
rect 23168 4868 23174 4870
rect 23230 4868 23254 4870
rect 23310 4868 23334 4870
rect 23390 4868 23414 4870
rect 23470 4868 23476 4870
rect 23168 4859 23476 4868
rect 22376 4616 22428 4622
rect 22376 4558 22428 4564
rect 22652 4616 22704 4622
rect 22652 4558 22704 4564
rect 23112 4276 23164 4282
rect 23112 4218 23164 4224
rect 23124 4078 23152 4218
rect 22376 4072 22428 4078
rect 22376 4014 22428 4020
rect 23112 4072 23164 4078
rect 23112 4014 23164 4020
rect 22100 4004 22152 4010
rect 22100 3946 22152 3952
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 22112 3738 22140 3946
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 22388 3194 22416 4014
rect 22652 4004 22704 4010
rect 22652 3946 22704 3952
rect 22376 3188 22428 3194
rect 22376 3130 22428 3136
rect 22664 3126 22692 3946
rect 23168 3836 23476 3845
rect 23168 3834 23174 3836
rect 23230 3834 23254 3836
rect 23310 3834 23334 3836
rect 23390 3834 23414 3836
rect 23470 3834 23476 3836
rect 23230 3782 23232 3834
rect 23412 3782 23414 3834
rect 23168 3780 23174 3782
rect 23230 3780 23254 3782
rect 23310 3780 23334 3782
rect 23390 3780 23414 3782
rect 23470 3780 23476 3782
rect 23168 3771 23476 3780
rect 23584 3738 23612 5170
rect 23664 5160 23716 5166
rect 23664 5102 23716 5108
rect 23572 3732 23624 3738
rect 23572 3674 23624 3680
rect 23676 3534 23704 5102
rect 23768 3738 23796 7822
rect 23860 7410 23888 8366
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23848 7404 23900 7410
rect 23848 7346 23900 7352
rect 23952 7002 23980 7822
rect 24044 7546 24072 8910
rect 24032 7540 24084 7546
rect 24032 7482 24084 7488
rect 24136 7410 24164 9318
rect 24216 9172 24268 9178
rect 24216 9114 24268 9120
rect 24228 9042 24256 9114
rect 24216 9036 24268 9042
rect 24216 8978 24268 8984
rect 24320 8480 24348 9318
rect 24872 9178 24900 9522
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24400 8492 24452 8498
rect 24320 8452 24400 8480
rect 24400 8434 24452 8440
rect 24308 8288 24360 8294
rect 24308 8230 24360 8236
rect 24216 7880 24268 7886
rect 24216 7822 24268 7828
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 24030 7032 24086 7041
rect 23940 6996 23992 7002
rect 24136 7002 24164 7142
rect 24030 6967 24086 6976
rect 24124 6996 24176 7002
rect 23940 6938 23992 6944
rect 24044 6934 24072 6967
rect 24124 6938 24176 6944
rect 24032 6928 24084 6934
rect 24032 6870 24084 6876
rect 24228 6322 24256 7822
rect 24320 7206 24348 8230
rect 24308 7200 24360 7206
rect 24308 7142 24360 7148
rect 24492 7200 24544 7206
rect 24492 7142 24544 7148
rect 24504 6866 24532 7142
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24216 6316 24268 6322
rect 24216 6258 24268 6264
rect 24688 6118 24716 6734
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 23848 6112 23900 6118
rect 23848 6054 23900 6060
rect 24492 6112 24544 6118
rect 24492 6054 24544 6060
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 23860 5710 23888 6054
rect 24504 5914 24532 6054
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 23848 5704 23900 5710
rect 23848 5646 23900 5652
rect 23860 4146 23888 5646
rect 24308 4480 24360 4486
rect 24308 4422 24360 4428
rect 24320 4146 24348 4422
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 24308 4140 24360 4146
rect 24308 4082 24360 4088
rect 23860 4026 23888 4082
rect 23860 3998 23980 4026
rect 23756 3732 23808 3738
rect 23756 3674 23808 3680
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 23848 3528 23900 3534
rect 23848 3470 23900 3476
rect 22652 3120 22704 3126
rect 22652 3062 22704 3068
rect 21548 3052 21600 3058
rect 21548 2994 21600 3000
rect 23676 2990 23704 3470
rect 23860 3126 23888 3470
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 21732 2984 21784 2990
rect 21732 2926 21784 2932
rect 23664 2984 23716 2990
rect 23664 2926 23716 2932
rect 21744 2854 21772 2926
rect 21732 2848 21784 2854
rect 21732 2790 21784 2796
rect 23168 2748 23476 2757
rect 23168 2746 23174 2748
rect 23230 2746 23254 2748
rect 23310 2746 23334 2748
rect 23390 2746 23414 2748
rect 23470 2746 23476 2748
rect 23230 2694 23232 2746
rect 23412 2694 23414 2746
rect 23168 2692 23174 2694
rect 23230 2692 23254 2694
rect 23310 2692 23334 2694
rect 23390 2692 23414 2694
rect 23470 2692 23476 2694
rect 23168 2683 23476 2692
rect 23676 2582 23704 2926
rect 23860 2854 23888 3062
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 23952 2774 23980 3998
rect 24124 4004 24176 4010
rect 24124 3946 24176 3952
rect 24136 3602 24164 3946
rect 24504 3942 24532 5850
rect 24780 4826 24808 6190
rect 24858 5808 24914 5817
rect 24964 5794 24992 10950
rect 25044 10600 25096 10606
rect 25044 10542 25096 10548
rect 25056 10266 25084 10542
rect 25044 10260 25096 10266
rect 25044 10202 25096 10208
rect 25148 10062 25176 11591
rect 25332 11286 25360 11630
rect 25320 11280 25372 11286
rect 25318 11248 25320 11257
rect 25372 11248 25374 11257
rect 25318 11183 25374 11192
rect 25504 11144 25556 11150
rect 25504 11086 25556 11092
rect 25320 11008 25372 11014
rect 25320 10950 25372 10956
rect 25332 10606 25360 10950
rect 25320 10600 25372 10606
rect 25320 10542 25372 10548
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25332 9994 25360 10542
rect 25320 9988 25372 9994
rect 25320 9930 25372 9936
rect 25044 9920 25096 9926
rect 25044 9862 25096 9868
rect 25056 9489 25084 9862
rect 25412 9512 25464 9518
rect 25042 9480 25098 9489
rect 25412 9454 25464 9460
rect 25042 9415 25098 9424
rect 25424 9178 25452 9454
rect 25412 9172 25464 9178
rect 25412 9114 25464 9120
rect 25412 8560 25464 8566
rect 25412 8502 25464 8508
rect 25320 8424 25372 8430
rect 25320 8366 25372 8372
rect 25332 7857 25360 8366
rect 25318 7848 25374 7857
rect 25318 7783 25374 7792
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25332 7546 25360 7686
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25320 7336 25372 7342
rect 25320 7278 25372 7284
rect 25134 7168 25190 7177
rect 25134 7103 25190 7112
rect 24914 5766 24992 5794
rect 24858 5743 24914 5752
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 24676 4820 24728 4826
rect 24676 4762 24728 4768
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 24688 4706 24716 4762
rect 24872 4706 24900 5646
rect 25044 5228 25096 5234
rect 25044 5170 25096 5176
rect 25056 4758 25084 5170
rect 24688 4678 24900 4706
rect 25044 4752 25096 4758
rect 25044 4694 25096 4700
rect 25148 4690 25176 7103
rect 25332 7041 25360 7278
rect 25318 7032 25374 7041
rect 25318 6967 25374 6976
rect 25320 5160 25372 5166
rect 25320 5102 25372 5108
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 24676 4480 24728 4486
rect 25044 4480 25096 4486
rect 24676 4422 24728 4428
rect 24872 4440 25044 4468
rect 24688 4146 24716 4422
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 24400 3936 24452 3942
rect 24400 3878 24452 3884
rect 24492 3936 24544 3942
rect 24492 3878 24544 3884
rect 24124 3596 24176 3602
rect 24124 3538 24176 3544
rect 24412 3058 24440 3878
rect 24504 3602 24532 3878
rect 24492 3596 24544 3602
rect 24492 3538 24544 3544
rect 24400 3052 24452 3058
rect 24400 2994 24452 3000
rect 24124 2848 24176 2854
rect 24124 2790 24176 2796
rect 23952 2746 24072 2774
rect 23664 2576 23716 2582
rect 23584 2536 23664 2564
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 21928 2281 21956 2382
rect 21914 2272 21970 2281
rect 21914 2207 21970 2216
rect 22020 2106 22048 2382
rect 23480 2372 23532 2378
rect 23480 2314 23532 2320
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 21456 2100 21508 2106
rect 21456 2042 21508 2048
rect 22008 2100 22060 2106
rect 22008 2042 22060 2048
rect 21468 1970 21496 2042
rect 21456 1964 21508 1970
rect 21456 1906 21508 1912
rect 22744 1896 22796 1902
rect 22744 1838 22796 1844
rect 22928 1896 22980 1902
rect 22928 1838 22980 1844
rect 22756 1562 22784 1838
rect 22836 1760 22888 1766
rect 22836 1702 22888 1708
rect 22744 1556 22796 1562
rect 22744 1498 22796 1504
rect 22848 1358 22876 1702
rect 22836 1352 22888 1358
rect 22836 1294 22888 1300
rect 21916 1216 21968 1222
rect 21916 1158 21968 1164
rect 21928 882 21956 1158
rect 21916 876 21968 882
rect 21916 818 21968 824
rect 22192 808 22244 814
rect 22006 776 22062 785
rect 20456 678 20484 734
rect 21364 740 21416 746
rect 22192 750 22244 756
rect 22006 711 22062 720
rect 21364 682 21416 688
rect 22020 678 22048 711
rect 22204 678 22232 750
rect 20444 672 20496 678
rect 20444 614 20496 620
rect 22008 672 22060 678
rect 22008 614 22060 620
rect 22192 672 22244 678
rect 22192 614 22244 620
rect 22112 474 22232 490
rect 19156 468 19208 474
rect 19156 410 19208 416
rect 19524 468 19576 474
rect 19524 410 19576 416
rect 22100 468 22232 474
rect 22152 462 22232 468
rect 22100 410 22152 416
rect 22204 338 22232 462
rect 22940 406 22968 1838
rect 23032 882 23060 2246
rect 23492 2038 23520 2314
rect 23480 2032 23532 2038
rect 23480 1974 23532 1980
rect 23492 1902 23520 1974
rect 23296 1896 23348 1902
rect 23294 1864 23296 1873
rect 23480 1896 23532 1902
rect 23348 1864 23350 1873
rect 23480 1838 23532 1844
rect 23294 1799 23350 1808
rect 23168 1660 23476 1669
rect 23168 1658 23174 1660
rect 23230 1658 23254 1660
rect 23310 1658 23334 1660
rect 23390 1658 23414 1660
rect 23470 1658 23476 1660
rect 23230 1606 23232 1658
rect 23412 1606 23414 1658
rect 23168 1604 23174 1606
rect 23230 1604 23254 1606
rect 23310 1604 23334 1606
rect 23390 1604 23414 1606
rect 23470 1604 23476 1606
rect 23168 1595 23476 1604
rect 23584 1544 23612 2536
rect 23664 2518 23716 2524
rect 24044 2514 24072 2746
rect 23756 2508 23808 2514
rect 23756 2450 23808 2456
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 23664 1760 23716 1766
rect 23664 1702 23716 1708
rect 23492 1516 23612 1544
rect 23492 1358 23520 1516
rect 23572 1420 23624 1426
rect 23572 1362 23624 1368
rect 23480 1352 23532 1358
rect 23480 1294 23532 1300
rect 23480 1012 23532 1018
rect 23480 954 23532 960
rect 23492 921 23520 954
rect 23478 912 23534 921
rect 23020 876 23072 882
rect 23584 882 23612 1362
rect 23478 847 23534 856
rect 23572 876 23624 882
rect 23020 818 23072 824
rect 23572 818 23624 824
rect 23676 678 23704 1702
rect 23664 672 23716 678
rect 23664 614 23716 620
rect 23168 572 23476 581
rect 23168 570 23174 572
rect 23230 570 23254 572
rect 23310 570 23334 572
rect 23390 570 23414 572
rect 23470 570 23476 572
rect 23230 518 23232 570
rect 23412 518 23414 570
rect 23168 516 23174 518
rect 23230 516 23254 518
rect 23310 516 23334 518
rect 23390 516 23414 518
rect 23470 516 23476 518
rect 23168 507 23476 516
rect 22928 400 22980 406
rect 22928 342 22980 348
rect 22100 332 22152 338
rect 22100 274 22152 280
rect 22192 332 22244 338
rect 22192 274 22244 280
rect 22112 134 22140 274
rect 23768 202 23796 2450
rect 23940 1828 23992 1834
rect 23940 1770 23992 1776
rect 23952 1358 23980 1770
rect 24032 1420 24084 1426
rect 24136 1408 24164 2790
rect 24504 2774 24532 3538
rect 24676 3392 24728 3398
rect 24676 3334 24728 3340
rect 24504 2746 24624 2774
rect 24308 2440 24360 2446
rect 24492 2440 24544 2446
rect 24360 2400 24440 2428
rect 24308 2382 24360 2388
rect 24308 2304 24360 2310
rect 24308 2246 24360 2252
rect 24216 1760 24268 1766
rect 24216 1702 24268 1708
rect 24084 1380 24164 1408
rect 24032 1362 24084 1368
rect 23940 1352 23992 1358
rect 23940 1294 23992 1300
rect 23848 1216 23900 1222
rect 23848 1158 23900 1164
rect 23860 814 23888 1158
rect 23848 808 23900 814
rect 23848 750 23900 756
rect 23938 776 23994 785
rect 24044 762 24072 1362
rect 23994 734 24072 762
rect 23938 711 23994 720
rect 23952 678 23980 711
rect 23940 672 23992 678
rect 23940 614 23992 620
rect 23756 196 23808 202
rect 23756 138 23808 144
rect 24228 134 24256 1702
rect 24320 474 24348 2246
rect 24412 1902 24440 2400
rect 24596 2428 24624 2746
rect 24688 2446 24716 3334
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 24544 2400 24624 2428
rect 24492 2382 24544 2388
rect 24400 1896 24452 1902
rect 24400 1838 24452 1844
rect 24412 1222 24440 1838
rect 24596 1766 24624 2400
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 24780 1970 24808 2994
rect 24872 2514 24900 4440
rect 25044 4422 25096 4428
rect 25148 4282 25176 4626
rect 25332 4622 25360 5102
rect 25424 4622 25452 8502
rect 25516 7936 25544 11086
rect 25688 10464 25740 10470
rect 25688 10406 25740 10412
rect 25700 10266 25728 10406
rect 25688 10260 25740 10266
rect 25688 10202 25740 10208
rect 25688 7948 25740 7954
rect 25516 7908 25688 7936
rect 25688 7890 25740 7896
rect 25504 7744 25556 7750
rect 25504 7686 25556 7692
rect 25596 7744 25648 7750
rect 25596 7686 25648 7692
rect 25320 4616 25372 4622
rect 25320 4558 25372 4564
rect 25412 4616 25464 4622
rect 25412 4558 25464 4564
rect 25516 4486 25544 7686
rect 25608 6866 25636 7686
rect 25596 6860 25648 6866
rect 25596 6802 25648 6808
rect 25596 6180 25648 6186
rect 25596 6122 25648 6128
rect 25608 5370 25636 6122
rect 25596 5364 25648 5370
rect 25596 5306 25648 5312
rect 25596 4752 25648 4758
rect 25596 4694 25648 4700
rect 25320 4480 25372 4486
rect 25320 4422 25372 4428
rect 25504 4480 25556 4486
rect 25504 4422 25556 4428
rect 25136 4276 25188 4282
rect 25136 4218 25188 4224
rect 25332 2774 25360 4422
rect 25412 3596 25464 3602
rect 25412 3538 25464 3544
rect 25424 3194 25452 3538
rect 25412 3188 25464 3194
rect 25412 3130 25464 3136
rect 25056 2746 25360 2774
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 25056 1970 25084 2746
rect 25608 2145 25636 4694
rect 25700 2990 25728 7890
rect 25792 3602 25820 12242
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 25884 11218 25912 12038
rect 26068 11898 26096 13330
rect 26436 12850 26464 13466
rect 26424 12844 26476 12850
rect 26424 12786 26476 12792
rect 26148 12776 26200 12782
rect 26148 12718 26200 12724
rect 26160 12617 26188 12718
rect 26332 12640 26384 12646
rect 26146 12608 26202 12617
rect 26332 12582 26384 12588
rect 26146 12543 26202 12552
rect 26160 12442 26188 12543
rect 26148 12436 26200 12442
rect 26148 12378 26200 12384
rect 26160 12306 26188 12378
rect 26148 12300 26200 12306
rect 26148 12242 26200 12248
rect 26056 11892 26108 11898
rect 26056 11834 26108 11840
rect 26240 11280 26292 11286
rect 26240 11222 26292 11228
rect 25872 11212 25924 11218
rect 25872 11154 25924 11160
rect 26148 11212 26200 11218
rect 26148 11154 26200 11160
rect 25870 10840 25926 10849
rect 25870 10775 25926 10784
rect 25964 10804 26016 10810
rect 25884 10266 25912 10775
rect 25964 10746 26016 10752
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 25976 9926 26004 10746
rect 26160 10606 26188 11154
rect 26252 10606 26280 11222
rect 26148 10600 26200 10606
rect 26148 10542 26200 10548
rect 26240 10600 26292 10606
rect 26240 10542 26292 10548
rect 26160 10130 26188 10542
rect 26148 10124 26200 10130
rect 26148 10066 26200 10072
rect 26252 10062 26280 10542
rect 26056 10056 26108 10062
rect 26240 10056 26292 10062
rect 26108 10004 26188 10010
rect 26056 9998 26188 10004
rect 26240 9998 26292 10004
rect 26068 9982 26188 9998
rect 25964 9920 26016 9926
rect 25964 9862 26016 9868
rect 25872 9444 25924 9450
rect 25872 9386 25924 9392
rect 25884 8634 25912 9386
rect 25976 9042 26004 9862
rect 26054 9616 26110 9625
rect 26054 9551 26110 9560
rect 26068 9518 26096 9551
rect 26056 9512 26108 9518
rect 26056 9454 26108 9460
rect 26068 9110 26096 9454
rect 26056 9104 26108 9110
rect 26056 9046 26108 9052
rect 25964 9036 26016 9042
rect 25964 8978 26016 8984
rect 25872 8628 25924 8634
rect 25872 8570 25924 8576
rect 25962 8392 26018 8401
rect 25962 8327 26018 8336
rect 25976 7886 26004 8327
rect 26160 7970 26188 9982
rect 26160 7942 26280 7970
rect 25872 7880 25924 7886
rect 25872 7822 25924 7828
rect 25964 7880 26016 7886
rect 25964 7822 26016 7828
rect 25884 7206 25912 7822
rect 26056 7336 26108 7342
rect 26056 7278 26108 7284
rect 25872 7200 25924 7206
rect 25872 7142 25924 7148
rect 25964 6860 26016 6866
rect 25964 6802 26016 6808
rect 25870 6760 25926 6769
rect 25870 6695 25872 6704
rect 25924 6695 25926 6704
rect 25872 6666 25924 6672
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 25884 5166 25912 5646
rect 25976 5302 26004 6802
rect 26068 6798 26096 7278
rect 26252 6882 26280 7942
rect 26160 6854 26280 6882
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26068 6254 26096 6734
rect 26056 6248 26108 6254
rect 26056 6190 26108 6196
rect 26056 5840 26108 5846
rect 26056 5782 26108 5788
rect 25964 5296 26016 5302
rect 25964 5238 26016 5244
rect 25872 5160 25924 5166
rect 25872 5102 25924 5108
rect 26068 4826 26096 5782
rect 26160 5710 26188 6854
rect 26240 6656 26292 6662
rect 26238 6624 26240 6633
rect 26292 6624 26294 6633
rect 26238 6559 26294 6568
rect 26344 5846 26372 12582
rect 26528 12481 26556 13824
rect 26620 13326 26648 14962
rect 26712 14822 26740 15302
rect 26790 15263 26846 15272
rect 26700 14816 26752 14822
rect 26700 14758 26752 14764
rect 26790 14512 26846 14521
rect 26896 14498 26924 16730
rect 26963 16348 27271 16357
rect 26963 16346 26969 16348
rect 27025 16346 27049 16348
rect 27105 16346 27129 16348
rect 27185 16346 27209 16348
rect 27265 16346 27271 16348
rect 27025 16294 27027 16346
rect 27207 16294 27209 16346
rect 26963 16292 26969 16294
rect 27025 16292 27049 16294
rect 27105 16292 27129 16294
rect 27185 16292 27209 16294
rect 27265 16292 27271 16294
rect 26963 16283 27271 16292
rect 26963 15260 27271 15269
rect 26963 15258 26969 15260
rect 27025 15258 27049 15260
rect 27105 15258 27129 15260
rect 27185 15258 27209 15260
rect 27265 15258 27271 15260
rect 27025 15206 27027 15258
rect 27207 15206 27209 15258
rect 26963 15204 26969 15206
rect 27025 15204 27049 15206
rect 27105 15204 27129 15206
rect 27185 15204 27209 15206
rect 27265 15204 27271 15206
rect 26963 15195 27271 15204
rect 26846 14470 26924 14498
rect 27356 14482 27384 19128
rect 27436 18148 27488 18154
rect 27436 18090 27488 18096
rect 27448 17202 27476 18090
rect 27436 17196 27488 17202
rect 27436 17138 27488 17144
rect 27448 16833 27476 17138
rect 27434 16824 27490 16833
rect 27434 16759 27490 16768
rect 27632 16658 27660 19207
rect 27712 18624 27764 18630
rect 27712 18566 27764 18572
rect 27724 18057 27752 18566
rect 27804 18148 27856 18154
rect 27804 18090 27856 18096
rect 27710 18048 27766 18057
rect 27710 17983 27766 17992
rect 27816 17542 27844 18090
rect 27804 17536 27856 17542
rect 27724 17496 27804 17524
rect 27724 17134 27752 17496
rect 27804 17478 27856 17484
rect 27712 17128 27764 17134
rect 27712 17070 27764 17076
rect 27804 16788 27856 16794
rect 27804 16730 27856 16736
rect 27436 16652 27488 16658
rect 27436 16594 27488 16600
rect 27620 16652 27672 16658
rect 27620 16594 27672 16600
rect 27448 15706 27476 16594
rect 27528 16584 27580 16590
rect 27528 16526 27580 16532
rect 27436 15700 27488 15706
rect 27436 15642 27488 15648
rect 27436 15564 27488 15570
rect 27436 15506 27488 15512
rect 27344 14476 27396 14482
rect 26790 14447 26846 14456
rect 26698 14104 26754 14113
rect 26698 14039 26754 14048
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26608 12776 26660 12782
rect 26608 12718 26660 12724
rect 26514 12472 26570 12481
rect 26514 12407 26570 12416
rect 26528 9674 26556 12407
rect 26620 12306 26648 12718
rect 26712 12646 26740 14039
rect 26804 13977 26832 14447
rect 27344 14418 27396 14424
rect 26884 14408 26936 14414
rect 26884 14350 26936 14356
rect 26790 13968 26846 13977
rect 26896 13938 26924 14350
rect 26963 14172 27271 14181
rect 26963 14170 26969 14172
rect 27025 14170 27049 14172
rect 27105 14170 27129 14172
rect 27185 14170 27209 14172
rect 27265 14170 27271 14172
rect 27025 14118 27027 14170
rect 27207 14118 27209 14170
rect 26963 14116 26969 14118
rect 27025 14116 27049 14118
rect 27105 14116 27129 14118
rect 27185 14116 27209 14118
rect 27265 14116 27271 14118
rect 26963 14107 27271 14116
rect 27448 14056 27476 15506
rect 27540 15094 27568 16526
rect 27618 15600 27674 15609
rect 27618 15535 27674 15544
rect 27528 15088 27580 15094
rect 27528 15030 27580 15036
rect 27632 14074 27660 15535
rect 27816 14770 27844 16730
rect 27894 16280 27950 16289
rect 27894 16215 27950 16224
rect 27908 16114 27936 16215
rect 27896 16108 27948 16114
rect 27896 16050 27948 16056
rect 27896 15904 27948 15910
rect 27896 15846 27948 15852
rect 27908 15162 27936 15846
rect 28000 15570 28028 22034
rect 31300 21956 31352 21962
rect 31300 21898 31352 21904
rect 29000 21616 29052 21622
rect 29000 21558 29052 21564
rect 28356 21548 28408 21554
rect 28356 21490 28408 21496
rect 28080 21412 28132 21418
rect 28080 21354 28132 21360
rect 27988 15564 28040 15570
rect 27988 15506 28040 15512
rect 27988 15428 28040 15434
rect 27988 15370 28040 15376
rect 27896 15156 27948 15162
rect 27896 15098 27948 15104
rect 27816 14742 27936 14770
rect 27804 14612 27856 14618
rect 27804 14554 27856 14560
rect 27712 14476 27764 14482
rect 27712 14418 27764 14424
rect 27172 14028 27476 14056
rect 27528 14068 27580 14074
rect 26790 13903 26846 13912
rect 26884 13932 26936 13938
rect 26884 13874 26936 13880
rect 27068 13932 27120 13938
rect 27172 13920 27200 14028
rect 27528 14010 27580 14016
rect 27620 14068 27672 14074
rect 27620 14010 27672 14016
rect 27540 13954 27568 14010
rect 27540 13938 27660 13954
rect 27120 13892 27200 13920
rect 27344 13932 27396 13938
rect 27068 13874 27120 13880
rect 27540 13932 27672 13938
rect 27540 13926 27620 13932
rect 27344 13874 27396 13880
rect 27620 13874 27672 13880
rect 26792 13728 26844 13734
rect 26792 13670 26844 13676
rect 26804 12850 26832 13670
rect 26896 12986 26924 13874
rect 27356 13138 27384 13874
rect 27436 13864 27488 13870
rect 27488 13824 27568 13852
rect 27436 13806 27488 13812
rect 27356 13110 27476 13138
rect 26963 13084 27271 13093
rect 26963 13082 26969 13084
rect 27025 13082 27049 13084
rect 27105 13082 27129 13084
rect 27185 13082 27209 13084
rect 27265 13082 27271 13084
rect 27025 13030 27027 13082
rect 27207 13030 27209 13082
rect 26963 13028 26969 13030
rect 27025 13028 27049 13030
rect 27105 13028 27129 13030
rect 27185 13028 27209 13030
rect 27265 13028 27271 13030
rect 26963 13019 27271 13028
rect 26884 12980 26936 12986
rect 26884 12922 26936 12928
rect 26792 12844 26844 12850
rect 26792 12786 26844 12792
rect 26700 12640 26752 12646
rect 26700 12582 26752 12588
rect 26712 12306 26740 12582
rect 26804 12434 26832 12786
rect 27160 12436 27212 12442
rect 26804 12406 27160 12434
rect 26804 12374 26832 12406
rect 27160 12378 27212 12384
rect 26792 12368 26844 12374
rect 26792 12310 26844 12316
rect 26884 12368 26936 12374
rect 26884 12310 26936 12316
rect 26608 12300 26660 12306
rect 26608 12242 26660 12248
rect 26700 12300 26752 12306
rect 26700 12242 26752 12248
rect 26896 12220 26924 12310
rect 26804 12192 26924 12220
rect 26804 11898 26832 12192
rect 26963 11996 27271 12005
rect 26963 11994 26969 11996
rect 27025 11994 27049 11996
rect 27105 11994 27129 11996
rect 27185 11994 27209 11996
rect 27265 11994 27271 11996
rect 27025 11942 27027 11994
rect 27207 11942 27209 11994
rect 26963 11940 26969 11942
rect 27025 11940 27049 11942
rect 27105 11940 27129 11942
rect 27185 11940 27209 11942
rect 27265 11940 27271 11942
rect 26963 11931 27271 11940
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 26620 11150 26648 11494
rect 26608 11144 26660 11150
rect 26608 11086 26660 11092
rect 26436 9646 26556 9674
rect 26436 8106 26464 9646
rect 26516 9036 26568 9042
rect 26516 8978 26568 8984
rect 26528 8634 26556 8978
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26620 8498 26648 11086
rect 26712 9926 26740 11698
rect 26700 9920 26752 9926
rect 26700 9862 26752 9868
rect 26700 9512 26752 9518
rect 26700 9454 26752 9460
rect 26712 9178 26740 9454
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26700 8968 26752 8974
rect 26700 8910 26752 8916
rect 26608 8492 26660 8498
rect 26608 8434 26660 8440
rect 26436 8078 26556 8106
rect 26528 7177 26556 8078
rect 26712 7954 26740 8910
rect 26804 8430 26832 11834
rect 27160 11688 27212 11694
rect 27158 11656 27160 11665
rect 27212 11656 27214 11665
rect 27158 11591 27214 11600
rect 27344 11144 27396 11150
rect 27344 11086 27396 11092
rect 26963 10908 27271 10917
rect 26963 10906 26969 10908
rect 27025 10906 27049 10908
rect 27105 10906 27129 10908
rect 27185 10906 27209 10908
rect 27265 10906 27271 10908
rect 27025 10854 27027 10906
rect 27207 10854 27209 10906
rect 26963 10852 26969 10854
rect 27025 10852 27049 10854
rect 27105 10852 27129 10854
rect 27185 10852 27209 10854
rect 27265 10852 27271 10854
rect 26963 10843 27271 10852
rect 26884 10056 26936 10062
rect 26884 9998 26936 10004
rect 26896 9722 26924 9998
rect 26963 9820 27271 9829
rect 26963 9818 26969 9820
rect 27025 9818 27049 9820
rect 27105 9818 27129 9820
rect 27185 9818 27209 9820
rect 27265 9818 27271 9820
rect 27025 9766 27027 9818
rect 27207 9766 27209 9818
rect 26963 9764 26969 9766
rect 27025 9764 27049 9766
rect 27105 9764 27129 9766
rect 27185 9764 27209 9766
rect 27265 9764 27271 9766
rect 26963 9755 27271 9764
rect 26884 9716 26936 9722
rect 26884 9658 26936 9664
rect 27356 9382 27384 11086
rect 26884 9376 26936 9382
rect 26884 9318 26936 9324
rect 27344 9376 27396 9382
rect 27344 9318 27396 9324
rect 26896 9178 26924 9318
rect 26884 9172 26936 9178
rect 26884 9114 26936 9120
rect 26884 8968 26936 8974
rect 26884 8910 26936 8916
rect 27344 8968 27396 8974
rect 27344 8910 27396 8916
rect 26792 8424 26844 8430
rect 26792 8366 26844 8372
rect 26700 7948 26752 7954
rect 26700 7890 26752 7896
rect 26514 7168 26570 7177
rect 26514 7103 26570 7112
rect 26516 6860 26568 6866
rect 26516 6802 26568 6808
rect 26528 6769 26556 6802
rect 26514 6760 26570 6769
rect 26514 6695 26570 6704
rect 26516 6656 26568 6662
rect 26516 6598 26568 6604
rect 26424 6180 26476 6186
rect 26424 6122 26476 6128
rect 26332 5840 26384 5846
rect 26332 5782 26384 5788
rect 26148 5704 26200 5710
rect 26148 5646 26200 5652
rect 26148 5568 26200 5574
rect 26148 5510 26200 5516
rect 26056 4820 26108 4826
rect 26056 4762 26108 4768
rect 26160 4146 26188 5510
rect 26148 4140 26200 4146
rect 26148 4082 26200 4088
rect 26240 4072 26292 4078
rect 26240 4014 26292 4020
rect 26056 3936 26108 3942
rect 26056 3878 26108 3884
rect 25780 3596 25832 3602
rect 25780 3538 25832 3544
rect 26068 3194 26096 3878
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 26056 3188 26108 3194
rect 26056 3130 26108 3136
rect 26160 3126 26188 3538
rect 26148 3120 26200 3126
rect 26148 3062 26200 3068
rect 26160 2990 26188 3062
rect 26252 2990 26280 4014
rect 26330 3088 26386 3097
rect 26330 3023 26386 3032
rect 25688 2984 25740 2990
rect 25688 2926 25740 2932
rect 26148 2984 26200 2990
rect 26148 2926 26200 2932
rect 26240 2984 26292 2990
rect 26240 2926 26292 2932
rect 26252 2446 26280 2926
rect 25688 2440 25740 2446
rect 25688 2382 25740 2388
rect 26240 2440 26292 2446
rect 26240 2382 26292 2388
rect 25594 2136 25650 2145
rect 25594 2071 25650 2080
rect 24768 1964 24820 1970
rect 24768 1906 24820 1912
rect 25044 1964 25096 1970
rect 25044 1906 25096 1912
rect 24584 1760 24636 1766
rect 24584 1702 24636 1708
rect 24492 1556 24544 1562
rect 24492 1498 24544 1504
rect 24400 1216 24452 1222
rect 24400 1158 24452 1164
rect 24504 678 24532 1498
rect 25594 1456 25650 1465
rect 25700 1426 25728 2382
rect 26344 2106 26372 3023
rect 26436 2582 26464 6122
rect 26528 3670 26556 6598
rect 26608 6248 26660 6254
rect 26608 6190 26660 6196
rect 26620 5302 26648 6190
rect 26712 5914 26740 7890
rect 26896 7546 26924 8910
rect 26963 8732 27271 8741
rect 26963 8730 26969 8732
rect 27025 8730 27049 8732
rect 27105 8730 27129 8732
rect 27185 8730 27209 8732
rect 27265 8730 27271 8732
rect 27025 8678 27027 8730
rect 27207 8678 27209 8730
rect 26963 8676 26969 8678
rect 27025 8676 27049 8678
rect 27105 8676 27129 8678
rect 27185 8676 27209 8678
rect 27265 8676 27271 8678
rect 26963 8667 27271 8676
rect 27356 8634 27384 8910
rect 27448 8634 27476 13110
rect 27540 11898 27568 13824
rect 27724 13734 27752 14418
rect 27816 13870 27844 14554
rect 27804 13864 27856 13870
rect 27804 13806 27856 13812
rect 27712 13728 27764 13734
rect 27712 13670 27764 13676
rect 27804 13524 27856 13530
rect 27908 13512 27936 14742
rect 28000 14385 28028 15370
rect 27986 14376 28042 14385
rect 27986 14311 28042 14320
rect 27988 14272 28040 14278
rect 27988 14214 28040 14220
rect 27856 13484 27936 13512
rect 27804 13466 27856 13472
rect 28000 13394 28028 14214
rect 28092 13433 28120 21354
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28172 16652 28224 16658
rect 28172 16594 28224 16600
rect 28184 15162 28212 16594
rect 28172 15156 28224 15162
rect 28172 15098 28224 15104
rect 28078 13424 28134 13433
rect 27988 13388 28040 13394
rect 28078 13359 28134 13368
rect 27988 13330 28040 13336
rect 27712 12980 27764 12986
rect 27712 12922 27764 12928
rect 27724 12306 27752 12922
rect 28092 12764 28120 13359
rect 27908 12736 28120 12764
rect 27712 12300 27764 12306
rect 27712 12242 27764 12248
rect 27528 11892 27580 11898
rect 27528 11834 27580 11840
rect 27908 11218 27936 12736
rect 28184 12714 28212 15098
rect 28276 13258 28304 18702
rect 28264 13252 28316 13258
rect 28264 13194 28316 13200
rect 28172 12708 28224 12714
rect 28172 12650 28224 12656
rect 27988 12640 28040 12646
rect 27988 12582 28040 12588
rect 28080 12640 28132 12646
rect 28080 12582 28132 12588
rect 28000 11898 28028 12582
rect 28092 12306 28120 12582
rect 28080 12300 28132 12306
rect 28080 12242 28132 12248
rect 28262 12200 28318 12209
rect 28262 12135 28318 12144
rect 27988 11892 28040 11898
rect 27988 11834 28040 11840
rect 27896 11212 27948 11218
rect 27896 11154 27948 11160
rect 27528 11144 27580 11150
rect 27528 11086 27580 11092
rect 27540 9178 27568 11086
rect 28080 11076 28132 11082
rect 28080 11018 28132 11024
rect 27712 10464 27764 10470
rect 27712 10406 27764 10412
rect 27724 9722 27752 10406
rect 27712 9716 27764 9722
rect 27712 9658 27764 9664
rect 27528 9172 27580 9178
rect 27528 9114 27580 9120
rect 27710 8936 27766 8945
rect 27710 8871 27766 8880
rect 27344 8628 27396 8634
rect 27344 8570 27396 8576
rect 27436 8628 27488 8634
rect 27436 8570 27488 8576
rect 27068 8492 27120 8498
rect 27068 8434 27120 8440
rect 27080 8090 27108 8434
rect 27068 8084 27120 8090
rect 27068 8026 27120 8032
rect 27436 7812 27488 7818
rect 27436 7754 27488 7760
rect 27344 7744 27396 7750
rect 27344 7686 27396 7692
rect 26963 7644 27271 7653
rect 26963 7642 26969 7644
rect 27025 7642 27049 7644
rect 27105 7642 27129 7644
rect 27185 7642 27209 7644
rect 27265 7642 27271 7644
rect 27025 7590 27027 7642
rect 27207 7590 27209 7642
rect 26963 7588 26969 7590
rect 27025 7588 27049 7590
rect 27105 7588 27129 7590
rect 27185 7588 27209 7590
rect 27265 7588 27271 7590
rect 26963 7579 27271 7588
rect 26884 7540 26936 7546
rect 26884 7482 26936 7488
rect 26792 7336 26844 7342
rect 26792 7278 26844 7284
rect 26804 7002 26832 7278
rect 26884 7200 26936 7206
rect 27252 7200 27304 7206
rect 26884 7142 26936 7148
rect 27250 7168 27252 7177
rect 27304 7168 27306 7177
rect 26792 6996 26844 7002
rect 26792 6938 26844 6944
rect 26896 6100 26924 7142
rect 27250 7103 27306 7112
rect 26963 6556 27271 6565
rect 26963 6554 26969 6556
rect 27025 6554 27049 6556
rect 27105 6554 27129 6556
rect 27185 6554 27209 6556
rect 27265 6554 27271 6556
rect 27025 6502 27027 6554
rect 27207 6502 27209 6554
rect 26963 6500 26969 6502
rect 27025 6500 27049 6502
rect 27105 6500 27129 6502
rect 27185 6500 27209 6502
rect 27265 6500 27271 6502
rect 26963 6491 27271 6500
rect 27066 6352 27122 6361
rect 27066 6287 27122 6296
rect 26976 6112 27028 6118
rect 26896 6072 26976 6100
rect 26976 6054 27028 6060
rect 26700 5908 26752 5914
rect 26700 5850 26752 5856
rect 27080 5846 27108 6287
rect 27356 6118 27384 7686
rect 27160 6112 27212 6118
rect 27160 6054 27212 6060
rect 27344 6112 27396 6118
rect 27344 6054 27396 6060
rect 27068 5840 27120 5846
rect 26974 5808 27030 5817
rect 27068 5782 27120 5788
rect 26974 5743 26976 5752
rect 27028 5743 27030 5752
rect 26976 5714 27028 5720
rect 26792 5636 26844 5642
rect 26792 5578 26844 5584
rect 26700 5568 26752 5574
rect 26700 5510 26752 5516
rect 26608 5296 26660 5302
rect 26608 5238 26660 5244
rect 26608 4684 26660 4690
rect 26608 4626 26660 4632
rect 26620 4593 26648 4626
rect 26606 4584 26662 4593
rect 26606 4519 26662 4528
rect 26516 3664 26568 3670
rect 26516 3606 26568 3612
rect 26620 2990 26648 4519
rect 26712 4026 26740 5510
rect 26804 4146 26832 5578
rect 26884 5568 26936 5574
rect 27172 5556 27200 6054
rect 27344 5704 27396 5710
rect 27344 5646 27396 5652
rect 27356 5556 27384 5646
rect 27172 5528 27384 5556
rect 26884 5510 26936 5516
rect 26792 4140 26844 4146
rect 26792 4082 26844 4088
rect 26712 3998 26832 4026
rect 26700 3936 26752 3942
rect 26700 3878 26752 3884
rect 26712 3670 26740 3878
rect 26700 3664 26752 3670
rect 26700 3606 26752 3612
rect 26608 2984 26660 2990
rect 26608 2926 26660 2932
rect 26712 2854 26740 3606
rect 26804 3058 26832 3998
rect 26792 3052 26844 3058
rect 26792 2994 26844 3000
rect 26700 2848 26752 2854
rect 26700 2790 26752 2796
rect 26712 2650 26740 2790
rect 26896 2774 26924 5510
rect 26963 5468 27271 5477
rect 26963 5466 26969 5468
rect 27025 5466 27049 5468
rect 27105 5466 27129 5468
rect 27185 5466 27209 5468
rect 27265 5466 27271 5468
rect 27025 5414 27027 5466
rect 27207 5414 27209 5466
rect 26963 5412 26969 5414
rect 27025 5412 27049 5414
rect 27105 5412 27129 5414
rect 27185 5412 27209 5414
rect 27265 5412 27271 5414
rect 26963 5403 27271 5412
rect 27356 5030 27384 5528
rect 27448 5166 27476 7754
rect 27620 6928 27672 6934
rect 27620 6870 27672 6876
rect 27528 6792 27580 6798
rect 27528 6734 27580 6740
rect 27540 5914 27568 6734
rect 27632 6458 27660 6870
rect 27620 6452 27672 6458
rect 27620 6394 27672 6400
rect 27528 5908 27580 5914
rect 27528 5850 27580 5856
rect 27436 5160 27488 5166
rect 27436 5102 27488 5108
rect 27344 5024 27396 5030
rect 27344 4966 27396 4972
rect 27436 5024 27488 5030
rect 27436 4966 27488 4972
rect 27356 4826 27384 4966
rect 27252 4820 27304 4826
rect 27252 4762 27304 4768
rect 27344 4820 27396 4826
rect 27344 4762 27396 4768
rect 27264 4554 27292 4762
rect 27448 4758 27476 4966
rect 27436 4752 27488 4758
rect 27436 4694 27488 4700
rect 27540 4690 27568 5850
rect 27724 4758 27752 8871
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 27816 7886 27844 8230
rect 27988 8084 28040 8090
rect 27988 8026 28040 8032
rect 27804 7880 27856 7886
rect 27804 7822 27856 7828
rect 27896 7880 27948 7886
rect 27896 7822 27948 7828
rect 27816 6798 27844 7822
rect 27908 7546 27936 7822
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 27896 7200 27948 7206
rect 27896 7142 27948 7148
rect 27908 6905 27936 7142
rect 28000 7002 28028 8026
rect 27988 6996 28040 7002
rect 27988 6938 28040 6944
rect 27894 6896 27950 6905
rect 27894 6831 27950 6840
rect 28092 6798 28120 11018
rect 28172 10464 28224 10470
rect 28172 10406 28224 10412
rect 28184 7886 28212 10406
rect 28276 10198 28304 12135
rect 28368 12102 28396 21490
rect 28448 21344 28500 21350
rect 28448 21286 28500 21292
rect 28460 17270 28488 21286
rect 28722 20904 28778 20913
rect 28722 20839 28778 20848
rect 28540 19848 28592 19854
rect 28540 19790 28592 19796
rect 28552 19242 28580 19790
rect 28540 19236 28592 19242
rect 28540 19178 28592 19184
rect 28448 17264 28500 17270
rect 28448 17206 28500 17212
rect 28552 16794 28580 19178
rect 28632 17264 28684 17270
rect 28632 17206 28684 17212
rect 28736 17218 28764 20839
rect 29012 20262 29040 21558
rect 30380 21480 30432 21486
rect 30380 21422 30432 21428
rect 30564 21480 30616 21486
rect 30564 21422 30616 21428
rect 30288 21412 30340 21418
rect 30288 21354 30340 21360
rect 29736 21344 29788 21350
rect 29736 21286 29788 21292
rect 30104 21344 30156 21350
rect 30104 21286 30156 21292
rect 29460 20936 29512 20942
rect 29460 20878 29512 20884
rect 29644 20936 29696 20942
rect 29644 20878 29696 20884
rect 29368 20596 29420 20602
rect 29368 20538 29420 20544
rect 29380 20398 29408 20538
rect 29092 20392 29144 20398
rect 29092 20334 29144 20340
rect 29276 20392 29328 20398
rect 29276 20334 29328 20340
rect 29368 20392 29420 20398
rect 29368 20334 29420 20340
rect 29000 20256 29052 20262
rect 29000 20198 29052 20204
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 28908 18148 28960 18154
rect 28908 18090 28960 18096
rect 28816 18080 28868 18086
rect 28816 18022 28868 18028
rect 28828 17338 28856 18022
rect 28920 17882 28948 18090
rect 28908 17876 28960 17882
rect 28908 17818 28960 17824
rect 28908 17740 28960 17746
rect 28908 17682 28960 17688
rect 28816 17332 28868 17338
rect 28816 17274 28868 17280
rect 28920 17270 28948 17682
rect 28908 17264 28960 17270
rect 28540 16788 28592 16794
rect 28540 16730 28592 16736
rect 28448 16584 28500 16590
rect 28644 16561 28672 17206
rect 28736 17190 28856 17218
rect 28908 17206 28960 17212
rect 28448 16526 28500 16532
rect 28630 16552 28686 16561
rect 28460 12986 28488 16526
rect 28630 16487 28686 16496
rect 28540 15496 28592 15502
rect 28540 15438 28592 15444
rect 28552 15162 28580 15438
rect 28540 15156 28592 15162
rect 28540 15098 28592 15104
rect 28448 12980 28500 12986
rect 28448 12922 28500 12928
rect 28356 12096 28408 12102
rect 28356 12038 28408 12044
rect 28448 11212 28500 11218
rect 28448 11154 28500 11160
rect 28264 10192 28316 10198
rect 28264 10134 28316 10140
rect 28460 10130 28488 11154
rect 28540 10464 28592 10470
rect 28540 10406 28592 10412
rect 28356 10124 28408 10130
rect 28356 10066 28408 10072
rect 28448 10124 28500 10130
rect 28448 10066 28500 10072
rect 28264 9920 28316 9926
rect 28264 9862 28316 9868
rect 28276 8498 28304 9862
rect 28368 9654 28396 10066
rect 28356 9648 28408 9654
rect 28356 9590 28408 9596
rect 28552 9586 28580 10406
rect 28540 9580 28592 9586
rect 28540 9522 28592 9528
rect 28552 8974 28580 9522
rect 28644 9042 28672 16487
rect 28722 16280 28778 16289
rect 28722 16215 28778 16224
rect 28736 16114 28764 16215
rect 28724 16108 28776 16114
rect 28724 16050 28776 16056
rect 28722 16008 28778 16017
rect 28722 15943 28724 15952
rect 28776 15943 28778 15952
rect 28724 15914 28776 15920
rect 28828 12986 28856 17190
rect 29012 16810 29040 19790
rect 29104 19242 29132 20334
rect 29184 19712 29236 19718
rect 29184 19654 29236 19660
rect 29196 19417 29224 19654
rect 29182 19408 29238 19417
rect 29182 19343 29238 19352
rect 29288 19310 29316 20334
rect 29380 19446 29408 20334
rect 29368 19440 29420 19446
rect 29368 19382 29420 19388
rect 29276 19304 29328 19310
rect 29276 19246 29328 19252
rect 29092 19236 29144 19242
rect 29092 19178 29144 19184
rect 29104 18086 29132 19178
rect 29184 18828 29236 18834
rect 29288 18816 29316 19246
rect 29380 18834 29408 19382
rect 29236 18788 29316 18816
rect 29368 18828 29420 18834
rect 29184 18770 29236 18776
rect 29368 18770 29420 18776
rect 29196 18222 29224 18770
rect 29276 18624 29328 18630
rect 29276 18566 29328 18572
rect 29184 18216 29236 18222
rect 29184 18158 29236 18164
rect 29092 18080 29144 18086
rect 29092 18022 29144 18028
rect 29104 17134 29132 18022
rect 29196 17746 29224 18158
rect 29184 17740 29236 17746
rect 29184 17682 29236 17688
rect 29196 17202 29224 17682
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 29092 17128 29144 17134
rect 29092 17070 29144 17076
rect 29012 16782 29224 16810
rect 29000 16652 29052 16658
rect 29000 16594 29052 16600
rect 28908 16448 28960 16454
rect 28908 16390 28960 16396
rect 28920 15094 28948 16390
rect 28908 15088 28960 15094
rect 28908 15030 28960 15036
rect 29012 14074 29040 16594
rect 29092 16176 29144 16182
rect 29092 16118 29144 16124
rect 29104 15065 29132 16118
rect 29090 15056 29146 15065
rect 29090 14991 29146 15000
rect 29104 14890 29132 14991
rect 29092 14884 29144 14890
rect 29092 14826 29144 14832
rect 29092 14272 29144 14278
rect 29092 14214 29144 14220
rect 29000 14068 29052 14074
rect 29000 14010 29052 14016
rect 28906 13968 28962 13977
rect 28906 13903 28962 13912
rect 28920 13410 28948 13903
rect 29104 13870 29132 14214
rect 29092 13864 29144 13870
rect 29092 13806 29144 13812
rect 29000 13728 29052 13734
rect 29000 13670 29052 13676
rect 29012 13530 29040 13670
rect 29000 13524 29052 13530
rect 29000 13466 29052 13472
rect 28920 13382 29132 13410
rect 29104 13326 29132 13382
rect 29092 13320 29144 13326
rect 29092 13262 29144 13268
rect 28908 13184 28960 13190
rect 28908 13126 28960 13132
rect 28816 12980 28868 12986
rect 28816 12922 28868 12928
rect 28724 12232 28776 12238
rect 28724 12174 28776 12180
rect 28816 12232 28868 12238
rect 28816 12174 28868 12180
rect 28736 11778 28764 12174
rect 28828 11898 28856 12174
rect 28816 11892 28868 11898
rect 28816 11834 28868 11840
rect 28736 11750 28856 11778
rect 28724 10532 28776 10538
rect 28724 10474 28776 10480
rect 28632 9036 28684 9042
rect 28632 8978 28684 8984
rect 28540 8968 28592 8974
rect 28540 8910 28592 8916
rect 28736 8498 28764 10474
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 28724 8492 28776 8498
rect 28724 8434 28776 8440
rect 28828 8090 28856 11750
rect 28920 11218 28948 13126
rect 29000 12776 29052 12782
rect 29000 12718 29052 12724
rect 29012 12238 29040 12718
rect 29000 12232 29052 12238
rect 29000 12174 29052 12180
rect 28908 11212 28960 11218
rect 28908 11154 28960 11160
rect 28908 10464 28960 10470
rect 28908 10406 28960 10412
rect 28920 9926 28948 10406
rect 28908 9920 28960 9926
rect 28908 9862 28960 9868
rect 28816 8084 28868 8090
rect 28816 8026 28868 8032
rect 28920 7970 28948 9862
rect 29000 9444 29052 9450
rect 29000 9386 29052 9392
rect 29012 8838 29040 9386
rect 29000 8832 29052 8838
rect 29000 8774 29052 8780
rect 28828 7942 28948 7970
rect 28172 7880 28224 7886
rect 28172 7822 28224 7828
rect 28264 7540 28316 7546
rect 28264 7482 28316 7488
rect 28276 7206 28304 7482
rect 28356 7404 28408 7410
rect 28408 7364 28488 7392
rect 28356 7346 28408 7352
rect 28264 7200 28316 7206
rect 28316 7160 28396 7188
rect 28264 7142 28316 7148
rect 27804 6792 27856 6798
rect 27804 6734 27856 6740
rect 28080 6792 28132 6798
rect 28080 6734 28132 6740
rect 28172 6384 28224 6390
rect 28170 6352 28172 6361
rect 28224 6352 28226 6361
rect 28170 6287 28226 6296
rect 27804 6112 27856 6118
rect 27804 6054 27856 6060
rect 27816 5778 27844 6054
rect 27804 5772 27856 5778
rect 27804 5714 27856 5720
rect 28172 5704 28224 5710
rect 28170 5672 28172 5681
rect 28224 5672 28226 5681
rect 28170 5607 28226 5616
rect 28172 5568 28224 5574
rect 28172 5510 28224 5516
rect 27896 5228 27948 5234
rect 27896 5170 27948 5176
rect 27712 4752 27764 4758
rect 27712 4694 27764 4700
rect 27344 4684 27396 4690
rect 27344 4626 27396 4632
rect 27528 4684 27580 4690
rect 27528 4626 27580 4632
rect 27252 4548 27304 4554
rect 27252 4490 27304 4496
rect 26963 4380 27271 4389
rect 26963 4378 26969 4380
rect 27025 4378 27049 4380
rect 27105 4378 27129 4380
rect 27185 4378 27209 4380
rect 27265 4378 27271 4380
rect 27025 4326 27027 4378
rect 27207 4326 27209 4378
rect 26963 4324 26969 4326
rect 27025 4324 27049 4326
rect 27105 4324 27129 4326
rect 27185 4324 27209 4326
rect 27265 4324 27271 4326
rect 26963 4315 27271 4324
rect 27356 4282 27384 4626
rect 27344 4276 27396 4282
rect 27344 4218 27396 4224
rect 27344 4072 27396 4078
rect 27344 4014 27396 4020
rect 27356 3738 27384 4014
rect 27540 3738 27568 4626
rect 27344 3732 27396 3738
rect 27344 3674 27396 3680
rect 27528 3732 27580 3738
rect 27528 3674 27580 3680
rect 27436 3664 27488 3670
rect 27436 3606 27488 3612
rect 26963 3292 27271 3301
rect 26963 3290 26969 3292
rect 27025 3290 27049 3292
rect 27105 3290 27129 3292
rect 27185 3290 27209 3292
rect 27265 3290 27271 3292
rect 27025 3238 27027 3290
rect 27207 3238 27209 3290
rect 26963 3236 26969 3238
rect 27025 3236 27049 3238
rect 27105 3236 27129 3238
rect 27185 3236 27209 3238
rect 27265 3236 27271 3238
rect 26963 3227 27271 3236
rect 27344 2848 27396 2854
rect 27344 2790 27396 2796
rect 26896 2746 27108 2774
rect 26700 2644 26752 2650
rect 26700 2586 26752 2592
rect 26424 2576 26476 2582
rect 26424 2518 26476 2524
rect 27080 2514 27108 2746
rect 27068 2508 27120 2514
rect 27068 2450 27120 2456
rect 26976 2440 27028 2446
rect 26896 2400 26976 2428
rect 26608 2304 26660 2310
rect 26608 2246 26660 2252
rect 26332 2100 26384 2106
rect 26332 2042 26384 2048
rect 26238 1864 26294 1873
rect 26294 1822 26372 1850
rect 26238 1799 26294 1808
rect 25594 1391 25596 1400
rect 25648 1391 25650 1400
rect 25688 1420 25740 1426
rect 25596 1362 25648 1368
rect 25688 1362 25740 1368
rect 24584 1352 24636 1358
rect 25700 1329 25728 1362
rect 24584 1294 24636 1300
rect 25686 1320 25742 1329
rect 24596 1018 24624 1294
rect 26344 1290 26372 1822
rect 26620 1426 26648 2246
rect 26896 1986 26924 2400
rect 26976 2382 27028 2388
rect 26963 2204 27271 2213
rect 26963 2202 26969 2204
rect 27025 2202 27049 2204
rect 27105 2202 27129 2204
rect 27185 2202 27209 2204
rect 27265 2202 27271 2204
rect 27025 2150 27027 2202
rect 27207 2150 27209 2202
rect 26963 2148 26969 2150
rect 27025 2148 27049 2150
rect 27105 2148 27129 2150
rect 27185 2148 27209 2150
rect 27265 2148 27271 2150
rect 26963 2139 27271 2148
rect 26896 1958 27016 1986
rect 27356 1970 27384 2790
rect 27448 2106 27476 3606
rect 27526 3496 27582 3505
rect 27526 3431 27582 3440
rect 27540 3074 27568 3431
rect 27540 3058 27660 3074
rect 27540 3052 27672 3058
rect 27540 3046 27620 3052
rect 27436 2100 27488 2106
rect 27436 2042 27488 2048
rect 26988 1902 27016 1958
rect 27344 1964 27396 1970
rect 27344 1906 27396 1912
rect 26976 1896 27028 1902
rect 26976 1838 27028 1844
rect 26988 1426 27016 1838
rect 27068 1760 27120 1766
rect 27120 1708 27292 1714
rect 27068 1702 27292 1708
rect 27080 1686 27292 1702
rect 27264 1562 27292 1686
rect 27252 1556 27304 1562
rect 27252 1498 27304 1504
rect 27448 1426 27476 2042
rect 27540 1766 27568 3046
rect 27620 2994 27672 3000
rect 27908 2106 27936 5170
rect 28080 3936 28132 3942
rect 28080 3878 28132 3884
rect 27896 2100 27948 2106
rect 27896 2042 27948 2048
rect 27804 1896 27856 1902
rect 27804 1838 27856 1844
rect 27528 1760 27580 1766
rect 27528 1702 27580 1708
rect 27712 1760 27764 1766
rect 27712 1702 27764 1708
rect 27540 1562 27568 1702
rect 27528 1556 27580 1562
rect 27528 1498 27580 1504
rect 26608 1420 26660 1426
rect 26608 1362 26660 1368
rect 26976 1420 27028 1426
rect 26976 1362 27028 1368
rect 27436 1420 27488 1426
rect 27436 1362 27488 1368
rect 25686 1255 25742 1264
rect 26332 1284 26384 1290
rect 26332 1226 26384 1232
rect 25686 1048 25742 1057
rect 24584 1012 24636 1018
rect 25686 983 25688 992
rect 24584 954 24636 960
rect 25740 983 25742 992
rect 25688 954 25740 960
rect 26344 814 26372 1226
rect 26700 1216 26752 1222
rect 26700 1158 26752 1164
rect 26884 1216 26936 1222
rect 26884 1158 26936 1164
rect 26712 1018 26740 1158
rect 26700 1012 26752 1018
rect 26700 954 26752 960
rect 26896 882 26924 1158
rect 26963 1116 27271 1125
rect 26963 1114 26969 1116
rect 27025 1114 27049 1116
rect 27105 1114 27129 1116
rect 27185 1114 27209 1116
rect 27265 1114 27271 1116
rect 27025 1062 27027 1114
rect 27207 1062 27209 1114
rect 26963 1060 26969 1062
rect 27025 1060 27049 1062
rect 27105 1060 27129 1062
rect 27185 1060 27209 1062
rect 27265 1060 27271 1062
rect 26963 1051 27271 1060
rect 27448 898 27476 1362
rect 26884 876 26936 882
rect 26884 818 26936 824
rect 27356 870 27476 898
rect 27356 814 27384 870
rect 26332 808 26384 814
rect 26332 750 26384 756
rect 27344 808 27396 814
rect 27344 750 27396 756
rect 27540 678 27568 1498
rect 27724 1358 27752 1702
rect 27816 1426 27844 1838
rect 27804 1420 27856 1426
rect 27804 1362 27856 1368
rect 28092 1358 28120 3878
rect 28184 1358 28212 5510
rect 28264 4820 28316 4826
rect 28264 4762 28316 4768
rect 28276 3738 28304 4762
rect 28264 3732 28316 3738
rect 28264 3674 28316 3680
rect 28368 3618 28396 7160
rect 28276 3590 28396 3618
rect 28276 2990 28304 3590
rect 28356 3528 28408 3534
rect 28356 3470 28408 3476
rect 28264 2984 28316 2990
rect 28368 2961 28396 3470
rect 28264 2926 28316 2932
rect 28354 2952 28410 2961
rect 28354 2887 28410 2896
rect 28460 2774 28488 7364
rect 28540 7200 28592 7206
rect 28540 7142 28592 7148
rect 28552 6322 28580 7142
rect 28540 6316 28592 6322
rect 28540 6258 28592 6264
rect 28632 6248 28684 6254
rect 28632 6190 28684 6196
rect 28644 5386 28672 6190
rect 28552 5358 28672 5386
rect 28552 4298 28580 5358
rect 28630 5264 28686 5273
rect 28630 5199 28686 5208
rect 28644 4468 28672 5199
rect 28828 4570 28856 7942
rect 28908 7472 28960 7478
rect 28908 7414 28960 7420
rect 28920 4690 28948 7414
rect 29012 7410 29040 8774
rect 29104 8430 29132 13262
rect 29196 12442 29224 16782
rect 29288 15706 29316 18566
rect 29380 18222 29408 18770
rect 29368 18216 29420 18222
rect 29368 18158 29420 18164
rect 29380 17270 29408 18158
rect 29368 17264 29420 17270
rect 29368 17206 29420 17212
rect 29368 16992 29420 16998
rect 29368 16934 29420 16940
rect 29380 16153 29408 16934
rect 29366 16144 29422 16153
rect 29366 16079 29422 16088
rect 29380 16046 29408 16079
rect 29368 16040 29420 16046
rect 29368 15982 29420 15988
rect 29368 15904 29420 15910
rect 29366 15872 29368 15881
rect 29420 15872 29422 15881
rect 29366 15807 29422 15816
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 29276 15360 29328 15366
rect 29274 15328 29276 15337
rect 29328 15328 29330 15337
rect 29274 15263 29330 15272
rect 29472 15042 29500 20878
rect 29552 19848 29604 19854
rect 29552 19790 29604 19796
rect 29288 15014 29500 15042
rect 29288 14618 29316 15014
rect 29368 14952 29420 14958
rect 29368 14894 29420 14900
rect 29276 14612 29328 14618
rect 29276 14554 29328 14560
rect 29276 14408 29328 14414
rect 29276 14350 29328 14356
rect 29184 12436 29236 12442
rect 29184 12378 29236 12384
rect 29288 11898 29316 14350
rect 29380 13530 29408 14894
rect 29564 14074 29592 19790
rect 29656 16794 29684 20878
rect 29748 18834 29776 21286
rect 29828 20256 29880 20262
rect 29828 20198 29880 20204
rect 29736 18828 29788 18834
rect 29736 18770 29788 18776
rect 29736 18624 29788 18630
rect 29736 18566 29788 18572
rect 29748 18086 29776 18566
rect 29736 18080 29788 18086
rect 29736 18022 29788 18028
rect 29748 17814 29776 18022
rect 29736 17808 29788 17814
rect 29736 17750 29788 17756
rect 29736 17332 29788 17338
rect 29736 17274 29788 17280
rect 29644 16788 29696 16794
rect 29644 16730 29696 16736
rect 29644 16040 29696 16046
rect 29642 16008 29644 16017
rect 29696 16008 29698 16017
rect 29642 15943 29698 15952
rect 29644 15904 29696 15910
rect 29644 15846 29696 15852
rect 29656 15745 29684 15846
rect 29642 15736 29698 15745
rect 29642 15671 29698 15680
rect 29644 15564 29696 15570
rect 29644 15506 29696 15512
rect 29656 15026 29684 15506
rect 29644 15020 29696 15026
rect 29644 14962 29696 14968
rect 29656 14278 29684 14962
rect 29748 14958 29776 17274
rect 29840 16046 29868 20198
rect 29920 19372 29972 19378
rect 29920 19314 29972 19320
rect 29828 16040 29880 16046
rect 29828 15982 29880 15988
rect 29736 14952 29788 14958
rect 29736 14894 29788 14900
rect 29644 14272 29696 14278
rect 29644 14214 29696 14220
rect 29552 14068 29604 14074
rect 29552 14010 29604 14016
rect 29840 13954 29868 15982
rect 29932 14346 29960 19314
rect 30012 19236 30064 19242
rect 30012 19178 30064 19184
rect 30024 16538 30052 19178
rect 30116 17610 30144 21286
rect 30196 20256 30248 20262
rect 30196 20198 30248 20204
rect 30208 20058 30236 20198
rect 30196 20052 30248 20058
rect 30196 19994 30248 20000
rect 30300 19718 30328 21354
rect 30288 19712 30340 19718
rect 30288 19654 30340 19660
rect 30300 19258 30328 19654
rect 30208 19230 30328 19258
rect 30208 18834 30236 19230
rect 30300 19174 30328 19230
rect 30288 19168 30340 19174
rect 30288 19110 30340 19116
rect 30196 18828 30248 18834
rect 30196 18770 30248 18776
rect 30208 18329 30236 18770
rect 30288 18624 30340 18630
rect 30288 18566 30340 18572
rect 30194 18320 30250 18329
rect 30194 18255 30250 18264
rect 30194 18184 30250 18193
rect 30194 18119 30250 18128
rect 30208 18086 30236 18119
rect 30196 18080 30248 18086
rect 30196 18022 30248 18028
rect 30104 17604 30156 17610
rect 30104 17546 30156 17552
rect 30208 16726 30236 18022
rect 30300 17066 30328 18566
rect 30392 18290 30420 21422
rect 30472 19236 30524 19242
rect 30472 19178 30524 19184
rect 30380 18284 30432 18290
rect 30380 18226 30432 18232
rect 30288 17060 30340 17066
rect 30288 17002 30340 17008
rect 30392 16794 30420 18226
rect 30484 17678 30512 19178
rect 30472 17672 30524 17678
rect 30470 17640 30472 17649
rect 30524 17640 30526 17649
rect 30470 17575 30526 17584
rect 30576 17338 30604 21422
rect 30758 21244 31066 21253
rect 30758 21242 30764 21244
rect 30820 21242 30844 21244
rect 30900 21242 30924 21244
rect 30980 21242 31004 21244
rect 31060 21242 31066 21244
rect 30820 21190 30822 21242
rect 31002 21190 31004 21242
rect 30758 21188 30764 21190
rect 30820 21188 30844 21190
rect 30900 21188 30924 21190
rect 30980 21188 31004 21190
rect 31060 21188 31066 21190
rect 30758 21179 31066 21188
rect 31208 20256 31260 20262
rect 31208 20198 31260 20204
rect 30758 20156 31066 20165
rect 30758 20154 30764 20156
rect 30820 20154 30844 20156
rect 30900 20154 30924 20156
rect 30980 20154 31004 20156
rect 31060 20154 31066 20156
rect 30820 20102 30822 20154
rect 31002 20102 31004 20154
rect 30758 20100 30764 20102
rect 30820 20100 30844 20102
rect 30900 20100 30924 20102
rect 30980 20100 31004 20102
rect 31060 20100 31066 20102
rect 30758 20091 31066 20100
rect 30656 19372 30708 19378
rect 30656 19314 30708 19320
rect 30564 17332 30616 17338
rect 30564 17274 30616 17280
rect 30472 17128 30524 17134
rect 30472 17070 30524 17076
rect 30380 16788 30432 16794
rect 30380 16730 30432 16736
rect 30196 16720 30248 16726
rect 30196 16662 30248 16668
rect 30024 16510 30144 16538
rect 30012 14952 30064 14958
rect 30010 14920 30012 14929
rect 30064 14920 30066 14929
rect 30010 14855 30066 14864
rect 29920 14340 29972 14346
rect 29920 14282 29972 14288
rect 30116 14074 30144 16510
rect 30392 16266 30420 16730
rect 30300 16238 30420 16266
rect 30196 16176 30248 16182
rect 30196 16118 30248 16124
rect 30208 14657 30236 16118
rect 30194 14648 30250 14657
rect 30194 14583 30250 14592
rect 30300 14074 30328 16238
rect 30378 16008 30434 16017
rect 30378 15943 30434 15952
rect 30392 15162 30420 15943
rect 30380 15156 30432 15162
rect 30380 15098 30432 15104
rect 30380 14816 30432 14822
rect 30380 14758 30432 14764
rect 30104 14068 30156 14074
rect 30104 14010 30156 14016
rect 30288 14068 30340 14074
rect 30288 14010 30340 14016
rect 29564 13926 29868 13954
rect 29920 14000 29972 14006
rect 29920 13942 29972 13948
rect 29368 13524 29420 13530
rect 29368 13466 29420 13472
rect 29564 13394 29592 13926
rect 29828 13864 29880 13870
rect 29656 13832 29828 13852
rect 29880 13832 29882 13841
rect 29656 13824 29826 13832
rect 29368 13388 29420 13394
rect 29368 13330 29420 13336
rect 29552 13388 29604 13394
rect 29552 13330 29604 13336
rect 29276 11892 29328 11898
rect 29276 11834 29328 11840
rect 29276 11756 29328 11762
rect 29276 11698 29328 11704
rect 29184 11552 29236 11558
rect 29184 11494 29236 11500
rect 29196 9518 29224 11494
rect 29288 10674 29316 11698
rect 29380 11354 29408 13330
rect 29552 12708 29604 12714
rect 29552 12650 29604 12656
rect 29564 12617 29592 12650
rect 29550 12608 29606 12617
rect 29550 12543 29606 12552
rect 29550 12472 29606 12481
rect 29550 12407 29606 12416
rect 29368 11348 29420 11354
rect 29368 11290 29420 11296
rect 29276 10668 29328 10674
rect 29276 10610 29328 10616
rect 29276 10464 29328 10470
rect 29276 10406 29328 10412
rect 29184 9512 29236 9518
rect 29184 9454 29236 9460
rect 29092 8424 29144 8430
rect 29092 8366 29144 8372
rect 29184 8288 29236 8294
rect 29184 8230 29236 8236
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 29196 7206 29224 8230
rect 29288 7954 29316 10406
rect 29460 9376 29512 9382
rect 29460 9318 29512 9324
rect 29276 7948 29328 7954
rect 29276 7890 29328 7896
rect 29368 7744 29420 7750
rect 29368 7686 29420 7692
rect 29184 7200 29236 7206
rect 29184 7142 29236 7148
rect 29276 7200 29328 7206
rect 29276 7142 29328 7148
rect 28998 6760 29054 6769
rect 28998 6695 29054 6704
rect 29012 5302 29040 6695
rect 29000 5296 29052 5302
rect 29000 5238 29052 5244
rect 29092 5092 29144 5098
rect 29092 5034 29144 5040
rect 29000 5024 29052 5030
rect 29000 4966 29052 4972
rect 28908 4684 28960 4690
rect 28908 4626 28960 4632
rect 28828 4542 28948 4570
rect 28644 4440 28856 4468
rect 28552 4270 28764 4298
rect 28630 4040 28686 4049
rect 28630 3975 28686 3984
rect 28644 3194 28672 3975
rect 28632 3188 28684 3194
rect 28632 3130 28684 3136
rect 28460 2746 28580 2774
rect 28264 2304 28316 2310
rect 28264 2246 28316 2252
rect 27712 1352 27764 1358
rect 27712 1294 27764 1300
rect 28080 1352 28132 1358
rect 28080 1294 28132 1300
rect 28172 1352 28224 1358
rect 28172 1294 28224 1300
rect 28276 882 28304 2246
rect 28552 1018 28580 2746
rect 28736 2106 28764 4270
rect 28828 2650 28856 4440
rect 28816 2644 28868 2650
rect 28816 2586 28868 2592
rect 28816 2508 28868 2514
rect 28816 2450 28868 2456
rect 28632 2100 28684 2106
rect 28632 2042 28684 2048
rect 28724 2100 28776 2106
rect 28724 2042 28776 2048
rect 28644 1562 28672 2042
rect 28828 1766 28856 2450
rect 28920 1902 28948 4542
rect 28908 1896 28960 1902
rect 28908 1838 28960 1844
rect 29012 1850 29040 4966
rect 29104 4282 29132 5034
rect 29092 4276 29144 4282
rect 29092 4218 29144 4224
rect 29196 2666 29224 7142
rect 29288 6798 29316 7142
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29276 6112 29328 6118
rect 29276 6054 29328 6060
rect 29104 2638 29224 2666
rect 29104 2582 29132 2638
rect 29092 2576 29144 2582
rect 29092 2518 29144 2524
rect 29090 2408 29146 2417
rect 29090 2343 29092 2352
rect 29144 2343 29146 2352
rect 29092 2314 29144 2320
rect 29184 2032 29236 2038
rect 29182 2000 29184 2009
rect 29236 2000 29238 2009
rect 29288 1970 29316 6054
rect 29380 5914 29408 7686
rect 29472 7478 29500 9318
rect 29564 8362 29592 12407
rect 29656 11626 29684 13824
rect 29826 13767 29882 13776
rect 29932 13308 29960 13942
rect 30392 13870 30420 14758
rect 30380 13864 30432 13870
rect 30208 13824 30380 13852
rect 30104 13796 30156 13802
rect 30104 13738 30156 13744
rect 29748 13280 29960 13308
rect 29748 11830 29776 13280
rect 29918 13152 29974 13161
rect 29918 13087 29974 13096
rect 29826 12880 29882 12889
rect 29826 12815 29882 12824
rect 29840 12782 29868 12815
rect 29932 12782 29960 13087
rect 30116 12918 30144 13738
rect 30104 12912 30156 12918
rect 30104 12854 30156 12860
rect 29828 12776 29880 12782
rect 29828 12718 29880 12724
rect 29920 12776 29972 12782
rect 29920 12718 29972 12724
rect 30010 12744 30066 12753
rect 30010 12679 30066 12688
rect 30024 12646 30052 12679
rect 30012 12640 30064 12646
rect 30012 12582 30064 12588
rect 30208 12434 30236 13824
rect 30380 13806 30432 13812
rect 30116 12406 30236 12434
rect 29736 11824 29788 11830
rect 29736 11766 29788 11772
rect 29644 11620 29696 11626
rect 29644 11562 29696 11568
rect 29920 11620 29972 11626
rect 29920 11562 29972 11568
rect 29932 10538 29960 11562
rect 30116 11558 30144 12406
rect 30378 12336 30434 12345
rect 30378 12271 30380 12280
rect 30432 12271 30434 12280
rect 30380 12242 30432 12248
rect 30104 11552 30156 11558
rect 30104 11494 30156 11500
rect 30012 11076 30064 11082
rect 30012 11018 30064 11024
rect 29920 10532 29972 10538
rect 29920 10474 29972 10480
rect 29644 10464 29696 10470
rect 29644 10406 29696 10412
rect 29552 8356 29604 8362
rect 29552 8298 29604 8304
rect 29460 7472 29512 7478
rect 29460 7414 29512 7420
rect 29368 5908 29420 5914
rect 29368 5850 29420 5856
rect 29366 5128 29422 5137
rect 29366 5063 29422 5072
rect 29380 2650 29408 5063
rect 29472 3194 29500 7414
rect 29460 3188 29512 3194
rect 29460 3130 29512 3136
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 29460 2576 29512 2582
rect 29460 2518 29512 2524
rect 29182 1935 29238 1944
rect 29276 1964 29328 1970
rect 29276 1906 29328 1912
rect 29012 1822 29132 1850
rect 28816 1760 28868 1766
rect 28816 1702 28868 1708
rect 28632 1556 28684 1562
rect 28632 1498 28684 1504
rect 28540 1012 28592 1018
rect 28540 954 28592 960
rect 29000 944 29052 950
rect 29000 886 29052 892
rect 28264 876 28316 882
rect 28264 818 28316 824
rect 29012 785 29040 886
rect 29104 882 29132 1822
rect 29472 1442 29500 2518
rect 29564 2446 29592 8298
rect 29656 6866 29684 10406
rect 29736 8356 29788 8362
rect 29736 8298 29788 8304
rect 29644 6860 29696 6866
rect 29644 6802 29696 6808
rect 29748 3482 29776 8298
rect 29828 7744 29880 7750
rect 29828 7686 29880 7692
rect 29840 3602 29868 7686
rect 29932 5166 29960 10474
rect 30024 9042 30052 11018
rect 30116 10470 30144 11494
rect 30104 10464 30156 10470
rect 30104 10406 30156 10412
rect 30116 9926 30144 10406
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 30484 9178 30512 17070
rect 30576 14618 30604 17274
rect 30668 15978 30696 19314
rect 30758 19068 31066 19077
rect 30758 19066 30764 19068
rect 30820 19066 30844 19068
rect 30900 19066 30924 19068
rect 30980 19066 31004 19068
rect 31060 19066 31066 19068
rect 30820 19014 30822 19066
rect 31002 19014 31004 19066
rect 30758 19012 30764 19014
rect 30820 19012 30844 19014
rect 30900 19012 30924 19014
rect 30980 19012 31004 19014
rect 31060 19012 31066 19014
rect 30758 19003 31066 19012
rect 30758 17980 31066 17989
rect 30758 17978 30764 17980
rect 30820 17978 30844 17980
rect 30900 17978 30924 17980
rect 30980 17978 31004 17980
rect 31060 17978 31066 17980
rect 30820 17926 30822 17978
rect 31002 17926 31004 17978
rect 30758 17924 30764 17926
rect 30820 17924 30844 17926
rect 30900 17924 30924 17926
rect 30980 17924 31004 17926
rect 31060 17924 31066 17926
rect 30758 17915 31066 17924
rect 31116 17060 31168 17066
rect 31116 17002 31168 17008
rect 30758 16892 31066 16901
rect 30758 16890 30764 16892
rect 30820 16890 30844 16892
rect 30900 16890 30924 16892
rect 30980 16890 31004 16892
rect 31060 16890 31066 16892
rect 30820 16838 30822 16890
rect 31002 16838 31004 16890
rect 30758 16836 30764 16838
rect 30820 16836 30844 16838
rect 30900 16836 30924 16838
rect 30980 16836 31004 16838
rect 31060 16836 31066 16838
rect 30758 16827 31066 16836
rect 30656 15972 30708 15978
rect 30656 15914 30708 15920
rect 30758 15804 31066 15813
rect 30758 15802 30764 15804
rect 30820 15802 30844 15804
rect 30900 15802 30924 15804
rect 30980 15802 31004 15804
rect 31060 15802 31066 15804
rect 30820 15750 30822 15802
rect 31002 15750 31004 15802
rect 30758 15748 30764 15750
rect 30820 15748 30844 15750
rect 30900 15748 30924 15750
rect 30980 15748 31004 15750
rect 31060 15748 31066 15750
rect 30758 15739 31066 15748
rect 30758 14716 31066 14725
rect 30758 14714 30764 14716
rect 30820 14714 30844 14716
rect 30900 14714 30924 14716
rect 30980 14714 31004 14716
rect 31060 14714 31066 14716
rect 30820 14662 30822 14714
rect 31002 14662 31004 14714
rect 30758 14660 30764 14662
rect 30820 14660 30844 14662
rect 30900 14660 30924 14662
rect 30980 14660 31004 14662
rect 31060 14660 31066 14662
rect 30758 14651 31066 14660
rect 30564 14612 30616 14618
rect 30564 14554 30616 14560
rect 30576 13734 30604 14554
rect 30656 14408 30708 14414
rect 30656 14350 30708 14356
rect 30564 13728 30616 13734
rect 30564 13670 30616 13676
rect 30472 9172 30524 9178
rect 30472 9114 30524 9120
rect 30012 9036 30064 9042
rect 30012 8978 30064 8984
rect 30012 8288 30064 8294
rect 30012 8230 30064 8236
rect 30024 7954 30052 8230
rect 30012 7948 30064 7954
rect 30012 7890 30064 7896
rect 29920 5160 29972 5166
rect 29920 5102 29972 5108
rect 29828 3596 29880 3602
rect 29828 3538 29880 3544
rect 29748 3454 29868 3482
rect 29736 3188 29788 3194
rect 29736 3130 29788 3136
rect 29748 2514 29776 3130
rect 29736 2508 29788 2514
rect 29736 2450 29788 2456
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 29380 1414 29500 1442
rect 29748 1426 29776 2450
rect 29736 1420 29788 1426
rect 29092 876 29144 882
rect 29092 818 29144 824
rect 29380 814 29408 1414
rect 29736 1362 29788 1368
rect 29458 1320 29514 1329
rect 29458 1255 29514 1264
rect 29472 1018 29500 1255
rect 29840 1222 29868 3454
rect 30024 1902 30052 7890
rect 30668 6866 30696 14350
rect 30758 13628 31066 13637
rect 30758 13626 30764 13628
rect 30820 13626 30844 13628
rect 30900 13626 30924 13628
rect 30980 13626 31004 13628
rect 31060 13626 31066 13628
rect 30820 13574 30822 13626
rect 31002 13574 31004 13626
rect 30758 13572 30764 13574
rect 30820 13572 30844 13574
rect 30900 13572 30924 13574
rect 30980 13572 31004 13574
rect 31060 13572 31066 13574
rect 30758 13563 31066 13572
rect 30758 12540 31066 12549
rect 30758 12538 30764 12540
rect 30820 12538 30844 12540
rect 30900 12538 30924 12540
rect 30980 12538 31004 12540
rect 31060 12538 31066 12540
rect 30820 12486 30822 12538
rect 31002 12486 31004 12538
rect 30758 12484 30764 12486
rect 30820 12484 30844 12486
rect 30900 12484 30924 12486
rect 30980 12484 31004 12486
rect 31060 12484 31066 12486
rect 30758 12475 31066 12484
rect 30758 11452 31066 11461
rect 30758 11450 30764 11452
rect 30820 11450 30844 11452
rect 30900 11450 30924 11452
rect 30980 11450 31004 11452
rect 31060 11450 31066 11452
rect 30820 11398 30822 11450
rect 31002 11398 31004 11450
rect 30758 11396 30764 11398
rect 30820 11396 30844 11398
rect 30900 11396 30924 11398
rect 30980 11396 31004 11398
rect 31060 11396 31066 11398
rect 30758 11387 31066 11396
rect 31128 11121 31156 17002
rect 31220 16250 31248 20198
rect 31208 16244 31260 16250
rect 31208 16186 31260 16192
rect 31208 14272 31260 14278
rect 31208 14214 31260 14220
rect 31114 11112 31170 11121
rect 31114 11047 31170 11056
rect 30758 10364 31066 10373
rect 30758 10362 30764 10364
rect 30820 10362 30844 10364
rect 30900 10362 30924 10364
rect 30980 10362 31004 10364
rect 31060 10362 31066 10364
rect 30820 10310 30822 10362
rect 31002 10310 31004 10362
rect 30758 10308 30764 10310
rect 30820 10308 30844 10310
rect 30900 10308 30924 10310
rect 30980 10308 31004 10310
rect 31060 10308 31066 10310
rect 30758 10299 31066 10308
rect 30758 9276 31066 9285
rect 30758 9274 30764 9276
rect 30820 9274 30844 9276
rect 30900 9274 30924 9276
rect 30980 9274 31004 9276
rect 31060 9274 31066 9276
rect 30820 9222 30822 9274
rect 31002 9222 31004 9274
rect 30758 9220 30764 9222
rect 30820 9220 30844 9222
rect 30900 9220 30924 9222
rect 30980 9220 31004 9222
rect 31060 9220 31066 9222
rect 30758 9211 31066 9220
rect 30758 8188 31066 8197
rect 30758 8186 30764 8188
rect 30820 8186 30844 8188
rect 30900 8186 30924 8188
rect 30980 8186 31004 8188
rect 31060 8186 31066 8188
rect 30820 8134 30822 8186
rect 31002 8134 31004 8186
rect 30758 8132 30764 8134
rect 30820 8132 30844 8134
rect 30900 8132 30924 8134
rect 30980 8132 31004 8134
rect 31060 8132 31066 8134
rect 30758 8123 31066 8132
rect 30758 7100 31066 7109
rect 30758 7098 30764 7100
rect 30820 7098 30844 7100
rect 30900 7098 30924 7100
rect 30980 7098 31004 7100
rect 31060 7098 31066 7100
rect 30820 7046 30822 7098
rect 31002 7046 31004 7098
rect 30758 7044 30764 7046
rect 30820 7044 30844 7046
rect 30900 7044 30924 7046
rect 30980 7044 31004 7046
rect 31060 7044 31066 7046
rect 30758 7035 31066 7044
rect 30656 6860 30708 6866
rect 30656 6802 30708 6808
rect 30758 6012 31066 6021
rect 30758 6010 30764 6012
rect 30820 6010 30844 6012
rect 30900 6010 30924 6012
rect 30980 6010 31004 6012
rect 31060 6010 31066 6012
rect 30820 5958 30822 6010
rect 31002 5958 31004 6010
rect 30758 5956 30764 5958
rect 30820 5956 30844 5958
rect 30900 5956 30924 5958
rect 30980 5956 31004 5958
rect 31060 5956 31066 5958
rect 30758 5947 31066 5956
rect 31220 5302 31248 14214
rect 31312 12986 31340 21898
rect 31390 17232 31446 17241
rect 31390 17167 31446 17176
rect 31404 14958 31432 17167
rect 31392 14952 31444 14958
rect 31392 14894 31444 14900
rect 31300 12980 31352 12986
rect 31300 12922 31352 12928
rect 31208 5296 31260 5302
rect 31208 5238 31260 5244
rect 30758 4924 31066 4933
rect 30758 4922 30764 4924
rect 30820 4922 30844 4924
rect 30900 4922 30924 4924
rect 30980 4922 31004 4924
rect 31060 4922 31066 4924
rect 30820 4870 30822 4922
rect 31002 4870 31004 4922
rect 30758 4868 30764 4870
rect 30820 4868 30844 4870
rect 30900 4868 30924 4870
rect 30980 4868 31004 4870
rect 31060 4868 31066 4870
rect 30758 4859 31066 4868
rect 30758 3836 31066 3845
rect 30758 3834 30764 3836
rect 30820 3834 30844 3836
rect 30900 3834 30924 3836
rect 30980 3834 31004 3836
rect 31060 3834 31066 3836
rect 30820 3782 30822 3834
rect 31002 3782 31004 3834
rect 30758 3780 30764 3782
rect 30820 3780 30844 3782
rect 30900 3780 30924 3782
rect 30980 3780 31004 3782
rect 31060 3780 31066 3782
rect 30758 3771 31066 3780
rect 30758 2748 31066 2757
rect 30758 2746 30764 2748
rect 30820 2746 30844 2748
rect 30900 2746 30924 2748
rect 30980 2746 31004 2748
rect 31060 2746 31066 2748
rect 30820 2694 30822 2746
rect 31002 2694 31004 2746
rect 30758 2692 30764 2694
rect 30820 2692 30844 2694
rect 30900 2692 30924 2694
rect 30980 2692 31004 2694
rect 31060 2692 31066 2694
rect 30758 2683 31066 2692
rect 30012 1896 30064 1902
rect 30012 1838 30064 1844
rect 30758 1660 31066 1669
rect 30758 1658 30764 1660
rect 30820 1658 30844 1660
rect 30900 1658 30924 1660
rect 30980 1658 31004 1660
rect 31060 1658 31066 1660
rect 30820 1606 30822 1658
rect 31002 1606 31004 1658
rect 30758 1604 30764 1606
rect 30820 1604 30844 1606
rect 30900 1604 30924 1606
rect 30980 1604 31004 1606
rect 31060 1604 31066 1606
rect 30758 1595 31066 1604
rect 29828 1216 29880 1222
rect 29828 1158 29880 1164
rect 29920 1216 29972 1222
rect 29920 1158 29972 1164
rect 29460 1012 29512 1018
rect 29460 954 29512 960
rect 29368 808 29420 814
rect 28998 776 29054 785
rect 29368 750 29420 756
rect 28998 711 29054 720
rect 24492 672 24544 678
rect 24492 614 24544 620
rect 27528 672 27580 678
rect 27528 614 27580 620
rect 24308 468 24360 474
rect 24308 410 24360 416
rect 29932 377 29960 1158
rect 30758 572 31066 581
rect 30758 570 30764 572
rect 30820 570 30844 572
rect 30900 570 30924 572
rect 30980 570 31004 572
rect 31060 570 31066 572
rect 30820 518 30822 570
rect 31002 518 31004 570
rect 30758 516 30764 518
rect 30820 516 30844 518
rect 30900 516 30924 518
rect 30980 516 31004 518
rect 31060 516 31066 518
rect 30758 507 31066 516
rect 29918 368 29974 377
rect 29918 303 29974 312
rect 22100 128 22152 134
rect 22100 70 22152 76
rect 24216 128 24268 134
rect 24216 70 24268 76
rect 3884 60 3936 66
rect 3884 2 3936 8
rect 16212 60 16264 66
rect 16212 2 16264 8
rect 18880 60 18932 66
rect 18880 2 18932 8
<< via2 >>
rect 2502 21936 2558 21992
rect 846 21528 902 21584
rect 4199 21786 4255 21788
rect 4279 21786 4335 21788
rect 4359 21786 4415 21788
rect 4439 21786 4495 21788
rect 4199 21734 4245 21786
rect 4245 21734 4255 21786
rect 4279 21734 4309 21786
rect 4309 21734 4321 21786
rect 4321 21734 4335 21786
rect 4359 21734 4373 21786
rect 4373 21734 4385 21786
rect 4385 21734 4415 21786
rect 4439 21734 4449 21786
rect 4449 21734 4495 21786
rect 4199 21732 4255 21734
rect 4279 21732 4335 21734
rect 4359 21732 4415 21734
rect 4439 21732 4495 21734
rect 1858 20984 1914 21040
rect 662 19760 718 19816
rect 1674 19352 1730 19408
rect 1122 17856 1178 17912
rect 1030 17720 1086 17776
rect 662 14456 718 14512
rect 1674 13812 1676 13832
rect 1676 13812 1728 13832
rect 1728 13812 1730 13832
rect 1674 13776 1730 13812
rect 2042 17040 2098 17096
rect 1950 13504 2006 13560
rect 1766 12552 1822 12608
rect 1950 12280 2006 12336
rect 2410 16632 2466 16688
rect 2226 15952 2282 16008
rect 2226 12688 2282 12744
rect 2134 11736 2190 11792
rect 2134 10668 2190 10704
rect 2134 10648 2136 10668
rect 2136 10648 2188 10668
rect 2188 10648 2190 10668
rect 1030 7792 1086 7848
rect 1122 6024 1178 6080
rect 938 4664 994 4720
rect 1122 1400 1178 1456
rect 1766 6740 1768 6760
rect 1768 6740 1820 6760
rect 1820 6740 1822 6760
rect 1766 6704 1822 6740
rect 2042 8064 2098 8120
rect 2594 16088 2650 16144
rect 3146 17856 3202 17912
rect 2594 8472 2650 8528
rect 2226 3712 2282 3768
rect 2962 15408 3018 15464
rect 3514 18400 3570 18456
rect 3330 17992 3386 18048
rect 3514 18264 3570 18320
rect 4066 20884 4068 20904
rect 4068 20884 4120 20904
rect 4120 20884 4122 20904
rect 4066 20848 4122 20884
rect 4199 20698 4255 20700
rect 4279 20698 4335 20700
rect 4359 20698 4415 20700
rect 4439 20698 4495 20700
rect 4199 20646 4245 20698
rect 4245 20646 4255 20698
rect 4279 20646 4309 20698
rect 4309 20646 4321 20698
rect 4321 20646 4335 20698
rect 4359 20646 4373 20698
rect 4373 20646 4385 20698
rect 4385 20646 4415 20698
rect 4439 20646 4449 20698
rect 4449 20646 4495 20698
rect 4199 20644 4255 20646
rect 4279 20644 4335 20646
rect 4359 20644 4415 20646
rect 4439 20644 4495 20646
rect 4710 20340 4712 20360
rect 4712 20340 4764 20360
rect 4764 20340 4766 20360
rect 4710 20304 4766 20340
rect 4199 19610 4255 19612
rect 4279 19610 4335 19612
rect 4359 19610 4415 19612
rect 4439 19610 4495 19612
rect 4199 19558 4245 19610
rect 4245 19558 4255 19610
rect 4279 19558 4309 19610
rect 4309 19558 4321 19610
rect 4321 19558 4335 19610
rect 4359 19558 4373 19610
rect 4373 19558 4385 19610
rect 4385 19558 4415 19610
rect 4439 19558 4449 19610
rect 4449 19558 4495 19610
rect 4199 19556 4255 19558
rect 4279 19556 4335 19558
rect 4359 19556 4415 19558
rect 4439 19556 4495 19558
rect 3606 14864 3662 14920
rect 2962 14320 3018 14376
rect 2870 11600 2926 11656
rect 3054 12844 3110 12880
rect 3054 12824 3056 12844
rect 3056 12824 3108 12844
rect 3108 12824 3110 12844
rect 2778 7248 2834 7304
rect 2962 8200 3018 8256
rect 2962 7404 3018 7440
rect 2962 7384 2964 7404
rect 2964 7384 3016 7404
rect 3016 7384 3018 7404
rect 2962 6840 3018 6896
rect 3606 13368 3662 13424
rect 3606 13232 3662 13288
rect 3790 18264 3846 18320
rect 4434 19216 4490 19272
rect 4342 18944 4398 19000
rect 4618 19080 4674 19136
rect 5078 22208 5134 22264
rect 11150 22244 11152 22264
rect 11152 22244 11204 22264
rect 11204 22244 11206 22264
rect 4250 18672 4306 18728
rect 4434 18672 4490 18728
rect 4802 18808 4858 18864
rect 4199 18522 4255 18524
rect 4279 18522 4335 18524
rect 4359 18522 4415 18524
rect 4439 18522 4495 18524
rect 4199 18470 4245 18522
rect 4245 18470 4255 18522
rect 4279 18470 4309 18522
rect 4309 18470 4321 18522
rect 4321 18470 4335 18522
rect 4359 18470 4373 18522
rect 4373 18470 4385 18522
rect 4385 18470 4415 18522
rect 4439 18470 4449 18522
rect 4449 18470 4495 18522
rect 4199 18468 4255 18470
rect 4279 18468 4335 18470
rect 4359 18468 4415 18470
rect 4439 18468 4495 18470
rect 5446 19352 5502 19408
rect 4526 18128 4582 18184
rect 4894 18128 4950 18184
rect 4526 17584 4582 17640
rect 4199 17434 4255 17436
rect 4279 17434 4335 17436
rect 4359 17434 4415 17436
rect 4439 17434 4495 17436
rect 4199 17382 4245 17434
rect 4245 17382 4255 17434
rect 4279 17382 4309 17434
rect 4309 17382 4321 17434
rect 4321 17382 4335 17434
rect 4359 17382 4373 17434
rect 4373 17382 4385 17434
rect 4385 17382 4415 17434
rect 4439 17382 4449 17434
rect 4449 17382 4495 17434
rect 4199 17380 4255 17382
rect 4279 17380 4335 17382
rect 4359 17380 4415 17382
rect 4439 17380 4495 17382
rect 3974 16632 4030 16688
rect 4199 16346 4255 16348
rect 4279 16346 4335 16348
rect 4359 16346 4415 16348
rect 4439 16346 4495 16348
rect 4199 16294 4245 16346
rect 4245 16294 4255 16346
rect 4279 16294 4309 16346
rect 4309 16294 4321 16346
rect 4321 16294 4335 16346
rect 4359 16294 4373 16346
rect 4373 16294 4385 16346
rect 4385 16294 4415 16346
rect 4439 16294 4449 16346
rect 4449 16294 4495 16346
rect 4199 16292 4255 16294
rect 4279 16292 4335 16294
rect 4359 16292 4415 16294
rect 4439 16292 4495 16294
rect 4199 15258 4255 15260
rect 4279 15258 4335 15260
rect 4359 15258 4415 15260
rect 4439 15258 4495 15260
rect 4199 15206 4245 15258
rect 4245 15206 4255 15258
rect 4279 15206 4309 15258
rect 4309 15206 4321 15258
rect 4321 15206 4335 15258
rect 4359 15206 4373 15258
rect 4373 15206 4385 15258
rect 4385 15206 4415 15258
rect 4439 15206 4449 15258
rect 4449 15206 4495 15258
rect 4199 15204 4255 15206
rect 4279 15204 4335 15206
rect 4359 15204 4415 15206
rect 4439 15204 4495 15206
rect 4158 14592 4214 14648
rect 4199 14170 4255 14172
rect 4279 14170 4335 14172
rect 4359 14170 4415 14172
rect 4439 14170 4495 14172
rect 4199 14118 4245 14170
rect 4245 14118 4255 14170
rect 4279 14118 4309 14170
rect 4309 14118 4321 14170
rect 4321 14118 4335 14170
rect 4359 14118 4373 14170
rect 4373 14118 4385 14170
rect 4385 14118 4415 14170
rect 4439 14118 4449 14170
rect 4449 14118 4495 14170
rect 4199 14116 4255 14118
rect 4279 14116 4335 14118
rect 4359 14116 4415 14118
rect 4439 14116 4495 14118
rect 4199 13082 4255 13084
rect 4279 13082 4335 13084
rect 4359 13082 4415 13084
rect 4439 13082 4495 13084
rect 4199 13030 4245 13082
rect 4245 13030 4255 13082
rect 4279 13030 4309 13082
rect 4309 13030 4321 13082
rect 4321 13030 4335 13082
rect 4359 13030 4373 13082
rect 4373 13030 4385 13082
rect 4385 13030 4415 13082
rect 4439 13030 4449 13082
rect 4449 13030 4495 13082
rect 4199 13028 4255 13030
rect 4279 13028 4335 13030
rect 4359 13028 4415 13030
rect 4439 13028 4495 13030
rect 4199 11994 4255 11996
rect 4279 11994 4335 11996
rect 4359 11994 4415 11996
rect 4439 11994 4495 11996
rect 4199 11942 4245 11994
rect 4245 11942 4255 11994
rect 4279 11942 4309 11994
rect 4309 11942 4321 11994
rect 4321 11942 4335 11994
rect 4359 11942 4373 11994
rect 4373 11942 4385 11994
rect 4385 11942 4415 11994
rect 4439 11942 4449 11994
rect 4449 11942 4495 11994
rect 4199 11940 4255 11942
rect 4279 11940 4335 11942
rect 4359 11940 4415 11942
rect 4439 11940 4495 11942
rect 3698 11192 3754 11248
rect 5262 18128 5318 18184
rect 5262 17992 5318 18048
rect 5170 17856 5226 17912
rect 5170 13912 5226 13968
rect 5078 13096 5134 13152
rect 4894 12960 4950 13016
rect 4199 10906 4255 10908
rect 4279 10906 4335 10908
rect 4359 10906 4415 10908
rect 4439 10906 4495 10908
rect 4199 10854 4245 10906
rect 4245 10854 4255 10906
rect 4279 10854 4309 10906
rect 4309 10854 4321 10906
rect 4321 10854 4335 10906
rect 4359 10854 4373 10906
rect 4373 10854 4385 10906
rect 4385 10854 4415 10906
rect 4439 10854 4449 10906
rect 4449 10854 4495 10906
rect 4199 10852 4255 10854
rect 4279 10852 4335 10854
rect 4359 10852 4415 10854
rect 4439 10852 4495 10854
rect 4199 9818 4255 9820
rect 4279 9818 4335 9820
rect 4359 9818 4415 9820
rect 4439 9818 4495 9820
rect 4199 9766 4245 9818
rect 4245 9766 4255 9818
rect 4279 9766 4309 9818
rect 4309 9766 4321 9818
rect 4321 9766 4335 9818
rect 4359 9766 4373 9818
rect 4373 9766 4385 9818
rect 4385 9766 4415 9818
rect 4439 9766 4449 9818
rect 4449 9766 4495 9818
rect 4199 9764 4255 9766
rect 4279 9764 4335 9766
rect 4359 9764 4415 9766
rect 4439 9764 4495 9766
rect 4986 9968 5042 10024
rect 3330 7948 3386 7984
rect 3330 7928 3332 7948
rect 3332 7928 3384 7948
rect 3384 7928 3386 7948
rect 3330 7792 3386 7848
rect 3238 4664 3294 4720
rect 3238 4528 3294 4584
rect 2686 3984 2742 4040
rect 2686 3712 2742 3768
rect 3422 5752 3478 5808
rect 4199 8730 4255 8732
rect 4279 8730 4335 8732
rect 4359 8730 4415 8732
rect 4439 8730 4495 8732
rect 4199 8678 4245 8730
rect 4245 8678 4255 8730
rect 4279 8678 4309 8730
rect 4309 8678 4321 8730
rect 4321 8678 4335 8730
rect 4359 8678 4373 8730
rect 4373 8678 4385 8730
rect 4385 8678 4415 8730
rect 4439 8678 4449 8730
rect 4449 8678 4495 8730
rect 4199 8676 4255 8678
rect 4279 8676 4335 8678
rect 4359 8676 4415 8678
rect 4439 8676 4495 8678
rect 4199 7642 4255 7644
rect 4279 7642 4335 7644
rect 4359 7642 4415 7644
rect 4439 7642 4495 7644
rect 4199 7590 4245 7642
rect 4245 7590 4255 7642
rect 4279 7590 4309 7642
rect 4309 7590 4321 7642
rect 4321 7590 4335 7642
rect 4359 7590 4373 7642
rect 4373 7590 4385 7642
rect 4385 7590 4415 7642
rect 4439 7590 4449 7642
rect 4449 7590 4495 7642
rect 4199 7588 4255 7590
rect 4279 7588 4335 7590
rect 4359 7588 4415 7590
rect 4439 7588 4495 7590
rect 4066 6840 4122 6896
rect 4199 6554 4255 6556
rect 4279 6554 4335 6556
rect 4359 6554 4415 6556
rect 4439 6554 4495 6556
rect 4199 6502 4245 6554
rect 4245 6502 4255 6554
rect 4279 6502 4309 6554
rect 4309 6502 4321 6554
rect 4321 6502 4335 6554
rect 4359 6502 4373 6554
rect 4373 6502 4385 6554
rect 4385 6502 4415 6554
rect 4439 6502 4449 6554
rect 4449 6502 4495 6554
rect 4199 6500 4255 6502
rect 4279 6500 4335 6502
rect 4359 6500 4415 6502
rect 4439 6500 4495 6502
rect 4199 5466 4255 5468
rect 4279 5466 4335 5468
rect 4359 5466 4415 5468
rect 4439 5466 4495 5468
rect 4199 5414 4245 5466
rect 4245 5414 4255 5466
rect 4279 5414 4309 5466
rect 4309 5414 4321 5466
rect 4321 5414 4335 5466
rect 4359 5414 4373 5466
rect 4373 5414 4385 5466
rect 4385 5414 4415 5466
rect 4439 5414 4449 5466
rect 4449 5414 4495 5466
rect 4199 5412 4255 5414
rect 4279 5412 4335 5414
rect 4359 5412 4415 5414
rect 4439 5412 4495 5414
rect 3330 2624 3386 2680
rect 3514 3848 3570 3904
rect 3514 3712 3570 3768
rect 3882 3984 3938 4040
rect 3974 3712 4030 3768
rect 4199 4378 4255 4380
rect 4279 4378 4335 4380
rect 4359 4378 4415 4380
rect 4439 4378 4495 4380
rect 4199 4326 4245 4378
rect 4245 4326 4255 4378
rect 4279 4326 4309 4378
rect 4309 4326 4321 4378
rect 4321 4326 4335 4378
rect 4359 4326 4373 4378
rect 4373 4326 4385 4378
rect 4385 4326 4415 4378
rect 4439 4326 4449 4378
rect 4449 4326 4495 4378
rect 4199 4324 4255 4326
rect 4279 4324 4335 4326
rect 4359 4324 4415 4326
rect 4439 4324 4495 4326
rect 4710 3848 4766 3904
rect 4986 6160 5042 6216
rect 11150 22208 11206 22244
rect 5814 19896 5870 19952
rect 5998 20576 6054 20632
rect 6550 20712 6606 20768
rect 5538 18400 5594 18456
rect 5998 19116 6000 19136
rect 6000 19116 6052 19136
rect 6052 19116 6054 19136
rect 5998 19080 6054 19116
rect 5538 18284 5594 18320
rect 5538 18264 5540 18284
rect 5540 18264 5592 18284
rect 5592 18264 5594 18284
rect 5446 17176 5502 17232
rect 5814 18672 5870 18728
rect 6734 19488 6790 19544
rect 6550 19352 6606 19408
rect 6090 18672 6146 18728
rect 5998 17992 6054 18048
rect 5906 17720 5962 17776
rect 5722 16360 5778 16416
rect 5906 14048 5962 14104
rect 5446 13776 5502 13832
rect 5722 12416 5778 12472
rect 6642 18808 6698 18864
rect 6918 19916 6974 19952
rect 6918 19896 6920 19916
rect 6920 19896 6972 19916
rect 6972 19896 6974 19916
rect 8574 21800 8630 21856
rect 10046 22072 10102 22128
rect 10966 22072 11022 22128
rect 8482 21256 8538 21312
rect 7994 21242 8050 21244
rect 8074 21242 8130 21244
rect 8154 21242 8210 21244
rect 8234 21242 8290 21244
rect 7994 21190 8040 21242
rect 8040 21190 8050 21242
rect 8074 21190 8104 21242
rect 8104 21190 8116 21242
rect 8116 21190 8130 21242
rect 8154 21190 8168 21242
rect 8168 21190 8180 21242
rect 8180 21190 8210 21242
rect 8234 21190 8244 21242
rect 8244 21190 8290 21242
rect 7994 21188 8050 21190
rect 8074 21188 8130 21190
rect 8154 21188 8210 21190
rect 8234 21188 8290 21190
rect 7286 19760 7342 19816
rect 8390 20168 8446 20224
rect 7994 20154 8050 20156
rect 8074 20154 8130 20156
rect 8154 20154 8210 20156
rect 8234 20154 8290 20156
rect 7994 20102 8040 20154
rect 8040 20102 8050 20154
rect 8074 20102 8104 20154
rect 8104 20102 8116 20154
rect 8116 20102 8130 20154
rect 8154 20102 8168 20154
rect 8168 20102 8180 20154
rect 8180 20102 8210 20154
rect 8234 20102 8244 20154
rect 8244 20102 8290 20154
rect 7994 20100 8050 20102
rect 8074 20100 8130 20102
rect 8154 20100 8210 20102
rect 8234 20100 8290 20102
rect 9310 21256 9366 21312
rect 8758 20984 8814 21040
rect 8850 20576 8906 20632
rect 6918 18536 6974 18592
rect 6918 18264 6974 18320
rect 7378 18264 7434 18320
rect 6826 17992 6882 18048
rect 6090 15136 6146 15192
rect 6642 15544 6698 15600
rect 6642 15272 6698 15328
rect 6550 15020 6606 15056
rect 6550 15000 6552 15020
rect 6552 15000 6604 15020
rect 6604 15000 6606 15020
rect 6274 14728 6330 14784
rect 6182 14184 6238 14240
rect 6550 14476 6606 14512
rect 6550 14456 6552 14476
rect 6552 14456 6604 14476
rect 6604 14456 6606 14476
rect 5354 8608 5410 8664
rect 5630 8880 5686 8936
rect 3698 3576 3754 3632
rect 3882 3440 3938 3496
rect 4199 3290 4255 3292
rect 4279 3290 4335 3292
rect 4359 3290 4415 3292
rect 4439 3290 4495 3292
rect 4199 3238 4245 3290
rect 4245 3238 4255 3290
rect 4279 3238 4309 3290
rect 4309 3238 4321 3290
rect 4321 3238 4335 3290
rect 4359 3238 4373 3290
rect 4373 3238 4385 3290
rect 4385 3238 4415 3290
rect 4439 3238 4449 3290
rect 4449 3238 4495 3290
rect 4199 3236 4255 3238
rect 4279 3236 4335 3238
rect 4359 3236 4415 3238
rect 4439 3236 4495 3238
rect 4526 3052 4582 3088
rect 4526 3032 4528 3052
rect 4528 3032 4580 3052
rect 4580 3032 4582 3052
rect 3698 2760 3754 2816
rect 4526 2508 4582 2544
rect 4526 2488 4528 2508
rect 4528 2488 4580 2508
rect 4580 2488 4582 2508
rect 4199 2202 4255 2204
rect 4279 2202 4335 2204
rect 4359 2202 4415 2204
rect 4439 2202 4495 2204
rect 4199 2150 4245 2202
rect 4245 2150 4255 2202
rect 4279 2150 4309 2202
rect 4309 2150 4321 2202
rect 4321 2150 4335 2202
rect 4359 2150 4373 2202
rect 4373 2150 4385 2202
rect 4385 2150 4415 2202
rect 4439 2150 4449 2202
rect 4449 2150 4495 2202
rect 4199 2148 4255 2150
rect 4279 2148 4335 2150
rect 4359 2148 4415 2150
rect 4439 2148 4495 2150
rect 5170 5344 5226 5400
rect 4986 3612 4988 3632
rect 4988 3612 5040 3632
rect 5040 3612 5042 3632
rect 4986 3576 5042 3612
rect 4250 1964 4306 2000
rect 4250 1944 4252 1964
rect 4252 1944 4304 1964
rect 4304 1944 4306 1964
rect 4618 1672 4674 1728
rect 4066 1300 4068 1320
rect 4068 1300 4120 1320
rect 4120 1300 4122 1320
rect 4066 1264 4122 1300
rect 4199 1114 4255 1116
rect 4279 1114 4335 1116
rect 4359 1114 4415 1116
rect 4439 1114 4495 1116
rect 4199 1062 4245 1114
rect 4245 1062 4255 1114
rect 4279 1062 4309 1114
rect 4309 1062 4321 1114
rect 4321 1062 4335 1114
rect 4359 1062 4373 1114
rect 4373 1062 4385 1114
rect 4385 1062 4415 1114
rect 4439 1062 4449 1114
rect 4449 1062 4495 1114
rect 4199 1060 4255 1062
rect 4279 1060 4335 1062
rect 4359 1060 4415 1062
rect 4439 1060 4495 1062
rect 5354 6432 5410 6488
rect 6734 14592 6790 14648
rect 7286 14728 7342 14784
rect 8206 19372 8262 19408
rect 8206 19352 8208 19372
rect 8208 19352 8260 19372
rect 8260 19352 8262 19372
rect 7562 18264 7618 18320
rect 7746 18536 7802 18592
rect 7470 17856 7526 17912
rect 7010 13776 7066 13832
rect 6734 13232 6790 13288
rect 6366 12416 6422 12472
rect 5538 6024 5594 6080
rect 5538 5072 5594 5128
rect 6182 7384 6238 7440
rect 7470 13504 7526 13560
rect 7102 12416 7158 12472
rect 7194 11620 7250 11656
rect 7194 11600 7196 11620
rect 7196 11600 7248 11620
rect 7248 11600 7250 11620
rect 7994 19066 8050 19068
rect 8074 19066 8130 19068
rect 8154 19066 8210 19068
rect 8234 19066 8290 19068
rect 7994 19014 8040 19066
rect 8040 19014 8050 19066
rect 8074 19014 8104 19066
rect 8104 19014 8116 19066
rect 8116 19014 8130 19066
rect 8154 19014 8168 19066
rect 8168 19014 8180 19066
rect 8180 19014 8210 19066
rect 8234 19014 8244 19066
rect 8244 19014 8290 19066
rect 7994 19012 8050 19014
rect 8074 19012 8130 19014
rect 8154 19012 8210 19014
rect 8234 19012 8290 19014
rect 8206 18572 8208 18592
rect 8208 18572 8260 18592
rect 8260 18572 8262 18592
rect 8206 18536 8262 18572
rect 7994 17978 8050 17980
rect 8074 17978 8130 17980
rect 8154 17978 8210 17980
rect 8234 17978 8290 17980
rect 7994 17926 8040 17978
rect 8040 17926 8050 17978
rect 8074 17926 8104 17978
rect 8104 17926 8116 17978
rect 8116 17926 8130 17978
rect 8154 17926 8168 17978
rect 8168 17926 8180 17978
rect 8180 17926 8210 17978
rect 8234 17926 8244 17978
rect 8244 17926 8290 17978
rect 7994 17924 8050 17926
rect 8074 17924 8130 17926
rect 8154 17924 8210 17926
rect 8234 17924 8290 17926
rect 7994 16890 8050 16892
rect 8074 16890 8130 16892
rect 8154 16890 8210 16892
rect 8234 16890 8290 16892
rect 7994 16838 8040 16890
rect 8040 16838 8050 16890
rect 8074 16838 8104 16890
rect 8104 16838 8116 16890
rect 8116 16838 8130 16890
rect 8154 16838 8168 16890
rect 8168 16838 8180 16890
rect 8180 16838 8210 16890
rect 8234 16838 8244 16890
rect 8244 16838 8290 16890
rect 7994 16836 8050 16838
rect 8074 16836 8130 16838
rect 8154 16836 8210 16838
rect 8234 16836 8290 16838
rect 8482 19660 8484 19680
rect 8484 19660 8536 19680
rect 8536 19660 8538 19680
rect 8482 19624 8538 19660
rect 9586 20440 9642 20496
rect 9034 20304 9090 20360
rect 9034 19488 9090 19544
rect 8482 16768 8538 16824
rect 8390 16496 8446 16552
rect 7994 15802 8050 15804
rect 8074 15802 8130 15804
rect 8154 15802 8210 15804
rect 8234 15802 8290 15804
rect 7994 15750 8040 15802
rect 8040 15750 8050 15802
rect 8074 15750 8104 15802
rect 8104 15750 8116 15802
rect 8116 15750 8130 15802
rect 8154 15750 8168 15802
rect 8168 15750 8180 15802
rect 8180 15750 8210 15802
rect 8234 15750 8244 15802
rect 8244 15750 8290 15802
rect 7994 15748 8050 15750
rect 8074 15748 8130 15750
rect 8154 15748 8210 15750
rect 8234 15748 8290 15750
rect 7994 14714 8050 14716
rect 8074 14714 8130 14716
rect 8154 14714 8210 14716
rect 8234 14714 8290 14716
rect 7994 14662 8040 14714
rect 8040 14662 8050 14714
rect 8074 14662 8104 14714
rect 8104 14662 8116 14714
rect 8116 14662 8130 14714
rect 8154 14662 8168 14714
rect 8168 14662 8180 14714
rect 8180 14662 8210 14714
rect 8234 14662 8244 14714
rect 8244 14662 8290 14714
rect 7994 14660 8050 14662
rect 8074 14660 8130 14662
rect 8154 14660 8210 14662
rect 8234 14660 8290 14662
rect 7994 13626 8050 13628
rect 8074 13626 8130 13628
rect 8154 13626 8210 13628
rect 8234 13626 8290 13628
rect 7994 13574 8040 13626
rect 8040 13574 8050 13626
rect 8074 13574 8104 13626
rect 8104 13574 8116 13626
rect 8116 13574 8130 13626
rect 8154 13574 8168 13626
rect 8168 13574 8180 13626
rect 8180 13574 8210 13626
rect 8234 13574 8244 13626
rect 8244 13574 8290 13626
rect 7994 13572 8050 13574
rect 8074 13572 8130 13574
rect 8154 13572 8210 13574
rect 8234 13572 8290 13574
rect 7654 12552 7710 12608
rect 7994 12538 8050 12540
rect 8074 12538 8130 12540
rect 8154 12538 8210 12540
rect 8234 12538 8290 12540
rect 7994 12486 8040 12538
rect 8040 12486 8050 12538
rect 8074 12486 8104 12538
rect 8104 12486 8116 12538
rect 8116 12486 8130 12538
rect 8154 12486 8168 12538
rect 8168 12486 8180 12538
rect 8180 12486 8210 12538
rect 8234 12486 8244 12538
rect 8244 12486 8290 12538
rect 7994 12484 8050 12486
rect 8074 12484 8130 12486
rect 8154 12484 8210 12486
rect 8234 12484 8290 12486
rect 8850 17720 8906 17776
rect 8850 17040 8906 17096
rect 8574 15136 8630 15192
rect 8758 14592 8814 14648
rect 8666 14048 8722 14104
rect 6918 8880 6974 8936
rect 6458 8064 6514 8120
rect 6274 7248 6330 7304
rect 6090 5788 6092 5808
rect 6092 5788 6144 5808
rect 6144 5788 6146 5808
rect 6090 5752 6146 5788
rect 6550 7404 6606 7440
rect 6550 7384 6552 7404
rect 6552 7384 6604 7404
rect 6604 7384 6606 7404
rect 6918 8608 6974 8664
rect 7470 9036 7526 9072
rect 7470 9016 7472 9036
rect 7472 9016 7524 9036
rect 7524 9016 7526 9036
rect 7010 8336 7066 8392
rect 6918 6840 6974 6896
rect 7994 11450 8050 11452
rect 8074 11450 8130 11452
rect 8154 11450 8210 11452
rect 8234 11450 8290 11452
rect 7994 11398 8040 11450
rect 8040 11398 8050 11450
rect 8074 11398 8104 11450
rect 8104 11398 8116 11450
rect 8116 11398 8130 11450
rect 8154 11398 8168 11450
rect 8168 11398 8180 11450
rect 8180 11398 8210 11450
rect 8234 11398 8244 11450
rect 8244 11398 8290 11450
rect 7994 11396 8050 11398
rect 8074 11396 8130 11398
rect 8154 11396 8210 11398
rect 8234 11396 8290 11398
rect 7994 10362 8050 10364
rect 8074 10362 8130 10364
rect 8154 10362 8210 10364
rect 8234 10362 8290 10364
rect 7994 10310 8040 10362
rect 8040 10310 8050 10362
rect 8074 10310 8104 10362
rect 8104 10310 8116 10362
rect 8116 10310 8130 10362
rect 8154 10310 8168 10362
rect 8168 10310 8180 10362
rect 8180 10310 8210 10362
rect 8234 10310 8244 10362
rect 8244 10310 8290 10362
rect 7994 10308 8050 10310
rect 8074 10308 8130 10310
rect 8154 10308 8210 10310
rect 8234 10308 8290 10310
rect 7994 9274 8050 9276
rect 8074 9274 8130 9276
rect 8154 9274 8210 9276
rect 8234 9274 8290 9276
rect 7994 9222 8040 9274
rect 8040 9222 8050 9274
rect 8074 9222 8104 9274
rect 8104 9222 8116 9274
rect 8116 9222 8130 9274
rect 8154 9222 8168 9274
rect 8168 9222 8180 9274
rect 8180 9222 8210 9274
rect 8234 9222 8244 9274
rect 8244 9222 8290 9274
rect 7994 9220 8050 9222
rect 8074 9220 8130 9222
rect 8154 9220 8210 9222
rect 8234 9220 8290 9222
rect 8942 14184 8998 14240
rect 9494 20168 9550 20224
rect 9218 19216 9274 19272
rect 9218 18128 9274 18184
rect 9218 17584 9274 17640
rect 10230 21936 10286 21992
rect 10966 21528 11022 21584
rect 10598 20984 10654 21040
rect 9586 18536 9642 18592
rect 9678 18400 9734 18456
rect 10322 18808 10378 18864
rect 9678 17448 9734 17504
rect 9218 16360 9274 16416
rect 9770 17040 9826 17096
rect 9494 16768 9550 16824
rect 9678 16632 9734 16688
rect 9494 16360 9550 16416
rect 9218 13776 9274 13832
rect 9034 12552 9090 12608
rect 9402 11736 9458 11792
rect 10506 16496 10562 16552
rect 10414 15408 10470 15464
rect 10322 14592 10378 14648
rect 10322 14476 10378 14512
rect 10322 14456 10324 14476
rect 10324 14456 10376 14476
rect 10376 14456 10378 14476
rect 10322 14184 10378 14240
rect 10414 13368 10470 13424
rect 10782 21256 10838 21312
rect 11789 21786 11845 21788
rect 11869 21786 11925 21788
rect 11949 21786 12005 21788
rect 12029 21786 12085 21788
rect 11789 21734 11835 21786
rect 11835 21734 11845 21786
rect 11869 21734 11899 21786
rect 11899 21734 11911 21786
rect 11911 21734 11925 21786
rect 11949 21734 11963 21786
rect 11963 21734 11975 21786
rect 11975 21734 12005 21786
rect 12029 21734 12039 21786
rect 12039 21734 12085 21786
rect 11789 21732 11845 21734
rect 11869 21732 11925 21734
rect 11949 21732 12005 21734
rect 12029 21732 12085 21734
rect 10966 20596 11022 20632
rect 10966 20576 10968 20596
rect 10968 20576 11020 20596
rect 11020 20576 11022 20596
rect 10690 19352 10746 19408
rect 10690 19252 10692 19272
rect 10692 19252 10744 19272
rect 10744 19252 10746 19272
rect 10690 19216 10746 19252
rect 10690 18028 10692 18048
rect 10692 18028 10744 18048
rect 10744 18028 10746 18048
rect 10690 17992 10746 18028
rect 11242 18808 11298 18864
rect 11058 17720 11114 17776
rect 10598 15136 10654 15192
rect 10782 16768 10838 16824
rect 11058 16904 11114 16960
rect 10782 15816 10838 15872
rect 11610 21292 11612 21312
rect 11612 21292 11664 21312
rect 11664 21292 11666 21312
rect 11610 21256 11666 21292
rect 11426 18944 11482 19000
rect 11150 16496 11206 16552
rect 11150 15680 11206 15736
rect 11058 15308 11060 15328
rect 11060 15308 11112 15328
rect 11112 15308 11114 15328
rect 11058 15272 11114 15308
rect 13818 21936 13874 21992
rect 12254 21528 12310 21584
rect 12162 20984 12218 21040
rect 11789 20698 11845 20700
rect 11869 20698 11925 20700
rect 11949 20698 12005 20700
rect 12029 20698 12085 20700
rect 11789 20646 11835 20698
rect 11835 20646 11845 20698
rect 11869 20646 11899 20698
rect 11899 20646 11911 20698
rect 11911 20646 11925 20698
rect 11949 20646 11963 20698
rect 11963 20646 11975 20698
rect 11975 20646 12005 20698
rect 12029 20646 12039 20698
rect 12039 20646 12085 20698
rect 11789 20644 11845 20646
rect 11869 20644 11925 20646
rect 11949 20644 12005 20646
rect 12029 20644 12085 20646
rect 11789 19610 11845 19612
rect 11869 19610 11925 19612
rect 11949 19610 12005 19612
rect 12029 19610 12085 19612
rect 11789 19558 11835 19610
rect 11835 19558 11845 19610
rect 11869 19558 11899 19610
rect 11899 19558 11911 19610
rect 11911 19558 11925 19610
rect 11949 19558 11963 19610
rect 11963 19558 11975 19610
rect 11975 19558 12005 19610
rect 12029 19558 12039 19610
rect 12039 19558 12085 19610
rect 11789 19556 11845 19558
rect 11869 19556 11925 19558
rect 11949 19556 12005 19558
rect 12029 19556 12085 19558
rect 11789 18522 11845 18524
rect 11869 18522 11925 18524
rect 11949 18522 12005 18524
rect 12029 18522 12085 18524
rect 11789 18470 11835 18522
rect 11835 18470 11845 18522
rect 11869 18470 11899 18522
rect 11899 18470 11911 18522
rect 11911 18470 11925 18522
rect 11949 18470 11963 18522
rect 11963 18470 11975 18522
rect 11975 18470 12005 18522
rect 12029 18470 12039 18522
rect 12039 18470 12085 18522
rect 11789 18468 11845 18470
rect 11869 18468 11925 18470
rect 11949 18468 12005 18470
rect 12029 18468 12085 18470
rect 11702 17856 11758 17912
rect 11789 17434 11845 17436
rect 11869 17434 11925 17436
rect 11949 17434 12005 17436
rect 12029 17434 12085 17436
rect 11789 17382 11835 17434
rect 11835 17382 11845 17434
rect 11869 17382 11899 17434
rect 11899 17382 11911 17434
rect 11911 17382 11925 17434
rect 11949 17382 11963 17434
rect 11963 17382 11975 17434
rect 11975 17382 12005 17434
rect 12029 17382 12039 17434
rect 12039 17382 12085 17434
rect 11789 17380 11845 17382
rect 11869 17380 11925 17382
rect 11949 17380 12005 17382
rect 12029 17380 12085 17382
rect 12254 17040 12310 17096
rect 10414 12180 10416 12200
rect 10416 12180 10468 12200
rect 10468 12180 10470 12200
rect 10414 12144 10470 12180
rect 9954 11192 10010 11248
rect 8574 9016 8630 9072
rect 8850 8508 8852 8528
rect 8852 8508 8904 8528
rect 8904 8508 8906 8528
rect 8850 8472 8906 8508
rect 9586 11056 9642 11112
rect 7654 8200 7710 8256
rect 7994 8186 8050 8188
rect 8074 8186 8130 8188
rect 8154 8186 8210 8188
rect 8234 8186 8290 8188
rect 7994 8134 8040 8186
rect 8040 8134 8050 8186
rect 8074 8134 8104 8186
rect 8104 8134 8116 8186
rect 8116 8134 8130 8186
rect 8154 8134 8168 8186
rect 8168 8134 8180 8186
rect 8180 8134 8210 8186
rect 8234 8134 8244 8186
rect 8244 8134 8290 8186
rect 7994 8132 8050 8134
rect 8074 8132 8130 8134
rect 8154 8132 8210 8134
rect 8234 8132 8290 8134
rect 8206 7828 8208 7848
rect 8208 7828 8260 7848
rect 8260 7828 8262 7848
rect 8206 7792 8262 7828
rect 7562 7268 7618 7304
rect 7562 7248 7564 7268
rect 7564 7248 7616 7268
rect 7616 7248 7618 7268
rect 7994 7098 8050 7100
rect 8074 7098 8130 7100
rect 8154 7098 8210 7100
rect 8234 7098 8290 7100
rect 7994 7046 8040 7098
rect 8040 7046 8050 7098
rect 8074 7046 8104 7098
rect 8104 7046 8116 7098
rect 8116 7046 8130 7098
rect 8154 7046 8168 7098
rect 8168 7046 8180 7098
rect 8180 7046 8210 7098
rect 8234 7046 8244 7098
rect 8244 7046 8290 7098
rect 7994 7044 8050 7046
rect 8074 7044 8130 7046
rect 8154 7044 8210 7046
rect 8234 7044 8290 7046
rect 7994 6010 8050 6012
rect 8074 6010 8130 6012
rect 8154 6010 8210 6012
rect 8234 6010 8290 6012
rect 7994 5958 8040 6010
rect 8040 5958 8050 6010
rect 8074 5958 8104 6010
rect 8104 5958 8116 6010
rect 8116 5958 8130 6010
rect 8154 5958 8168 6010
rect 8168 5958 8180 6010
rect 8180 5958 8210 6010
rect 8234 5958 8244 6010
rect 8244 5958 8290 6010
rect 7994 5956 8050 5958
rect 8074 5956 8130 5958
rect 8154 5956 8210 5958
rect 8234 5956 8290 5958
rect 6458 5616 6514 5672
rect 5906 3732 5962 3768
rect 5906 3712 5908 3732
rect 5908 3712 5960 3732
rect 5960 3712 5962 3732
rect 5170 2488 5226 2544
rect 5170 1400 5226 1456
rect 5354 2488 5410 2544
rect 5998 2916 6054 2952
rect 5998 2896 6000 2916
rect 6000 2896 6052 2916
rect 6052 2896 6054 2916
rect 5998 2644 6054 2680
rect 5998 2624 6000 2644
rect 6000 2624 6052 2644
rect 6052 2624 6054 2644
rect 5538 1944 5594 2000
rect 6826 5072 6882 5128
rect 7194 4528 7250 4584
rect 6918 3576 6974 3632
rect 6550 2760 6606 2816
rect 6550 1708 6552 1728
rect 6552 1708 6604 1728
rect 6604 1708 6606 1728
rect 6550 1672 6606 1708
rect 6734 1264 6790 1320
rect 6642 992 6698 1048
rect 4250 312 4306 368
rect 7994 4922 8050 4924
rect 8074 4922 8130 4924
rect 8154 4922 8210 4924
rect 8234 4922 8290 4924
rect 7994 4870 8040 4922
rect 8040 4870 8050 4922
rect 8074 4870 8104 4922
rect 8104 4870 8116 4922
rect 8116 4870 8130 4922
rect 8154 4870 8168 4922
rect 8168 4870 8180 4922
rect 8180 4870 8210 4922
rect 8234 4870 8244 4922
rect 8244 4870 8290 4922
rect 7994 4868 8050 4870
rect 8074 4868 8130 4870
rect 8154 4868 8210 4870
rect 8234 4868 8290 4870
rect 8206 4564 8208 4584
rect 8208 4564 8260 4584
rect 8260 4564 8262 4584
rect 8206 4528 8262 4564
rect 7994 3834 8050 3836
rect 8074 3834 8130 3836
rect 8154 3834 8210 3836
rect 8234 3834 8290 3836
rect 7994 3782 8040 3834
rect 8040 3782 8050 3834
rect 8074 3782 8104 3834
rect 8104 3782 8116 3834
rect 8116 3782 8130 3834
rect 8154 3782 8168 3834
rect 8168 3782 8180 3834
rect 8180 3782 8210 3834
rect 8234 3782 8244 3834
rect 8244 3782 8290 3834
rect 7994 3780 8050 3782
rect 8074 3780 8130 3782
rect 8154 3780 8210 3782
rect 8234 3780 8290 3782
rect 8850 5208 8906 5264
rect 8758 4664 8814 4720
rect 8666 4528 8722 4584
rect 8574 3984 8630 4040
rect 7994 2746 8050 2748
rect 8074 2746 8130 2748
rect 8154 2746 8210 2748
rect 8234 2746 8290 2748
rect 7994 2694 8040 2746
rect 8040 2694 8050 2746
rect 8074 2694 8104 2746
rect 8104 2694 8116 2746
rect 8116 2694 8130 2746
rect 8154 2694 8168 2746
rect 8168 2694 8180 2746
rect 8180 2694 8210 2746
rect 8234 2694 8244 2746
rect 8244 2694 8290 2746
rect 7994 2692 8050 2694
rect 8074 2692 8130 2694
rect 8154 2692 8210 2694
rect 8234 2692 8290 2694
rect 9126 7656 9182 7712
rect 9586 7656 9642 7712
rect 9126 6196 9128 6216
rect 9128 6196 9180 6216
rect 9180 6196 9182 6216
rect 9126 6160 9182 6196
rect 7994 1658 8050 1660
rect 8074 1658 8130 1660
rect 8154 1658 8210 1660
rect 8234 1658 8290 1660
rect 7994 1606 8040 1658
rect 8040 1606 8050 1658
rect 8074 1606 8104 1658
rect 8104 1606 8116 1658
rect 8116 1606 8130 1658
rect 8154 1606 8168 1658
rect 8168 1606 8180 1658
rect 8180 1606 8210 1658
rect 8234 1606 8244 1658
rect 8244 1606 8290 1658
rect 7994 1604 8050 1606
rect 8074 1604 8130 1606
rect 8154 1604 8210 1606
rect 8234 1604 8290 1606
rect 8298 1128 8354 1184
rect 9310 1128 9366 1184
rect 10230 6976 10286 7032
rect 11058 13640 11114 13696
rect 10874 12824 10930 12880
rect 10782 11736 10838 11792
rect 11058 12688 11114 12744
rect 12162 16396 12164 16416
rect 12164 16396 12216 16416
rect 12216 16396 12218 16416
rect 12162 16360 12218 16396
rect 11789 16346 11845 16348
rect 11869 16346 11925 16348
rect 11949 16346 12005 16348
rect 12029 16346 12085 16348
rect 11789 16294 11835 16346
rect 11835 16294 11845 16346
rect 11869 16294 11899 16346
rect 11899 16294 11911 16346
rect 11911 16294 11925 16346
rect 11949 16294 11963 16346
rect 11963 16294 11975 16346
rect 11975 16294 12005 16346
rect 12029 16294 12039 16346
rect 12039 16294 12085 16346
rect 11789 16292 11845 16294
rect 11869 16292 11925 16294
rect 11949 16292 12005 16294
rect 12029 16292 12085 16294
rect 12438 20848 12494 20904
rect 12806 17992 12862 18048
rect 12806 16788 12862 16824
rect 12806 16768 12808 16788
rect 12808 16768 12860 16788
rect 12860 16768 12862 16788
rect 11789 15258 11845 15260
rect 11869 15258 11925 15260
rect 11949 15258 12005 15260
rect 12029 15258 12085 15260
rect 11789 15206 11835 15258
rect 11835 15206 11845 15258
rect 11869 15206 11899 15258
rect 11899 15206 11911 15258
rect 11911 15206 11925 15258
rect 11949 15206 11963 15258
rect 11963 15206 11975 15258
rect 11975 15206 12005 15258
rect 12029 15206 12039 15258
rect 12039 15206 12085 15258
rect 11789 15204 11845 15206
rect 11869 15204 11925 15206
rect 11949 15204 12005 15206
rect 12029 15204 12085 15206
rect 11789 14170 11845 14172
rect 11869 14170 11925 14172
rect 11949 14170 12005 14172
rect 12029 14170 12085 14172
rect 11789 14118 11835 14170
rect 11835 14118 11845 14170
rect 11869 14118 11899 14170
rect 11899 14118 11911 14170
rect 11911 14118 11925 14170
rect 11949 14118 11963 14170
rect 11963 14118 11975 14170
rect 11975 14118 12005 14170
rect 12029 14118 12039 14170
rect 12039 14118 12085 14170
rect 11789 14116 11845 14118
rect 11869 14116 11925 14118
rect 11949 14116 12005 14118
rect 12029 14116 12085 14118
rect 11978 13912 12034 13968
rect 11978 13776 12034 13832
rect 11242 12960 11298 13016
rect 11058 11600 11114 11656
rect 10874 11328 10930 11384
rect 10782 10376 10838 10432
rect 11610 12960 11666 13016
rect 11794 13232 11850 13288
rect 11789 13082 11845 13084
rect 11869 13082 11925 13084
rect 11949 13082 12005 13084
rect 12029 13082 12085 13084
rect 11789 13030 11835 13082
rect 11835 13030 11845 13082
rect 11869 13030 11899 13082
rect 11899 13030 11911 13082
rect 11911 13030 11925 13082
rect 11949 13030 11963 13082
rect 11963 13030 11975 13082
rect 11975 13030 12005 13082
rect 12029 13030 12039 13082
rect 12039 13030 12085 13082
rect 11789 13028 11845 13030
rect 11869 13028 11925 13030
rect 11949 13028 12005 13030
rect 12029 13028 12085 13030
rect 13082 18264 13138 18320
rect 13818 21256 13874 21312
rect 14094 21392 14150 21448
rect 19338 22092 19394 22128
rect 19338 22072 19340 22092
rect 19340 22072 19392 22092
rect 19392 22072 19394 22092
rect 22466 22072 22522 22128
rect 14278 19352 14334 19408
rect 13450 18808 13506 18864
rect 13634 18148 13690 18184
rect 13634 18128 13636 18148
rect 13636 18128 13688 18148
rect 13688 18128 13690 18148
rect 13358 17720 13414 17776
rect 13634 17176 13690 17232
rect 13634 16496 13690 16552
rect 13174 16360 13230 16416
rect 13082 15036 13084 15056
rect 13084 15036 13136 15056
rect 13136 15036 13138 15056
rect 13082 15000 13138 15036
rect 12714 14456 12770 14512
rect 12438 13096 12494 13152
rect 11794 12552 11850 12608
rect 12346 12416 12402 12472
rect 11978 12280 12034 12336
rect 11610 12144 11666 12200
rect 11789 11994 11845 11996
rect 11869 11994 11925 11996
rect 11949 11994 12005 11996
rect 12029 11994 12085 11996
rect 11789 11942 11835 11994
rect 11835 11942 11845 11994
rect 11869 11942 11899 11994
rect 11899 11942 11911 11994
rect 11911 11942 11925 11994
rect 11949 11942 11963 11994
rect 11963 11942 11975 11994
rect 11975 11942 12005 11994
rect 12029 11942 12039 11994
rect 12039 11942 12085 11994
rect 11789 11940 11845 11942
rect 11869 11940 11925 11942
rect 11949 11940 12005 11942
rect 12029 11940 12085 11942
rect 11978 11736 12034 11792
rect 13082 14184 13138 14240
rect 14002 16904 14058 16960
rect 13818 15816 13874 15872
rect 13450 15544 13506 15600
rect 14554 19760 14610 19816
rect 15584 21242 15640 21244
rect 15664 21242 15720 21244
rect 15744 21242 15800 21244
rect 15824 21242 15880 21244
rect 15584 21190 15630 21242
rect 15630 21190 15640 21242
rect 15664 21190 15694 21242
rect 15694 21190 15706 21242
rect 15706 21190 15720 21242
rect 15744 21190 15758 21242
rect 15758 21190 15770 21242
rect 15770 21190 15800 21242
rect 15824 21190 15834 21242
rect 15834 21190 15880 21242
rect 15584 21188 15640 21190
rect 15664 21188 15720 21190
rect 15744 21188 15800 21190
rect 15824 21188 15880 21190
rect 15198 20596 15254 20632
rect 15198 20576 15200 20596
rect 15200 20576 15252 20596
rect 15252 20576 15254 20596
rect 13450 13948 13452 13968
rect 13452 13948 13504 13968
rect 13504 13948 13506 13968
rect 12898 13368 12954 13424
rect 12714 12280 12770 12336
rect 12346 11872 12402 11928
rect 12438 11756 12494 11792
rect 12438 11736 12440 11756
rect 12440 11736 12492 11756
rect 12492 11736 12494 11756
rect 13450 13912 13506 13948
rect 13358 13776 13414 13832
rect 13818 13232 13874 13288
rect 13818 13096 13874 13152
rect 13174 11872 13230 11928
rect 11789 10906 11845 10908
rect 11869 10906 11925 10908
rect 11949 10906 12005 10908
rect 12029 10906 12085 10908
rect 11789 10854 11835 10906
rect 11835 10854 11845 10906
rect 11869 10854 11899 10906
rect 11899 10854 11911 10906
rect 11911 10854 11925 10906
rect 11949 10854 11963 10906
rect 11963 10854 11975 10906
rect 11975 10854 12005 10906
rect 12029 10854 12039 10906
rect 12039 10854 12085 10906
rect 11789 10852 11845 10854
rect 11869 10852 11925 10854
rect 11949 10852 12005 10854
rect 12029 10852 12085 10854
rect 11426 10240 11482 10296
rect 11242 9152 11298 9208
rect 10506 6568 10562 6624
rect 10874 6704 10930 6760
rect 10782 6024 10838 6080
rect 10322 5480 10378 5536
rect 7994 570 8050 572
rect 8074 570 8130 572
rect 8154 570 8210 572
rect 8234 570 8290 572
rect 7994 518 8040 570
rect 8040 518 8050 570
rect 8074 518 8104 570
rect 8104 518 8116 570
rect 8116 518 8130 570
rect 8154 518 8168 570
rect 8168 518 8180 570
rect 8180 518 8210 570
rect 8234 518 8244 570
rect 8244 518 8290 570
rect 7994 516 8050 518
rect 8074 516 8130 518
rect 8154 516 8210 518
rect 8234 516 8290 518
rect 11150 7248 11206 7304
rect 11789 9818 11845 9820
rect 11869 9818 11925 9820
rect 11949 9818 12005 9820
rect 12029 9818 12085 9820
rect 11789 9766 11835 9818
rect 11835 9766 11845 9818
rect 11869 9766 11899 9818
rect 11899 9766 11911 9818
rect 11911 9766 11925 9818
rect 11949 9766 11963 9818
rect 11963 9766 11975 9818
rect 11975 9766 12005 9818
rect 12029 9766 12039 9818
rect 12039 9766 12085 9818
rect 11789 9764 11845 9766
rect 11869 9764 11925 9766
rect 11949 9764 12005 9766
rect 12029 9764 12085 9766
rect 12346 10920 12402 10976
rect 12254 10240 12310 10296
rect 12806 11056 12862 11112
rect 12622 10376 12678 10432
rect 13266 10376 13322 10432
rect 12162 9152 12218 9208
rect 11789 8730 11845 8732
rect 11869 8730 11925 8732
rect 11949 8730 12005 8732
rect 12029 8730 12085 8732
rect 11789 8678 11835 8730
rect 11835 8678 11845 8730
rect 11869 8678 11899 8730
rect 11899 8678 11911 8730
rect 11911 8678 11925 8730
rect 11949 8678 11963 8730
rect 11963 8678 11975 8730
rect 11975 8678 12005 8730
rect 12029 8678 12039 8730
rect 12039 8678 12085 8730
rect 11789 8676 11845 8678
rect 11869 8676 11925 8678
rect 11949 8676 12005 8678
rect 12029 8676 12085 8678
rect 11789 7642 11845 7644
rect 11869 7642 11925 7644
rect 11949 7642 12005 7644
rect 12029 7642 12085 7644
rect 11789 7590 11835 7642
rect 11835 7590 11845 7642
rect 11869 7590 11899 7642
rect 11899 7590 11911 7642
rect 11911 7590 11925 7642
rect 11949 7590 11963 7642
rect 11963 7590 11975 7642
rect 11975 7590 12005 7642
rect 12029 7590 12039 7642
rect 12039 7590 12085 7642
rect 11789 7588 11845 7590
rect 11869 7588 11925 7590
rect 11949 7588 12005 7590
rect 12029 7588 12085 7590
rect 11518 6860 11574 6896
rect 11518 6840 11520 6860
rect 11520 6840 11572 6860
rect 11572 6840 11574 6860
rect 10874 5208 10930 5264
rect 10966 2760 11022 2816
rect 11610 6432 11666 6488
rect 11426 6196 11428 6216
rect 11428 6196 11480 6216
rect 11480 6196 11482 6216
rect 11426 6160 11482 6196
rect 11610 6160 11666 6216
rect 11789 6554 11845 6556
rect 11869 6554 11925 6556
rect 11949 6554 12005 6556
rect 12029 6554 12085 6556
rect 11789 6502 11835 6554
rect 11835 6502 11845 6554
rect 11869 6502 11899 6554
rect 11899 6502 11911 6554
rect 11911 6502 11925 6554
rect 11949 6502 11963 6554
rect 11963 6502 11975 6554
rect 11975 6502 12005 6554
rect 12029 6502 12039 6554
rect 12039 6502 12085 6554
rect 11789 6500 11845 6502
rect 11869 6500 11925 6502
rect 11949 6500 12005 6502
rect 12029 6500 12085 6502
rect 12898 7248 12954 7304
rect 13082 6976 13138 7032
rect 14002 12300 14058 12336
rect 14002 12280 14004 12300
rect 14004 12280 14056 12300
rect 14056 12280 14058 12300
rect 13818 10920 13874 10976
rect 11702 5888 11758 5944
rect 11789 5466 11845 5468
rect 11869 5466 11925 5468
rect 11949 5466 12005 5468
rect 12029 5466 12085 5468
rect 11789 5414 11835 5466
rect 11835 5414 11845 5466
rect 11869 5414 11899 5466
rect 11899 5414 11911 5466
rect 11911 5414 11925 5466
rect 11949 5414 11963 5466
rect 11963 5414 11975 5466
rect 11975 5414 12005 5466
rect 12029 5414 12039 5466
rect 12039 5414 12085 5466
rect 11789 5412 11845 5414
rect 11869 5412 11925 5414
rect 11949 5412 12005 5414
rect 12029 5412 12085 5414
rect 11426 2624 11482 2680
rect 11789 4378 11845 4380
rect 11869 4378 11925 4380
rect 11949 4378 12005 4380
rect 12029 4378 12085 4380
rect 11789 4326 11835 4378
rect 11835 4326 11845 4378
rect 11869 4326 11899 4378
rect 11899 4326 11911 4378
rect 11911 4326 11925 4378
rect 11949 4326 11963 4378
rect 11963 4326 11975 4378
rect 11975 4326 12005 4378
rect 12029 4326 12039 4378
rect 12039 4326 12085 4378
rect 11789 4324 11845 4326
rect 11869 4324 11925 4326
rect 11949 4324 12005 4326
rect 12029 4324 12085 4326
rect 12254 4256 12310 4312
rect 11789 3290 11845 3292
rect 11869 3290 11925 3292
rect 11949 3290 12005 3292
rect 12029 3290 12085 3292
rect 11789 3238 11835 3290
rect 11835 3238 11845 3290
rect 11869 3238 11899 3290
rect 11899 3238 11911 3290
rect 11911 3238 11925 3290
rect 11949 3238 11963 3290
rect 11963 3238 11975 3290
rect 11975 3238 12005 3290
rect 12029 3238 12039 3290
rect 12039 3238 12085 3290
rect 11789 3236 11845 3238
rect 11869 3236 11925 3238
rect 11949 3236 12005 3238
rect 12029 3236 12085 3238
rect 11794 2760 11850 2816
rect 13542 6976 13598 7032
rect 13358 6568 13414 6624
rect 14094 11756 14150 11792
rect 14094 11736 14096 11756
rect 14096 11736 14148 11756
rect 14148 11736 14150 11756
rect 15584 20154 15640 20156
rect 15664 20154 15720 20156
rect 15744 20154 15800 20156
rect 15824 20154 15880 20156
rect 15584 20102 15630 20154
rect 15630 20102 15640 20154
rect 15664 20102 15694 20154
rect 15694 20102 15706 20154
rect 15706 20102 15720 20154
rect 15744 20102 15758 20154
rect 15758 20102 15770 20154
rect 15770 20102 15800 20154
rect 15824 20102 15834 20154
rect 15834 20102 15880 20154
rect 15584 20100 15640 20102
rect 15664 20100 15720 20102
rect 15744 20100 15800 20102
rect 15824 20100 15880 20102
rect 16762 20848 16818 20904
rect 16578 20440 16634 20496
rect 15584 19066 15640 19068
rect 15664 19066 15720 19068
rect 15744 19066 15800 19068
rect 15824 19066 15880 19068
rect 15584 19014 15630 19066
rect 15630 19014 15640 19066
rect 15664 19014 15694 19066
rect 15694 19014 15706 19066
rect 15706 19014 15720 19066
rect 15744 19014 15758 19066
rect 15758 19014 15770 19066
rect 15770 19014 15800 19066
rect 15824 19014 15834 19066
rect 15834 19014 15880 19066
rect 15584 19012 15640 19014
rect 15664 19012 15720 19014
rect 15744 19012 15800 19014
rect 15824 19012 15880 19014
rect 16118 19216 16174 19272
rect 15584 17978 15640 17980
rect 15664 17978 15720 17980
rect 15744 17978 15800 17980
rect 15824 17978 15880 17980
rect 15584 17926 15630 17978
rect 15630 17926 15640 17978
rect 15664 17926 15694 17978
rect 15694 17926 15706 17978
rect 15706 17926 15720 17978
rect 15744 17926 15758 17978
rect 15758 17926 15770 17978
rect 15770 17926 15800 17978
rect 15824 17926 15834 17978
rect 15834 17926 15880 17978
rect 15584 17924 15640 17926
rect 15664 17924 15720 17926
rect 15744 17924 15800 17926
rect 15824 17924 15880 17926
rect 15014 16632 15070 16688
rect 16486 19216 16542 19272
rect 16394 17992 16450 18048
rect 15584 16890 15640 16892
rect 15664 16890 15720 16892
rect 15744 16890 15800 16892
rect 15824 16890 15880 16892
rect 15584 16838 15630 16890
rect 15630 16838 15640 16890
rect 15664 16838 15694 16890
rect 15694 16838 15706 16890
rect 15706 16838 15720 16890
rect 15744 16838 15758 16890
rect 15758 16838 15770 16890
rect 15770 16838 15800 16890
rect 15824 16838 15834 16890
rect 15834 16838 15880 16890
rect 15584 16836 15640 16838
rect 15664 16836 15720 16838
rect 15744 16836 15800 16838
rect 15824 16836 15880 16838
rect 14830 14864 14886 14920
rect 15584 15802 15640 15804
rect 15664 15802 15720 15804
rect 15744 15802 15800 15804
rect 15824 15802 15880 15804
rect 15584 15750 15630 15802
rect 15630 15750 15640 15802
rect 15664 15750 15694 15802
rect 15694 15750 15706 15802
rect 15706 15750 15720 15802
rect 15744 15750 15758 15802
rect 15758 15750 15770 15802
rect 15770 15750 15800 15802
rect 15824 15750 15834 15802
rect 15834 15750 15880 15802
rect 15584 15748 15640 15750
rect 15664 15748 15720 15750
rect 15744 15748 15800 15750
rect 15824 15748 15880 15750
rect 15584 14714 15640 14716
rect 15664 14714 15720 14716
rect 15744 14714 15800 14716
rect 15824 14714 15880 14716
rect 15584 14662 15630 14714
rect 15630 14662 15640 14714
rect 15664 14662 15694 14714
rect 15694 14662 15706 14714
rect 15706 14662 15720 14714
rect 15744 14662 15758 14714
rect 15758 14662 15770 14714
rect 15770 14662 15800 14714
rect 15824 14662 15834 14714
rect 15834 14662 15880 14714
rect 15584 14660 15640 14662
rect 15664 14660 15720 14662
rect 15744 14660 15800 14662
rect 15824 14660 15880 14662
rect 15658 13776 15714 13832
rect 15584 13626 15640 13628
rect 15664 13626 15720 13628
rect 15744 13626 15800 13628
rect 15824 13626 15880 13628
rect 15584 13574 15630 13626
rect 15630 13574 15640 13626
rect 15664 13574 15694 13626
rect 15694 13574 15706 13626
rect 15706 13574 15720 13626
rect 15744 13574 15758 13626
rect 15758 13574 15770 13626
rect 15770 13574 15800 13626
rect 15824 13574 15834 13626
rect 15834 13574 15880 13626
rect 15584 13572 15640 13574
rect 15664 13572 15720 13574
rect 15744 13572 15800 13574
rect 15824 13572 15880 13574
rect 14554 11328 14610 11384
rect 13910 7284 13912 7304
rect 13912 7284 13964 7304
rect 13964 7284 13966 7304
rect 13910 7248 13966 7284
rect 13542 5616 13598 5672
rect 14462 7792 14518 7848
rect 15584 12538 15640 12540
rect 15664 12538 15720 12540
rect 15744 12538 15800 12540
rect 15824 12538 15880 12540
rect 15584 12486 15630 12538
rect 15630 12486 15640 12538
rect 15664 12486 15694 12538
rect 15694 12486 15706 12538
rect 15706 12486 15720 12538
rect 15744 12486 15758 12538
rect 15758 12486 15770 12538
rect 15770 12486 15800 12538
rect 15824 12486 15834 12538
rect 15834 12486 15880 12538
rect 15584 12484 15640 12486
rect 15664 12484 15720 12486
rect 15744 12484 15800 12486
rect 15824 12484 15880 12486
rect 15584 11450 15640 11452
rect 15664 11450 15720 11452
rect 15744 11450 15800 11452
rect 15824 11450 15880 11452
rect 15584 11398 15630 11450
rect 15630 11398 15640 11450
rect 15664 11398 15694 11450
rect 15694 11398 15706 11450
rect 15706 11398 15720 11450
rect 15744 11398 15758 11450
rect 15758 11398 15770 11450
rect 15770 11398 15800 11450
rect 15824 11398 15834 11450
rect 15834 11398 15880 11450
rect 15584 11396 15640 11398
rect 15664 11396 15720 11398
rect 15744 11396 15800 11398
rect 15824 11396 15880 11398
rect 15750 11076 15806 11112
rect 15750 11056 15752 11076
rect 15752 11056 15804 11076
rect 15804 11056 15806 11076
rect 15584 10362 15640 10364
rect 15664 10362 15720 10364
rect 15744 10362 15800 10364
rect 15824 10362 15880 10364
rect 15584 10310 15630 10362
rect 15630 10310 15640 10362
rect 15664 10310 15694 10362
rect 15694 10310 15706 10362
rect 15706 10310 15720 10362
rect 15744 10310 15758 10362
rect 15758 10310 15770 10362
rect 15770 10310 15800 10362
rect 15824 10310 15834 10362
rect 15834 10310 15880 10362
rect 15584 10308 15640 10310
rect 15664 10308 15720 10310
rect 15744 10308 15800 10310
rect 15824 10308 15880 10310
rect 15106 7284 15108 7304
rect 15108 7284 15160 7304
rect 15160 7284 15162 7304
rect 13910 3440 13966 3496
rect 15106 7248 15162 7284
rect 15290 6976 15346 7032
rect 15290 6432 15346 6488
rect 15584 9274 15640 9276
rect 15664 9274 15720 9276
rect 15744 9274 15800 9276
rect 15824 9274 15880 9276
rect 15584 9222 15630 9274
rect 15630 9222 15640 9274
rect 15664 9222 15694 9274
rect 15694 9222 15706 9274
rect 15706 9222 15720 9274
rect 15744 9222 15758 9274
rect 15758 9222 15770 9274
rect 15770 9222 15800 9274
rect 15824 9222 15834 9274
rect 15834 9222 15880 9274
rect 15584 9220 15640 9222
rect 15664 9220 15720 9222
rect 15744 9220 15800 9222
rect 15824 9220 15880 9222
rect 16302 14220 16304 14240
rect 16304 14220 16356 14240
rect 16356 14220 16358 14240
rect 16302 14184 16358 14220
rect 16854 16516 16910 16552
rect 16854 16496 16856 16516
rect 16856 16496 16908 16516
rect 16908 16496 16910 16516
rect 17958 21528 18014 21584
rect 18234 18808 18290 18864
rect 17958 18672 18014 18728
rect 18234 16360 18290 16416
rect 17038 15408 17094 15464
rect 16946 15000 17002 15056
rect 16578 14592 16634 14648
rect 15584 8186 15640 8188
rect 15664 8186 15720 8188
rect 15744 8186 15800 8188
rect 15824 8186 15880 8188
rect 15584 8134 15630 8186
rect 15630 8134 15640 8186
rect 15664 8134 15694 8186
rect 15694 8134 15706 8186
rect 15706 8134 15720 8186
rect 15744 8134 15758 8186
rect 15758 8134 15770 8186
rect 15770 8134 15800 8186
rect 15824 8134 15834 8186
rect 15834 8134 15880 8186
rect 15584 8132 15640 8134
rect 15664 8132 15720 8134
rect 15744 8132 15800 8134
rect 15824 8132 15880 8134
rect 15584 7098 15640 7100
rect 15664 7098 15720 7100
rect 15744 7098 15800 7100
rect 15824 7098 15880 7100
rect 15584 7046 15630 7098
rect 15630 7046 15640 7098
rect 15664 7046 15694 7098
rect 15694 7046 15706 7098
rect 15706 7046 15720 7098
rect 15744 7046 15758 7098
rect 15758 7046 15770 7098
rect 15770 7046 15800 7098
rect 15824 7046 15834 7098
rect 15834 7046 15880 7098
rect 15584 7044 15640 7046
rect 15664 7044 15720 7046
rect 15744 7044 15800 7046
rect 15824 7044 15880 7046
rect 15750 6704 15806 6760
rect 15934 6296 15990 6352
rect 15290 6024 15346 6080
rect 15198 4528 15254 4584
rect 14922 4020 14924 4040
rect 14924 4020 14976 4040
rect 14976 4020 14978 4040
rect 14922 3984 14978 4020
rect 14094 3440 14150 3496
rect 14830 3440 14886 3496
rect 15584 6010 15640 6012
rect 15664 6010 15720 6012
rect 15744 6010 15800 6012
rect 15824 6010 15880 6012
rect 15584 5958 15630 6010
rect 15630 5958 15640 6010
rect 15664 5958 15694 6010
rect 15694 5958 15706 6010
rect 15706 5958 15720 6010
rect 15744 5958 15758 6010
rect 15758 5958 15770 6010
rect 15770 5958 15800 6010
rect 15824 5958 15834 6010
rect 15834 5958 15880 6010
rect 15584 5956 15640 5958
rect 15664 5956 15720 5958
rect 15744 5956 15800 5958
rect 15824 5956 15880 5958
rect 16118 7928 16174 7984
rect 16670 11056 16726 11112
rect 16578 10668 16634 10704
rect 16578 10648 16580 10668
rect 16580 10648 16632 10668
rect 16632 10648 16634 10668
rect 16118 6296 16174 6352
rect 16302 6860 16358 6896
rect 16578 10104 16634 10160
rect 17314 15544 17370 15600
rect 18970 18808 19026 18864
rect 17682 15272 17738 15328
rect 18142 15564 18198 15600
rect 18142 15544 18144 15564
rect 18144 15544 18196 15564
rect 18196 15544 18198 15564
rect 17774 14864 17830 14920
rect 17498 14456 17554 14512
rect 17590 13368 17646 13424
rect 19379 21786 19435 21788
rect 19459 21786 19515 21788
rect 19539 21786 19595 21788
rect 19619 21786 19675 21788
rect 19379 21734 19425 21786
rect 19425 21734 19435 21786
rect 19459 21734 19489 21786
rect 19489 21734 19501 21786
rect 19501 21734 19515 21786
rect 19539 21734 19553 21786
rect 19553 21734 19565 21786
rect 19565 21734 19595 21786
rect 19619 21734 19629 21786
rect 19629 21734 19675 21786
rect 19379 21732 19435 21734
rect 19459 21732 19515 21734
rect 19539 21732 19595 21734
rect 19619 21732 19675 21734
rect 19379 20698 19435 20700
rect 19459 20698 19515 20700
rect 19539 20698 19595 20700
rect 19619 20698 19675 20700
rect 19379 20646 19425 20698
rect 19425 20646 19435 20698
rect 19459 20646 19489 20698
rect 19489 20646 19501 20698
rect 19501 20646 19515 20698
rect 19539 20646 19553 20698
rect 19553 20646 19565 20698
rect 19565 20646 19595 20698
rect 19619 20646 19629 20698
rect 19629 20646 19675 20698
rect 19379 20644 19435 20646
rect 19459 20644 19515 20646
rect 19539 20644 19595 20646
rect 19619 20644 19675 20646
rect 20350 21664 20406 21720
rect 22006 21548 22062 21584
rect 22006 21528 22008 21548
rect 22008 21528 22060 21548
rect 22060 21528 22062 21548
rect 19890 20576 19946 20632
rect 19379 19610 19435 19612
rect 19459 19610 19515 19612
rect 19539 19610 19595 19612
rect 19619 19610 19675 19612
rect 19379 19558 19425 19610
rect 19425 19558 19435 19610
rect 19459 19558 19489 19610
rect 19489 19558 19501 19610
rect 19501 19558 19515 19610
rect 19539 19558 19553 19610
rect 19553 19558 19565 19610
rect 19565 19558 19595 19610
rect 19619 19558 19629 19610
rect 19629 19558 19675 19610
rect 19379 19556 19435 19558
rect 19459 19556 19515 19558
rect 19539 19556 19595 19558
rect 19619 19556 19675 19558
rect 18878 15272 18934 15328
rect 19379 18522 19435 18524
rect 19459 18522 19515 18524
rect 19539 18522 19595 18524
rect 19619 18522 19675 18524
rect 19379 18470 19425 18522
rect 19425 18470 19435 18522
rect 19459 18470 19489 18522
rect 19489 18470 19501 18522
rect 19501 18470 19515 18522
rect 19539 18470 19553 18522
rect 19553 18470 19565 18522
rect 19565 18470 19595 18522
rect 19619 18470 19629 18522
rect 19629 18470 19675 18522
rect 19379 18468 19435 18470
rect 19459 18468 19515 18470
rect 19539 18468 19595 18470
rect 19619 18468 19675 18470
rect 19379 17434 19435 17436
rect 19459 17434 19515 17436
rect 19539 17434 19595 17436
rect 19619 17434 19675 17436
rect 19379 17382 19425 17434
rect 19425 17382 19435 17434
rect 19459 17382 19489 17434
rect 19489 17382 19501 17434
rect 19501 17382 19515 17434
rect 19539 17382 19553 17434
rect 19553 17382 19565 17434
rect 19565 17382 19595 17434
rect 19619 17382 19629 17434
rect 19629 17382 19675 17434
rect 19379 17380 19435 17382
rect 19459 17380 19515 17382
rect 19539 17380 19595 17382
rect 19619 17380 19675 17382
rect 19522 16904 19578 16960
rect 19379 16346 19435 16348
rect 19459 16346 19515 16348
rect 19539 16346 19595 16348
rect 19619 16346 19675 16348
rect 19379 16294 19425 16346
rect 19425 16294 19435 16346
rect 19459 16294 19489 16346
rect 19489 16294 19501 16346
rect 19501 16294 19515 16346
rect 19539 16294 19553 16346
rect 19553 16294 19565 16346
rect 19565 16294 19595 16346
rect 19619 16294 19629 16346
rect 19629 16294 19675 16346
rect 19379 16292 19435 16294
rect 19459 16292 19515 16294
rect 19539 16292 19595 16294
rect 19619 16292 19675 16294
rect 19379 15258 19435 15260
rect 19459 15258 19515 15260
rect 19539 15258 19595 15260
rect 19619 15258 19675 15260
rect 19379 15206 19425 15258
rect 19425 15206 19435 15258
rect 19459 15206 19489 15258
rect 19489 15206 19501 15258
rect 19501 15206 19515 15258
rect 19539 15206 19553 15258
rect 19553 15206 19565 15258
rect 19565 15206 19595 15258
rect 19619 15206 19629 15258
rect 19629 15206 19675 15258
rect 19379 15204 19435 15206
rect 19459 15204 19515 15206
rect 19539 15204 19595 15206
rect 19619 15204 19675 15206
rect 19798 15136 19854 15192
rect 19154 13812 19156 13832
rect 19156 13812 19208 13832
rect 19208 13812 19210 13832
rect 17682 12144 17738 12200
rect 16762 9968 16818 10024
rect 16302 6840 16304 6860
rect 16304 6840 16356 6860
rect 16356 6840 16358 6860
rect 16486 6704 16542 6760
rect 16210 5752 16266 5808
rect 17038 6568 17094 6624
rect 16026 5344 16082 5400
rect 15584 4922 15640 4924
rect 15664 4922 15720 4924
rect 15744 4922 15800 4924
rect 15824 4922 15880 4924
rect 15584 4870 15630 4922
rect 15630 4870 15640 4922
rect 15664 4870 15694 4922
rect 15694 4870 15706 4922
rect 15706 4870 15720 4922
rect 15744 4870 15758 4922
rect 15758 4870 15770 4922
rect 15770 4870 15800 4922
rect 15824 4870 15834 4922
rect 15834 4870 15880 4922
rect 15584 4868 15640 4870
rect 15664 4868 15720 4870
rect 15744 4868 15800 4870
rect 15824 4868 15880 4870
rect 15584 3834 15640 3836
rect 15664 3834 15720 3836
rect 15744 3834 15800 3836
rect 15824 3834 15880 3836
rect 15584 3782 15630 3834
rect 15630 3782 15640 3834
rect 15664 3782 15694 3834
rect 15694 3782 15706 3834
rect 15706 3782 15720 3834
rect 15744 3782 15758 3834
rect 15758 3782 15770 3834
rect 15770 3782 15800 3834
rect 15824 3782 15834 3834
rect 15834 3782 15880 3834
rect 15584 3780 15640 3782
rect 15664 3780 15720 3782
rect 15744 3780 15800 3782
rect 15824 3780 15880 3782
rect 16302 4392 16358 4448
rect 12254 2624 12310 2680
rect 11886 2352 11942 2408
rect 11789 2202 11845 2204
rect 11869 2202 11925 2204
rect 11949 2202 12005 2204
rect 12029 2202 12085 2204
rect 11789 2150 11835 2202
rect 11835 2150 11845 2202
rect 11869 2150 11899 2202
rect 11899 2150 11911 2202
rect 11911 2150 11925 2202
rect 11949 2150 11963 2202
rect 11963 2150 11975 2202
rect 11975 2150 12005 2202
rect 12029 2150 12039 2202
rect 12039 2150 12085 2202
rect 11789 2148 11845 2150
rect 11869 2148 11925 2150
rect 11949 2148 12005 2150
rect 12029 2148 12085 2150
rect 12438 2352 12494 2408
rect 11426 992 11482 1048
rect 11789 1114 11845 1116
rect 11869 1114 11925 1116
rect 11949 1114 12005 1116
rect 12029 1114 12085 1116
rect 11789 1062 11835 1114
rect 11835 1062 11845 1114
rect 11869 1062 11899 1114
rect 11899 1062 11911 1114
rect 11911 1062 11925 1114
rect 11949 1062 11963 1114
rect 11963 1062 11975 1114
rect 11975 1062 12005 1114
rect 12029 1062 12039 1114
rect 12039 1062 12085 1114
rect 11789 1060 11845 1062
rect 11869 1060 11925 1062
rect 11949 1060 12005 1062
rect 12029 1060 12085 1062
rect 11794 876 11850 912
rect 11794 856 11796 876
rect 11796 856 11848 876
rect 11848 856 11850 876
rect 15584 2746 15640 2748
rect 15664 2746 15720 2748
rect 15744 2746 15800 2748
rect 15824 2746 15880 2748
rect 15584 2694 15630 2746
rect 15630 2694 15640 2746
rect 15664 2694 15694 2746
rect 15694 2694 15706 2746
rect 15706 2694 15720 2746
rect 15744 2694 15758 2746
rect 15758 2694 15770 2746
rect 15770 2694 15800 2746
rect 15824 2694 15834 2746
rect 15834 2694 15880 2746
rect 15584 2692 15640 2694
rect 15664 2692 15720 2694
rect 15744 2692 15800 2694
rect 15824 2692 15880 2694
rect 15584 1658 15640 1660
rect 15664 1658 15720 1660
rect 15744 1658 15800 1660
rect 15824 1658 15880 1660
rect 15584 1606 15630 1658
rect 15630 1606 15640 1658
rect 15664 1606 15694 1658
rect 15694 1606 15706 1658
rect 15706 1606 15720 1658
rect 15744 1606 15758 1658
rect 15758 1606 15770 1658
rect 15770 1606 15800 1658
rect 15824 1606 15834 1658
rect 15834 1606 15880 1658
rect 15584 1604 15640 1606
rect 15664 1604 15720 1606
rect 15744 1604 15800 1606
rect 15824 1604 15880 1606
rect 15584 570 15640 572
rect 15664 570 15720 572
rect 15744 570 15800 572
rect 15824 570 15880 572
rect 15584 518 15630 570
rect 15630 518 15640 570
rect 15664 518 15694 570
rect 15694 518 15706 570
rect 15706 518 15720 570
rect 15744 518 15758 570
rect 15758 518 15770 570
rect 15770 518 15800 570
rect 15824 518 15834 570
rect 15834 518 15880 570
rect 15584 516 15640 518
rect 15664 516 15720 518
rect 15744 516 15800 518
rect 15824 516 15880 518
rect 16302 2796 16304 2816
rect 16304 2796 16356 2816
rect 16356 2796 16358 2816
rect 16302 2760 16358 2796
rect 17498 6432 17554 6488
rect 19154 13776 19210 13812
rect 19706 14728 19762 14784
rect 19614 14592 19670 14648
rect 19379 14170 19435 14172
rect 19459 14170 19515 14172
rect 19539 14170 19595 14172
rect 19619 14170 19675 14172
rect 19379 14118 19425 14170
rect 19425 14118 19435 14170
rect 19459 14118 19489 14170
rect 19489 14118 19501 14170
rect 19501 14118 19515 14170
rect 19539 14118 19553 14170
rect 19553 14118 19565 14170
rect 19565 14118 19595 14170
rect 19619 14118 19629 14170
rect 19629 14118 19675 14170
rect 19379 14116 19435 14118
rect 19459 14116 19515 14118
rect 19539 14116 19595 14118
rect 19619 14116 19675 14118
rect 19522 13948 19524 13968
rect 19524 13948 19576 13968
rect 19576 13948 19578 13968
rect 19522 13912 19578 13948
rect 18970 12416 19026 12472
rect 19982 17720 20038 17776
rect 22006 19624 22062 19680
rect 21178 18264 21234 18320
rect 21270 17720 21326 17776
rect 20534 16360 20590 16416
rect 23570 21836 23572 21856
rect 23572 21836 23624 21856
rect 23624 21836 23626 21856
rect 23570 21800 23626 21836
rect 23202 21428 23204 21448
rect 23204 21428 23256 21448
rect 23256 21428 23258 21448
rect 23202 21392 23258 21428
rect 22558 20304 22614 20360
rect 22466 19660 22468 19680
rect 22468 19660 22520 19680
rect 22520 19660 22522 19680
rect 22466 19624 22522 19660
rect 22190 18400 22246 18456
rect 22098 16940 22100 16960
rect 22100 16940 22152 16960
rect 22152 16940 22154 16960
rect 22098 16904 22154 16940
rect 21546 16632 21602 16688
rect 20810 15852 20812 15872
rect 20812 15852 20864 15872
rect 20864 15852 20866 15872
rect 20810 15816 20866 15852
rect 20442 14864 20498 14920
rect 20166 14184 20222 14240
rect 19890 14048 19946 14104
rect 19379 13082 19435 13084
rect 19459 13082 19515 13084
rect 19539 13082 19595 13084
rect 19619 13082 19675 13084
rect 19379 13030 19425 13082
rect 19425 13030 19435 13082
rect 19459 13030 19489 13082
rect 19489 13030 19501 13082
rect 19501 13030 19515 13082
rect 19539 13030 19553 13082
rect 19553 13030 19565 13082
rect 19565 13030 19595 13082
rect 19619 13030 19629 13082
rect 19629 13030 19675 13082
rect 19379 13028 19435 13030
rect 19459 13028 19515 13030
rect 19539 13028 19595 13030
rect 19619 13028 19675 13030
rect 19379 11994 19435 11996
rect 19459 11994 19515 11996
rect 19539 11994 19595 11996
rect 19619 11994 19675 11996
rect 19379 11942 19425 11994
rect 19425 11942 19435 11994
rect 19459 11942 19489 11994
rect 19489 11942 19501 11994
rect 19501 11942 19515 11994
rect 19539 11942 19553 11994
rect 19553 11942 19565 11994
rect 19565 11942 19595 11994
rect 19619 11942 19629 11994
rect 19629 11942 19675 11994
rect 19379 11940 19435 11942
rect 19459 11940 19515 11942
rect 19539 11940 19595 11942
rect 19619 11940 19675 11942
rect 21362 15408 21418 15464
rect 20626 13776 20682 13832
rect 21914 16224 21970 16280
rect 22926 19080 22982 19136
rect 23174 21242 23230 21244
rect 23254 21242 23310 21244
rect 23334 21242 23390 21244
rect 23414 21242 23470 21244
rect 23174 21190 23220 21242
rect 23220 21190 23230 21242
rect 23254 21190 23284 21242
rect 23284 21190 23296 21242
rect 23296 21190 23310 21242
rect 23334 21190 23348 21242
rect 23348 21190 23360 21242
rect 23360 21190 23390 21242
rect 23414 21190 23424 21242
rect 23424 21190 23470 21242
rect 23174 21188 23230 21190
rect 23254 21188 23310 21190
rect 23334 21188 23390 21190
rect 23414 21188 23470 21190
rect 23174 20154 23230 20156
rect 23254 20154 23310 20156
rect 23334 20154 23390 20156
rect 23414 20154 23470 20156
rect 23174 20102 23220 20154
rect 23220 20102 23230 20154
rect 23254 20102 23284 20154
rect 23284 20102 23296 20154
rect 23296 20102 23310 20154
rect 23334 20102 23348 20154
rect 23348 20102 23360 20154
rect 23360 20102 23390 20154
rect 23414 20102 23424 20154
rect 23424 20102 23470 20154
rect 23174 20100 23230 20102
rect 23254 20100 23310 20102
rect 23334 20100 23390 20102
rect 23414 20100 23470 20102
rect 23110 19896 23166 19952
rect 23174 19066 23230 19068
rect 23254 19066 23310 19068
rect 23334 19066 23390 19068
rect 23414 19066 23470 19068
rect 23174 19014 23220 19066
rect 23220 19014 23230 19066
rect 23254 19014 23284 19066
rect 23284 19014 23296 19066
rect 23296 19014 23310 19066
rect 23334 19014 23348 19066
rect 23348 19014 23360 19066
rect 23360 19014 23390 19066
rect 23414 19014 23424 19066
rect 23424 19014 23470 19066
rect 23174 19012 23230 19014
rect 23254 19012 23310 19014
rect 23334 19012 23390 19014
rect 23414 19012 23470 19014
rect 23478 18808 23534 18864
rect 23018 17992 23074 18048
rect 23174 17978 23230 17980
rect 23254 17978 23310 17980
rect 23334 17978 23390 17980
rect 23414 17978 23470 17980
rect 23174 17926 23220 17978
rect 23220 17926 23230 17978
rect 23254 17926 23284 17978
rect 23284 17926 23296 17978
rect 23296 17926 23310 17978
rect 23334 17926 23348 17978
rect 23348 17926 23360 17978
rect 23360 17926 23390 17978
rect 23414 17926 23424 17978
rect 23424 17926 23470 17978
rect 23174 17924 23230 17926
rect 23254 17924 23310 17926
rect 23334 17924 23390 17926
rect 23414 17924 23470 17926
rect 22926 17040 22982 17096
rect 21822 15816 21878 15872
rect 21270 13132 21272 13152
rect 21272 13132 21324 13152
rect 21324 13132 21326 13152
rect 21270 13096 21326 13132
rect 21178 12416 21234 12472
rect 22006 15544 22062 15600
rect 23478 17740 23534 17776
rect 23478 17720 23480 17740
rect 23480 17720 23532 17740
rect 23532 17720 23534 17740
rect 23846 20576 23902 20632
rect 23938 19916 23994 19952
rect 23938 19896 23940 19916
rect 23940 19896 23992 19916
rect 23992 19896 23994 19916
rect 24214 21664 24270 21720
rect 24030 19080 24086 19136
rect 23846 18536 23902 18592
rect 23294 17448 23350 17504
rect 23386 17212 23388 17232
rect 23388 17212 23440 17232
rect 23440 17212 23442 17232
rect 23386 17176 23442 17212
rect 23174 16890 23230 16892
rect 23254 16890 23310 16892
rect 23334 16890 23390 16892
rect 23414 16890 23470 16892
rect 23174 16838 23220 16890
rect 23220 16838 23230 16890
rect 23254 16838 23284 16890
rect 23284 16838 23296 16890
rect 23296 16838 23310 16890
rect 23334 16838 23348 16890
rect 23348 16838 23360 16890
rect 23360 16838 23390 16890
rect 23414 16838 23424 16890
rect 23424 16838 23470 16890
rect 23174 16836 23230 16838
rect 23254 16836 23310 16838
rect 23334 16836 23390 16838
rect 23414 16836 23470 16838
rect 23478 16632 23534 16688
rect 22374 14728 22430 14784
rect 23174 15802 23230 15804
rect 23254 15802 23310 15804
rect 23334 15802 23390 15804
rect 23414 15802 23470 15804
rect 23174 15750 23220 15802
rect 23220 15750 23230 15802
rect 23254 15750 23284 15802
rect 23284 15750 23296 15802
rect 23296 15750 23310 15802
rect 23334 15750 23348 15802
rect 23348 15750 23360 15802
rect 23360 15750 23390 15802
rect 23414 15750 23424 15802
rect 23424 15750 23470 15802
rect 23174 15748 23230 15750
rect 23254 15748 23310 15750
rect 23334 15748 23390 15750
rect 23414 15748 23470 15750
rect 23846 16652 23902 16688
rect 23846 16632 23848 16652
rect 23848 16632 23900 16652
rect 23900 16632 23902 16652
rect 24122 17176 24178 17232
rect 24490 21548 24546 21584
rect 24490 21528 24492 21548
rect 24492 21528 24544 21548
rect 24544 21528 24546 21548
rect 25134 21120 25190 21176
rect 25410 20848 25466 20904
rect 26969 21786 27025 21788
rect 27049 21786 27105 21788
rect 27129 21786 27185 21788
rect 27209 21786 27265 21788
rect 26969 21734 27015 21786
rect 27015 21734 27025 21786
rect 27049 21734 27079 21786
rect 27079 21734 27091 21786
rect 27091 21734 27105 21786
rect 27129 21734 27143 21786
rect 27143 21734 27155 21786
rect 27155 21734 27185 21786
rect 27209 21734 27219 21786
rect 27219 21734 27265 21786
rect 26969 21732 27025 21734
rect 27049 21732 27105 21734
rect 27129 21732 27185 21734
rect 27209 21732 27265 21734
rect 25870 21664 25926 21720
rect 25778 21392 25834 21448
rect 24490 17856 24546 17912
rect 23938 16396 23940 16416
rect 23940 16396 23992 16416
rect 23992 16396 23994 16416
rect 23938 16360 23994 16396
rect 23846 15680 23902 15736
rect 23174 14714 23230 14716
rect 23254 14714 23310 14716
rect 23334 14714 23390 14716
rect 23414 14714 23470 14716
rect 23174 14662 23220 14714
rect 23220 14662 23230 14714
rect 23254 14662 23284 14714
rect 23284 14662 23296 14714
rect 23296 14662 23310 14714
rect 23334 14662 23348 14714
rect 23348 14662 23360 14714
rect 23360 14662 23390 14714
rect 23414 14662 23424 14714
rect 23424 14662 23470 14714
rect 23174 14660 23230 14662
rect 23254 14660 23310 14662
rect 23334 14660 23390 14662
rect 23414 14660 23470 14662
rect 23110 14456 23166 14512
rect 24030 14728 24086 14784
rect 23938 14476 23994 14512
rect 23938 14456 23940 14476
rect 23940 14456 23992 14476
rect 23992 14456 23994 14476
rect 23174 13626 23230 13628
rect 23254 13626 23310 13628
rect 23334 13626 23390 13628
rect 23414 13626 23470 13628
rect 23174 13574 23220 13626
rect 23220 13574 23230 13626
rect 23254 13574 23284 13626
rect 23284 13574 23296 13626
rect 23296 13574 23310 13626
rect 23334 13574 23348 13626
rect 23348 13574 23360 13626
rect 23360 13574 23390 13626
rect 23414 13574 23424 13626
rect 23424 13574 23470 13626
rect 23174 13572 23230 13574
rect 23254 13572 23310 13574
rect 23334 13572 23390 13574
rect 23414 13572 23470 13574
rect 22006 13368 22062 13424
rect 21546 12144 21602 12200
rect 19798 11192 19854 11248
rect 19379 10906 19435 10908
rect 19459 10906 19515 10908
rect 19539 10906 19595 10908
rect 19619 10906 19675 10908
rect 19379 10854 19425 10906
rect 19425 10854 19435 10906
rect 19459 10854 19489 10906
rect 19489 10854 19501 10906
rect 19501 10854 19515 10906
rect 19539 10854 19553 10906
rect 19553 10854 19565 10906
rect 19565 10854 19595 10906
rect 19619 10854 19629 10906
rect 19629 10854 19675 10906
rect 19379 10852 19435 10854
rect 19459 10852 19515 10854
rect 19539 10852 19595 10854
rect 19619 10852 19675 10854
rect 19982 11056 20038 11112
rect 20442 10512 20498 10568
rect 18510 8880 18566 8936
rect 19379 9818 19435 9820
rect 19459 9818 19515 9820
rect 19539 9818 19595 9820
rect 19619 9818 19675 9820
rect 19379 9766 19425 9818
rect 19425 9766 19435 9818
rect 19459 9766 19489 9818
rect 19489 9766 19501 9818
rect 19501 9766 19515 9818
rect 19539 9766 19553 9818
rect 19553 9766 19565 9818
rect 19565 9766 19595 9818
rect 19619 9766 19629 9818
rect 19629 9766 19675 9818
rect 19379 9764 19435 9766
rect 19459 9764 19515 9766
rect 19539 9764 19595 9766
rect 19619 9764 19675 9766
rect 18050 8356 18106 8392
rect 18050 8336 18052 8356
rect 18052 8336 18104 8356
rect 18104 8336 18106 8356
rect 17958 7520 18014 7576
rect 17958 7420 17960 7440
rect 17960 7420 18012 7440
rect 18012 7420 18014 7440
rect 17958 7384 18014 7420
rect 17774 5208 17830 5264
rect 17590 5072 17646 5128
rect 17498 4664 17554 4720
rect 16762 3440 16818 3496
rect 18602 7284 18604 7304
rect 18604 7284 18656 7304
rect 18656 7284 18658 7304
rect 18602 7248 18658 7284
rect 19379 8730 19435 8732
rect 19459 8730 19515 8732
rect 19539 8730 19595 8732
rect 19619 8730 19675 8732
rect 19379 8678 19425 8730
rect 19425 8678 19435 8730
rect 19459 8678 19489 8730
rect 19489 8678 19501 8730
rect 19501 8678 19515 8730
rect 19539 8678 19553 8730
rect 19553 8678 19565 8730
rect 19565 8678 19595 8730
rect 19619 8678 19629 8730
rect 19629 8678 19675 8730
rect 19379 8676 19435 8678
rect 19459 8676 19515 8678
rect 19539 8676 19595 8678
rect 19619 8676 19675 8678
rect 19246 8336 19302 8392
rect 19379 7642 19435 7644
rect 19459 7642 19515 7644
rect 19539 7642 19595 7644
rect 19619 7642 19675 7644
rect 19379 7590 19425 7642
rect 19425 7590 19435 7642
rect 19459 7590 19489 7642
rect 19489 7590 19501 7642
rect 19501 7590 19515 7642
rect 19539 7590 19553 7642
rect 19553 7590 19565 7642
rect 19565 7590 19595 7642
rect 19619 7590 19629 7642
rect 19629 7590 19675 7642
rect 19379 7588 19435 7590
rect 19459 7588 19515 7590
rect 19539 7588 19595 7590
rect 19619 7588 19675 7590
rect 21914 12960 21970 13016
rect 23294 12724 23296 12744
rect 23296 12724 23348 12744
rect 23348 12724 23350 12744
rect 23294 12688 23350 12724
rect 24490 16224 24546 16280
rect 25502 20304 25558 20360
rect 24950 19216 25006 19272
rect 25502 17992 25558 18048
rect 24122 13912 24178 13968
rect 24766 13640 24822 13696
rect 23174 12538 23230 12540
rect 23254 12538 23310 12540
rect 23334 12538 23390 12540
rect 23414 12538 23470 12540
rect 23174 12486 23220 12538
rect 23220 12486 23230 12538
rect 23254 12486 23284 12538
rect 23284 12486 23296 12538
rect 23296 12486 23310 12538
rect 23334 12486 23348 12538
rect 23348 12486 23360 12538
rect 23360 12486 23390 12538
rect 23414 12486 23424 12538
rect 23424 12486 23470 12538
rect 23174 12484 23230 12486
rect 23254 12484 23310 12486
rect 23334 12484 23390 12486
rect 23414 12484 23470 12486
rect 24306 12960 24362 13016
rect 22466 11212 22522 11248
rect 22466 11192 22468 11212
rect 22468 11192 22520 11212
rect 22520 11192 22522 11212
rect 21362 10784 21418 10840
rect 20902 7248 20958 7304
rect 20718 6860 20774 6896
rect 20718 6840 20720 6860
rect 20720 6840 20772 6860
rect 20772 6840 20774 6860
rect 19379 6554 19435 6556
rect 19459 6554 19515 6556
rect 19539 6554 19595 6556
rect 19619 6554 19675 6556
rect 19379 6502 19425 6554
rect 19425 6502 19435 6554
rect 19459 6502 19489 6554
rect 19489 6502 19501 6554
rect 19501 6502 19515 6554
rect 19539 6502 19553 6554
rect 19553 6502 19565 6554
rect 19565 6502 19595 6554
rect 19619 6502 19629 6554
rect 19629 6502 19675 6554
rect 19379 6500 19435 6502
rect 19459 6500 19515 6502
rect 19539 6500 19595 6502
rect 19619 6500 19675 6502
rect 19379 5466 19435 5468
rect 19459 5466 19515 5468
rect 19539 5466 19595 5468
rect 19619 5466 19675 5468
rect 19379 5414 19425 5466
rect 19425 5414 19435 5466
rect 19459 5414 19489 5466
rect 19489 5414 19501 5466
rect 19501 5414 19515 5466
rect 19539 5414 19553 5466
rect 19553 5414 19565 5466
rect 19565 5414 19595 5466
rect 19619 5414 19629 5466
rect 19629 5414 19675 5466
rect 19379 5412 19435 5414
rect 19459 5412 19515 5414
rect 19539 5412 19595 5414
rect 19619 5412 19675 5414
rect 19154 4392 19210 4448
rect 19379 4378 19435 4380
rect 19459 4378 19515 4380
rect 19539 4378 19595 4380
rect 19619 4378 19675 4380
rect 19379 4326 19425 4378
rect 19425 4326 19435 4378
rect 19459 4326 19489 4378
rect 19489 4326 19501 4378
rect 19501 4326 19515 4378
rect 19539 4326 19553 4378
rect 19553 4326 19565 4378
rect 19565 4326 19595 4378
rect 19619 4326 19629 4378
rect 19629 4326 19675 4378
rect 19379 4324 19435 4326
rect 19459 4324 19515 4326
rect 19539 4324 19595 4326
rect 19619 4324 19675 4326
rect 19379 3290 19435 3292
rect 19459 3290 19515 3292
rect 19539 3290 19595 3292
rect 19619 3290 19675 3292
rect 19379 3238 19425 3290
rect 19425 3238 19435 3290
rect 19459 3238 19489 3290
rect 19489 3238 19501 3290
rect 19501 3238 19515 3290
rect 19539 3238 19553 3290
rect 19553 3238 19565 3290
rect 19565 3238 19595 3290
rect 19619 3238 19629 3290
rect 19629 3238 19675 3290
rect 19379 3236 19435 3238
rect 19459 3236 19515 3238
rect 19539 3236 19595 3238
rect 19619 3236 19675 3238
rect 19706 3032 19762 3088
rect 21362 7792 21418 7848
rect 17958 1828 18014 1864
rect 17958 1808 17960 1828
rect 17960 1808 18012 1828
rect 18012 1808 18014 1828
rect 19379 2202 19435 2204
rect 19459 2202 19515 2204
rect 19539 2202 19595 2204
rect 19619 2202 19675 2204
rect 19379 2150 19425 2202
rect 19425 2150 19435 2202
rect 19459 2150 19489 2202
rect 19489 2150 19501 2202
rect 19501 2150 19515 2202
rect 19539 2150 19553 2202
rect 19553 2150 19565 2202
rect 19565 2150 19595 2202
rect 19619 2150 19629 2202
rect 19629 2150 19675 2202
rect 19379 2148 19435 2150
rect 19459 2148 19515 2150
rect 19539 2148 19595 2150
rect 19619 2148 19675 2150
rect 19062 1808 19118 1864
rect 18234 1264 18290 1320
rect 18878 1264 18934 1320
rect 19430 1400 19486 1456
rect 19379 1114 19435 1116
rect 19459 1114 19515 1116
rect 19539 1114 19595 1116
rect 19619 1114 19675 1116
rect 19379 1062 19425 1114
rect 19425 1062 19435 1114
rect 19459 1062 19489 1114
rect 19489 1062 19501 1114
rect 19501 1062 19515 1114
rect 19539 1062 19553 1114
rect 19553 1062 19565 1114
rect 19565 1062 19595 1114
rect 19619 1062 19629 1114
rect 19629 1062 19675 1114
rect 19379 1060 19435 1062
rect 19459 1060 19515 1062
rect 19539 1060 19595 1062
rect 19619 1060 19675 1062
rect 21086 2760 21142 2816
rect 20626 2252 20628 2272
rect 20628 2252 20680 2272
rect 20680 2252 20682 2272
rect 20626 2216 20682 2252
rect 20718 1828 20774 1864
rect 20902 2080 20958 2136
rect 20718 1808 20720 1828
rect 20720 1808 20772 1828
rect 20772 1808 20774 1828
rect 20718 1012 20774 1048
rect 20718 992 20720 1012
rect 20720 992 20772 1012
rect 20772 992 20774 1012
rect 23294 11636 23296 11656
rect 23296 11636 23348 11656
rect 23348 11636 23350 11656
rect 23294 11600 23350 11636
rect 23174 11450 23230 11452
rect 23254 11450 23310 11452
rect 23334 11450 23390 11452
rect 23414 11450 23470 11452
rect 23174 11398 23220 11450
rect 23220 11398 23230 11450
rect 23254 11398 23284 11450
rect 23284 11398 23296 11450
rect 23296 11398 23310 11450
rect 23334 11398 23348 11450
rect 23348 11398 23360 11450
rect 23360 11398 23390 11450
rect 23414 11398 23424 11450
rect 23424 11398 23470 11450
rect 23174 11396 23230 11398
rect 23254 11396 23310 11398
rect 23334 11396 23390 11398
rect 23414 11396 23470 11398
rect 22926 10648 22982 10704
rect 24490 11600 24546 11656
rect 26238 19080 26294 19136
rect 25870 17484 25872 17504
rect 25872 17484 25924 17504
rect 25924 17484 25926 17504
rect 25870 17448 25926 17484
rect 25778 15136 25834 15192
rect 25686 14864 25742 14920
rect 26606 19216 26662 19272
rect 25962 15680 26018 15736
rect 26238 15816 26294 15872
rect 26146 14864 26202 14920
rect 26606 18300 26608 18320
rect 26608 18300 26660 18320
rect 26660 18300 26662 18320
rect 26606 18264 26662 18300
rect 26606 17176 26662 17232
rect 26969 20698 27025 20700
rect 27049 20698 27105 20700
rect 27129 20698 27185 20700
rect 27209 20698 27265 20700
rect 26969 20646 27015 20698
rect 27015 20646 27025 20698
rect 27049 20646 27079 20698
rect 27079 20646 27091 20698
rect 27091 20646 27105 20698
rect 27129 20646 27143 20698
rect 27143 20646 27155 20698
rect 27155 20646 27185 20698
rect 27209 20646 27219 20698
rect 27219 20646 27265 20698
rect 26969 20644 27025 20646
rect 27049 20644 27105 20646
rect 27129 20644 27185 20646
rect 27209 20644 27265 20646
rect 26969 19610 27025 19612
rect 27049 19610 27105 19612
rect 27129 19610 27185 19612
rect 27209 19610 27265 19612
rect 26969 19558 27015 19610
rect 27015 19558 27025 19610
rect 27049 19558 27079 19610
rect 27079 19558 27091 19610
rect 27091 19558 27105 19610
rect 27129 19558 27143 19610
rect 27143 19558 27155 19610
rect 27155 19558 27185 19610
rect 27209 19558 27219 19610
rect 27219 19558 27265 19610
rect 26969 19556 27025 19558
rect 27049 19556 27105 19558
rect 27129 19556 27185 19558
rect 27209 19556 27265 19558
rect 26974 19252 26976 19272
rect 26976 19252 27028 19272
rect 27028 19252 27030 19272
rect 26974 19216 27030 19252
rect 27618 19216 27674 19272
rect 26969 18522 27025 18524
rect 27049 18522 27105 18524
rect 27129 18522 27185 18524
rect 27209 18522 27265 18524
rect 26969 18470 27015 18522
rect 27015 18470 27025 18522
rect 27049 18470 27079 18522
rect 27079 18470 27091 18522
rect 27091 18470 27105 18522
rect 27129 18470 27143 18522
rect 27143 18470 27155 18522
rect 27155 18470 27185 18522
rect 27209 18470 27219 18522
rect 27219 18470 27265 18522
rect 26969 18468 27025 18470
rect 27049 18468 27105 18470
rect 27129 18468 27185 18470
rect 27209 18468 27265 18470
rect 27066 17876 27122 17912
rect 27066 17856 27068 17876
rect 27068 17856 27120 17876
rect 27120 17856 27122 17876
rect 26969 17434 27025 17436
rect 27049 17434 27105 17436
rect 27129 17434 27185 17436
rect 27209 17434 27265 17436
rect 26969 17382 27015 17434
rect 27015 17382 27025 17434
rect 27049 17382 27079 17434
rect 27079 17382 27091 17434
rect 27091 17382 27105 17434
rect 27129 17382 27143 17434
rect 27143 17382 27155 17434
rect 27155 17382 27185 17434
rect 27209 17382 27219 17434
rect 27219 17382 27265 17434
rect 26969 17380 27025 17382
rect 27049 17380 27105 17382
rect 27129 17380 27185 17382
rect 27209 17380 27265 17382
rect 26698 17040 26754 17096
rect 26606 16632 26662 16688
rect 26790 15680 26846 15736
rect 26514 14320 26570 14376
rect 25134 11600 25190 11656
rect 24214 10648 24270 10704
rect 24214 10548 24216 10568
rect 24216 10548 24268 10568
rect 24268 10548 24270 10568
rect 23174 10362 23230 10364
rect 23254 10362 23310 10364
rect 23334 10362 23390 10364
rect 23414 10362 23470 10364
rect 23174 10310 23220 10362
rect 23220 10310 23230 10362
rect 23254 10310 23284 10362
rect 23284 10310 23296 10362
rect 23296 10310 23310 10362
rect 23334 10310 23348 10362
rect 23348 10310 23360 10362
rect 23360 10310 23390 10362
rect 23414 10310 23424 10362
rect 23424 10310 23470 10362
rect 23174 10308 23230 10310
rect 23254 10308 23310 10310
rect 23334 10308 23390 10310
rect 23414 10308 23470 10310
rect 24214 10512 24270 10548
rect 24122 9460 24124 9480
rect 24124 9460 24176 9480
rect 24176 9460 24178 9480
rect 24122 9424 24178 9460
rect 23174 9274 23230 9276
rect 23254 9274 23310 9276
rect 23334 9274 23390 9276
rect 23414 9274 23470 9276
rect 23174 9222 23220 9274
rect 23220 9222 23230 9274
rect 23254 9222 23284 9274
rect 23284 9222 23296 9274
rect 23296 9222 23310 9274
rect 23334 9222 23348 9274
rect 23348 9222 23360 9274
rect 23360 9222 23390 9274
rect 23414 9222 23424 9274
rect 23424 9222 23470 9274
rect 23174 9220 23230 9222
rect 23254 9220 23310 9222
rect 23334 9220 23390 9222
rect 23414 9220 23470 9222
rect 24766 9580 24822 9616
rect 24766 9560 24768 9580
rect 24768 9560 24820 9580
rect 24820 9560 24822 9580
rect 23174 8186 23230 8188
rect 23254 8186 23310 8188
rect 23334 8186 23390 8188
rect 23414 8186 23470 8188
rect 23174 8134 23220 8186
rect 23220 8134 23230 8186
rect 23254 8134 23284 8186
rect 23284 8134 23296 8186
rect 23296 8134 23310 8186
rect 23334 8134 23348 8186
rect 23348 8134 23360 8186
rect 23360 8134 23390 8186
rect 23414 8134 23424 8186
rect 23424 8134 23470 8186
rect 23174 8132 23230 8134
rect 23254 8132 23310 8134
rect 23334 8132 23390 8134
rect 23414 8132 23470 8134
rect 22650 6704 22706 6760
rect 23174 7098 23230 7100
rect 23254 7098 23310 7100
rect 23334 7098 23390 7100
rect 23414 7098 23470 7100
rect 23174 7046 23220 7098
rect 23220 7046 23230 7098
rect 23254 7046 23284 7098
rect 23284 7046 23296 7098
rect 23296 7046 23310 7098
rect 23334 7046 23348 7098
rect 23348 7046 23360 7098
rect 23360 7046 23390 7098
rect 23414 7046 23424 7098
rect 23424 7046 23470 7098
rect 23174 7044 23230 7046
rect 23254 7044 23310 7046
rect 23334 7044 23390 7046
rect 23414 7044 23470 7046
rect 23386 6316 23442 6352
rect 23386 6296 23388 6316
rect 23388 6296 23440 6316
rect 23440 6296 23442 6316
rect 21638 4528 21694 4584
rect 22374 5616 22430 5672
rect 23174 6010 23230 6012
rect 23254 6010 23310 6012
rect 23334 6010 23390 6012
rect 23414 6010 23470 6012
rect 23174 5958 23220 6010
rect 23220 5958 23230 6010
rect 23254 5958 23284 6010
rect 23284 5958 23296 6010
rect 23296 5958 23310 6010
rect 23334 5958 23348 6010
rect 23348 5958 23360 6010
rect 23360 5958 23390 6010
rect 23414 5958 23424 6010
rect 23424 5958 23470 6010
rect 23174 5956 23230 5958
rect 23254 5956 23310 5958
rect 23334 5956 23390 5958
rect 23414 5956 23470 5958
rect 23386 5752 23442 5808
rect 23174 4922 23230 4924
rect 23254 4922 23310 4924
rect 23334 4922 23390 4924
rect 23414 4922 23470 4924
rect 23174 4870 23220 4922
rect 23220 4870 23230 4922
rect 23254 4870 23284 4922
rect 23284 4870 23296 4922
rect 23296 4870 23310 4922
rect 23334 4870 23348 4922
rect 23348 4870 23360 4922
rect 23360 4870 23390 4922
rect 23414 4870 23424 4922
rect 23424 4870 23470 4922
rect 23174 4868 23230 4870
rect 23254 4868 23310 4870
rect 23334 4868 23390 4870
rect 23414 4868 23470 4870
rect 23174 3834 23230 3836
rect 23254 3834 23310 3836
rect 23334 3834 23390 3836
rect 23414 3834 23470 3836
rect 23174 3782 23220 3834
rect 23220 3782 23230 3834
rect 23254 3782 23284 3834
rect 23284 3782 23296 3834
rect 23296 3782 23310 3834
rect 23334 3782 23348 3834
rect 23348 3782 23360 3834
rect 23360 3782 23390 3834
rect 23414 3782 23424 3834
rect 23424 3782 23470 3834
rect 23174 3780 23230 3782
rect 23254 3780 23310 3782
rect 23334 3780 23390 3782
rect 23414 3780 23470 3782
rect 24030 6976 24086 7032
rect 23174 2746 23230 2748
rect 23254 2746 23310 2748
rect 23334 2746 23390 2748
rect 23414 2746 23470 2748
rect 23174 2694 23220 2746
rect 23220 2694 23230 2746
rect 23254 2694 23284 2746
rect 23284 2694 23296 2746
rect 23296 2694 23310 2746
rect 23334 2694 23348 2746
rect 23348 2694 23360 2746
rect 23360 2694 23390 2746
rect 23414 2694 23424 2746
rect 23424 2694 23470 2746
rect 23174 2692 23230 2694
rect 23254 2692 23310 2694
rect 23334 2692 23390 2694
rect 23414 2692 23470 2694
rect 24858 5752 24914 5808
rect 25318 11228 25320 11248
rect 25320 11228 25372 11248
rect 25372 11228 25374 11248
rect 25318 11192 25374 11228
rect 25042 9424 25098 9480
rect 25318 7792 25374 7848
rect 25134 7112 25190 7168
rect 25318 6976 25374 7032
rect 21914 2216 21970 2272
rect 22006 720 22062 776
rect 23294 1844 23296 1864
rect 23296 1844 23348 1864
rect 23348 1844 23350 1864
rect 23294 1808 23350 1844
rect 23174 1658 23230 1660
rect 23254 1658 23310 1660
rect 23334 1658 23390 1660
rect 23414 1658 23470 1660
rect 23174 1606 23220 1658
rect 23220 1606 23230 1658
rect 23254 1606 23284 1658
rect 23284 1606 23296 1658
rect 23296 1606 23310 1658
rect 23334 1606 23348 1658
rect 23348 1606 23360 1658
rect 23360 1606 23390 1658
rect 23414 1606 23424 1658
rect 23424 1606 23470 1658
rect 23174 1604 23230 1606
rect 23254 1604 23310 1606
rect 23334 1604 23390 1606
rect 23414 1604 23470 1606
rect 23478 856 23534 912
rect 23174 570 23230 572
rect 23254 570 23310 572
rect 23334 570 23390 572
rect 23414 570 23470 572
rect 23174 518 23220 570
rect 23220 518 23230 570
rect 23254 518 23284 570
rect 23284 518 23296 570
rect 23296 518 23310 570
rect 23334 518 23348 570
rect 23348 518 23360 570
rect 23360 518 23390 570
rect 23414 518 23424 570
rect 23424 518 23470 570
rect 23174 516 23230 518
rect 23254 516 23310 518
rect 23334 516 23390 518
rect 23414 516 23470 518
rect 23938 720 23994 776
rect 26146 12552 26202 12608
rect 25870 10784 25926 10840
rect 26054 9560 26110 9616
rect 25962 8336 26018 8392
rect 25870 6724 25926 6760
rect 25870 6704 25872 6724
rect 25872 6704 25924 6724
rect 25924 6704 25926 6724
rect 26238 6604 26240 6624
rect 26240 6604 26292 6624
rect 26292 6604 26294 6624
rect 26238 6568 26294 6604
rect 26790 15272 26846 15328
rect 26790 14456 26846 14512
rect 26969 16346 27025 16348
rect 27049 16346 27105 16348
rect 27129 16346 27185 16348
rect 27209 16346 27265 16348
rect 26969 16294 27015 16346
rect 27015 16294 27025 16346
rect 27049 16294 27079 16346
rect 27079 16294 27091 16346
rect 27091 16294 27105 16346
rect 27129 16294 27143 16346
rect 27143 16294 27155 16346
rect 27155 16294 27185 16346
rect 27209 16294 27219 16346
rect 27219 16294 27265 16346
rect 26969 16292 27025 16294
rect 27049 16292 27105 16294
rect 27129 16292 27185 16294
rect 27209 16292 27265 16294
rect 26969 15258 27025 15260
rect 27049 15258 27105 15260
rect 27129 15258 27185 15260
rect 27209 15258 27265 15260
rect 26969 15206 27015 15258
rect 27015 15206 27025 15258
rect 27049 15206 27079 15258
rect 27079 15206 27091 15258
rect 27091 15206 27105 15258
rect 27129 15206 27143 15258
rect 27143 15206 27155 15258
rect 27155 15206 27185 15258
rect 27209 15206 27219 15258
rect 27219 15206 27265 15258
rect 26969 15204 27025 15206
rect 27049 15204 27105 15206
rect 27129 15204 27185 15206
rect 27209 15204 27265 15206
rect 27434 16768 27490 16824
rect 27710 17992 27766 18048
rect 26698 14048 26754 14104
rect 26514 12416 26570 12472
rect 26790 13912 26846 13968
rect 26969 14170 27025 14172
rect 27049 14170 27105 14172
rect 27129 14170 27185 14172
rect 27209 14170 27265 14172
rect 26969 14118 27015 14170
rect 27015 14118 27025 14170
rect 27049 14118 27079 14170
rect 27079 14118 27091 14170
rect 27091 14118 27105 14170
rect 27129 14118 27143 14170
rect 27143 14118 27155 14170
rect 27155 14118 27185 14170
rect 27209 14118 27219 14170
rect 27219 14118 27265 14170
rect 26969 14116 27025 14118
rect 27049 14116 27105 14118
rect 27129 14116 27185 14118
rect 27209 14116 27265 14118
rect 27618 15544 27674 15600
rect 27894 16224 27950 16280
rect 26969 13082 27025 13084
rect 27049 13082 27105 13084
rect 27129 13082 27185 13084
rect 27209 13082 27265 13084
rect 26969 13030 27015 13082
rect 27015 13030 27025 13082
rect 27049 13030 27079 13082
rect 27079 13030 27091 13082
rect 27091 13030 27105 13082
rect 27129 13030 27143 13082
rect 27143 13030 27155 13082
rect 27155 13030 27185 13082
rect 27209 13030 27219 13082
rect 27219 13030 27265 13082
rect 26969 13028 27025 13030
rect 27049 13028 27105 13030
rect 27129 13028 27185 13030
rect 27209 13028 27265 13030
rect 26969 11994 27025 11996
rect 27049 11994 27105 11996
rect 27129 11994 27185 11996
rect 27209 11994 27265 11996
rect 26969 11942 27015 11994
rect 27015 11942 27025 11994
rect 27049 11942 27079 11994
rect 27079 11942 27091 11994
rect 27091 11942 27105 11994
rect 27129 11942 27143 11994
rect 27143 11942 27155 11994
rect 27155 11942 27185 11994
rect 27209 11942 27219 11994
rect 27219 11942 27265 11994
rect 26969 11940 27025 11942
rect 27049 11940 27105 11942
rect 27129 11940 27185 11942
rect 27209 11940 27265 11942
rect 27158 11636 27160 11656
rect 27160 11636 27212 11656
rect 27212 11636 27214 11656
rect 27158 11600 27214 11636
rect 26969 10906 27025 10908
rect 27049 10906 27105 10908
rect 27129 10906 27185 10908
rect 27209 10906 27265 10908
rect 26969 10854 27015 10906
rect 27015 10854 27025 10906
rect 27049 10854 27079 10906
rect 27079 10854 27091 10906
rect 27091 10854 27105 10906
rect 27129 10854 27143 10906
rect 27143 10854 27155 10906
rect 27155 10854 27185 10906
rect 27209 10854 27219 10906
rect 27219 10854 27265 10906
rect 26969 10852 27025 10854
rect 27049 10852 27105 10854
rect 27129 10852 27185 10854
rect 27209 10852 27265 10854
rect 26969 9818 27025 9820
rect 27049 9818 27105 9820
rect 27129 9818 27185 9820
rect 27209 9818 27265 9820
rect 26969 9766 27015 9818
rect 27015 9766 27025 9818
rect 27049 9766 27079 9818
rect 27079 9766 27091 9818
rect 27091 9766 27105 9818
rect 27129 9766 27143 9818
rect 27143 9766 27155 9818
rect 27155 9766 27185 9818
rect 27209 9766 27219 9818
rect 27219 9766 27265 9818
rect 26969 9764 27025 9766
rect 27049 9764 27105 9766
rect 27129 9764 27185 9766
rect 27209 9764 27265 9766
rect 26514 7112 26570 7168
rect 26514 6704 26570 6760
rect 26330 3032 26386 3088
rect 25594 2080 25650 2136
rect 25594 1420 25650 1456
rect 26969 8730 27025 8732
rect 27049 8730 27105 8732
rect 27129 8730 27185 8732
rect 27209 8730 27265 8732
rect 26969 8678 27015 8730
rect 27015 8678 27025 8730
rect 27049 8678 27079 8730
rect 27079 8678 27091 8730
rect 27091 8678 27105 8730
rect 27129 8678 27143 8730
rect 27143 8678 27155 8730
rect 27155 8678 27185 8730
rect 27209 8678 27219 8730
rect 27219 8678 27265 8730
rect 26969 8676 27025 8678
rect 27049 8676 27105 8678
rect 27129 8676 27185 8678
rect 27209 8676 27265 8678
rect 27986 14320 28042 14376
rect 28078 13368 28134 13424
rect 28262 12144 28318 12200
rect 27710 8880 27766 8936
rect 26969 7642 27025 7644
rect 27049 7642 27105 7644
rect 27129 7642 27185 7644
rect 27209 7642 27265 7644
rect 26969 7590 27015 7642
rect 27015 7590 27025 7642
rect 27049 7590 27079 7642
rect 27079 7590 27091 7642
rect 27091 7590 27105 7642
rect 27129 7590 27143 7642
rect 27143 7590 27155 7642
rect 27155 7590 27185 7642
rect 27209 7590 27219 7642
rect 27219 7590 27265 7642
rect 26969 7588 27025 7590
rect 27049 7588 27105 7590
rect 27129 7588 27185 7590
rect 27209 7588 27265 7590
rect 27250 7148 27252 7168
rect 27252 7148 27304 7168
rect 27304 7148 27306 7168
rect 27250 7112 27306 7148
rect 26969 6554 27025 6556
rect 27049 6554 27105 6556
rect 27129 6554 27185 6556
rect 27209 6554 27265 6556
rect 26969 6502 27015 6554
rect 27015 6502 27025 6554
rect 27049 6502 27079 6554
rect 27079 6502 27091 6554
rect 27091 6502 27105 6554
rect 27129 6502 27143 6554
rect 27143 6502 27155 6554
rect 27155 6502 27185 6554
rect 27209 6502 27219 6554
rect 27219 6502 27265 6554
rect 26969 6500 27025 6502
rect 27049 6500 27105 6502
rect 27129 6500 27185 6502
rect 27209 6500 27265 6502
rect 27066 6296 27122 6352
rect 26974 5772 27030 5808
rect 26974 5752 26976 5772
rect 26976 5752 27028 5772
rect 27028 5752 27030 5772
rect 26606 4528 26662 4584
rect 26969 5466 27025 5468
rect 27049 5466 27105 5468
rect 27129 5466 27185 5468
rect 27209 5466 27265 5468
rect 26969 5414 27015 5466
rect 27015 5414 27025 5466
rect 27049 5414 27079 5466
rect 27079 5414 27091 5466
rect 27091 5414 27105 5466
rect 27129 5414 27143 5466
rect 27143 5414 27155 5466
rect 27155 5414 27185 5466
rect 27209 5414 27219 5466
rect 27219 5414 27265 5466
rect 26969 5412 27025 5414
rect 27049 5412 27105 5414
rect 27129 5412 27185 5414
rect 27209 5412 27265 5414
rect 27894 6840 27950 6896
rect 28722 20848 28778 20904
rect 28630 16496 28686 16552
rect 28722 16224 28778 16280
rect 28722 15972 28778 16008
rect 28722 15952 28724 15972
rect 28724 15952 28776 15972
rect 28776 15952 28778 15972
rect 29182 19352 29238 19408
rect 29090 15000 29146 15056
rect 28906 13912 28962 13968
rect 28170 6332 28172 6352
rect 28172 6332 28224 6352
rect 28224 6332 28226 6352
rect 28170 6296 28226 6332
rect 28170 5652 28172 5672
rect 28172 5652 28224 5672
rect 28224 5652 28226 5672
rect 28170 5616 28226 5652
rect 26969 4378 27025 4380
rect 27049 4378 27105 4380
rect 27129 4378 27185 4380
rect 27209 4378 27265 4380
rect 26969 4326 27015 4378
rect 27015 4326 27025 4378
rect 27049 4326 27079 4378
rect 27079 4326 27091 4378
rect 27091 4326 27105 4378
rect 27129 4326 27143 4378
rect 27143 4326 27155 4378
rect 27155 4326 27185 4378
rect 27209 4326 27219 4378
rect 27219 4326 27265 4378
rect 26969 4324 27025 4326
rect 27049 4324 27105 4326
rect 27129 4324 27185 4326
rect 27209 4324 27265 4326
rect 26969 3290 27025 3292
rect 27049 3290 27105 3292
rect 27129 3290 27185 3292
rect 27209 3290 27265 3292
rect 26969 3238 27015 3290
rect 27015 3238 27025 3290
rect 27049 3238 27079 3290
rect 27079 3238 27091 3290
rect 27091 3238 27105 3290
rect 27129 3238 27143 3290
rect 27143 3238 27155 3290
rect 27155 3238 27185 3290
rect 27209 3238 27219 3290
rect 27219 3238 27265 3290
rect 26969 3236 27025 3238
rect 27049 3236 27105 3238
rect 27129 3236 27185 3238
rect 27209 3236 27265 3238
rect 26238 1808 26294 1864
rect 25594 1400 25596 1420
rect 25596 1400 25648 1420
rect 25648 1400 25650 1420
rect 25686 1264 25742 1320
rect 26969 2202 27025 2204
rect 27049 2202 27105 2204
rect 27129 2202 27185 2204
rect 27209 2202 27265 2204
rect 26969 2150 27015 2202
rect 27015 2150 27025 2202
rect 27049 2150 27079 2202
rect 27079 2150 27091 2202
rect 27091 2150 27105 2202
rect 27129 2150 27143 2202
rect 27143 2150 27155 2202
rect 27155 2150 27185 2202
rect 27209 2150 27219 2202
rect 27219 2150 27265 2202
rect 26969 2148 27025 2150
rect 27049 2148 27105 2150
rect 27129 2148 27185 2150
rect 27209 2148 27265 2150
rect 27526 3440 27582 3496
rect 25686 1012 25742 1048
rect 25686 992 25688 1012
rect 25688 992 25740 1012
rect 25740 992 25742 1012
rect 26969 1114 27025 1116
rect 27049 1114 27105 1116
rect 27129 1114 27185 1116
rect 27209 1114 27265 1116
rect 26969 1062 27015 1114
rect 27015 1062 27025 1114
rect 27049 1062 27079 1114
rect 27079 1062 27091 1114
rect 27091 1062 27105 1114
rect 27129 1062 27143 1114
rect 27143 1062 27155 1114
rect 27155 1062 27185 1114
rect 27209 1062 27219 1114
rect 27219 1062 27265 1114
rect 26969 1060 27025 1062
rect 27049 1060 27105 1062
rect 27129 1060 27185 1062
rect 27209 1060 27265 1062
rect 28354 2896 28410 2952
rect 28630 5208 28686 5264
rect 29366 16088 29422 16144
rect 29366 15852 29368 15872
rect 29368 15852 29420 15872
rect 29420 15852 29422 15872
rect 29366 15816 29422 15852
rect 29274 15308 29276 15328
rect 29276 15308 29328 15328
rect 29328 15308 29330 15328
rect 29274 15272 29330 15308
rect 29642 15988 29644 16008
rect 29644 15988 29696 16008
rect 29696 15988 29698 16008
rect 29642 15952 29698 15988
rect 29642 15680 29698 15736
rect 30194 18264 30250 18320
rect 30194 18128 30250 18184
rect 30470 17620 30472 17640
rect 30472 17620 30524 17640
rect 30524 17620 30526 17640
rect 30470 17584 30526 17620
rect 30764 21242 30820 21244
rect 30844 21242 30900 21244
rect 30924 21242 30980 21244
rect 31004 21242 31060 21244
rect 30764 21190 30810 21242
rect 30810 21190 30820 21242
rect 30844 21190 30874 21242
rect 30874 21190 30886 21242
rect 30886 21190 30900 21242
rect 30924 21190 30938 21242
rect 30938 21190 30950 21242
rect 30950 21190 30980 21242
rect 31004 21190 31014 21242
rect 31014 21190 31060 21242
rect 30764 21188 30820 21190
rect 30844 21188 30900 21190
rect 30924 21188 30980 21190
rect 31004 21188 31060 21190
rect 30764 20154 30820 20156
rect 30844 20154 30900 20156
rect 30924 20154 30980 20156
rect 31004 20154 31060 20156
rect 30764 20102 30810 20154
rect 30810 20102 30820 20154
rect 30844 20102 30874 20154
rect 30874 20102 30886 20154
rect 30886 20102 30900 20154
rect 30924 20102 30938 20154
rect 30938 20102 30950 20154
rect 30950 20102 30980 20154
rect 31004 20102 31014 20154
rect 31014 20102 31060 20154
rect 30764 20100 30820 20102
rect 30844 20100 30900 20102
rect 30924 20100 30980 20102
rect 31004 20100 31060 20102
rect 30010 14900 30012 14920
rect 30012 14900 30064 14920
rect 30064 14900 30066 14920
rect 30010 14864 30066 14900
rect 30194 14592 30250 14648
rect 30378 15952 30434 16008
rect 29550 12552 29606 12608
rect 29550 12416 29606 12472
rect 28998 6704 29054 6760
rect 28630 3984 28686 4040
rect 29090 2372 29146 2408
rect 29090 2352 29092 2372
rect 29092 2352 29144 2372
rect 29144 2352 29146 2372
rect 29182 1980 29184 2000
rect 29184 1980 29236 2000
rect 29236 1980 29238 2000
rect 29182 1944 29238 1980
rect 29826 13812 29828 13832
rect 29828 13812 29880 13832
rect 29880 13812 29882 13832
rect 29826 13776 29882 13812
rect 29918 13096 29974 13152
rect 29826 12824 29882 12880
rect 30010 12688 30066 12744
rect 30378 12300 30434 12336
rect 30378 12280 30380 12300
rect 30380 12280 30432 12300
rect 30432 12280 30434 12300
rect 29366 5072 29422 5128
rect 30764 19066 30820 19068
rect 30844 19066 30900 19068
rect 30924 19066 30980 19068
rect 31004 19066 31060 19068
rect 30764 19014 30810 19066
rect 30810 19014 30820 19066
rect 30844 19014 30874 19066
rect 30874 19014 30886 19066
rect 30886 19014 30900 19066
rect 30924 19014 30938 19066
rect 30938 19014 30950 19066
rect 30950 19014 30980 19066
rect 31004 19014 31014 19066
rect 31014 19014 31060 19066
rect 30764 19012 30820 19014
rect 30844 19012 30900 19014
rect 30924 19012 30980 19014
rect 31004 19012 31060 19014
rect 30764 17978 30820 17980
rect 30844 17978 30900 17980
rect 30924 17978 30980 17980
rect 31004 17978 31060 17980
rect 30764 17926 30810 17978
rect 30810 17926 30820 17978
rect 30844 17926 30874 17978
rect 30874 17926 30886 17978
rect 30886 17926 30900 17978
rect 30924 17926 30938 17978
rect 30938 17926 30950 17978
rect 30950 17926 30980 17978
rect 31004 17926 31014 17978
rect 31014 17926 31060 17978
rect 30764 17924 30820 17926
rect 30844 17924 30900 17926
rect 30924 17924 30980 17926
rect 31004 17924 31060 17926
rect 30764 16890 30820 16892
rect 30844 16890 30900 16892
rect 30924 16890 30980 16892
rect 31004 16890 31060 16892
rect 30764 16838 30810 16890
rect 30810 16838 30820 16890
rect 30844 16838 30874 16890
rect 30874 16838 30886 16890
rect 30886 16838 30900 16890
rect 30924 16838 30938 16890
rect 30938 16838 30950 16890
rect 30950 16838 30980 16890
rect 31004 16838 31014 16890
rect 31014 16838 31060 16890
rect 30764 16836 30820 16838
rect 30844 16836 30900 16838
rect 30924 16836 30980 16838
rect 31004 16836 31060 16838
rect 30764 15802 30820 15804
rect 30844 15802 30900 15804
rect 30924 15802 30980 15804
rect 31004 15802 31060 15804
rect 30764 15750 30810 15802
rect 30810 15750 30820 15802
rect 30844 15750 30874 15802
rect 30874 15750 30886 15802
rect 30886 15750 30900 15802
rect 30924 15750 30938 15802
rect 30938 15750 30950 15802
rect 30950 15750 30980 15802
rect 31004 15750 31014 15802
rect 31014 15750 31060 15802
rect 30764 15748 30820 15750
rect 30844 15748 30900 15750
rect 30924 15748 30980 15750
rect 31004 15748 31060 15750
rect 30764 14714 30820 14716
rect 30844 14714 30900 14716
rect 30924 14714 30980 14716
rect 31004 14714 31060 14716
rect 30764 14662 30810 14714
rect 30810 14662 30820 14714
rect 30844 14662 30874 14714
rect 30874 14662 30886 14714
rect 30886 14662 30900 14714
rect 30924 14662 30938 14714
rect 30938 14662 30950 14714
rect 30950 14662 30980 14714
rect 31004 14662 31014 14714
rect 31014 14662 31060 14714
rect 30764 14660 30820 14662
rect 30844 14660 30900 14662
rect 30924 14660 30980 14662
rect 31004 14660 31060 14662
rect 29458 1264 29514 1320
rect 30764 13626 30820 13628
rect 30844 13626 30900 13628
rect 30924 13626 30980 13628
rect 31004 13626 31060 13628
rect 30764 13574 30810 13626
rect 30810 13574 30820 13626
rect 30844 13574 30874 13626
rect 30874 13574 30886 13626
rect 30886 13574 30900 13626
rect 30924 13574 30938 13626
rect 30938 13574 30950 13626
rect 30950 13574 30980 13626
rect 31004 13574 31014 13626
rect 31014 13574 31060 13626
rect 30764 13572 30820 13574
rect 30844 13572 30900 13574
rect 30924 13572 30980 13574
rect 31004 13572 31060 13574
rect 30764 12538 30820 12540
rect 30844 12538 30900 12540
rect 30924 12538 30980 12540
rect 31004 12538 31060 12540
rect 30764 12486 30810 12538
rect 30810 12486 30820 12538
rect 30844 12486 30874 12538
rect 30874 12486 30886 12538
rect 30886 12486 30900 12538
rect 30924 12486 30938 12538
rect 30938 12486 30950 12538
rect 30950 12486 30980 12538
rect 31004 12486 31014 12538
rect 31014 12486 31060 12538
rect 30764 12484 30820 12486
rect 30844 12484 30900 12486
rect 30924 12484 30980 12486
rect 31004 12484 31060 12486
rect 30764 11450 30820 11452
rect 30844 11450 30900 11452
rect 30924 11450 30980 11452
rect 31004 11450 31060 11452
rect 30764 11398 30810 11450
rect 30810 11398 30820 11450
rect 30844 11398 30874 11450
rect 30874 11398 30886 11450
rect 30886 11398 30900 11450
rect 30924 11398 30938 11450
rect 30938 11398 30950 11450
rect 30950 11398 30980 11450
rect 31004 11398 31014 11450
rect 31014 11398 31060 11450
rect 30764 11396 30820 11398
rect 30844 11396 30900 11398
rect 30924 11396 30980 11398
rect 31004 11396 31060 11398
rect 31114 11056 31170 11112
rect 30764 10362 30820 10364
rect 30844 10362 30900 10364
rect 30924 10362 30980 10364
rect 31004 10362 31060 10364
rect 30764 10310 30810 10362
rect 30810 10310 30820 10362
rect 30844 10310 30874 10362
rect 30874 10310 30886 10362
rect 30886 10310 30900 10362
rect 30924 10310 30938 10362
rect 30938 10310 30950 10362
rect 30950 10310 30980 10362
rect 31004 10310 31014 10362
rect 31014 10310 31060 10362
rect 30764 10308 30820 10310
rect 30844 10308 30900 10310
rect 30924 10308 30980 10310
rect 31004 10308 31060 10310
rect 30764 9274 30820 9276
rect 30844 9274 30900 9276
rect 30924 9274 30980 9276
rect 31004 9274 31060 9276
rect 30764 9222 30810 9274
rect 30810 9222 30820 9274
rect 30844 9222 30874 9274
rect 30874 9222 30886 9274
rect 30886 9222 30900 9274
rect 30924 9222 30938 9274
rect 30938 9222 30950 9274
rect 30950 9222 30980 9274
rect 31004 9222 31014 9274
rect 31014 9222 31060 9274
rect 30764 9220 30820 9222
rect 30844 9220 30900 9222
rect 30924 9220 30980 9222
rect 31004 9220 31060 9222
rect 30764 8186 30820 8188
rect 30844 8186 30900 8188
rect 30924 8186 30980 8188
rect 31004 8186 31060 8188
rect 30764 8134 30810 8186
rect 30810 8134 30820 8186
rect 30844 8134 30874 8186
rect 30874 8134 30886 8186
rect 30886 8134 30900 8186
rect 30924 8134 30938 8186
rect 30938 8134 30950 8186
rect 30950 8134 30980 8186
rect 31004 8134 31014 8186
rect 31014 8134 31060 8186
rect 30764 8132 30820 8134
rect 30844 8132 30900 8134
rect 30924 8132 30980 8134
rect 31004 8132 31060 8134
rect 30764 7098 30820 7100
rect 30844 7098 30900 7100
rect 30924 7098 30980 7100
rect 31004 7098 31060 7100
rect 30764 7046 30810 7098
rect 30810 7046 30820 7098
rect 30844 7046 30874 7098
rect 30874 7046 30886 7098
rect 30886 7046 30900 7098
rect 30924 7046 30938 7098
rect 30938 7046 30950 7098
rect 30950 7046 30980 7098
rect 31004 7046 31014 7098
rect 31014 7046 31060 7098
rect 30764 7044 30820 7046
rect 30844 7044 30900 7046
rect 30924 7044 30980 7046
rect 31004 7044 31060 7046
rect 30764 6010 30820 6012
rect 30844 6010 30900 6012
rect 30924 6010 30980 6012
rect 31004 6010 31060 6012
rect 30764 5958 30810 6010
rect 30810 5958 30820 6010
rect 30844 5958 30874 6010
rect 30874 5958 30886 6010
rect 30886 5958 30900 6010
rect 30924 5958 30938 6010
rect 30938 5958 30950 6010
rect 30950 5958 30980 6010
rect 31004 5958 31014 6010
rect 31014 5958 31060 6010
rect 30764 5956 30820 5958
rect 30844 5956 30900 5958
rect 30924 5956 30980 5958
rect 31004 5956 31060 5958
rect 31390 17176 31446 17232
rect 30764 4922 30820 4924
rect 30844 4922 30900 4924
rect 30924 4922 30980 4924
rect 31004 4922 31060 4924
rect 30764 4870 30810 4922
rect 30810 4870 30820 4922
rect 30844 4870 30874 4922
rect 30874 4870 30886 4922
rect 30886 4870 30900 4922
rect 30924 4870 30938 4922
rect 30938 4870 30950 4922
rect 30950 4870 30980 4922
rect 31004 4870 31014 4922
rect 31014 4870 31060 4922
rect 30764 4868 30820 4870
rect 30844 4868 30900 4870
rect 30924 4868 30980 4870
rect 31004 4868 31060 4870
rect 30764 3834 30820 3836
rect 30844 3834 30900 3836
rect 30924 3834 30980 3836
rect 31004 3834 31060 3836
rect 30764 3782 30810 3834
rect 30810 3782 30820 3834
rect 30844 3782 30874 3834
rect 30874 3782 30886 3834
rect 30886 3782 30900 3834
rect 30924 3782 30938 3834
rect 30938 3782 30950 3834
rect 30950 3782 30980 3834
rect 31004 3782 31014 3834
rect 31014 3782 31060 3834
rect 30764 3780 30820 3782
rect 30844 3780 30900 3782
rect 30924 3780 30980 3782
rect 31004 3780 31060 3782
rect 30764 2746 30820 2748
rect 30844 2746 30900 2748
rect 30924 2746 30980 2748
rect 31004 2746 31060 2748
rect 30764 2694 30810 2746
rect 30810 2694 30820 2746
rect 30844 2694 30874 2746
rect 30874 2694 30886 2746
rect 30886 2694 30900 2746
rect 30924 2694 30938 2746
rect 30938 2694 30950 2746
rect 30950 2694 30980 2746
rect 31004 2694 31014 2746
rect 31014 2694 31060 2746
rect 30764 2692 30820 2694
rect 30844 2692 30900 2694
rect 30924 2692 30980 2694
rect 31004 2692 31060 2694
rect 30764 1658 30820 1660
rect 30844 1658 30900 1660
rect 30924 1658 30980 1660
rect 31004 1658 31060 1660
rect 30764 1606 30810 1658
rect 30810 1606 30820 1658
rect 30844 1606 30874 1658
rect 30874 1606 30886 1658
rect 30886 1606 30900 1658
rect 30924 1606 30938 1658
rect 30938 1606 30950 1658
rect 30950 1606 30980 1658
rect 31004 1606 31014 1658
rect 31014 1606 31060 1658
rect 30764 1604 30820 1606
rect 30844 1604 30900 1606
rect 30924 1604 30980 1606
rect 31004 1604 31060 1606
rect 28998 720 29054 776
rect 30764 570 30820 572
rect 30844 570 30900 572
rect 30924 570 30980 572
rect 31004 570 31060 572
rect 30764 518 30810 570
rect 30810 518 30820 570
rect 30844 518 30874 570
rect 30874 518 30886 570
rect 30886 518 30900 570
rect 30924 518 30938 570
rect 30938 518 30950 570
rect 30950 518 30980 570
rect 31004 518 31014 570
rect 31014 518 31060 570
rect 30764 516 30820 518
rect 30844 516 30900 518
rect 30924 516 30980 518
rect 31004 516 31060 518
rect 29918 312 29974 368
<< metal3 >>
rect 5073 22266 5139 22269
rect 11145 22266 11211 22269
rect 5073 22264 11211 22266
rect 5073 22208 5078 22264
rect 5134 22208 11150 22264
rect 11206 22208 11211 22264
rect 5073 22206 11211 22208
rect 5073 22203 5139 22206
rect 11145 22203 11211 22206
rect 10041 22130 10107 22133
rect 10174 22130 10180 22132
rect 10041 22128 10180 22130
rect 10041 22072 10046 22128
rect 10102 22072 10180 22128
rect 10041 22070 10180 22072
rect 10041 22067 10107 22070
rect 10174 22068 10180 22070
rect 10244 22068 10250 22132
rect 10961 22130 11027 22133
rect 14406 22130 14412 22132
rect 10961 22128 14412 22130
rect 10961 22072 10966 22128
rect 11022 22072 14412 22128
rect 10961 22070 14412 22072
rect 10961 22067 11027 22070
rect 14406 22068 14412 22070
rect 14476 22068 14482 22132
rect 19333 22130 19399 22133
rect 22461 22130 22527 22133
rect 19333 22128 22527 22130
rect 19333 22072 19338 22128
rect 19394 22072 22466 22128
rect 22522 22072 22527 22128
rect 19333 22070 22527 22072
rect 19333 22067 19399 22070
rect 22461 22067 22527 22070
rect 2497 21994 2563 21997
rect 8702 21994 8708 21996
rect 2497 21992 8708 21994
rect 2497 21936 2502 21992
rect 2558 21936 8708 21992
rect 2497 21934 8708 21936
rect 2497 21931 2563 21934
rect 8702 21932 8708 21934
rect 8772 21932 8778 21996
rect 10225 21994 10291 21997
rect 13813 21996 13879 21997
rect 12566 21994 12572 21996
rect 10225 21992 12572 21994
rect 10225 21936 10230 21992
rect 10286 21936 12572 21992
rect 10225 21934 12572 21936
rect 10225 21931 10291 21934
rect 12566 21932 12572 21934
rect 12636 21932 12642 21996
rect 13813 21992 13860 21996
rect 13924 21994 13930 21996
rect 13813 21936 13818 21992
rect 13813 21932 13860 21936
rect 13924 21934 13970 21994
rect 13924 21932 13930 21934
rect 13813 21931 13879 21932
rect 8569 21858 8635 21861
rect 23565 21860 23631 21861
rect 9254 21858 9260 21860
rect 8569 21856 9260 21858
rect 8569 21800 8574 21856
rect 8630 21800 9260 21856
rect 8569 21798 9260 21800
rect 8569 21795 8635 21798
rect 9254 21796 9260 21798
rect 9324 21796 9330 21860
rect 23565 21858 23612 21860
rect 23520 21856 23612 21858
rect 23520 21800 23570 21856
rect 23520 21798 23612 21800
rect 23565 21796 23612 21798
rect 23676 21796 23682 21860
rect 23565 21795 23631 21796
rect 4189 21792 4505 21793
rect 4189 21728 4195 21792
rect 4259 21728 4275 21792
rect 4339 21728 4355 21792
rect 4419 21728 4435 21792
rect 4499 21728 4505 21792
rect 4189 21727 4505 21728
rect 11779 21792 12095 21793
rect 11779 21728 11785 21792
rect 11849 21728 11865 21792
rect 11929 21728 11945 21792
rect 12009 21728 12025 21792
rect 12089 21728 12095 21792
rect 11779 21727 12095 21728
rect 19369 21792 19685 21793
rect 19369 21728 19375 21792
rect 19439 21728 19455 21792
rect 19519 21728 19535 21792
rect 19599 21728 19615 21792
rect 19679 21728 19685 21792
rect 19369 21727 19685 21728
rect 26959 21792 27275 21793
rect 26959 21728 26965 21792
rect 27029 21728 27045 21792
rect 27109 21728 27125 21792
rect 27189 21728 27205 21792
rect 27269 21728 27275 21792
rect 26959 21727 27275 21728
rect 20345 21722 20411 21725
rect 24209 21722 24275 21725
rect 25865 21722 25931 21725
rect 20345 21720 25931 21722
rect 20345 21664 20350 21720
rect 20406 21664 24214 21720
rect 24270 21664 25870 21720
rect 25926 21664 25931 21720
rect 20345 21662 25931 21664
rect 20345 21659 20411 21662
rect 24209 21659 24275 21662
rect 25865 21659 25931 21662
rect 841 21586 907 21589
rect 10961 21586 11027 21589
rect 12249 21588 12315 21589
rect 11462 21586 11468 21588
rect 841 21584 2790 21586
rect 841 21528 846 21584
rect 902 21528 2790 21584
rect 841 21526 2790 21528
rect 841 21523 907 21526
rect 2730 21450 2790 21526
rect 10961 21584 11468 21586
rect 10961 21528 10966 21584
rect 11022 21528 11468 21584
rect 10961 21526 11468 21528
rect 10961 21523 11027 21526
rect 11462 21524 11468 21526
rect 11532 21524 11538 21588
rect 12198 21586 12204 21588
rect 12158 21526 12204 21586
rect 12268 21584 12315 21588
rect 12310 21528 12315 21584
rect 12198 21524 12204 21526
rect 12268 21524 12315 21528
rect 16982 21524 16988 21588
rect 17052 21586 17058 21588
rect 17953 21586 18019 21589
rect 17052 21584 18019 21586
rect 17052 21528 17958 21584
rect 18014 21528 18019 21584
rect 17052 21526 18019 21528
rect 17052 21524 17058 21526
rect 12249 21523 12315 21524
rect 17953 21523 18019 21526
rect 22001 21586 22067 21589
rect 24485 21586 24551 21589
rect 22001 21584 24551 21586
rect 22001 21528 22006 21584
rect 22062 21528 24490 21584
rect 24546 21528 24551 21584
rect 22001 21526 24551 21528
rect 22001 21523 22067 21526
rect 24485 21523 24551 21526
rect 14089 21450 14155 21453
rect 2730 21448 14155 21450
rect 2730 21392 14094 21448
rect 14150 21392 14155 21448
rect 2730 21390 14155 21392
rect 14089 21387 14155 21390
rect 23197 21450 23263 21453
rect 25773 21450 25839 21453
rect 23197 21448 25839 21450
rect 23197 21392 23202 21448
rect 23258 21392 25778 21448
rect 25834 21392 25839 21448
rect 23197 21390 25839 21392
rect 23197 21387 23263 21390
rect 25773 21387 25839 21390
rect 8477 21314 8543 21317
rect 9305 21314 9371 21317
rect 8477 21312 9371 21314
rect 8477 21256 8482 21312
rect 8538 21256 9310 21312
rect 9366 21256 9371 21312
rect 8477 21254 9371 21256
rect 8477 21251 8543 21254
rect 9305 21251 9371 21254
rect 10777 21314 10843 21317
rect 11605 21314 11671 21317
rect 10777 21312 11671 21314
rect 10777 21256 10782 21312
rect 10838 21256 11610 21312
rect 11666 21256 11671 21312
rect 10777 21254 11671 21256
rect 10777 21251 10843 21254
rect 11605 21251 11671 21254
rect 13118 21252 13124 21316
rect 13188 21314 13194 21316
rect 13813 21314 13879 21317
rect 13188 21312 13879 21314
rect 13188 21256 13818 21312
rect 13874 21256 13879 21312
rect 13188 21254 13879 21256
rect 13188 21252 13194 21254
rect 13813 21251 13879 21254
rect 7984 21248 8300 21249
rect 7984 21184 7990 21248
rect 8054 21184 8070 21248
rect 8134 21184 8150 21248
rect 8214 21184 8230 21248
rect 8294 21184 8300 21248
rect 7984 21183 8300 21184
rect 15574 21248 15890 21249
rect 15574 21184 15580 21248
rect 15644 21184 15660 21248
rect 15724 21184 15740 21248
rect 15804 21184 15820 21248
rect 15884 21184 15890 21248
rect 15574 21183 15890 21184
rect 23164 21248 23480 21249
rect 23164 21184 23170 21248
rect 23234 21184 23250 21248
rect 23314 21184 23330 21248
rect 23394 21184 23410 21248
rect 23474 21184 23480 21248
rect 23164 21183 23480 21184
rect 30754 21248 31070 21249
rect 30754 21184 30760 21248
rect 30824 21184 30840 21248
rect 30904 21184 30920 21248
rect 30984 21184 31000 21248
rect 31064 21184 31070 21248
rect 30754 21183 31070 21184
rect 11278 21178 11284 21180
rect 8526 21118 11284 21178
rect 1853 21042 1919 21045
rect 8526 21042 8586 21118
rect 11278 21116 11284 21118
rect 11348 21116 11354 21180
rect 25129 21178 25195 21181
rect 26366 21178 26372 21180
rect 25129 21176 26372 21178
rect 25129 21120 25134 21176
rect 25190 21120 26372 21176
rect 25129 21118 26372 21120
rect 25129 21115 25195 21118
rect 26366 21116 26372 21118
rect 26436 21116 26442 21180
rect 1853 21040 8586 21042
rect 1853 20984 1858 21040
rect 1914 20984 8586 21040
rect 1853 20982 8586 20984
rect 8753 21042 8819 21045
rect 10593 21042 10659 21045
rect 8753 21040 10659 21042
rect 8753 20984 8758 21040
rect 8814 20984 10598 21040
rect 10654 20984 10659 21040
rect 8753 20982 10659 20984
rect 1853 20979 1919 20982
rect 8753 20979 8819 20982
rect 10593 20979 10659 20982
rect 12157 21042 12223 21045
rect 12157 21040 12266 21042
rect 12157 20984 12162 21040
rect 12218 20984 12266 21040
rect 12157 20979 12266 20984
rect 4061 20906 4127 20909
rect 11094 20906 11100 20908
rect 4061 20904 11100 20906
rect 4061 20848 4066 20904
rect 4122 20848 11100 20904
rect 4061 20846 11100 20848
rect 4061 20843 4127 20846
rect 11094 20844 11100 20846
rect 11164 20844 11170 20908
rect 12206 20906 12266 20979
rect 12433 20906 12499 20909
rect 12206 20904 12499 20906
rect 12206 20848 12438 20904
rect 12494 20848 12499 20904
rect 12206 20846 12499 20848
rect 12433 20843 12499 20846
rect 16757 20906 16823 20909
rect 23606 20906 23612 20908
rect 16757 20904 23612 20906
rect 16757 20848 16762 20904
rect 16818 20848 23612 20904
rect 16757 20846 23612 20848
rect 16757 20843 16823 20846
rect 23606 20844 23612 20846
rect 23676 20844 23682 20908
rect 25405 20906 25471 20909
rect 28717 20906 28783 20909
rect 25405 20904 28783 20906
rect 25405 20848 25410 20904
rect 25466 20848 28722 20904
rect 28778 20848 28783 20904
rect 25405 20846 28783 20848
rect 25405 20843 25471 20846
rect 28717 20843 28783 20846
rect 6545 20770 6611 20773
rect 8886 20770 8892 20772
rect 6545 20768 8892 20770
rect 6545 20712 6550 20768
rect 6606 20712 8892 20768
rect 6545 20710 8892 20712
rect 6545 20707 6611 20710
rect 8886 20708 8892 20710
rect 8956 20708 8962 20772
rect 4189 20704 4505 20705
rect 4189 20640 4195 20704
rect 4259 20640 4275 20704
rect 4339 20640 4355 20704
rect 4419 20640 4435 20704
rect 4499 20640 4505 20704
rect 4189 20639 4505 20640
rect 11779 20704 12095 20705
rect 11779 20640 11785 20704
rect 11849 20640 11865 20704
rect 11929 20640 11945 20704
rect 12009 20640 12025 20704
rect 12089 20640 12095 20704
rect 11779 20639 12095 20640
rect 19369 20704 19685 20705
rect 19369 20640 19375 20704
rect 19439 20640 19455 20704
rect 19519 20640 19535 20704
rect 19599 20640 19615 20704
rect 19679 20640 19685 20704
rect 19369 20639 19685 20640
rect 26959 20704 27275 20705
rect 26959 20640 26965 20704
rect 27029 20640 27045 20704
rect 27109 20640 27125 20704
rect 27189 20640 27205 20704
rect 27269 20640 27275 20704
rect 26959 20639 27275 20640
rect 5993 20634 6059 20637
rect 8845 20634 8911 20637
rect 10961 20636 11027 20637
rect 10910 20634 10916 20636
rect 5993 20632 8911 20634
rect 5993 20576 5998 20632
rect 6054 20576 8850 20632
rect 8906 20576 8911 20632
rect 5993 20574 8911 20576
rect 10870 20574 10916 20634
rect 10980 20632 11027 20636
rect 11022 20576 11027 20632
rect 5993 20571 6059 20574
rect 8845 20571 8911 20574
rect 10910 20572 10916 20574
rect 10980 20572 11027 20576
rect 13670 20572 13676 20636
rect 13740 20634 13746 20636
rect 15193 20634 15259 20637
rect 13740 20632 15259 20634
rect 13740 20576 15198 20632
rect 15254 20576 15259 20632
rect 13740 20574 15259 20576
rect 13740 20572 13746 20574
rect 10961 20571 11027 20572
rect 15193 20571 15259 20574
rect 19885 20634 19951 20637
rect 23841 20634 23907 20637
rect 19885 20632 23907 20634
rect 19885 20576 19890 20632
rect 19946 20576 23846 20632
rect 23902 20576 23907 20632
rect 19885 20574 23907 20576
rect 19885 20571 19951 20574
rect 23841 20571 23907 20574
rect 9581 20498 9647 20501
rect 9806 20498 9812 20500
rect 9581 20496 9812 20498
rect 9581 20440 9586 20496
rect 9642 20440 9812 20496
rect 9581 20438 9812 20440
rect 9581 20435 9647 20438
rect 9806 20436 9812 20438
rect 9876 20436 9882 20500
rect 16062 20436 16068 20500
rect 16132 20498 16138 20500
rect 16573 20498 16639 20501
rect 16132 20496 16639 20498
rect 16132 20440 16578 20496
rect 16634 20440 16639 20496
rect 16132 20438 16639 20440
rect 16132 20436 16138 20438
rect 16573 20435 16639 20438
rect 4705 20362 4771 20365
rect 9029 20362 9095 20365
rect 4705 20360 9095 20362
rect 4705 20304 4710 20360
rect 4766 20304 9034 20360
rect 9090 20304 9095 20360
rect 4705 20302 9095 20304
rect 4705 20299 4771 20302
rect 9029 20299 9095 20302
rect 22553 20362 22619 20365
rect 25497 20362 25563 20365
rect 22553 20360 25563 20362
rect 22553 20304 22558 20360
rect 22614 20304 25502 20360
rect 25558 20304 25563 20360
rect 22553 20302 25563 20304
rect 22553 20299 22619 20302
rect 25497 20299 25563 20302
rect 8385 20226 8451 20229
rect 9489 20226 9555 20229
rect 8385 20224 9555 20226
rect 8385 20168 8390 20224
rect 8446 20168 9494 20224
rect 9550 20168 9555 20224
rect 8385 20166 9555 20168
rect 8385 20163 8451 20166
rect 9489 20163 9555 20166
rect 7984 20160 8300 20161
rect 7984 20096 7990 20160
rect 8054 20096 8070 20160
rect 8134 20096 8150 20160
rect 8214 20096 8230 20160
rect 8294 20096 8300 20160
rect 7984 20095 8300 20096
rect 15574 20160 15890 20161
rect 15574 20096 15580 20160
rect 15644 20096 15660 20160
rect 15724 20096 15740 20160
rect 15804 20096 15820 20160
rect 15884 20096 15890 20160
rect 15574 20095 15890 20096
rect 23164 20160 23480 20161
rect 23164 20096 23170 20160
rect 23234 20096 23250 20160
rect 23314 20096 23330 20160
rect 23394 20096 23410 20160
rect 23474 20096 23480 20160
rect 23164 20095 23480 20096
rect 30754 20160 31070 20161
rect 30754 20096 30760 20160
rect 30824 20096 30840 20160
rect 30904 20096 30920 20160
rect 30984 20096 31000 20160
rect 31064 20096 31070 20160
rect 30754 20095 31070 20096
rect 5809 19954 5875 19957
rect 6913 19954 6979 19957
rect 5809 19952 6979 19954
rect 5809 19896 5814 19952
rect 5870 19896 6918 19952
rect 6974 19896 6979 19952
rect 5809 19894 6979 19896
rect 5809 19891 5875 19894
rect 6913 19891 6979 19894
rect 23105 19954 23171 19957
rect 23933 19954 23999 19957
rect 23105 19952 23999 19954
rect 23105 19896 23110 19952
rect 23166 19896 23938 19952
rect 23994 19896 23999 19952
rect 23105 19894 23999 19896
rect 23105 19891 23171 19894
rect 23933 19891 23999 19894
rect 657 19818 723 19821
rect 7281 19818 7347 19821
rect 14549 19818 14615 19821
rect 657 19816 7114 19818
rect 657 19760 662 19816
rect 718 19760 7114 19816
rect 657 19758 7114 19760
rect 657 19755 723 19758
rect 7054 19682 7114 19758
rect 7281 19816 14615 19818
rect 7281 19760 7286 19816
rect 7342 19760 14554 19816
rect 14610 19760 14615 19816
rect 7281 19758 14615 19760
rect 7281 19755 7347 19758
rect 14549 19755 14615 19758
rect 8477 19682 8543 19685
rect 7054 19680 8543 19682
rect 7054 19624 8482 19680
rect 8538 19624 8543 19680
rect 7054 19622 8543 19624
rect 8477 19619 8543 19622
rect 22001 19682 22067 19685
rect 22461 19682 22527 19685
rect 22001 19680 22527 19682
rect 22001 19624 22006 19680
rect 22062 19624 22466 19680
rect 22522 19624 22527 19680
rect 22001 19622 22527 19624
rect 22001 19619 22067 19622
rect 22461 19619 22527 19622
rect 4189 19616 4505 19617
rect 4189 19552 4195 19616
rect 4259 19552 4275 19616
rect 4339 19552 4355 19616
rect 4419 19552 4435 19616
rect 4499 19552 4505 19616
rect 4189 19551 4505 19552
rect 11779 19616 12095 19617
rect 11779 19552 11785 19616
rect 11849 19552 11865 19616
rect 11929 19552 11945 19616
rect 12009 19552 12025 19616
rect 12089 19552 12095 19616
rect 11779 19551 12095 19552
rect 19369 19616 19685 19617
rect 19369 19552 19375 19616
rect 19439 19552 19455 19616
rect 19519 19552 19535 19616
rect 19599 19552 19615 19616
rect 19679 19552 19685 19616
rect 19369 19551 19685 19552
rect 26959 19616 27275 19617
rect 26959 19552 26965 19616
rect 27029 19552 27045 19616
rect 27109 19552 27125 19616
rect 27189 19552 27205 19616
rect 27269 19552 27275 19616
rect 26959 19551 27275 19552
rect 6729 19546 6795 19549
rect 9029 19546 9095 19549
rect 6729 19544 9095 19546
rect 6729 19488 6734 19544
rect 6790 19488 9034 19544
rect 9090 19488 9095 19544
rect 6729 19486 9095 19488
rect 6729 19483 6795 19486
rect 9029 19483 9095 19486
rect 1669 19410 1735 19413
rect 5441 19410 5507 19413
rect 1669 19408 5507 19410
rect 1669 19352 1674 19408
rect 1730 19352 5446 19408
rect 5502 19352 5507 19408
rect 1669 19350 5507 19352
rect 1669 19347 1735 19350
rect 5441 19347 5507 19350
rect 6545 19410 6611 19413
rect 6678 19410 6684 19412
rect 6545 19408 6684 19410
rect 6545 19352 6550 19408
rect 6606 19352 6684 19408
rect 6545 19350 6684 19352
rect 6545 19347 6611 19350
rect 6678 19348 6684 19350
rect 6748 19348 6754 19412
rect 8201 19410 8267 19413
rect 10685 19410 10751 19413
rect 14273 19410 14339 19413
rect 29177 19410 29243 19413
rect 8201 19408 9506 19410
rect 8201 19352 8206 19408
rect 8262 19352 9506 19408
rect 8201 19350 9506 19352
rect 8201 19347 8267 19350
rect 4429 19274 4495 19277
rect 9213 19274 9279 19277
rect 4429 19272 9279 19274
rect 4429 19216 4434 19272
rect 4490 19216 9218 19272
rect 9274 19216 9279 19272
rect 4429 19214 9279 19216
rect 9446 19274 9506 19350
rect 10685 19408 14339 19410
rect 10685 19352 10690 19408
rect 10746 19352 14278 19408
rect 14334 19352 14339 19408
rect 10685 19350 14339 19352
rect 10685 19347 10751 19350
rect 14273 19347 14339 19350
rect 23430 19408 29243 19410
rect 23430 19352 29182 19408
rect 29238 19352 29243 19408
rect 23430 19350 29243 19352
rect 10685 19274 10751 19277
rect 9446 19272 10751 19274
rect 9446 19216 10690 19272
rect 10746 19216 10751 19272
rect 9446 19214 10751 19216
rect 4429 19211 4495 19214
rect 9213 19211 9279 19214
rect 10685 19211 10751 19214
rect 15326 19212 15332 19276
rect 15396 19274 15402 19276
rect 16113 19274 16179 19277
rect 16481 19276 16547 19277
rect 15396 19272 16179 19274
rect 15396 19216 16118 19272
rect 16174 19216 16179 19272
rect 15396 19214 16179 19216
rect 15396 19212 15402 19214
rect 16113 19211 16179 19214
rect 16430 19212 16436 19276
rect 16500 19274 16547 19276
rect 23430 19274 23490 19350
rect 29177 19347 29243 19350
rect 16500 19272 16592 19274
rect 16542 19216 16592 19272
rect 16500 19214 16592 19216
rect 22878 19214 23490 19274
rect 24945 19274 25011 19277
rect 26601 19274 26667 19277
rect 24945 19272 26667 19274
rect 24945 19216 24950 19272
rect 25006 19216 26606 19272
rect 26662 19216 26667 19272
rect 24945 19214 26667 19216
rect 16500 19212 16547 19214
rect 16481 19211 16547 19212
rect 22878 19141 22938 19214
rect 24945 19211 25011 19214
rect 26601 19211 26667 19214
rect 26969 19274 27035 19277
rect 27613 19274 27679 19277
rect 26969 19272 27679 19274
rect 26969 19216 26974 19272
rect 27030 19216 27618 19272
rect 27674 19216 27679 19272
rect 26969 19214 27679 19216
rect 26969 19211 27035 19214
rect 27613 19211 27679 19214
rect 4613 19138 4679 19141
rect 5993 19138 6059 19141
rect 4613 19136 6059 19138
rect 4613 19080 4618 19136
rect 4674 19080 5998 19136
rect 6054 19080 6059 19136
rect 4613 19078 6059 19080
rect 22878 19136 22987 19141
rect 22878 19080 22926 19136
rect 22982 19080 22987 19136
rect 22878 19078 22987 19080
rect 4613 19075 4679 19078
rect 5993 19075 6059 19078
rect 22921 19075 22987 19078
rect 24025 19138 24091 19141
rect 26233 19138 26299 19141
rect 24025 19136 26299 19138
rect 24025 19080 24030 19136
rect 24086 19080 26238 19136
rect 26294 19080 26299 19136
rect 24025 19078 26299 19080
rect 24025 19075 24091 19078
rect 26233 19075 26299 19078
rect 7984 19072 8300 19073
rect 7984 19008 7990 19072
rect 8054 19008 8070 19072
rect 8134 19008 8150 19072
rect 8214 19008 8230 19072
rect 8294 19008 8300 19072
rect 7984 19007 8300 19008
rect 15574 19072 15890 19073
rect 15574 19008 15580 19072
rect 15644 19008 15660 19072
rect 15724 19008 15740 19072
rect 15804 19008 15820 19072
rect 15884 19008 15890 19072
rect 15574 19007 15890 19008
rect 23164 19072 23480 19073
rect 23164 19008 23170 19072
rect 23234 19008 23250 19072
rect 23314 19008 23330 19072
rect 23394 19008 23410 19072
rect 23474 19008 23480 19072
rect 23164 19007 23480 19008
rect 30754 19072 31070 19073
rect 30754 19008 30760 19072
rect 30824 19008 30840 19072
rect 30904 19008 30920 19072
rect 30984 19008 31000 19072
rect 31064 19008 31070 19072
rect 30754 19007 31070 19008
rect 3734 18940 3740 19004
rect 3804 19002 3810 19004
rect 4337 19002 4403 19005
rect 11421 19002 11487 19005
rect 3804 19000 4403 19002
rect 3804 18944 4342 19000
rect 4398 18944 4403 19000
rect 3804 18942 4403 18944
rect 3804 18940 3810 18942
rect 4337 18939 4403 18942
rect 4662 18942 7252 19002
rect 4662 18866 4722 18942
rect 4294 18806 4722 18866
rect 4797 18866 4863 18869
rect 6637 18866 6703 18869
rect 4797 18864 6703 18866
rect 4797 18808 4802 18864
rect 4858 18808 6642 18864
rect 6698 18808 6703 18864
rect 4797 18806 6703 18808
rect 7192 18866 7252 18942
rect 11421 19000 13692 19002
rect 11421 18944 11426 19000
rect 11482 18944 13692 19000
rect 11421 18942 13692 18944
rect 11421 18939 11487 18942
rect 10317 18866 10383 18869
rect 11237 18866 11303 18869
rect 13445 18866 13511 18869
rect 7192 18864 13511 18866
rect 7192 18808 10322 18864
rect 10378 18808 11242 18864
rect 11298 18808 13450 18864
rect 13506 18808 13511 18864
rect 7192 18806 13511 18808
rect 13632 18866 13692 18942
rect 18229 18866 18295 18869
rect 13632 18864 18295 18866
rect 13632 18808 18234 18864
rect 18290 18808 18295 18864
rect 13632 18806 18295 18808
rect 4294 18733 4354 18806
rect 4797 18803 4863 18806
rect 6637 18803 6703 18806
rect 10317 18803 10383 18806
rect 11237 18803 11303 18806
rect 13445 18803 13511 18806
rect 18229 18803 18295 18806
rect 18965 18866 19031 18869
rect 23473 18866 23539 18869
rect 24710 18866 24716 18868
rect 18965 18864 22110 18866
rect 18965 18808 18970 18864
rect 19026 18808 22110 18864
rect 18965 18806 22110 18808
rect 18965 18803 19031 18806
rect 4245 18728 4354 18733
rect 4245 18672 4250 18728
rect 4306 18672 4354 18728
rect 4245 18670 4354 18672
rect 4429 18730 4495 18733
rect 5809 18730 5875 18733
rect 4429 18728 5875 18730
rect 4429 18672 4434 18728
rect 4490 18672 5814 18728
rect 5870 18672 5875 18728
rect 4429 18670 5875 18672
rect 4245 18667 4311 18670
rect 4429 18667 4495 18670
rect 5809 18667 5875 18670
rect 6085 18730 6151 18733
rect 10358 18730 10364 18732
rect 6085 18728 10364 18730
rect 6085 18672 6090 18728
rect 6146 18672 10364 18728
rect 6085 18670 10364 18672
rect 6085 18667 6151 18670
rect 10358 18668 10364 18670
rect 10428 18730 10434 18732
rect 17953 18730 18019 18733
rect 10428 18728 18019 18730
rect 10428 18672 17958 18728
rect 18014 18672 18019 18728
rect 10428 18670 18019 18672
rect 22050 18730 22110 18806
rect 23473 18864 24716 18866
rect 23473 18808 23478 18864
rect 23534 18808 24716 18864
rect 23473 18806 24716 18808
rect 23473 18803 23539 18806
rect 24710 18804 24716 18806
rect 24780 18804 24786 18868
rect 25262 18730 25268 18732
rect 22050 18670 25268 18730
rect 10428 18668 10434 18670
rect 17953 18667 18019 18670
rect 25262 18668 25268 18670
rect 25332 18668 25338 18732
rect 6913 18594 6979 18597
rect 4662 18592 6979 18594
rect 4662 18536 6918 18592
rect 6974 18536 6979 18592
rect 4662 18534 6979 18536
rect 4189 18528 4505 18529
rect 4189 18464 4195 18528
rect 4259 18464 4275 18528
rect 4339 18464 4355 18528
rect 4419 18464 4435 18528
rect 4499 18464 4505 18528
rect 4189 18463 4505 18464
rect 3509 18458 3575 18461
rect 3374 18456 3575 18458
rect 3374 18400 3514 18456
rect 3570 18400 3575 18456
rect 3374 18398 3575 18400
rect 3374 18186 3434 18398
rect 3509 18395 3575 18398
rect 3509 18322 3575 18325
rect 3785 18322 3851 18325
rect 4662 18322 4722 18534
rect 6913 18531 6979 18534
rect 7741 18596 7807 18597
rect 7741 18592 7788 18596
rect 7852 18594 7858 18596
rect 8201 18594 8267 18597
rect 9581 18594 9647 18597
rect 7741 18536 7746 18592
rect 7741 18532 7788 18536
rect 7852 18534 7898 18594
rect 8201 18592 9647 18594
rect 8201 18536 8206 18592
rect 8262 18536 9586 18592
rect 9642 18536 9647 18592
rect 8201 18534 9647 18536
rect 7852 18532 7858 18534
rect 7741 18531 7807 18532
rect 8201 18531 8267 18534
rect 9581 18531 9647 18534
rect 23841 18594 23907 18597
rect 26182 18594 26188 18596
rect 23841 18592 26188 18594
rect 23841 18536 23846 18592
rect 23902 18536 26188 18592
rect 23841 18534 26188 18536
rect 23841 18531 23907 18534
rect 26182 18532 26188 18534
rect 26252 18532 26258 18596
rect 11779 18528 12095 18529
rect 11779 18464 11785 18528
rect 11849 18464 11865 18528
rect 11929 18464 11945 18528
rect 12009 18464 12025 18528
rect 12089 18464 12095 18528
rect 11779 18463 12095 18464
rect 19369 18528 19685 18529
rect 19369 18464 19375 18528
rect 19439 18464 19455 18528
rect 19519 18464 19535 18528
rect 19599 18464 19615 18528
rect 19679 18464 19685 18528
rect 19369 18463 19685 18464
rect 26959 18528 27275 18529
rect 26959 18464 26965 18528
rect 27029 18464 27045 18528
rect 27109 18464 27125 18528
rect 27189 18464 27205 18528
rect 27269 18464 27275 18528
rect 26959 18463 27275 18464
rect 5533 18458 5599 18461
rect 9673 18458 9739 18461
rect 5533 18456 9739 18458
rect 5533 18400 5538 18456
rect 5594 18400 9678 18456
rect 9734 18400 9739 18456
rect 5533 18398 9739 18400
rect 5533 18395 5599 18398
rect 9673 18395 9739 18398
rect 22185 18458 22251 18461
rect 25814 18458 25820 18460
rect 22185 18456 25820 18458
rect 22185 18400 22190 18456
rect 22246 18400 25820 18456
rect 22185 18398 25820 18400
rect 22185 18395 22251 18398
rect 25814 18396 25820 18398
rect 25884 18396 25890 18460
rect 3509 18320 4722 18322
rect 3509 18264 3514 18320
rect 3570 18264 3790 18320
rect 3846 18264 4722 18320
rect 3509 18262 4722 18264
rect 5533 18322 5599 18325
rect 6913 18322 6979 18325
rect 5533 18320 6979 18322
rect 5533 18264 5538 18320
rect 5594 18264 6918 18320
rect 6974 18264 6979 18320
rect 5533 18262 6979 18264
rect 3509 18259 3575 18262
rect 3785 18259 3851 18262
rect 5533 18259 5599 18262
rect 6913 18259 6979 18262
rect 7046 18260 7052 18324
rect 7116 18322 7122 18324
rect 7373 18322 7439 18325
rect 7116 18320 7439 18322
rect 7116 18264 7378 18320
rect 7434 18264 7439 18320
rect 7116 18262 7439 18264
rect 7116 18260 7122 18262
rect 7373 18259 7439 18262
rect 7557 18322 7623 18325
rect 10726 18322 10732 18324
rect 7557 18320 10732 18322
rect 7557 18264 7562 18320
rect 7618 18264 10732 18320
rect 7557 18262 10732 18264
rect 7557 18259 7623 18262
rect 10726 18260 10732 18262
rect 10796 18322 10802 18324
rect 13077 18322 13143 18325
rect 10796 18320 13143 18322
rect 10796 18264 13082 18320
rect 13138 18264 13143 18320
rect 10796 18262 13143 18264
rect 10796 18260 10802 18262
rect 13077 18259 13143 18262
rect 21173 18322 21239 18325
rect 26601 18322 26667 18325
rect 21173 18320 26667 18322
rect 21173 18264 21178 18320
rect 21234 18264 26606 18320
rect 26662 18264 26667 18320
rect 21173 18262 26667 18264
rect 21173 18259 21239 18262
rect 26601 18259 26667 18262
rect 30046 18260 30052 18324
rect 30116 18322 30122 18324
rect 30189 18322 30255 18325
rect 30116 18320 30255 18322
rect 30116 18264 30194 18320
rect 30250 18264 30255 18320
rect 30116 18262 30255 18264
rect 30116 18260 30122 18262
rect 30189 18259 30255 18262
rect 4521 18186 4587 18189
rect 3374 18184 4587 18186
rect 3374 18128 4526 18184
rect 4582 18128 4587 18184
rect 3374 18126 4587 18128
rect 4521 18123 4587 18126
rect 4654 18124 4660 18188
rect 4724 18186 4730 18188
rect 4889 18186 4955 18189
rect 4724 18184 4955 18186
rect 4724 18128 4894 18184
rect 4950 18128 4955 18184
rect 4724 18126 4955 18128
rect 4724 18124 4730 18126
rect 4889 18123 4955 18126
rect 5257 18186 5323 18189
rect 9213 18186 9279 18189
rect 5257 18184 9279 18186
rect 5257 18128 5262 18184
rect 5318 18128 9218 18184
rect 9274 18128 9279 18184
rect 5257 18126 9279 18128
rect 5257 18123 5323 18126
rect 9213 18123 9279 18126
rect 13486 18124 13492 18188
rect 13556 18186 13562 18188
rect 13629 18186 13695 18189
rect 30189 18186 30255 18189
rect 13556 18184 30255 18186
rect 13556 18128 13634 18184
rect 13690 18128 30194 18184
rect 30250 18128 30255 18184
rect 13556 18126 30255 18128
rect 13556 18124 13562 18126
rect 13629 18123 13695 18126
rect 30189 18123 30255 18126
rect 3325 18050 3391 18053
rect 3918 18050 3924 18052
rect 3325 18048 3924 18050
rect 3325 17992 3330 18048
rect 3386 17992 3924 18048
rect 3325 17990 3924 17992
rect 3325 17987 3391 17990
rect 3918 17988 3924 17990
rect 3988 17988 3994 18052
rect 4838 17988 4844 18052
rect 4908 18050 4914 18052
rect 5257 18050 5323 18053
rect 5993 18052 6059 18053
rect 5390 18050 5396 18052
rect 4908 17990 5090 18050
rect 4908 17988 4914 17990
rect 1117 17914 1183 17917
rect 3141 17914 3207 17917
rect 1117 17912 3207 17914
rect 1117 17856 1122 17912
rect 1178 17856 3146 17912
rect 3202 17856 3207 17912
rect 1117 17854 3207 17856
rect 5030 17914 5090 17990
rect 5257 18048 5396 18050
rect 5257 17992 5262 18048
rect 5318 17992 5396 18048
rect 5257 17990 5396 17992
rect 5257 17987 5323 17990
rect 5390 17988 5396 17990
rect 5460 17988 5466 18052
rect 5942 18050 5948 18052
rect 5902 17990 5948 18050
rect 6012 18048 6059 18052
rect 6054 17992 6059 18048
rect 5942 17988 5948 17990
rect 6012 17988 6059 17992
rect 5993 17987 6059 17988
rect 6821 18050 6887 18053
rect 7782 18050 7788 18052
rect 6821 18048 7788 18050
rect 6821 17992 6826 18048
rect 6882 17992 7788 18048
rect 6821 17990 7788 17992
rect 6821 17987 6887 17990
rect 7782 17988 7788 17990
rect 7852 17988 7858 18052
rect 10685 18050 10751 18053
rect 12801 18050 12867 18053
rect 10685 18048 12867 18050
rect 10685 17992 10690 18048
rect 10746 17992 12806 18048
rect 12862 17992 12867 18048
rect 10685 17990 12867 17992
rect 10685 17987 10751 17990
rect 12801 17987 12867 17990
rect 16389 18050 16455 18053
rect 23013 18050 23079 18053
rect 16389 18048 23079 18050
rect 16389 17992 16394 18048
rect 16450 17992 23018 18048
rect 23074 17992 23079 18048
rect 16389 17990 23079 17992
rect 16389 17987 16455 17990
rect 23013 17987 23079 17990
rect 25497 18050 25563 18053
rect 27705 18050 27771 18053
rect 25497 18048 27771 18050
rect 25497 17992 25502 18048
rect 25558 17992 27710 18048
rect 27766 17992 27771 18048
rect 25497 17990 27771 17992
rect 25497 17987 25563 17990
rect 27705 17987 27771 17990
rect 7984 17984 8300 17985
rect 7984 17920 7990 17984
rect 8054 17920 8070 17984
rect 8134 17920 8150 17984
rect 8214 17920 8230 17984
rect 8294 17920 8300 17984
rect 7984 17919 8300 17920
rect 15574 17984 15890 17985
rect 15574 17920 15580 17984
rect 15644 17920 15660 17984
rect 15724 17920 15740 17984
rect 15804 17920 15820 17984
rect 15884 17920 15890 17984
rect 15574 17919 15890 17920
rect 23164 17984 23480 17985
rect 23164 17920 23170 17984
rect 23234 17920 23250 17984
rect 23314 17920 23330 17984
rect 23394 17920 23410 17984
rect 23474 17920 23480 17984
rect 23164 17919 23480 17920
rect 30754 17984 31070 17985
rect 30754 17920 30760 17984
rect 30824 17920 30840 17984
rect 30904 17920 30920 17984
rect 30984 17920 31000 17984
rect 31064 17920 31070 17984
rect 30754 17919 31070 17920
rect 5165 17914 5231 17917
rect 7465 17914 7531 17917
rect 11697 17916 11763 17917
rect 11646 17914 11652 17916
rect 5030 17912 5231 17914
rect 5030 17856 5170 17912
rect 5226 17856 5231 17912
rect 5030 17854 5231 17856
rect 1117 17851 1183 17854
rect 3141 17851 3207 17854
rect 5165 17851 5231 17854
rect 5398 17912 7531 17914
rect 5398 17856 7470 17912
rect 7526 17856 7531 17912
rect 5398 17854 7531 17856
rect 11606 17854 11652 17914
rect 11716 17912 11763 17916
rect 11758 17856 11763 17912
rect 1025 17778 1091 17781
rect 5398 17778 5458 17854
rect 7465 17851 7531 17854
rect 11646 17852 11652 17854
rect 11716 17852 11763 17856
rect 11697 17851 11763 17852
rect 24485 17914 24551 17917
rect 27061 17914 27127 17917
rect 24485 17912 27127 17914
rect 24485 17856 24490 17912
rect 24546 17856 27066 17912
rect 27122 17856 27127 17912
rect 24485 17854 27127 17856
rect 24485 17851 24551 17854
rect 27061 17851 27127 17854
rect 1025 17776 5458 17778
rect 1025 17720 1030 17776
rect 1086 17720 5458 17776
rect 1025 17718 5458 17720
rect 5901 17778 5967 17781
rect 8845 17778 8911 17781
rect 11053 17778 11119 17781
rect 13353 17778 13419 17781
rect 5901 17776 8724 17778
rect 5901 17720 5906 17776
rect 5962 17720 8724 17776
rect 5901 17718 8724 17720
rect 1025 17715 1091 17718
rect 5901 17715 5967 17718
rect 4521 17642 4587 17645
rect 4521 17640 8586 17642
rect 4521 17584 4526 17640
rect 4582 17584 8586 17640
rect 4521 17582 8586 17584
rect 4521 17579 4587 17582
rect 8526 17508 8586 17582
rect 8518 17444 8524 17508
rect 8588 17444 8594 17508
rect 8664 17506 8724 17718
rect 8845 17776 13419 17778
rect 8845 17720 8850 17776
rect 8906 17720 11058 17776
rect 11114 17720 13358 17776
rect 13414 17720 13419 17776
rect 8845 17718 13419 17720
rect 8845 17715 8911 17718
rect 11053 17715 11119 17718
rect 13353 17715 13419 17718
rect 19977 17778 20043 17781
rect 21265 17778 21331 17781
rect 19977 17776 21331 17778
rect 19977 17720 19982 17776
rect 20038 17720 21270 17776
rect 21326 17720 21331 17776
rect 19977 17718 21331 17720
rect 19977 17715 20043 17718
rect 21265 17715 21331 17718
rect 23473 17778 23539 17781
rect 23606 17778 23612 17780
rect 23473 17776 23612 17778
rect 23473 17720 23478 17776
rect 23534 17720 23612 17776
rect 23473 17718 23612 17720
rect 23473 17715 23539 17718
rect 23606 17716 23612 17718
rect 23676 17716 23682 17780
rect 9213 17642 9279 17645
rect 30465 17642 30531 17645
rect 9213 17640 30531 17642
rect 9213 17584 9218 17640
rect 9274 17584 30470 17640
rect 30526 17584 30531 17640
rect 9213 17582 30531 17584
rect 9213 17579 9279 17582
rect 30465 17579 30531 17582
rect 9673 17506 9739 17509
rect 8664 17504 9739 17506
rect 8664 17448 9678 17504
rect 9734 17448 9739 17504
rect 8664 17446 9739 17448
rect 9673 17443 9739 17446
rect 23289 17506 23355 17509
rect 25865 17506 25931 17509
rect 23289 17504 25931 17506
rect 23289 17448 23294 17504
rect 23350 17448 25870 17504
rect 25926 17448 25931 17504
rect 23289 17446 25931 17448
rect 23289 17443 23355 17446
rect 25865 17443 25931 17446
rect 4189 17440 4505 17441
rect 4189 17376 4195 17440
rect 4259 17376 4275 17440
rect 4339 17376 4355 17440
rect 4419 17376 4435 17440
rect 4499 17376 4505 17440
rect 4189 17375 4505 17376
rect 11779 17440 12095 17441
rect 11779 17376 11785 17440
rect 11849 17376 11865 17440
rect 11929 17376 11945 17440
rect 12009 17376 12025 17440
rect 12089 17376 12095 17440
rect 11779 17375 12095 17376
rect 19369 17440 19685 17441
rect 19369 17376 19375 17440
rect 19439 17376 19455 17440
rect 19519 17376 19535 17440
rect 19599 17376 19615 17440
rect 19679 17376 19685 17440
rect 19369 17375 19685 17376
rect 26959 17440 27275 17441
rect 26959 17376 26965 17440
rect 27029 17376 27045 17440
rect 27109 17376 27125 17440
rect 27189 17376 27205 17440
rect 27269 17376 27275 17440
rect 26959 17375 27275 17376
rect 10542 17370 10548 17372
rect 5214 17310 10548 17370
rect 5214 17234 5274 17310
rect 10542 17308 10548 17310
rect 10612 17308 10618 17372
rect 2730 17174 5274 17234
rect 5441 17234 5507 17237
rect 11462 17234 11468 17236
rect 5441 17232 11468 17234
rect 5441 17176 5446 17232
rect 5502 17176 11468 17232
rect 5441 17174 11468 17176
rect 2037 17098 2103 17101
rect 2730 17098 2790 17174
rect 5441 17171 5507 17174
rect 11462 17172 11468 17174
rect 11532 17172 11538 17236
rect 13629 17234 13695 17237
rect 23381 17234 23447 17237
rect 13629 17232 23447 17234
rect 13629 17176 13634 17232
rect 13690 17176 23386 17232
rect 23442 17176 23447 17232
rect 13629 17174 23447 17176
rect 13629 17171 13695 17174
rect 23381 17171 23447 17174
rect 24117 17234 24183 17237
rect 26601 17234 26667 17237
rect 31385 17234 31451 17237
rect 24117 17232 31451 17234
rect 24117 17176 24122 17232
rect 24178 17176 26606 17232
rect 26662 17176 31390 17232
rect 31446 17176 31451 17232
rect 24117 17174 31451 17176
rect 24117 17171 24183 17174
rect 26601 17171 26667 17174
rect 31385 17171 31451 17174
rect 8845 17098 8911 17101
rect 2037 17096 2790 17098
rect 2037 17040 2042 17096
rect 2098 17040 2790 17096
rect 2037 17038 2790 17040
rect 7790 17096 8911 17098
rect 7790 17040 8850 17096
rect 8906 17040 8911 17096
rect 7790 17038 8911 17040
rect 2037 17035 2103 17038
rect 7790 16962 7850 17038
rect 8845 17035 8911 17038
rect 9765 17098 9831 17101
rect 12249 17098 12315 17101
rect 9765 17096 12315 17098
rect 9765 17040 9770 17096
rect 9826 17040 12254 17096
rect 12310 17040 12315 17096
rect 9765 17038 12315 17040
rect 9765 17035 9831 17038
rect 12249 17035 12315 17038
rect 22921 17098 22987 17101
rect 26693 17098 26759 17101
rect 22921 17096 26759 17098
rect 22921 17040 22926 17096
rect 22982 17040 26698 17096
rect 26754 17040 26759 17096
rect 22921 17038 26759 17040
rect 22921 17035 22987 17038
rect 26693 17035 26759 17038
rect 2730 16902 7850 16962
rect 11053 16962 11119 16965
rect 13997 16962 14063 16965
rect 11053 16960 14063 16962
rect 11053 16904 11058 16960
rect 11114 16904 14002 16960
rect 14058 16904 14063 16960
rect 11053 16902 14063 16904
rect 2405 16690 2471 16693
rect 2730 16690 2790 16902
rect 11053 16899 11119 16902
rect 13997 16899 14063 16902
rect 19517 16962 19583 16965
rect 22093 16962 22159 16965
rect 19517 16960 22159 16962
rect 19517 16904 19522 16960
rect 19578 16904 22098 16960
rect 22154 16904 22159 16960
rect 19517 16902 22159 16904
rect 19517 16899 19583 16902
rect 22093 16899 22159 16902
rect 7984 16896 8300 16897
rect 7984 16832 7990 16896
rect 8054 16832 8070 16896
rect 8134 16832 8150 16896
rect 8214 16832 8230 16896
rect 8294 16832 8300 16896
rect 7984 16831 8300 16832
rect 15574 16896 15890 16897
rect 15574 16832 15580 16896
rect 15644 16832 15660 16896
rect 15724 16832 15740 16896
rect 15804 16832 15820 16896
rect 15884 16832 15890 16896
rect 15574 16831 15890 16832
rect 23164 16896 23480 16897
rect 23164 16832 23170 16896
rect 23234 16832 23250 16896
rect 23314 16832 23330 16896
rect 23394 16832 23410 16896
rect 23474 16832 23480 16896
rect 23164 16831 23480 16832
rect 30754 16896 31070 16897
rect 30754 16832 30760 16896
rect 30824 16832 30840 16896
rect 30904 16832 30920 16896
rect 30984 16832 31000 16896
rect 31064 16832 31070 16896
rect 30754 16831 31070 16832
rect 8477 16826 8543 16829
rect 9489 16826 9555 16829
rect 8477 16824 9555 16826
rect 8477 16768 8482 16824
rect 8538 16768 9494 16824
rect 9550 16768 9555 16824
rect 8477 16766 9555 16768
rect 8477 16763 8543 16766
rect 9489 16763 9555 16766
rect 10777 16826 10843 16829
rect 12801 16826 12867 16829
rect 27429 16826 27495 16829
rect 10777 16824 12867 16826
rect 10777 16768 10782 16824
rect 10838 16768 12806 16824
rect 12862 16768 12867 16824
rect 10777 16766 12867 16768
rect 10777 16763 10843 16766
rect 12801 16763 12867 16766
rect 23614 16824 27495 16826
rect 23614 16768 27434 16824
rect 27490 16768 27495 16824
rect 23614 16766 27495 16768
rect 2405 16688 2790 16690
rect 2405 16632 2410 16688
rect 2466 16632 2790 16688
rect 2405 16630 2790 16632
rect 3969 16690 4035 16693
rect 9673 16690 9739 16693
rect 3969 16688 9739 16690
rect 3969 16632 3974 16688
rect 4030 16632 9678 16688
rect 9734 16632 9739 16688
rect 3969 16630 9739 16632
rect 2405 16627 2471 16630
rect 3969 16627 4035 16630
rect 9673 16627 9739 16630
rect 15009 16690 15075 16693
rect 21541 16690 21607 16693
rect 15009 16688 21607 16690
rect 15009 16632 15014 16688
rect 15070 16632 21546 16688
rect 21602 16632 21607 16688
rect 15009 16630 21607 16632
rect 15009 16627 15075 16630
rect 21541 16627 21607 16630
rect 23473 16690 23539 16693
rect 23614 16690 23674 16766
rect 27429 16763 27495 16766
rect 23473 16688 23674 16690
rect 23473 16632 23478 16688
rect 23534 16632 23674 16688
rect 23473 16630 23674 16632
rect 23841 16690 23907 16693
rect 26601 16690 26667 16693
rect 23841 16688 26667 16690
rect 23841 16632 23846 16688
rect 23902 16632 26606 16688
rect 26662 16632 26667 16688
rect 23841 16630 26667 16632
rect 23473 16627 23539 16630
rect 23841 16627 23907 16630
rect 26601 16627 26667 16630
rect 8385 16554 8451 16557
rect 10501 16554 10567 16557
rect 8385 16552 10567 16554
rect 8385 16496 8390 16552
rect 8446 16496 10506 16552
rect 10562 16496 10567 16552
rect 8385 16494 10567 16496
rect 8385 16491 8451 16494
rect 10501 16491 10567 16494
rect 11145 16554 11211 16557
rect 13629 16554 13695 16557
rect 11145 16552 13695 16554
rect 11145 16496 11150 16552
rect 11206 16496 13634 16552
rect 13690 16496 13695 16552
rect 11145 16494 13695 16496
rect 11145 16491 11211 16494
rect 13629 16491 13695 16494
rect 16849 16554 16915 16557
rect 28625 16554 28691 16557
rect 16849 16552 28691 16554
rect 16849 16496 16854 16552
rect 16910 16496 28630 16552
rect 28686 16496 28691 16552
rect 16849 16494 28691 16496
rect 16849 16491 16915 16494
rect 28625 16491 28691 16494
rect 5717 16418 5783 16421
rect 9213 16418 9279 16421
rect 9489 16418 9555 16421
rect 5717 16416 9555 16418
rect 5717 16360 5722 16416
rect 5778 16360 9218 16416
rect 9274 16360 9494 16416
rect 9550 16360 9555 16416
rect 5717 16358 9555 16360
rect 5717 16355 5783 16358
rect 9213 16355 9279 16358
rect 9489 16355 9555 16358
rect 12157 16418 12223 16421
rect 13169 16418 13235 16421
rect 18229 16418 18295 16421
rect 12157 16416 18295 16418
rect 12157 16360 12162 16416
rect 12218 16360 13174 16416
rect 13230 16360 18234 16416
rect 18290 16360 18295 16416
rect 12157 16358 18295 16360
rect 12157 16355 12223 16358
rect 13169 16355 13235 16358
rect 18229 16355 18295 16358
rect 20529 16418 20595 16421
rect 23933 16418 23999 16421
rect 20529 16416 23999 16418
rect 20529 16360 20534 16416
rect 20590 16360 23938 16416
rect 23994 16360 23999 16416
rect 20529 16358 23999 16360
rect 20529 16355 20595 16358
rect 23933 16355 23999 16358
rect 4189 16352 4505 16353
rect 4189 16288 4195 16352
rect 4259 16288 4275 16352
rect 4339 16288 4355 16352
rect 4419 16288 4435 16352
rect 4499 16288 4505 16352
rect 4189 16287 4505 16288
rect 11779 16352 12095 16353
rect 11779 16288 11785 16352
rect 11849 16288 11865 16352
rect 11929 16288 11945 16352
rect 12009 16288 12025 16352
rect 12089 16288 12095 16352
rect 11779 16287 12095 16288
rect 19369 16352 19685 16353
rect 19369 16288 19375 16352
rect 19439 16288 19455 16352
rect 19519 16288 19535 16352
rect 19599 16288 19615 16352
rect 19679 16288 19685 16352
rect 19369 16287 19685 16288
rect 26959 16352 27275 16353
rect 26959 16288 26965 16352
rect 27029 16288 27045 16352
rect 27109 16288 27125 16352
rect 27189 16288 27205 16352
rect 27269 16288 27275 16352
rect 26959 16287 27275 16288
rect 21909 16282 21975 16285
rect 24485 16282 24551 16285
rect 21909 16280 24551 16282
rect 21909 16224 21914 16280
rect 21970 16224 24490 16280
rect 24546 16224 24551 16280
rect 21909 16222 24551 16224
rect 21909 16219 21975 16222
rect 24485 16219 24551 16222
rect 27889 16282 27955 16285
rect 28717 16282 28783 16285
rect 27889 16280 28783 16282
rect 27889 16224 27894 16280
rect 27950 16224 28722 16280
rect 28778 16224 28783 16280
rect 27889 16222 28783 16224
rect 27889 16219 27955 16222
rect 28717 16219 28783 16222
rect 2589 16146 2655 16149
rect 29361 16146 29427 16149
rect 2589 16144 29427 16146
rect 2589 16088 2594 16144
rect 2650 16088 29366 16144
rect 29422 16088 29427 16144
rect 2589 16086 29427 16088
rect 2589 16083 2655 16086
rect 29361 16083 29427 16086
rect 2221 16010 2287 16013
rect 28717 16010 28783 16013
rect 2221 16008 28783 16010
rect 2221 15952 2226 16008
rect 2282 15952 28722 16008
rect 28778 15952 28783 16008
rect 2221 15950 28783 15952
rect 2221 15947 2287 15950
rect 28717 15947 28783 15950
rect 29637 16010 29703 16013
rect 30373 16010 30439 16013
rect 29637 16008 30439 16010
rect 29637 15952 29642 16008
rect 29698 15952 30378 16008
rect 30434 15952 30439 16008
rect 29637 15950 30439 15952
rect 29637 15947 29703 15950
rect 30373 15947 30439 15950
rect 10777 15874 10843 15877
rect 13813 15874 13879 15877
rect 10777 15872 13879 15874
rect 10777 15816 10782 15872
rect 10838 15816 13818 15872
rect 13874 15816 13879 15872
rect 10777 15814 13879 15816
rect 10777 15811 10843 15814
rect 13813 15811 13879 15814
rect 20805 15874 20871 15877
rect 21817 15874 21883 15877
rect 20805 15872 21883 15874
rect 20805 15816 20810 15872
rect 20866 15816 21822 15872
rect 21878 15816 21883 15872
rect 20805 15814 21883 15816
rect 20805 15811 20871 15814
rect 21817 15811 21883 15814
rect 26233 15874 26299 15877
rect 29361 15874 29427 15877
rect 26233 15872 29427 15874
rect 26233 15816 26238 15872
rect 26294 15816 29366 15872
rect 29422 15816 29427 15872
rect 26233 15814 29427 15816
rect 26233 15811 26299 15814
rect 29361 15811 29427 15814
rect 7984 15808 8300 15809
rect 7984 15744 7990 15808
rect 8054 15744 8070 15808
rect 8134 15744 8150 15808
rect 8214 15744 8230 15808
rect 8294 15744 8300 15808
rect 7984 15743 8300 15744
rect 15574 15808 15890 15809
rect 15574 15744 15580 15808
rect 15644 15744 15660 15808
rect 15724 15744 15740 15808
rect 15804 15744 15820 15808
rect 15884 15744 15890 15808
rect 15574 15743 15890 15744
rect 23164 15808 23480 15809
rect 23164 15744 23170 15808
rect 23234 15744 23250 15808
rect 23314 15744 23330 15808
rect 23394 15744 23410 15808
rect 23474 15744 23480 15808
rect 23164 15743 23480 15744
rect 30754 15808 31070 15809
rect 30754 15744 30760 15808
rect 30824 15744 30840 15808
rect 30904 15744 30920 15808
rect 30984 15744 31000 15808
rect 31064 15744 31070 15808
rect 30754 15743 31070 15744
rect 9622 15676 9628 15740
rect 9692 15738 9698 15740
rect 11145 15738 11211 15741
rect 9692 15736 11211 15738
rect 9692 15680 11150 15736
rect 11206 15680 11211 15736
rect 9692 15678 11211 15680
rect 9692 15676 9698 15678
rect 11145 15675 11211 15678
rect 23841 15738 23907 15741
rect 25957 15738 26023 15741
rect 23841 15736 26023 15738
rect 23841 15680 23846 15736
rect 23902 15680 25962 15736
rect 26018 15680 26023 15736
rect 23841 15678 26023 15680
rect 23841 15675 23907 15678
rect 25957 15675 26023 15678
rect 26785 15738 26851 15741
rect 29637 15738 29703 15741
rect 26785 15736 29703 15738
rect 26785 15680 26790 15736
rect 26846 15680 29642 15736
rect 29698 15680 29703 15736
rect 26785 15678 29703 15680
rect 26785 15675 26851 15678
rect 29637 15675 29703 15678
rect 6637 15602 6703 15605
rect 13445 15602 13511 15605
rect 6637 15600 13511 15602
rect 6637 15544 6642 15600
rect 6698 15544 13450 15600
rect 13506 15544 13511 15600
rect 6637 15542 13511 15544
rect 6637 15539 6703 15542
rect 13445 15539 13511 15542
rect 17309 15602 17375 15605
rect 18137 15602 18203 15605
rect 17309 15600 18203 15602
rect 17309 15544 17314 15600
rect 17370 15544 18142 15600
rect 18198 15544 18203 15600
rect 17309 15542 18203 15544
rect 17309 15539 17375 15542
rect 18137 15539 18203 15542
rect 22001 15602 22067 15605
rect 27613 15602 27679 15605
rect 22001 15600 27679 15602
rect 22001 15544 22006 15600
rect 22062 15544 27618 15600
rect 27674 15544 27679 15600
rect 22001 15542 27679 15544
rect 22001 15539 22067 15542
rect 27613 15539 27679 15542
rect 2957 15466 3023 15469
rect 10409 15466 10475 15469
rect 2957 15464 10475 15466
rect 2957 15408 2962 15464
rect 3018 15408 10414 15464
rect 10470 15408 10475 15464
rect 2957 15406 10475 15408
rect 2957 15403 3023 15406
rect 10409 15403 10475 15406
rect 17033 15466 17099 15469
rect 21357 15466 21423 15469
rect 24158 15466 24164 15468
rect 17033 15464 19810 15466
rect 17033 15408 17038 15464
rect 17094 15408 19810 15464
rect 17033 15406 19810 15408
rect 17033 15403 17099 15406
rect 6637 15330 6703 15333
rect 11053 15330 11119 15333
rect 6637 15328 11119 15330
rect 6637 15272 6642 15328
rect 6698 15272 11058 15328
rect 11114 15272 11119 15328
rect 6637 15270 11119 15272
rect 6637 15267 6703 15270
rect 11053 15267 11119 15270
rect 17677 15330 17743 15333
rect 18873 15330 18939 15333
rect 17677 15328 18939 15330
rect 17677 15272 17682 15328
rect 17738 15272 18878 15328
rect 18934 15272 18939 15328
rect 17677 15270 18939 15272
rect 19750 15330 19810 15406
rect 21357 15464 24164 15466
rect 21357 15408 21362 15464
rect 21418 15408 24164 15464
rect 21357 15406 24164 15408
rect 21357 15403 21423 15406
rect 24158 15404 24164 15406
rect 24228 15404 24234 15468
rect 26006 15406 27538 15466
rect 26006 15330 26066 15406
rect 19750 15270 26066 15330
rect 17677 15267 17743 15270
rect 18873 15267 18939 15270
rect 26366 15268 26372 15332
rect 26436 15330 26442 15332
rect 26785 15330 26851 15333
rect 26436 15328 26851 15330
rect 26436 15272 26790 15328
rect 26846 15272 26851 15328
rect 26436 15270 26851 15272
rect 27478 15330 27538 15406
rect 29269 15330 29335 15333
rect 27478 15328 29335 15330
rect 27478 15272 29274 15328
rect 29330 15272 29335 15328
rect 27478 15270 29335 15272
rect 26436 15268 26442 15270
rect 26785 15267 26851 15270
rect 29269 15267 29335 15270
rect 4189 15264 4505 15265
rect 4189 15200 4195 15264
rect 4259 15200 4275 15264
rect 4339 15200 4355 15264
rect 4419 15200 4435 15264
rect 4499 15200 4505 15264
rect 4189 15199 4505 15200
rect 11779 15264 12095 15265
rect 11779 15200 11785 15264
rect 11849 15200 11865 15264
rect 11929 15200 11945 15264
rect 12009 15200 12025 15264
rect 12089 15200 12095 15264
rect 11779 15199 12095 15200
rect 19369 15264 19685 15265
rect 19369 15200 19375 15264
rect 19439 15200 19455 15264
rect 19519 15200 19535 15264
rect 19599 15200 19615 15264
rect 19679 15200 19685 15264
rect 19369 15199 19685 15200
rect 26959 15264 27275 15265
rect 26959 15200 26965 15264
rect 27029 15200 27045 15264
rect 27109 15200 27125 15264
rect 27189 15200 27205 15264
rect 27269 15200 27275 15264
rect 26959 15199 27275 15200
rect 6085 15194 6151 15197
rect 8569 15194 8635 15197
rect 10593 15196 10659 15197
rect 6085 15192 8635 15194
rect 6085 15136 6090 15192
rect 6146 15136 8574 15192
rect 8630 15136 8635 15192
rect 6085 15134 8635 15136
rect 6085 15131 6151 15134
rect 8569 15131 8635 15134
rect 10542 15132 10548 15196
rect 10612 15194 10659 15196
rect 19793 15194 19859 15197
rect 25773 15194 25839 15197
rect 10612 15192 10704 15194
rect 10654 15136 10704 15192
rect 10612 15134 10704 15136
rect 19793 15192 25839 15194
rect 19793 15136 19798 15192
rect 19854 15136 25778 15192
rect 25834 15136 25839 15192
rect 19793 15134 25839 15136
rect 10612 15132 10659 15134
rect 10593 15131 10659 15132
rect 19793 15131 19859 15134
rect 25773 15131 25839 15134
rect 6545 15058 6611 15061
rect 13077 15058 13143 15061
rect 6545 15056 13143 15058
rect 6545 15000 6550 15056
rect 6606 15000 13082 15056
rect 13138 15000 13143 15056
rect 6545 14998 13143 15000
rect 6545 14995 6611 14998
rect 13077 14995 13143 14998
rect 16941 15058 17007 15061
rect 29085 15058 29151 15061
rect 16941 15056 29151 15058
rect 16941 15000 16946 15056
rect 17002 15000 29090 15056
rect 29146 15000 29151 15056
rect 16941 14998 29151 15000
rect 16941 14995 17007 14998
rect 29085 14995 29151 14998
rect 3601 14922 3667 14925
rect 12198 14922 12204 14924
rect 3601 14920 12204 14922
rect 3601 14864 3606 14920
rect 3662 14864 12204 14920
rect 3601 14862 12204 14864
rect 3601 14859 3667 14862
rect 12198 14860 12204 14862
rect 12268 14860 12274 14924
rect 14825 14922 14891 14925
rect 17769 14922 17835 14925
rect 14825 14920 17835 14922
rect 14825 14864 14830 14920
rect 14886 14864 17774 14920
rect 17830 14864 17835 14920
rect 14825 14862 17835 14864
rect 14825 14859 14891 14862
rect 17769 14859 17835 14862
rect 20437 14922 20503 14925
rect 25681 14922 25747 14925
rect 20437 14920 25747 14922
rect 20437 14864 20442 14920
rect 20498 14864 25686 14920
rect 25742 14864 25747 14920
rect 20437 14862 25747 14864
rect 20437 14859 20503 14862
rect 25681 14859 25747 14862
rect 26141 14922 26207 14925
rect 29494 14922 29500 14924
rect 26141 14920 29500 14922
rect 26141 14864 26146 14920
rect 26202 14864 29500 14920
rect 26141 14862 29500 14864
rect 26141 14859 26207 14862
rect 29494 14860 29500 14862
rect 29564 14922 29570 14924
rect 30005 14922 30071 14925
rect 29564 14920 30071 14922
rect 29564 14864 30010 14920
rect 30066 14864 30071 14920
rect 29564 14862 30071 14864
rect 29564 14860 29570 14862
rect 30005 14859 30071 14862
rect 6269 14786 6335 14789
rect 7281 14786 7347 14789
rect 6269 14784 7347 14786
rect 6269 14728 6274 14784
rect 6330 14728 7286 14784
rect 7342 14728 7347 14784
rect 6269 14726 7347 14728
rect 6269 14723 6335 14726
rect 7281 14723 7347 14726
rect 19701 14786 19767 14789
rect 22369 14786 22435 14789
rect 19701 14784 22435 14786
rect 19701 14728 19706 14784
rect 19762 14728 22374 14784
rect 22430 14728 22435 14784
rect 19701 14726 22435 14728
rect 19701 14723 19767 14726
rect 22369 14723 22435 14726
rect 24025 14786 24091 14789
rect 26144 14786 26204 14859
rect 24025 14784 26204 14786
rect 24025 14728 24030 14784
rect 24086 14728 26204 14784
rect 24025 14726 26204 14728
rect 24025 14723 24091 14726
rect 7984 14720 8300 14721
rect 7984 14656 7990 14720
rect 8054 14656 8070 14720
rect 8134 14656 8150 14720
rect 8214 14656 8230 14720
rect 8294 14656 8300 14720
rect 7984 14655 8300 14656
rect 15574 14720 15890 14721
rect 15574 14656 15580 14720
rect 15644 14656 15660 14720
rect 15724 14656 15740 14720
rect 15804 14656 15820 14720
rect 15884 14656 15890 14720
rect 15574 14655 15890 14656
rect 23164 14720 23480 14721
rect 23164 14656 23170 14720
rect 23234 14656 23250 14720
rect 23314 14656 23330 14720
rect 23394 14656 23410 14720
rect 23474 14656 23480 14720
rect 23164 14655 23480 14656
rect 30754 14720 31070 14721
rect 30754 14656 30760 14720
rect 30824 14656 30840 14720
rect 30904 14656 30920 14720
rect 30984 14656 31000 14720
rect 31064 14656 31070 14720
rect 30754 14655 31070 14656
rect 4153 14650 4219 14653
rect 6729 14650 6795 14653
rect 4153 14648 6795 14650
rect 4153 14592 4158 14648
rect 4214 14592 6734 14648
rect 6790 14592 6795 14648
rect 4153 14590 6795 14592
rect 4153 14587 4219 14590
rect 6729 14587 6795 14590
rect 8753 14650 8819 14653
rect 10317 14650 10383 14653
rect 16573 14650 16639 14653
rect 19609 14650 19675 14653
rect 30189 14650 30255 14653
rect 8753 14648 12634 14650
rect 8753 14592 8758 14648
rect 8814 14592 10322 14648
rect 10378 14592 12634 14648
rect 8753 14590 12634 14592
rect 8753 14587 8819 14590
rect 10317 14587 10383 14590
rect 657 14514 723 14517
rect 6545 14514 6611 14517
rect 10317 14514 10383 14517
rect 657 14512 10383 14514
rect 657 14456 662 14512
rect 718 14456 6550 14512
rect 6606 14456 10322 14512
rect 10378 14456 10383 14512
rect 657 14454 10383 14456
rect 12574 14514 12634 14590
rect 16573 14648 19675 14650
rect 16573 14592 16578 14648
rect 16634 14592 19614 14648
rect 19670 14592 19675 14648
rect 16573 14590 19675 14592
rect 16573 14587 16639 14590
rect 19609 14587 19675 14590
rect 23614 14648 30255 14650
rect 23614 14592 30194 14648
rect 30250 14592 30255 14648
rect 23614 14590 30255 14592
rect 12709 14514 12775 14517
rect 12574 14512 12775 14514
rect 12574 14456 12714 14512
rect 12770 14456 12775 14512
rect 12574 14454 12775 14456
rect 657 14451 723 14454
rect 6545 14451 6611 14454
rect 10317 14451 10383 14454
rect 12709 14451 12775 14454
rect 17493 14514 17559 14517
rect 23105 14514 23171 14517
rect 17493 14512 23171 14514
rect 17493 14456 17498 14512
rect 17554 14456 23110 14512
rect 23166 14456 23171 14512
rect 17493 14454 23171 14456
rect 17493 14451 17559 14454
rect 23105 14451 23171 14454
rect 2957 14378 3023 14381
rect 23614 14378 23674 14590
rect 30189 14587 30255 14590
rect 23933 14514 23999 14517
rect 26785 14514 26851 14517
rect 2957 14376 23674 14378
rect 2957 14320 2962 14376
rect 3018 14320 23674 14376
rect 2957 14318 23674 14320
rect 23798 14512 26851 14514
rect 23798 14456 23938 14512
rect 23994 14456 26790 14512
rect 26846 14456 26851 14512
rect 23798 14454 26851 14456
rect 2957 14315 3023 14318
rect 6177 14242 6243 14245
rect 8937 14242 9003 14245
rect 10317 14244 10383 14245
rect 10317 14242 10364 14244
rect 6177 14240 9003 14242
rect 6177 14184 6182 14240
rect 6238 14184 8942 14240
rect 8998 14184 9003 14240
rect 6177 14182 9003 14184
rect 10272 14240 10364 14242
rect 10272 14184 10322 14240
rect 10272 14182 10364 14184
rect 6177 14179 6243 14182
rect 8937 14179 9003 14182
rect 10317 14180 10364 14182
rect 10428 14180 10434 14244
rect 12198 14180 12204 14244
rect 12268 14180 12274 14244
rect 13077 14242 13143 14245
rect 16297 14242 16363 14245
rect 13077 14240 16363 14242
rect 13077 14184 13082 14240
rect 13138 14184 16302 14240
rect 16358 14184 16363 14240
rect 13077 14182 16363 14184
rect 10317 14179 10383 14180
rect 4189 14176 4505 14177
rect 4189 14112 4195 14176
rect 4259 14112 4275 14176
rect 4339 14112 4355 14176
rect 4419 14112 4435 14176
rect 4499 14112 4505 14176
rect 4189 14111 4505 14112
rect 11779 14176 12095 14177
rect 11779 14112 11785 14176
rect 11849 14112 11865 14176
rect 11929 14112 11945 14176
rect 12009 14112 12025 14176
rect 12089 14112 12095 14176
rect 11779 14111 12095 14112
rect 5901 14106 5967 14109
rect 8661 14106 8727 14109
rect 5901 14104 8727 14106
rect 5901 14048 5906 14104
rect 5962 14048 8666 14104
rect 8722 14048 8727 14104
rect 5901 14046 8727 14048
rect 5901 14043 5967 14046
rect 8661 14043 8727 14046
rect 5165 13970 5231 13973
rect 11973 13970 12039 13973
rect 5165 13968 12039 13970
rect 5165 13912 5170 13968
rect 5226 13912 11978 13968
rect 12034 13912 12039 13968
rect 5165 13910 12039 13912
rect 5165 13907 5231 13910
rect 11973 13907 12039 13910
rect 1669 13836 1735 13837
rect 1669 13832 1716 13836
rect 1780 13834 1786 13836
rect 5441 13834 5507 13837
rect 7005 13834 7071 13837
rect 9213 13834 9279 13837
rect 1669 13776 1674 13832
rect 1669 13772 1716 13776
rect 1780 13774 1826 13834
rect 5441 13832 7071 13834
rect 5441 13776 5446 13832
rect 5502 13776 7010 13832
rect 7066 13776 7071 13832
rect 5441 13774 7071 13776
rect 1780 13772 1786 13774
rect 1669 13771 1735 13772
rect 5441 13771 5507 13774
rect 7005 13771 7071 13774
rect 7790 13832 9279 13834
rect 7790 13776 9218 13832
rect 9274 13776 9279 13832
rect 7790 13774 9279 13776
rect 6494 13636 6500 13700
rect 6564 13698 6570 13700
rect 7790 13698 7850 13774
rect 9213 13771 9279 13774
rect 11094 13772 11100 13836
rect 11164 13834 11170 13836
rect 11973 13834 12039 13837
rect 11164 13832 12039 13834
rect 11164 13776 11978 13832
rect 12034 13776 12039 13832
rect 11164 13774 12039 13776
rect 12206 13834 12266 14180
rect 13077 14179 13143 14182
rect 16297 14179 16363 14182
rect 20161 14242 20227 14245
rect 23798 14242 23858 14454
rect 23933 14451 23999 14454
rect 26785 14451 26851 14454
rect 26509 14378 26575 14381
rect 27981 14378 28047 14381
rect 26509 14376 28047 14378
rect 26509 14320 26514 14376
rect 26570 14320 27986 14376
rect 28042 14320 28047 14376
rect 26509 14318 28047 14320
rect 26509 14315 26575 14318
rect 27981 14315 28047 14318
rect 20161 14240 23858 14242
rect 20161 14184 20166 14240
rect 20222 14184 23858 14240
rect 20161 14182 23858 14184
rect 20161 14179 20227 14182
rect 19369 14176 19685 14177
rect 19369 14112 19375 14176
rect 19439 14112 19455 14176
rect 19519 14112 19535 14176
rect 19599 14112 19615 14176
rect 19679 14112 19685 14176
rect 19369 14111 19685 14112
rect 26959 14176 27275 14177
rect 26959 14112 26965 14176
rect 27029 14112 27045 14176
rect 27109 14112 27125 14176
rect 27189 14112 27205 14176
rect 27269 14112 27275 14176
rect 26959 14111 27275 14112
rect 19885 14106 19951 14109
rect 26693 14106 26759 14109
rect 19885 14104 26759 14106
rect 19885 14048 19890 14104
rect 19946 14048 26698 14104
rect 26754 14048 26759 14104
rect 19885 14046 26759 14048
rect 19885 14043 19951 14046
rect 26693 14043 26759 14046
rect 13445 13970 13511 13973
rect 19517 13970 19583 13973
rect 24117 13970 24183 13973
rect 13445 13968 13554 13970
rect 13445 13912 13450 13968
rect 13506 13912 13554 13968
rect 13445 13907 13554 13912
rect 19517 13968 24183 13970
rect 19517 13912 19522 13968
rect 19578 13912 24122 13968
rect 24178 13912 24183 13968
rect 19517 13910 24183 13912
rect 19517 13907 19583 13910
rect 24117 13907 24183 13910
rect 26785 13970 26851 13973
rect 28901 13970 28967 13973
rect 26785 13968 28967 13970
rect 26785 13912 26790 13968
rect 26846 13912 28906 13968
rect 28962 13912 28967 13968
rect 26785 13910 28967 13912
rect 26785 13907 26851 13910
rect 28901 13907 28967 13910
rect 13353 13834 13419 13837
rect 12206 13832 13419 13834
rect 12206 13776 13358 13832
rect 13414 13776 13419 13832
rect 12206 13774 13419 13776
rect 11164 13772 11170 13774
rect 11973 13771 12039 13774
rect 13353 13771 13419 13774
rect 6564 13638 7850 13698
rect 11053 13698 11119 13701
rect 13494 13698 13554 13907
rect 15653 13834 15719 13837
rect 19149 13834 19215 13837
rect 15653 13832 19215 13834
rect 15653 13776 15658 13832
rect 15714 13776 19154 13832
rect 19210 13776 19215 13832
rect 15653 13774 19215 13776
rect 15653 13771 15719 13774
rect 19149 13771 19215 13774
rect 20621 13834 20687 13837
rect 29821 13834 29887 13837
rect 30046 13834 30052 13836
rect 20621 13832 23674 13834
rect 20621 13776 20626 13832
rect 20682 13776 23674 13832
rect 20621 13774 23674 13776
rect 20621 13771 20687 13774
rect 11053 13696 13554 13698
rect 11053 13640 11058 13696
rect 11114 13640 13554 13696
rect 11053 13638 13554 13640
rect 23614 13698 23674 13774
rect 29821 13832 30052 13834
rect 29821 13776 29826 13832
rect 29882 13776 30052 13832
rect 29821 13774 30052 13776
rect 29821 13771 29887 13774
rect 30046 13772 30052 13774
rect 30116 13772 30122 13836
rect 24761 13698 24827 13701
rect 23614 13696 24827 13698
rect 23614 13640 24766 13696
rect 24822 13640 24827 13696
rect 23614 13638 24827 13640
rect 6564 13636 6570 13638
rect 11053 13635 11119 13638
rect 24761 13635 24827 13638
rect 7984 13632 8300 13633
rect 7984 13568 7990 13632
rect 8054 13568 8070 13632
rect 8134 13568 8150 13632
rect 8214 13568 8230 13632
rect 8294 13568 8300 13632
rect 7984 13567 8300 13568
rect 15574 13632 15890 13633
rect 15574 13568 15580 13632
rect 15644 13568 15660 13632
rect 15724 13568 15740 13632
rect 15804 13568 15820 13632
rect 15884 13568 15890 13632
rect 15574 13567 15890 13568
rect 23164 13632 23480 13633
rect 23164 13568 23170 13632
rect 23234 13568 23250 13632
rect 23314 13568 23330 13632
rect 23394 13568 23410 13632
rect 23474 13568 23480 13632
rect 23164 13567 23480 13568
rect 30754 13632 31070 13633
rect 30754 13568 30760 13632
rect 30824 13568 30840 13632
rect 30904 13568 30920 13632
rect 30984 13568 31000 13632
rect 31064 13568 31070 13632
rect 30754 13567 31070 13568
rect 1945 13562 2011 13565
rect 7465 13562 7531 13565
rect 1945 13560 7531 13562
rect 1945 13504 1950 13560
rect 2006 13504 7470 13560
rect 7526 13504 7531 13560
rect 1945 13502 7531 13504
rect 1945 13499 2011 13502
rect 7465 13499 7531 13502
rect 8518 13500 8524 13564
rect 8588 13562 8594 13564
rect 8588 13502 15026 13562
rect 8588 13500 8594 13502
rect 3601 13426 3667 13429
rect 10409 13426 10475 13429
rect 3601 13424 10475 13426
rect 3601 13368 3606 13424
rect 3662 13368 10414 13424
rect 10470 13368 10475 13424
rect 3601 13366 10475 13368
rect 3601 13363 3667 13366
rect 10409 13363 10475 13366
rect 10550 13366 12082 13426
rect 3601 13290 3667 13293
rect 6729 13290 6795 13293
rect 3601 13288 6795 13290
rect 3601 13232 3606 13288
rect 3662 13232 6734 13288
rect 6790 13232 6795 13288
rect 3601 13230 6795 13232
rect 3601 13227 3667 13230
rect 6729 13227 6795 13230
rect 7598 13228 7604 13292
rect 7668 13290 7674 13292
rect 10550 13290 10610 13366
rect 11789 13290 11855 13293
rect 7668 13230 10610 13290
rect 11654 13288 11855 13290
rect 11654 13232 11794 13288
rect 11850 13232 11855 13288
rect 11654 13230 11855 13232
rect 12022 13290 12082 13366
rect 12382 13364 12388 13428
rect 12452 13426 12458 13428
rect 12893 13426 12959 13429
rect 12452 13424 12959 13426
rect 12452 13368 12898 13424
rect 12954 13368 12959 13424
rect 12452 13366 12959 13368
rect 14966 13426 15026 13502
rect 17585 13426 17651 13429
rect 14966 13424 17651 13426
rect 14966 13368 17590 13424
rect 17646 13368 17651 13424
rect 14966 13366 17651 13368
rect 12452 13364 12458 13366
rect 12893 13363 12959 13366
rect 17585 13363 17651 13366
rect 22001 13426 22067 13429
rect 28073 13426 28139 13429
rect 22001 13424 28139 13426
rect 22001 13368 22006 13424
rect 22062 13368 28078 13424
rect 28134 13368 28139 13424
rect 22001 13366 28139 13368
rect 22001 13363 22067 13366
rect 28073 13363 28139 13366
rect 13813 13290 13879 13293
rect 12022 13288 13879 13290
rect 12022 13232 13818 13288
rect 13874 13232 13879 13288
rect 12022 13230 13879 13232
rect 7668 13228 7674 13230
rect 5073 13154 5139 13157
rect 11654 13154 11714 13230
rect 11789 13227 11855 13230
rect 13813 13227 13879 13230
rect 22502 13228 22508 13292
rect 22572 13290 22578 13292
rect 22572 13230 27538 13290
rect 22572 13228 22578 13230
rect 5073 13152 11714 13154
rect 5073 13096 5078 13152
rect 5134 13096 11714 13152
rect 5073 13094 11714 13096
rect 12433 13154 12499 13157
rect 13813 13154 13879 13157
rect 12433 13152 13879 13154
rect 12433 13096 12438 13152
rect 12494 13096 13818 13152
rect 13874 13096 13879 13152
rect 12433 13094 13879 13096
rect 5073 13091 5139 13094
rect 12433 13091 12499 13094
rect 13813 13091 13879 13094
rect 21265 13154 21331 13157
rect 26366 13154 26372 13156
rect 21265 13152 26372 13154
rect 21265 13096 21270 13152
rect 21326 13096 26372 13152
rect 21265 13094 26372 13096
rect 21265 13091 21331 13094
rect 26366 13092 26372 13094
rect 26436 13092 26442 13156
rect 27478 13154 27538 13230
rect 29913 13154 29979 13157
rect 27478 13152 29979 13154
rect 27478 13096 29918 13152
rect 29974 13096 29979 13152
rect 27478 13094 29979 13096
rect 29913 13091 29979 13094
rect 4189 13088 4505 13089
rect 4189 13024 4195 13088
rect 4259 13024 4275 13088
rect 4339 13024 4355 13088
rect 4419 13024 4435 13088
rect 4499 13024 4505 13088
rect 4189 13023 4505 13024
rect 11779 13088 12095 13089
rect 11779 13024 11785 13088
rect 11849 13024 11865 13088
rect 11929 13024 11945 13088
rect 12009 13024 12025 13088
rect 12089 13024 12095 13088
rect 11779 13023 12095 13024
rect 19369 13088 19685 13089
rect 19369 13024 19375 13088
rect 19439 13024 19455 13088
rect 19519 13024 19535 13088
rect 19599 13024 19615 13088
rect 19679 13024 19685 13088
rect 19369 13023 19685 13024
rect 26959 13088 27275 13089
rect 26959 13024 26965 13088
rect 27029 13024 27045 13088
rect 27109 13024 27125 13088
rect 27189 13024 27205 13088
rect 27269 13024 27275 13088
rect 26959 13023 27275 13024
rect 4889 13018 4955 13021
rect 11237 13020 11303 13021
rect 4889 13016 11116 13018
rect 4889 12960 4894 13016
rect 4950 12960 11116 13016
rect 4889 12958 11116 12960
rect 4889 12955 4955 12958
rect 3049 12882 3115 12885
rect 10869 12882 10935 12885
rect 3049 12880 10935 12882
rect 3049 12824 3054 12880
rect 3110 12824 10874 12880
rect 10930 12824 10935 12880
rect 3049 12822 10935 12824
rect 11056 12882 11116 12958
rect 11237 13016 11284 13020
rect 11348 13018 11354 13020
rect 11237 12960 11242 13016
rect 11237 12956 11284 12960
rect 11348 12958 11394 13018
rect 11348 12956 11354 12958
rect 11462 12956 11468 13020
rect 11532 13018 11538 13020
rect 11605 13018 11671 13021
rect 11532 13016 11671 13018
rect 11532 12960 11610 13016
rect 11666 12960 11671 13016
rect 11532 12958 11671 12960
rect 11532 12956 11538 12958
rect 11237 12955 11303 12956
rect 11605 12955 11671 12958
rect 12382 12956 12388 13020
rect 12452 12956 12458 13020
rect 21909 13018 21975 13021
rect 24301 13018 24367 13021
rect 21909 13016 24367 13018
rect 21909 12960 21914 13016
rect 21970 12960 24306 13016
rect 24362 12960 24367 13016
rect 21909 12958 24367 12960
rect 12390 12882 12450 12956
rect 21909 12955 21975 12958
rect 24301 12955 24367 12958
rect 11056 12822 12450 12882
rect 3049 12819 3115 12822
rect 10869 12819 10935 12822
rect 21950 12820 21956 12884
rect 22020 12882 22026 12884
rect 29821 12882 29887 12885
rect 22020 12880 29887 12882
rect 22020 12824 29826 12880
rect 29882 12824 29887 12880
rect 22020 12822 29887 12824
rect 22020 12820 22026 12822
rect 29821 12819 29887 12822
rect 2221 12746 2287 12749
rect 11053 12746 11119 12749
rect 2221 12744 11119 12746
rect 2221 12688 2226 12744
rect 2282 12688 11058 12744
rect 11114 12688 11119 12744
rect 2221 12686 11119 12688
rect 2221 12683 2287 12686
rect 11053 12683 11119 12686
rect 23289 12746 23355 12749
rect 23289 12744 23674 12746
rect 23289 12688 23294 12744
rect 23350 12688 23674 12744
rect 23289 12686 23674 12688
rect 23289 12683 23355 12686
rect 1761 12610 1827 12613
rect 7649 12610 7715 12613
rect 1761 12608 7715 12610
rect 1761 12552 1766 12608
rect 1822 12552 7654 12608
rect 7710 12552 7715 12608
rect 1761 12550 7715 12552
rect 1761 12547 1827 12550
rect 7649 12547 7715 12550
rect 9029 12610 9095 12613
rect 11789 12610 11855 12613
rect 9029 12608 11855 12610
rect 9029 12552 9034 12608
rect 9090 12552 11794 12608
rect 11850 12552 11855 12608
rect 9029 12550 11855 12552
rect 9029 12547 9095 12550
rect 11789 12547 11855 12550
rect 7984 12544 8300 12545
rect 7984 12480 7990 12544
rect 8054 12480 8070 12544
rect 8134 12480 8150 12544
rect 8214 12480 8230 12544
rect 8294 12480 8300 12544
rect 7984 12479 8300 12480
rect 15574 12544 15890 12545
rect 15574 12480 15580 12544
rect 15644 12480 15660 12544
rect 15724 12480 15740 12544
rect 15804 12480 15820 12544
rect 15884 12480 15890 12544
rect 15574 12479 15890 12480
rect 23164 12544 23480 12545
rect 23164 12480 23170 12544
rect 23234 12480 23250 12544
rect 23314 12480 23330 12544
rect 23394 12480 23410 12544
rect 23474 12480 23480 12544
rect 23164 12479 23480 12480
rect 3734 12412 3740 12476
rect 3804 12474 3810 12476
rect 5717 12474 5783 12477
rect 3804 12472 5783 12474
rect 3804 12416 5722 12472
rect 5778 12416 5783 12472
rect 3804 12414 5783 12416
rect 3804 12412 3810 12414
rect 5717 12411 5783 12414
rect 6361 12474 6427 12477
rect 7097 12474 7163 12477
rect 12341 12474 12407 12477
rect 13486 12474 13492 12476
rect 6361 12472 7163 12474
rect 6361 12416 6366 12472
rect 6422 12416 7102 12472
rect 7158 12416 7163 12472
rect 6361 12414 7163 12416
rect 6361 12411 6427 12414
rect 7097 12411 7163 12414
rect 8710 12472 13492 12474
rect 8710 12416 12346 12472
rect 12402 12416 13492 12472
rect 8710 12414 13492 12416
rect 1945 12338 2011 12341
rect 8710 12338 8770 12414
rect 12341 12411 12407 12414
rect 13486 12412 13492 12414
rect 13556 12412 13562 12476
rect 18965 12474 19031 12477
rect 21173 12474 21239 12477
rect 18965 12472 21239 12474
rect 18965 12416 18970 12472
rect 19026 12416 21178 12472
rect 21234 12416 21239 12472
rect 18965 12414 21239 12416
rect 23614 12474 23674 12686
rect 26182 12684 26188 12748
rect 26252 12746 26258 12748
rect 30005 12746 30071 12749
rect 26252 12744 30071 12746
rect 26252 12688 30010 12744
rect 30066 12688 30071 12744
rect 26252 12686 30071 12688
rect 26252 12684 26258 12686
rect 30005 12683 30071 12686
rect 26141 12610 26207 12613
rect 29545 12610 29611 12613
rect 26141 12608 29611 12610
rect 26141 12552 26146 12608
rect 26202 12552 29550 12608
rect 29606 12552 29611 12608
rect 26141 12550 29611 12552
rect 26141 12547 26207 12550
rect 29545 12547 29611 12550
rect 30754 12544 31070 12545
rect 30754 12480 30760 12544
rect 30824 12480 30840 12544
rect 30904 12480 30920 12544
rect 30984 12480 31000 12544
rect 31064 12480 31070 12544
rect 30754 12479 31070 12480
rect 26509 12474 26575 12477
rect 29545 12476 29611 12477
rect 29494 12474 29500 12476
rect 23614 12472 26575 12474
rect 23614 12416 26514 12472
rect 26570 12416 26575 12472
rect 23614 12414 26575 12416
rect 29454 12414 29500 12474
rect 29564 12472 29611 12476
rect 29606 12416 29611 12472
rect 18965 12411 19031 12414
rect 21173 12411 21239 12414
rect 26509 12411 26575 12414
rect 29494 12412 29500 12414
rect 29564 12412 29611 12416
rect 29545 12411 29611 12412
rect 1945 12336 8770 12338
rect 1945 12280 1950 12336
rect 2006 12280 8770 12336
rect 1945 12278 8770 12280
rect 1945 12275 2011 12278
rect 8886 12276 8892 12340
rect 8956 12338 8962 12340
rect 11973 12338 12039 12341
rect 8956 12336 12039 12338
rect 8956 12280 11978 12336
rect 12034 12280 12039 12336
rect 8956 12278 12039 12280
rect 8956 12276 8962 12278
rect 11973 12275 12039 12278
rect 12709 12338 12775 12341
rect 13997 12338 14063 12341
rect 12709 12336 14063 12338
rect 12709 12280 12714 12336
rect 12770 12280 14002 12336
rect 14058 12280 14063 12336
rect 12709 12278 14063 12280
rect 12709 12275 12775 12278
rect 13997 12275 14063 12278
rect 22870 12276 22876 12340
rect 22940 12338 22946 12340
rect 30373 12338 30439 12341
rect 22940 12336 30439 12338
rect 22940 12280 30378 12336
rect 30434 12280 30439 12336
rect 22940 12278 30439 12280
rect 22940 12276 22946 12278
rect 30373 12275 30439 12278
rect 6678 12140 6684 12204
rect 6748 12202 6754 12204
rect 10409 12202 10475 12205
rect 6748 12200 10475 12202
rect 6748 12144 10414 12200
rect 10470 12144 10475 12200
rect 6748 12142 10475 12144
rect 6748 12140 6754 12142
rect 10409 12139 10475 12142
rect 11605 12202 11671 12205
rect 17677 12202 17743 12205
rect 11605 12200 17743 12202
rect 11605 12144 11610 12200
rect 11666 12144 17682 12200
rect 17738 12144 17743 12200
rect 11605 12142 17743 12144
rect 11605 12139 11671 12142
rect 17677 12139 17743 12142
rect 21541 12202 21607 12205
rect 28257 12202 28323 12205
rect 21541 12200 28323 12202
rect 21541 12144 21546 12200
rect 21602 12144 28262 12200
rect 28318 12144 28323 12200
rect 21541 12142 28323 12144
rect 21541 12139 21607 12142
rect 28257 12139 28323 12142
rect 4189 12000 4505 12001
rect 4189 11936 4195 12000
rect 4259 11936 4275 12000
rect 4339 11936 4355 12000
rect 4419 11936 4435 12000
rect 4499 11936 4505 12000
rect 4189 11935 4505 11936
rect 11779 12000 12095 12001
rect 11779 11936 11785 12000
rect 11849 11936 11865 12000
rect 11929 11936 11945 12000
rect 12009 11936 12025 12000
rect 12089 11936 12095 12000
rect 11779 11935 12095 11936
rect 19369 12000 19685 12001
rect 19369 11936 19375 12000
rect 19439 11936 19455 12000
rect 19519 11936 19535 12000
rect 19599 11936 19615 12000
rect 19679 11936 19685 12000
rect 19369 11935 19685 11936
rect 26959 12000 27275 12001
rect 26959 11936 26965 12000
rect 27029 11936 27045 12000
rect 27109 11936 27125 12000
rect 27189 11936 27205 12000
rect 27269 11936 27275 12000
rect 26959 11935 27275 11936
rect 12341 11930 12407 11933
rect 13169 11930 13235 11933
rect 12341 11928 13235 11930
rect 12341 11872 12346 11928
rect 12402 11872 13174 11928
rect 13230 11872 13235 11928
rect 12341 11870 13235 11872
rect 12341 11867 12407 11870
rect 13169 11867 13235 11870
rect 2129 11794 2195 11797
rect 9397 11794 9463 11797
rect 10777 11796 10843 11797
rect 2129 11792 9463 11794
rect 2129 11736 2134 11792
rect 2190 11736 9402 11792
rect 9458 11736 9463 11792
rect 2129 11734 9463 11736
rect 2129 11731 2195 11734
rect 9397 11731 9463 11734
rect 10726 11732 10732 11796
rect 10796 11794 10843 11796
rect 10796 11792 10888 11794
rect 10838 11736 10888 11792
rect 10796 11734 10888 11736
rect 10796 11732 10843 11734
rect 11646 11732 11652 11796
rect 11716 11794 11722 11796
rect 11973 11794 12039 11797
rect 11716 11792 12039 11794
rect 11716 11736 11978 11792
rect 12034 11736 12039 11792
rect 11716 11734 12039 11736
rect 11716 11732 11722 11734
rect 10777 11731 10843 11732
rect 11973 11731 12039 11734
rect 12433 11794 12499 11797
rect 14089 11794 14155 11797
rect 12433 11792 14155 11794
rect 12433 11736 12438 11792
rect 12494 11736 14094 11792
rect 14150 11736 14155 11792
rect 12433 11734 14155 11736
rect 12433 11731 12499 11734
rect 14089 11731 14155 11734
rect 2865 11658 2931 11661
rect 7189 11658 7255 11661
rect 2865 11656 7255 11658
rect 2865 11600 2870 11656
rect 2926 11600 7194 11656
rect 7250 11600 7255 11656
rect 2865 11598 7255 11600
rect 2865 11595 2931 11598
rect 7189 11595 7255 11598
rect 7782 11596 7788 11660
rect 7852 11658 7858 11660
rect 11053 11658 11119 11661
rect 7852 11656 11119 11658
rect 7852 11600 11058 11656
rect 11114 11600 11119 11656
rect 7852 11598 11119 11600
rect 7852 11596 7858 11598
rect 11053 11595 11119 11598
rect 23289 11658 23355 11661
rect 24485 11658 24551 11661
rect 23289 11656 24551 11658
rect 23289 11600 23294 11656
rect 23350 11600 24490 11656
rect 24546 11600 24551 11656
rect 23289 11598 24551 11600
rect 23289 11595 23355 11598
rect 24485 11595 24551 11598
rect 25129 11658 25195 11661
rect 27153 11658 27219 11661
rect 25129 11656 27219 11658
rect 25129 11600 25134 11656
rect 25190 11600 27158 11656
rect 27214 11600 27219 11656
rect 25129 11598 27219 11600
rect 25129 11595 25195 11598
rect 27153 11595 27219 11598
rect 7984 11456 8300 11457
rect 7984 11392 7990 11456
rect 8054 11392 8070 11456
rect 8134 11392 8150 11456
rect 8214 11392 8230 11456
rect 8294 11392 8300 11456
rect 7984 11391 8300 11392
rect 15574 11456 15890 11457
rect 15574 11392 15580 11456
rect 15644 11392 15660 11456
rect 15724 11392 15740 11456
rect 15804 11392 15820 11456
rect 15884 11392 15890 11456
rect 15574 11391 15890 11392
rect 23164 11456 23480 11457
rect 23164 11392 23170 11456
rect 23234 11392 23250 11456
rect 23314 11392 23330 11456
rect 23394 11392 23410 11456
rect 23474 11392 23480 11456
rect 23164 11391 23480 11392
rect 30754 11456 31070 11457
rect 30754 11392 30760 11456
rect 30824 11392 30840 11456
rect 30904 11392 30920 11456
rect 30984 11392 31000 11456
rect 31064 11392 31070 11456
rect 30754 11391 31070 11392
rect 10869 11386 10935 11389
rect 14549 11386 14615 11389
rect 10869 11384 14615 11386
rect 10869 11328 10874 11384
rect 10930 11328 14554 11384
rect 14610 11328 14615 11384
rect 10869 11326 14615 11328
rect 10869 11323 10935 11326
rect 14549 11323 14615 11326
rect 3693 11250 3759 11253
rect 9949 11250 10015 11253
rect 19793 11250 19859 11253
rect 3693 11248 19859 11250
rect 3693 11192 3698 11248
rect 3754 11192 9954 11248
rect 10010 11192 19798 11248
rect 19854 11192 19859 11248
rect 3693 11190 19859 11192
rect 3693 11187 3759 11190
rect 9949 11187 10015 11190
rect 19793 11187 19859 11190
rect 22461 11250 22527 11253
rect 25313 11250 25379 11253
rect 22461 11248 25379 11250
rect 22461 11192 22466 11248
rect 22522 11192 25318 11248
rect 25374 11192 25379 11248
rect 22461 11190 25379 11192
rect 22461 11187 22527 11190
rect 25313 11187 25379 11190
rect 9581 11114 9647 11117
rect 12801 11114 12867 11117
rect 9581 11112 12867 11114
rect 9581 11056 9586 11112
rect 9642 11056 12806 11112
rect 12862 11056 12867 11112
rect 9581 11054 12867 11056
rect 9581 11051 9647 11054
rect 12801 11051 12867 11054
rect 15142 11052 15148 11116
rect 15212 11114 15218 11116
rect 15745 11114 15811 11117
rect 15212 11112 15811 11114
rect 15212 11056 15750 11112
rect 15806 11056 15811 11112
rect 15212 11054 15811 11056
rect 15212 11052 15218 11054
rect 15745 11051 15811 11054
rect 16665 11114 16731 11117
rect 19977 11114 20043 11117
rect 31109 11114 31175 11117
rect 16665 11112 31175 11114
rect 16665 11056 16670 11112
rect 16726 11056 19982 11112
rect 20038 11056 31114 11112
rect 31170 11056 31175 11112
rect 16665 11054 31175 11056
rect 16665 11051 16731 11054
rect 19977 11051 20043 11054
rect 31109 11051 31175 11054
rect 12341 10978 12407 10981
rect 13813 10978 13879 10981
rect 12341 10976 13879 10978
rect 12341 10920 12346 10976
rect 12402 10920 13818 10976
rect 13874 10920 13879 10976
rect 12341 10918 13879 10920
rect 12341 10915 12407 10918
rect 13813 10915 13879 10918
rect 4189 10912 4505 10913
rect 4189 10848 4195 10912
rect 4259 10848 4275 10912
rect 4339 10848 4355 10912
rect 4419 10848 4435 10912
rect 4499 10848 4505 10912
rect 4189 10847 4505 10848
rect 11779 10912 12095 10913
rect 11779 10848 11785 10912
rect 11849 10848 11865 10912
rect 11929 10848 11945 10912
rect 12009 10848 12025 10912
rect 12089 10848 12095 10912
rect 11779 10847 12095 10848
rect 19369 10912 19685 10913
rect 19369 10848 19375 10912
rect 19439 10848 19455 10912
rect 19519 10848 19535 10912
rect 19599 10848 19615 10912
rect 19679 10848 19685 10912
rect 19369 10847 19685 10848
rect 26959 10912 27275 10913
rect 26959 10848 26965 10912
rect 27029 10848 27045 10912
rect 27109 10848 27125 10912
rect 27189 10848 27205 10912
rect 27269 10848 27275 10912
rect 26959 10847 27275 10848
rect 21357 10842 21423 10845
rect 25865 10842 25931 10845
rect 21357 10840 25931 10842
rect 21357 10784 21362 10840
rect 21418 10784 25870 10840
rect 25926 10784 25931 10840
rect 21357 10782 25931 10784
rect 21357 10779 21423 10782
rect 25865 10779 25931 10782
rect 2129 10706 2195 10709
rect 9622 10706 9628 10708
rect 2129 10704 9628 10706
rect 2129 10648 2134 10704
rect 2190 10648 9628 10704
rect 2129 10646 9628 10648
rect 2129 10643 2195 10646
rect 9622 10644 9628 10646
rect 9692 10644 9698 10708
rect 16573 10706 16639 10709
rect 12390 10704 16639 10706
rect 12390 10648 16578 10704
rect 16634 10648 16639 10704
rect 12390 10646 16639 10648
rect 5574 10508 5580 10572
rect 5644 10570 5650 10572
rect 12390 10570 12450 10646
rect 16573 10643 16639 10646
rect 22921 10706 22987 10709
rect 24209 10706 24275 10709
rect 22921 10704 24275 10706
rect 22921 10648 22926 10704
rect 22982 10648 24214 10704
rect 24270 10648 24275 10704
rect 22921 10646 24275 10648
rect 22921 10643 22987 10646
rect 24209 10643 24275 10646
rect 5644 10510 12450 10570
rect 20437 10570 20503 10573
rect 24209 10570 24275 10573
rect 20437 10568 24275 10570
rect 20437 10512 20442 10568
rect 20498 10512 24214 10568
rect 24270 10512 24275 10568
rect 20437 10510 24275 10512
rect 5644 10508 5650 10510
rect 20437 10507 20503 10510
rect 24209 10507 24275 10510
rect 10777 10434 10843 10437
rect 12617 10434 12683 10437
rect 13261 10434 13327 10437
rect 10777 10432 13327 10434
rect 10777 10376 10782 10432
rect 10838 10376 12622 10432
rect 12678 10376 13266 10432
rect 13322 10376 13327 10432
rect 10777 10374 13327 10376
rect 10777 10371 10843 10374
rect 12617 10371 12683 10374
rect 13261 10371 13327 10374
rect 7984 10368 8300 10369
rect 7984 10304 7990 10368
rect 8054 10304 8070 10368
rect 8134 10304 8150 10368
rect 8214 10304 8230 10368
rect 8294 10304 8300 10368
rect 7984 10303 8300 10304
rect 15574 10368 15890 10369
rect 15574 10304 15580 10368
rect 15644 10304 15660 10368
rect 15724 10304 15740 10368
rect 15804 10304 15820 10368
rect 15884 10304 15890 10368
rect 15574 10303 15890 10304
rect 23164 10368 23480 10369
rect 23164 10304 23170 10368
rect 23234 10304 23250 10368
rect 23314 10304 23330 10368
rect 23394 10304 23410 10368
rect 23474 10304 23480 10368
rect 23164 10303 23480 10304
rect 30754 10368 31070 10369
rect 30754 10304 30760 10368
rect 30824 10304 30840 10368
rect 30904 10304 30920 10368
rect 30984 10304 31000 10368
rect 31064 10304 31070 10368
rect 30754 10303 31070 10304
rect 11421 10298 11487 10301
rect 12249 10298 12315 10301
rect 11421 10296 12315 10298
rect 11421 10240 11426 10296
rect 11482 10240 12254 10296
rect 12310 10240 12315 10296
rect 11421 10238 12315 10240
rect 11421 10235 11487 10238
rect 12249 10235 12315 10238
rect 3918 10100 3924 10164
rect 3988 10162 3994 10164
rect 16573 10162 16639 10165
rect 3988 10160 16639 10162
rect 3988 10104 16578 10160
rect 16634 10104 16639 10160
rect 3988 10102 16639 10104
rect 3988 10100 3994 10102
rect 16573 10099 16639 10102
rect 4981 10026 5047 10029
rect 16757 10026 16823 10029
rect 4981 10024 16823 10026
rect 4981 9968 4986 10024
rect 5042 9968 16762 10024
rect 16818 9968 16823 10024
rect 4981 9966 16823 9968
rect 4981 9963 5047 9966
rect 16757 9963 16823 9966
rect 4189 9824 4505 9825
rect 4189 9760 4195 9824
rect 4259 9760 4275 9824
rect 4339 9760 4355 9824
rect 4419 9760 4435 9824
rect 4499 9760 4505 9824
rect 4189 9759 4505 9760
rect 11779 9824 12095 9825
rect 11779 9760 11785 9824
rect 11849 9760 11865 9824
rect 11929 9760 11945 9824
rect 12009 9760 12025 9824
rect 12089 9760 12095 9824
rect 11779 9759 12095 9760
rect 19369 9824 19685 9825
rect 19369 9760 19375 9824
rect 19439 9760 19455 9824
rect 19519 9760 19535 9824
rect 19599 9760 19615 9824
rect 19679 9760 19685 9824
rect 19369 9759 19685 9760
rect 26959 9824 27275 9825
rect 26959 9760 26965 9824
rect 27029 9760 27045 9824
rect 27109 9760 27125 9824
rect 27189 9760 27205 9824
rect 27269 9760 27275 9824
rect 26959 9759 27275 9760
rect 24761 9618 24827 9621
rect 26049 9618 26115 9621
rect 24761 9616 26115 9618
rect 24761 9560 24766 9616
rect 24822 9560 26054 9616
rect 26110 9560 26115 9616
rect 24761 9558 26115 9560
rect 24761 9555 24827 9558
rect 26049 9555 26115 9558
rect 24117 9482 24183 9485
rect 25037 9482 25103 9485
rect 24117 9480 25103 9482
rect 24117 9424 24122 9480
rect 24178 9424 25042 9480
rect 25098 9424 25103 9480
rect 24117 9422 25103 9424
rect 24117 9419 24183 9422
rect 25037 9419 25103 9422
rect 7984 9280 8300 9281
rect 7984 9216 7990 9280
rect 8054 9216 8070 9280
rect 8134 9216 8150 9280
rect 8214 9216 8230 9280
rect 8294 9216 8300 9280
rect 7984 9215 8300 9216
rect 15574 9280 15890 9281
rect 15574 9216 15580 9280
rect 15644 9216 15660 9280
rect 15724 9216 15740 9280
rect 15804 9216 15820 9280
rect 15884 9216 15890 9280
rect 15574 9215 15890 9216
rect 23164 9280 23480 9281
rect 23164 9216 23170 9280
rect 23234 9216 23250 9280
rect 23314 9216 23330 9280
rect 23394 9216 23410 9280
rect 23474 9216 23480 9280
rect 23164 9215 23480 9216
rect 30754 9280 31070 9281
rect 30754 9216 30760 9280
rect 30824 9216 30840 9280
rect 30904 9216 30920 9280
rect 30984 9216 31000 9280
rect 31064 9216 31070 9280
rect 30754 9215 31070 9216
rect 11237 9210 11303 9213
rect 12157 9210 12223 9213
rect 11237 9208 12223 9210
rect 11237 9152 11242 9208
rect 11298 9152 12162 9208
rect 12218 9152 12223 9208
rect 11237 9150 12223 9152
rect 11237 9147 11303 9150
rect 12157 9147 12223 9150
rect 7465 9074 7531 9077
rect 8569 9074 8635 9077
rect 7465 9072 8635 9074
rect 7465 9016 7470 9072
rect 7526 9016 8574 9072
rect 8630 9016 8635 9072
rect 7465 9014 8635 9016
rect 7465 9011 7531 9014
rect 8569 9011 8635 9014
rect 5625 8938 5691 8941
rect 6913 8938 6979 8941
rect 5625 8936 6979 8938
rect 5625 8880 5630 8936
rect 5686 8880 6918 8936
rect 6974 8880 6979 8936
rect 5625 8878 6979 8880
rect 5625 8875 5691 8878
rect 6913 8875 6979 8878
rect 18505 8938 18571 8941
rect 27705 8938 27771 8941
rect 18505 8936 27771 8938
rect 18505 8880 18510 8936
rect 18566 8880 27710 8936
rect 27766 8880 27771 8936
rect 18505 8878 27771 8880
rect 18505 8875 18571 8878
rect 27705 8875 27771 8878
rect 4189 8736 4505 8737
rect 4189 8672 4195 8736
rect 4259 8672 4275 8736
rect 4339 8672 4355 8736
rect 4419 8672 4435 8736
rect 4499 8672 4505 8736
rect 4189 8671 4505 8672
rect 11779 8736 12095 8737
rect 11779 8672 11785 8736
rect 11849 8672 11865 8736
rect 11929 8672 11945 8736
rect 12009 8672 12025 8736
rect 12089 8672 12095 8736
rect 11779 8671 12095 8672
rect 19369 8736 19685 8737
rect 19369 8672 19375 8736
rect 19439 8672 19455 8736
rect 19519 8672 19535 8736
rect 19599 8672 19615 8736
rect 19679 8672 19685 8736
rect 19369 8671 19685 8672
rect 26959 8736 27275 8737
rect 26959 8672 26965 8736
rect 27029 8672 27045 8736
rect 27109 8672 27125 8736
rect 27189 8672 27205 8736
rect 27269 8672 27275 8736
rect 26959 8671 27275 8672
rect 5349 8666 5415 8669
rect 6913 8666 6979 8669
rect 5349 8664 6979 8666
rect 5349 8608 5354 8664
rect 5410 8608 6918 8664
rect 6974 8608 6979 8664
rect 5349 8606 6979 8608
rect 5349 8603 5415 8606
rect 6913 8603 6979 8606
rect 2589 8530 2655 8533
rect 8845 8530 8911 8533
rect 2589 8528 8911 8530
rect 2589 8472 2594 8528
rect 2650 8472 8850 8528
rect 8906 8472 8911 8528
rect 2589 8470 8911 8472
rect 2589 8467 2655 8470
rect 8845 8467 8911 8470
rect 7005 8394 7071 8397
rect 18045 8394 18111 8397
rect 7005 8392 18111 8394
rect 7005 8336 7010 8392
rect 7066 8336 18050 8392
rect 18106 8336 18111 8392
rect 7005 8334 18111 8336
rect 7005 8331 7071 8334
rect 18045 8331 18111 8334
rect 19241 8394 19307 8397
rect 25957 8394 26023 8397
rect 19241 8392 26023 8394
rect 19241 8336 19246 8392
rect 19302 8336 25962 8392
rect 26018 8336 26023 8392
rect 19241 8334 26023 8336
rect 19241 8331 19307 8334
rect 25957 8331 26023 8334
rect 2957 8258 3023 8261
rect 7649 8258 7715 8261
rect 2957 8256 7715 8258
rect 2957 8200 2962 8256
rect 3018 8200 7654 8256
rect 7710 8200 7715 8256
rect 2957 8198 7715 8200
rect 2957 8195 3023 8198
rect 7649 8195 7715 8198
rect 7984 8192 8300 8193
rect 7984 8128 7990 8192
rect 8054 8128 8070 8192
rect 8134 8128 8150 8192
rect 8214 8128 8230 8192
rect 8294 8128 8300 8192
rect 7984 8127 8300 8128
rect 15574 8192 15890 8193
rect 15574 8128 15580 8192
rect 15644 8128 15660 8192
rect 15724 8128 15740 8192
rect 15804 8128 15820 8192
rect 15884 8128 15890 8192
rect 15574 8127 15890 8128
rect 23164 8192 23480 8193
rect 23164 8128 23170 8192
rect 23234 8128 23250 8192
rect 23314 8128 23330 8192
rect 23394 8128 23410 8192
rect 23474 8128 23480 8192
rect 23164 8127 23480 8128
rect 30754 8192 31070 8193
rect 30754 8128 30760 8192
rect 30824 8128 30840 8192
rect 30904 8128 30920 8192
rect 30984 8128 31000 8192
rect 31064 8128 31070 8192
rect 30754 8127 31070 8128
rect 2037 8122 2103 8125
rect 6453 8122 6519 8125
rect 2037 8120 6519 8122
rect 2037 8064 2042 8120
rect 2098 8064 6458 8120
rect 6514 8064 6519 8120
rect 2037 8062 6519 8064
rect 2037 8059 2103 8062
rect 6453 8059 6519 8062
rect 3325 7986 3391 7989
rect 16113 7986 16179 7989
rect 3325 7984 16179 7986
rect 3325 7928 3330 7984
rect 3386 7928 16118 7984
rect 16174 7928 16179 7984
rect 3325 7926 16179 7928
rect 3325 7923 3391 7926
rect 16113 7923 16179 7926
rect 1025 7850 1091 7853
rect 3325 7850 3391 7853
rect 1025 7848 3391 7850
rect 1025 7792 1030 7848
rect 1086 7792 3330 7848
rect 3386 7792 3391 7848
rect 1025 7790 3391 7792
rect 1025 7787 1091 7790
rect 3325 7787 3391 7790
rect 8201 7850 8267 7853
rect 14457 7850 14523 7853
rect 8201 7848 14523 7850
rect 8201 7792 8206 7848
rect 8262 7792 14462 7848
rect 14518 7792 14523 7848
rect 8201 7790 14523 7792
rect 8201 7787 8267 7790
rect 14457 7787 14523 7790
rect 21357 7850 21423 7853
rect 25313 7850 25379 7853
rect 21357 7848 25379 7850
rect 21357 7792 21362 7848
rect 21418 7792 25318 7848
rect 25374 7792 25379 7848
rect 21357 7790 25379 7792
rect 21357 7787 21423 7790
rect 25313 7787 25379 7790
rect 9121 7714 9187 7717
rect 9581 7714 9647 7717
rect 9121 7712 9647 7714
rect 9121 7656 9126 7712
rect 9182 7656 9586 7712
rect 9642 7656 9647 7712
rect 9121 7654 9647 7656
rect 9121 7651 9187 7654
rect 9581 7651 9647 7654
rect 4189 7648 4505 7649
rect 4189 7584 4195 7648
rect 4259 7584 4275 7648
rect 4339 7584 4355 7648
rect 4419 7584 4435 7648
rect 4499 7584 4505 7648
rect 4189 7583 4505 7584
rect 11779 7648 12095 7649
rect 11779 7584 11785 7648
rect 11849 7584 11865 7648
rect 11929 7584 11945 7648
rect 12009 7584 12025 7648
rect 12089 7584 12095 7648
rect 11779 7583 12095 7584
rect 19369 7648 19685 7649
rect 19369 7584 19375 7648
rect 19439 7584 19455 7648
rect 19519 7584 19535 7648
rect 19599 7584 19615 7648
rect 19679 7584 19685 7648
rect 19369 7583 19685 7584
rect 26959 7648 27275 7649
rect 26959 7584 26965 7648
rect 27029 7584 27045 7648
rect 27109 7584 27125 7648
rect 27189 7584 27205 7648
rect 27269 7584 27275 7648
rect 26959 7583 27275 7584
rect 17953 7580 18019 7581
rect 17902 7578 17908 7580
rect 17862 7518 17908 7578
rect 17972 7576 18019 7580
rect 18014 7520 18019 7576
rect 17902 7516 17908 7518
rect 17972 7516 18019 7520
rect 17953 7515 18019 7516
rect 2957 7442 3023 7445
rect 6177 7442 6243 7445
rect 2957 7440 6243 7442
rect 2957 7384 2962 7440
rect 3018 7384 6182 7440
rect 6238 7384 6243 7440
rect 2957 7382 6243 7384
rect 2957 7379 3023 7382
rect 6177 7379 6243 7382
rect 6545 7442 6611 7445
rect 17953 7442 18019 7445
rect 6545 7440 18019 7442
rect 6545 7384 6550 7440
rect 6606 7384 17958 7440
rect 18014 7384 18019 7440
rect 6545 7382 18019 7384
rect 6545 7379 6611 7382
rect 17953 7379 18019 7382
rect 2773 7306 2839 7309
rect 6269 7306 6335 7309
rect 7557 7306 7623 7309
rect 2773 7304 2882 7306
rect 2773 7248 2778 7304
rect 2834 7248 2882 7304
rect 2773 7243 2882 7248
rect 6269 7304 7623 7306
rect 6269 7248 6274 7304
rect 6330 7248 7562 7304
rect 7618 7248 7623 7304
rect 6269 7246 7623 7248
rect 6269 7243 6335 7246
rect 7557 7243 7623 7246
rect 11145 7306 11211 7309
rect 12893 7306 12959 7309
rect 11145 7304 12959 7306
rect 11145 7248 11150 7304
rect 11206 7248 12898 7304
rect 12954 7248 12959 7304
rect 11145 7246 12959 7248
rect 11145 7243 11211 7246
rect 12893 7243 12959 7246
rect 13905 7306 13971 7309
rect 15101 7306 15167 7309
rect 13905 7304 15167 7306
rect 13905 7248 13910 7304
rect 13966 7248 15106 7304
rect 15162 7248 15167 7304
rect 13905 7246 15167 7248
rect 13905 7243 13971 7246
rect 15101 7243 15167 7246
rect 18597 7306 18663 7309
rect 20897 7306 20963 7309
rect 18597 7304 20963 7306
rect 18597 7248 18602 7304
rect 18658 7248 20902 7304
rect 20958 7248 20963 7304
rect 18597 7246 20963 7248
rect 18597 7243 18663 7246
rect 20897 7243 20963 7246
rect 2822 6898 2882 7243
rect 25129 7170 25195 7173
rect 26509 7170 26575 7173
rect 27245 7170 27311 7173
rect 25129 7168 27311 7170
rect 25129 7112 25134 7168
rect 25190 7112 26514 7168
rect 26570 7112 27250 7168
rect 27306 7112 27311 7168
rect 25129 7110 27311 7112
rect 25129 7107 25195 7110
rect 26509 7107 26575 7110
rect 27245 7107 27311 7110
rect 7984 7104 8300 7105
rect 7984 7040 7990 7104
rect 8054 7040 8070 7104
rect 8134 7040 8150 7104
rect 8214 7040 8230 7104
rect 8294 7040 8300 7104
rect 7984 7039 8300 7040
rect 15574 7104 15890 7105
rect 15574 7040 15580 7104
rect 15644 7040 15660 7104
rect 15724 7040 15740 7104
rect 15804 7040 15820 7104
rect 15884 7040 15890 7104
rect 15574 7039 15890 7040
rect 23164 7104 23480 7105
rect 23164 7040 23170 7104
rect 23234 7040 23250 7104
rect 23314 7040 23330 7104
rect 23394 7040 23410 7104
rect 23474 7040 23480 7104
rect 23164 7039 23480 7040
rect 30754 7104 31070 7105
rect 30754 7040 30760 7104
rect 30824 7040 30840 7104
rect 30904 7040 30920 7104
rect 30984 7040 31000 7104
rect 31064 7040 31070 7104
rect 30754 7039 31070 7040
rect 10225 7034 10291 7037
rect 13077 7034 13143 7037
rect 10225 7032 13143 7034
rect 10225 6976 10230 7032
rect 10286 6976 13082 7032
rect 13138 6976 13143 7032
rect 10225 6974 13143 6976
rect 10225 6971 10291 6974
rect 13077 6971 13143 6974
rect 13537 7034 13603 7037
rect 15285 7034 15351 7037
rect 13537 7032 15351 7034
rect 13537 6976 13542 7032
rect 13598 6976 15290 7032
rect 15346 6976 15351 7032
rect 13537 6974 15351 6976
rect 13537 6971 13603 6974
rect 15285 6971 15351 6974
rect 24025 7034 24091 7037
rect 25313 7034 25379 7037
rect 24025 7032 25379 7034
rect 24025 6976 24030 7032
rect 24086 6976 25318 7032
rect 25374 6976 25379 7032
rect 24025 6974 25379 6976
rect 24025 6971 24091 6974
rect 25313 6971 25379 6974
rect 2957 6898 3023 6901
rect 2822 6896 3023 6898
rect 2822 6840 2962 6896
rect 3018 6840 3023 6896
rect 2822 6838 3023 6840
rect 2957 6835 3023 6838
rect 4061 6898 4127 6901
rect 6913 6898 6979 6901
rect 4061 6896 6979 6898
rect 4061 6840 4066 6896
rect 4122 6840 6918 6896
rect 6974 6840 6979 6896
rect 4061 6838 6979 6840
rect 4061 6835 4127 6838
rect 6913 6835 6979 6838
rect 11513 6898 11579 6901
rect 16297 6898 16363 6901
rect 11513 6896 16363 6898
rect 11513 6840 11518 6896
rect 11574 6840 16302 6896
rect 16358 6840 16363 6896
rect 11513 6838 16363 6840
rect 11513 6835 11579 6838
rect 16297 6835 16363 6838
rect 20713 6898 20779 6901
rect 27889 6898 27955 6901
rect 20713 6896 27955 6898
rect 20713 6840 20718 6896
rect 20774 6840 27894 6896
rect 27950 6840 27955 6896
rect 20713 6838 27955 6840
rect 20713 6835 20779 6838
rect 27889 6835 27955 6838
rect 1761 6762 1827 6765
rect 10869 6762 10935 6765
rect 15745 6762 15811 6765
rect 1761 6760 10935 6762
rect 1761 6704 1766 6760
rect 1822 6704 10874 6760
rect 10930 6704 10935 6760
rect 1761 6702 10935 6704
rect 1761 6699 1827 6702
rect 10869 6699 10935 6702
rect 11654 6760 15811 6762
rect 11654 6704 15750 6760
rect 15806 6704 15811 6760
rect 11654 6702 15811 6704
rect 10501 6626 10567 6629
rect 11654 6626 11714 6702
rect 15745 6699 15811 6702
rect 16481 6762 16547 6765
rect 22645 6762 22711 6765
rect 25865 6762 25931 6765
rect 16481 6760 22110 6762
rect 16481 6704 16486 6760
rect 16542 6704 22110 6760
rect 16481 6702 22110 6704
rect 16481 6699 16547 6702
rect 10501 6624 11714 6626
rect 10501 6568 10506 6624
rect 10562 6568 11714 6624
rect 10501 6566 11714 6568
rect 13353 6626 13419 6629
rect 17033 6626 17099 6629
rect 13353 6624 17099 6626
rect 13353 6568 13358 6624
rect 13414 6568 17038 6624
rect 17094 6568 17099 6624
rect 13353 6566 17099 6568
rect 22050 6626 22110 6702
rect 22645 6760 25931 6762
rect 22645 6704 22650 6760
rect 22706 6704 25870 6760
rect 25926 6704 25931 6760
rect 22645 6702 25931 6704
rect 22645 6699 22711 6702
rect 25865 6699 25931 6702
rect 26509 6762 26575 6765
rect 28993 6762 29059 6765
rect 26509 6760 29059 6762
rect 26509 6704 26514 6760
rect 26570 6704 28998 6760
rect 29054 6704 29059 6760
rect 26509 6702 29059 6704
rect 26509 6699 26575 6702
rect 28993 6699 29059 6702
rect 26233 6626 26299 6629
rect 22050 6624 26299 6626
rect 22050 6568 26238 6624
rect 26294 6568 26299 6624
rect 22050 6566 26299 6568
rect 10501 6563 10567 6566
rect 13353 6563 13419 6566
rect 17033 6563 17099 6566
rect 26233 6563 26299 6566
rect 4189 6560 4505 6561
rect 4189 6496 4195 6560
rect 4259 6496 4275 6560
rect 4339 6496 4355 6560
rect 4419 6496 4435 6560
rect 4499 6496 4505 6560
rect 4189 6495 4505 6496
rect 11779 6560 12095 6561
rect 11779 6496 11785 6560
rect 11849 6496 11865 6560
rect 11929 6496 11945 6560
rect 12009 6496 12025 6560
rect 12089 6496 12095 6560
rect 11779 6495 12095 6496
rect 19369 6560 19685 6561
rect 19369 6496 19375 6560
rect 19439 6496 19455 6560
rect 19519 6496 19535 6560
rect 19599 6496 19615 6560
rect 19679 6496 19685 6560
rect 19369 6495 19685 6496
rect 26959 6560 27275 6561
rect 26959 6496 26965 6560
rect 27029 6496 27045 6560
rect 27109 6496 27125 6560
rect 27189 6496 27205 6560
rect 27269 6496 27275 6560
rect 26959 6495 27275 6496
rect 5349 6490 5415 6493
rect 11605 6490 11671 6493
rect 5349 6488 11671 6490
rect 5349 6432 5354 6488
rect 5410 6432 11610 6488
rect 11666 6432 11671 6488
rect 5349 6430 11671 6432
rect 5349 6427 5415 6430
rect 11605 6427 11671 6430
rect 15285 6490 15351 6493
rect 17493 6490 17559 6493
rect 15285 6488 17559 6490
rect 15285 6432 15290 6488
rect 15346 6432 17498 6488
rect 17554 6432 17559 6488
rect 15285 6430 17559 6432
rect 15285 6427 15351 6430
rect 17493 6427 17559 6430
rect 1710 6292 1716 6356
rect 1780 6354 1786 6356
rect 15929 6354 15995 6357
rect 16113 6354 16179 6357
rect 23381 6354 23447 6357
rect 1780 6352 15995 6354
rect 1780 6296 15934 6352
rect 15990 6296 15995 6352
rect 1780 6294 15995 6296
rect 1780 6292 1786 6294
rect 15929 6291 15995 6294
rect 16070 6352 23447 6354
rect 16070 6296 16118 6352
rect 16174 6296 23386 6352
rect 23442 6296 23447 6352
rect 16070 6294 23447 6296
rect 16070 6291 16179 6294
rect 23381 6291 23447 6294
rect 27061 6354 27127 6357
rect 28165 6354 28231 6357
rect 27061 6352 28231 6354
rect 27061 6296 27066 6352
rect 27122 6296 28170 6352
rect 28226 6296 28231 6352
rect 27061 6294 28231 6296
rect 27061 6291 27127 6294
rect 28165 6291 28231 6294
rect 4981 6218 5047 6221
rect 9121 6218 9187 6221
rect 11421 6218 11487 6221
rect 4981 6216 8586 6218
rect 4981 6160 4986 6216
rect 5042 6160 8586 6216
rect 4981 6158 8586 6160
rect 4981 6155 5047 6158
rect 1117 6082 1183 6085
rect 5533 6082 5599 6085
rect 1117 6080 5599 6082
rect 1117 6024 1122 6080
rect 1178 6024 5538 6080
rect 5594 6024 5599 6080
rect 1117 6022 5599 6024
rect 8526 6082 8586 6158
rect 9121 6216 11487 6218
rect 9121 6160 9126 6216
rect 9182 6160 11426 6216
rect 11482 6160 11487 6216
rect 9121 6158 11487 6160
rect 9121 6155 9187 6158
rect 11421 6155 11487 6158
rect 11605 6218 11671 6221
rect 16070 6218 16130 6291
rect 11605 6216 16130 6218
rect 11605 6160 11610 6216
rect 11666 6160 16130 6216
rect 11605 6158 16130 6160
rect 11605 6155 11671 6158
rect 10777 6082 10843 6085
rect 15285 6082 15351 6085
rect 8526 6022 9690 6082
rect 1117 6019 1183 6022
rect 5533 6019 5599 6022
rect 7984 6016 8300 6017
rect 7984 5952 7990 6016
rect 8054 5952 8070 6016
rect 8134 5952 8150 6016
rect 8214 5952 8230 6016
rect 8294 5952 8300 6016
rect 7984 5951 8300 5952
rect 9630 5946 9690 6022
rect 10777 6080 15351 6082
rect 10777 6024 10782 6080
rect 10838 6024 15290 6080
rect 15346 6024 15351 6080
rect 10777 6022 15351 6024
rect 10777 6019 10843 6022
rect 15285 6019 15351 6022
rect 15574 6016 15890 6017
rect 15574 5952 15580 6016
rect 15644 5952 15660 6016
rect 15724 5952 15740 6016
rect 15804 5952 15820 6016
rect 15884 5952 15890 6016
rect 15574 5951 15890 5952
rect 23164 6016 23480 6017
rect 23164 5952 23170 6016
rect 23234 5952 23250 6016
rect 23314 5952 23330 6016
rect 23394 5952 23410 6016
rect 23474 5952 23480 6016
rect 23164 5951 23480 5952
rect 30754 6016 31070 6017
rect 30754 5952 30760 6016
rect 30824 5952 30840 6016
rect 30904 5952 30920 6016
rect 30984 5952 31000 6016
rect 31064 5952 31070 6016
rect 30754 5951 31070 5952
rect 11697 5946 11763 5949
rect 9630 5944 11763 5946
rect 9630 5888 11702 5944
rect 11758 5888 11763 5944
rect 9630 5886 11763 5888
rect 11697 5883 11763 5886
rect 3417 5810 3483 5813
rect 6085 5810 6151 5813
rect 16205 5810 16271 5813
rect 3417 5808 16271 5810
rect 3417 5752 3422 5808
rect 3478 5752 6090 5808
rect 6146 5752 16210 5808
rect 16266 5752 16271 5808
rect 3417 5750 16271 5752
rect 3417 5747 3483 5750
rect 6085 5747 6151 5750
rect 16205 5747 16271 5750
rect 23381 5810 23447 5813
rect 24853 5810 24919 5813
rect 26969 5810 27035 5813
rect 23381 5808 27035 5810
rect 23381 5752 23386 5808
rect 23442 5752 24858 5808
rect 24914 5752 26974 5808
rect 27030 5752 27035 5808
rect 23381 5750 27035 5752
rect 23381 5747 23447 5750
rect 24853 5747 24919 5750
rect 26969 5747 27035 5750
rect 6453 5674 6519 5677
rect 13537 5674 13603 5677
rect 6453 5672 13603 5674
rect 6453 5616 6458 5672
rect 6514 5616 13542 5672
rect 13598 5616 13603 5672
rect 6453 5614 13603 5616
rect 6453 5611 6519 5614
rect 13537 5611 13603 5614
rect 22369 5674 22435 5677
rect 28165 5674 28231 5677
rect 22369 5672 28231 5674
rect 22369 5616 22374 5672
rect 22430 5616 28170 5672
rect 28226 5616 28231 5672
rect 22369 5614 28231 5616
rect 22369 5611 22435 5614
rect 28165 5611 28231 5614
rect 6678 5476 6684 5540
rect 6748 5538 6754 5540
rect 10317 5538 10383 5541
rect 6748 5536 10383 5538
rect 6748 5480 10322 5536
rect 10378 5480 10383 5536
rect 6748 5478 10383 5480
rect 6748 5476 6754 5478
rect 10317 5475 10383 5478
rect 4189 5472 4505 5473
rect 4189 5408 4195 5472
rect 4259 5408 4275 5472
rect 4339 5408 4355 5472
rect 4419 5408 4435 5472
rect 4499 5408 4505 5472
rect 4189 5407 4505 5408
rect 11779 5472 12095 5473
rect 11779 5408 11785 5472
rect 11849 5408 11865 5472
rect 11929 5408 11945 5472
rect 12009 5408 12025 5472
rect 12089 5408 12095 5472
rect 11779 5407 12095 5408
rect 19369 5472 19685 5473
rect 19369 5408 19375 5472
rect 19439 5408 19455 5472
rect 19519 5408 19535 5472
rect 19599 5408 19615 5472
rect 19679 5408 19685 5472
rect 19369 5407 19685 5408
rect 26959 5472 27275 5473
rect 26959 5408 26965 5472
rect 27029 5408 27045 5472
rect 27109 5408 27125 5472
rect 27189 5408 27205 5472
rect 27269 5408 27275 5472
rect 26959 5407 27275 5408
rect 5165 5402 5231 5405
rect 16021 5402 16087 5405
rect 5165 5400 11714 5402
rect 5165 5344 5170 5400
rect 5226 5344 11714 5400
rect 5165 5342 11714 5344
rect 5165 5339 5231 5342
rect 8845 5266 8911 5269
rect 10869 5266 10935 5269
rect 8845 5264 10935 5266
rect 8845 5208 8850 5264
rect 8906 5208 10874 5264
rect 10930 5208 10935 5264
rect 8845 5206 10935 5208
rect 11654 5266 11714 5342
rect 12206 5400 16087 5402
rect 12206 5344 16026 5400
rect 16082 5344 16087 5400
rect 12206 5342 16087 5344
rect 12206 5266 12266 5342
rect 16021 5339 16087 5342
rect 11654 5206 12266 5266
rect 17769 5266 17835 5269
rect 28625 5266 28691 5269
rect 17769 5264 28691 5266
rect 17769 5208 17774 5264
rect 17830 5208 28630 5264
rect 28686 5208 28691 5264
rect 17769 5206 28691 5208
rect 8845 5203 8911 5206
rect 10869 5203 10935 5206
rect 17769 5203 17835 5206
rect 28625 5203 28691 5206
rect 5533 5130 5599 5133
rect 6821 5130 6887 5133
rect 5533 5128 6887 5130
rect 5533 5072 5538 5128
rect 5594 5072 6826 5128
rect 6882 5072 6887 5128
rect 5533 5070 6887 5072
rect 5533 5067 5599 5070
rect 6821 5067 6887 5070
rect 17585 5130 17651 5133
rect 29361 5130 29427 5133
rect 17585 5128 29427 5130
rect 17585 5072 17590 5128
rect 17646 5072 29366 5128
rect 29422 5072 29427 5128
rect 17585 5070 29427 5072
rect 17585 5067 17651 5070
rect 29361 5067 29427 5070
rect 7984 4928 8300 4929
rect 7984 4864 7990 4928
rect 8054 4864 8070 4928
rect 8134 4864 8150 4928
rect 8214 4864 8230 4928
rect 8294 4864 8300 4928
rect 7984 4863 8300 4864
rect 15574 4928 15890 4929
rect 15574 4864 15580 4928
rect 15644 4864 15660 4928
rect 15724 4864 15740 4928
rect 15804 4864 15820 4928
rect 15884 4864 15890 4928
rect 15574 4863 15890 4864
rect 23164 4928 23480 4929
rect 23164 4864 23170 4928
rect 23234 4864 23250 4928
rect 23314 4864 23330 4928
rect 23394 4864 23410 4928
rect 23474 4864 23480 4928
rect 23164 4863 23480 4864
rect 30754 4928 31070 4929
rect 30754 4864 30760 4928
rect 30824 4864 30840 4928
rect 30904 4864 30920 4928
rect 30984 4864 31000 4928
rect 31064 4864 31070 4928
rect 30754 4863 31070 4864
rect 933 4722 999 4725
rect 3233 4722 3299 4725
rect 8753 4722 8819 4725
rect 933 4720 8819 4722
rect 933 4664 938 4720
rect 994 4664 3238 4720
rect 3294 4664 8758 4720
rect 8814 4664 8819 4720
rect 933 4662 8819 4664
rect 933 4659 999 4662
rect 3233 4659 3299 4662
rect 8753 4659 8819 4662
rect 17493 4722 17559 4725
rect 23790 4722 23796 4724
rect 17493 4720 23796 4722
rect 17493 4664 17498 4720
rect 17554 4664 23796 4720
rect 17493 4662 23796 4664
rect 17493 4659 17559 4662
rect 23790 4660 23796 4662
rect 23860 4660 23866 4724
rect 3233 4586 3299 4589
rect 7189 4586 7255 4589
rect 8201 4586 8267 4589
rect 3233 4584 8267 4586
rect 3233 4528 3238 4584
rect 3294 4528 7194 4584
rect 7250 4528 8206 4584
rect 8262 4528 8267 4584
rect 3233 4526 8267 4528
rect 3233 4523 3299 4526
rect 7189 4523 7255 4526
rect 8201 4523 8267 4526
rect 8661 4586 8727 4589
rect 15193 4586 15259 4589
rect 8661 4584 15259 4586
rect 8661 4528 8666 4584
rect 8722 4528 15198 4584
rect 15254 4528 15259 4584
rect 8661 4526 15259 4528
rect 8661 4523 8727 4526
rect 15193 4523 15259 4526
rect 21633 4586 21699 4589
rect 26601 4586 26667 4589
rect 21633 4584 26667 4586
rect 21633 4528 21638 4584
rect 21694 4528 26606 4584
rect 26662 4528 26667 4584
rect 21633 4526 26667 4528
rect 21633 4523 21699 4526
rect 26601 4523 26667 4526
rect 16297 4450 16363 4453
rect 19149 4450 19215 4453
rect 16297 4448 19215 4450
rect 16297 4392 16302 4448
rect 16358 4392 19154 4448
rect 19210 4392 19215 4448
rect 16297 4390 19215 4392
rect 16297 4387 16363 4390
rect 19149 4387 19215 4390
rect 4189 4384 4505 4385
rect 4189 4320 4195 4384
rect 4259 4320 4275 4384
rect 4339 4320 4355 4384
rect 4419 4320 4435 4384
rect 4499 4320 4505 4384
rect 4189 4319 4505 4320
rect 11779 4384 12095 4385
rect 11779 4320 11785 4384
rect 11849 4320 11865 4384
rect 11929 4320 11945 4384
rect 12009 4320 12025 4384
rect 12089 4320 12095 4384
rect 11779 4319 12095 4320
rect 19369 4384 19685 4385
rect 19369 4320 19375 4384
rect 19439 4320 19455 4384
rect 19519 4320 19535 4384
rect 19599 4320 19615 4384
rect 19679 4320 19685 4384
rect 19369 4319 19685 4320
rect 26959 4384 27275 4385
rect 26959 4320 26965 4384
rect 27029 4320 27045 4384
rect 27109 4320 27125 4384
rect 27189 4320 27205 4384
rect 27269 4320 27275 4384
rect 26959 4319 27275 4320
rect 12249 4314 12315 4317
rect 17902 4314 17908 4316
rect 12249 4312 17908 4314
rect 12249 4256 12254 4312
rect 12310 4256 17908 4312
rect 12249 4254 17908 4256
rect 12249 4251 12315 4254
rect 17902 4252 17908 4254
rect 17972 4252 17978 4316
rect 2681 4042 2747 4045
rect 3877 4042 3943 4045
rect 8569 4042 8635 4045
rect 2681 4040 8635 4042
rect 2681 3984 2686 4040
rect 2742 3984 3882 4040
rect 3938 3984 8574 4040
rect 8630 3984 8635 4040
rect 2681 3982 8635 3984
rect 2681 3979 2747 3982
rect 3877 3979 3943 3982
rect 8569 3979 8635 3982
rect 14917 4042 14983 4045
rect 28625 4042 28691 4045
rect 14917 4040 28691 4042
rect 14917 3984 14922 4040
rect 14978 3984 28630 4040
rect 28686 3984 28691 4040
rect 14917 3982 28691 3984
rect 14917 3979 14983 3982
rect 28625 3979 28691 3982
rect 3509 3906 3575 3909
rect 4705 3906 4771 3909
rect 3509 3904 4771 3906
rect 3509 3848 3514 3904
rect 3570 3848 4710 3904
rect 4766 3848 4771 3904
rect 3509 3846 4771 3848
rect 3509 3843 3575 3846
rect 4705 3843 4771 3846
rect 7984 3840 8300 3841
rect 7984 3776 7990 3840
rect 8054 3776 8070 3840
rect 8134 3776 8150 3840
rect 8214 3776 8230 3840
rect 8294 3776 8300 3840
rect 7984 3775 8300 3776
rect 15574 3840 15890 3841
rect 15574 3776 15580 3840
rect 15644 3776 15660 3840
rect 15724 3776 15740 3840
rect 15804 3776 15820 3840
rect 15884 3776 15890 3840
rect 15574 3775 15890 3776
rect 23164 3840 23480 3841
rect 23164 3776 23170 3840
rect 23234 3776 23250 3840
rect 23314 3776 23330 3840
rect 23394 3776 23410 3840
rect 23474 3776 23480 3840
rect 23164 3775 23480 3776
rect 30754 3840 31070 3841
rect 30754 3776 30760 3840
rect 30824 3776 30840 3840
rect 30904 3776 30920 3840
rect 30984 3776 31000 3840
rect 31064 3776 31070 3840
rect 30754 3775 31070 3776
rect 2221 3770 2287 3773
rect 2681 3770 2747 3773
rect 2221 3768 2747 3770
rect 2221 3712 2226 3768
rect 2282 3712 2686 3768
rect 2742 3712 2747 3768
rect 2221 3710 2747 3712
rect 2221 3707 2287 3710
rect 2681 3707 2747 3710
rect 3509 3770 3575 3773
rect 3969 3770 4035 3773
rect 5901 3770 5967 3773
rect 3509 3768 5967 3770
rect 3509 3712 3514 3768
rect 3570 3712 3974 3768
rect 4030 3712 5906 3768
rect 5962 3712 5967 3768
rect 3509 3710 5967 3712
rect 3509 3707 3575 3710
rect 3969 3707 4035 3710
rect 5901 3707 5967 3710
rect 3693 3634 3759 3637
rect 4981 3634 5047 3637
rect 6913 3634 6979 3637
rect 3693 3632 6979 3634
rect 3693 3576 3698 3632
rect 3754 3576 4986 3632
rect 5042 3576 6918 3632
rect 6974 3576 6979 3632
rect 3693 3574 6979 3576
rect 3693 3571 3759 3574
rect 4981 3571 5047 3574
rect 6913 3571 6979 3574
rect 3877 3498 3943 3501
rect 13905 3498 13971 3501
rect 3877 3496 13971 3498
rect 3877 3440 3882 3496
rect 3938 3440 13910 3496
rect 13966 3440 13971 3496
rect 3877 3438 13971 3440
rect 3877 3435 3943 3438
rect 13905 3435 13971 3438
rect 14089 3498 14155 3501
rect 14825 3498 14891 3501
rect 16757 3498 16823 3501
rect 27521 3498 27587 3501
rect 14089 3496 27587 3498
rect 14089 3440 14094 3496
rect 14150 3440 14830 3496
rect 14886 3440 16762 3496
rect 16818 3440 27526 3496
rect 27582 3440 27587 3496
rect 14089 3438 27587 3440
rect 14089 3435 14155 3438
rect 14825 3435 14891 3438
rect 16757 3435 16823 3438
rect 27521 3435 27587 3438
rect 4189 3296 4505 3297
rect 4189 3232 4195 3296
rect 4259 3232 4275 3296
rect 4339 3232 4355 3296
rect 4419 3232 4435 3296
rect 4499 3232 4505 3296
rect 4189 3231 4505 3232
rect 11779 3296 12095 3297
rect 11779 3232 11785 3296
rect 11849 3232 11865 3296
rect 11929 3232 11945 3296
rect 12009 3232 12025 3296
rect 12089 3232 12095 3296
rect 11779 3231 12095 3232
rect 19369 3296 19685 3297
rect 19369 3232 19375 3296
rect 19439 3232 19455 3296
rect 19519 3232 19535 3296
rect 19599 3232 19615 3296
rect 19679 3232 19685 3296
rect 19369 3231 19685 3232
rect 26959 3296 27275 3297
rect 26959 3232 26965 3296
rect 27029 3232 27045 3296
rect 27109 3232 27125 3296
rect 27189 3232 27205 3296
rect 27269 3232 27275 3296
rect 26959 3231 27275 3232
rect 4521 3090 4587 3093
rect 15142 3090 15148 3092
rect 4521 3088 15148 3090
rect 4521 3032 4526 3088
rect 4582 3032 15148 3088
rect 4521 3030 15148 3032
rect 4521 3027 4587 3030
rect 15142 3028 15148 3030
rect 15212 3028 15218 3092
rect 19701 3090 19767 3093
rect 26325 3090 26391 3093
rect 19701 3088 26391 3090
rect 19701 3032 19706 3088
rect 19762 3032 26330 3088
rect 26386 3032 26391 3088
rect 19701 3030 26391 3032
rect 19701 3027 19767 3030
rect 26325 3027 26391 3030
rect 5993 2954 6059 2957
rect 28349 2954 28415 2957
rect 5993 2952 28415 2954
rect 5993 2896 5998 2952
rect 6054 2896 28354 2952
rect 28410 2896 28415 2952
rect 5993 2894 28415 2896
rect 5993 2891 6059 2894
rect 28349 2891 28415 2894
rect 3693 2818 3759 2821
rect 6545 2818 6611 2821
rect 3693 2816 6611 2818
rect 3693 2760 3698 2816
rect 3754 2760 6550 2816
rect 6606 2760 6611 2816
rect 3693 2758 6611 2760
rect 3693 2755 3759 2758
rect 6545 2755 6611 2758
rect 10961 2818 11027 2821
rect 11789 2818 11855 2821
rect 10961 2816 11855 2818
rect 10961 2760 10966 2816
rect 11022 2760 11794 2816
rect 11850 2760 11855 2816
rect 10961 2758 11855 2760
rect 10961 2755 11027 2758
rect 11789 2755 11855 2758
rect 16297 2818 16363 2821
rect 21081 2818 21147 2821
rect 16297 2816 21147 2818
rect 16297 2760 16302 2816
rect 16358 2760 21086 2816
rect 21142 2760 21147 2816
rect 16297 2758 21147 2760
rect 16297 2755 16363 2758
rect 21081 2755 21147 2758
rect 7984 2752 8300 2753
rect 7984 2688 7990 2752
rect 8054 2688 8070 2752
rect 8134 2688 8150 2752
rect 8214 2688 8230 2752
rect 8294 2688 8300 2752
rect 7984 2687 8300 2688
rect 15574 2752 15890 2753
rect 15574 2688 15580 2752
rect 15644 2688 15660 2752
rect 15724 2688 15740 2752
rect 15804 2688 15820 2752
rect 15884 2688 15890 2752
rect 15574 2687 15890 2688
rect 23164 2752 23480 2753
rect 23164 2688 23170 2752
rect 23234 2688 23250 2752
rect 23314 2688 23330 2752
rect 23394 2688 23410 2752
rect 23474 2688 23480 2752
rect 23164 2687 23480 2688
rect 30754 2752 31070 2753
rect 30754 2688 30760 2752
rect 30824 2688 30840 2752
rect 30904 2688 30920 2752
rect 30984 2688 31000 2752
rect 31064 2688 31070 2752
rect 30754 2687 31070 2688
rect 3325 2682 3391 2685
rect 5993 2682 6059 2685
rect 3325 2680 6059 2682
rect 3325 2624 3330 2680
rect 3386 2624 5998 2680
rect 6054 2624 6059 2680
rect 3325 2622 6059 2624
rect 3325 2619 3391 2622
rect 5993 2619 6059 2622
rect 11421 2682 11487 2685
rect 12249 2682 12315 2685
rect 11421 2680 12315 2682
rect 11421 2624 11426 2680
rect 11482 2624 12254 2680
rect 12310 2624 12315 2680
rect 11421 2622 12315 2624
rect 11421 2619 11487 2622
rect 12249 2619 12315 2622
rect 4521 2546 4587 2549
rect 5165 2546 5231 2549
rect 4521 2544 5231 2546
rect 4521 2488 4526 2544
rect 4582 2488 5170 2544
rect 5226 2488 5231 2544
rect 4521 2486 5231 2488
rect 4521 2483 4587 2486
rect 5165 2483 5231 2486
rect 5349 2546 5415 2549
rect 24710 2546 24716 2548
rect 5349 2544 24716 2546
rect 5349 2488 5354 2544
rect 5410 2488 24716 2544
rect 5349 2486 24716 2488
rect 5349 2483 5415 2486
rect 24710 2484 24716 2486
rect 24780 2484 24786 2548
rect 11881 2410 11947 2413
rect 12433 2410 12499 2413
rect 11881 2408 12499 2410
rect 11881 2352 11886 2408
rect 11942 2352 12438 2408
rect 12494 2352 12499 2408
rect 11881 2350 12499 2352
rect 11881 2347 11947 2350
rect 12433 2347 12499 2350
rect 15142 2348 15148 2412
rect 15212 2410 15218 2412
rect 29085 2410 29151 2413
rect 15212 2408 29151 2410
rect 15212 2352 29090 2408
rect 29146 2352 29151 2408
rect 15212 2350 29151 2352
rect 15212 2348 15218 2350
rect 29085 2347 29151 2350
rect 20621 2274 20687 2277
rect 21909 2274 21975 2277
rect 20621 2272 21975 2274
rect 20621 2216 20626 2272
rect 20682 2216 21914 2272
rect 21970 2216 21975 2272
rect 20621 2214 21975 2216
rect 20621 2211 20687 2214
rect 21909 2211 21975 2214
rect 4189 2208 4505 2209
rect 4189 2144 4195 2208
rect 4259 2144 4275 2208
rect 4339 2144 4355 2208
rect 4419 2144 4435 2208
rect 4499 2144 4505 2208
rect 4189 2143 4505 2144
rect 11779 2208 12095 2209
rect 11779 2144 11785 2208
rect 11849 2144 11865 2208
rect 11929 2144 11945 2208
rect 12009 2144 12025 2208
rect 12089 2144 12095 2208
rect 11779 2143 12095 2144
rect 19369 2208 19685 2209
rect 19369 2144 19375 2208
rect 19439 2144 19455 2208
rect 19519 2144 19535 2208
rect 19599 2144 19615 2208
rect 19679 2144 19685 2208
rect 19369 2143 19685 2144
rect 26959 2208 27275 2209
rect 26959 2144 26965 2208
rect 27029 2144 27045 2208
rect 27109 2144 27125 2208
rect 27189 2144 27205 2208
rect 27269 2144 27275 2208
rect 26959 2143 27275 2144
rect 20897 2138 20963 2141
rect 25589 2138 25655 2141
rect 20897 2136 25655 2138
rect 20897 2080 20902 2136
rect 20958 2080 25594 2136
rect 25650 2080 25655 2136
rect 20897 2078 25655 2080
rect 20897 2075 20963 2078
rect 25589 2075 25655 2078
rect 4245 2002 4311 2005
rect 5533 2004 5599 2005
rect 5533 2002 5580 2004
rect 4245 2000 5274 2002
rect 4245 1944 4250 2000
rect 4306 1944 5274 2000
rect 4245 1942 5274 1944
rect 5488 2000 5580 2002
rect 5488 1944 5538 2000
rect 5488 1942 5580 1944
rect 4245 1939 4311 1942
rect 5214 1866 5274 1942
rect 5533 1940 5580 1942
rect 5644 1940 5650 2004
rect 29177 2002 29243 2005
rect 12390 2000 29243 2002
rect 12390 1944 29182 2000
rect 29238 1944 29243 2000
rect 12390 1942 29243 1944
rect 5533 1939 5599 1940
rect 12390 1866 12450 1942
rect 29177 1939 29243 1942
rect 5214 1806 12450 1866
rect 17953 1866 18019 1869
rect 19057 1866 19123 1869
rect 17953 1864 19123 1866
rect 17953 1808 17958 1864
rect 18014 1808 19062 1864
rect 19118 1808 19123 1864
rect 17953 1806 19123 1808
rect 17953 1803 18019 1806
rect 19057 1803 19123 1806
rect 20713 1866 20779 1869
rect 23289 1866 23355 1869
rect 26233 1866 26299 1869
rect 20713 1864 26299 1866
rect 20713 1808 20718 1864
rect 20774 1808 23294 1864
rect 23350 1808 26238 1864
rect 26294 1808 26299 1864
rect 20713 1806 26299 1808
rect 20713 1803 20779 1806
rect 23289 1803 23355 1806
rect 26233 1803 26299 1806
rect 4613 1730 4679 1733
rect 6545 1730 6611 1733
rect 4613 1728 6611 1730
rect 4613 1672 4618 1728
rect 4674 1672 6550 1728
rect 6606 1672 6611 1728
rect 4613 1670 6611 1672
rect 4613 1667 4679 1670
rect 6545 1667 6611 1670
rect 7984 1664 8300 1665
rect 7984 1600 7990 1664
rect 8054 1600 8070 1664
rect 8134 1600 8150 1664
rect 8214 1600 8230 1664
rect 8294 1600 8300 1664
rect 7984 1599 8300 1600
rect 15574 1664 15890 1665
rect 15574 1600 15580 1664
rect 15644 1600 15660 1664
rect 15724 1600 15740 1664
rect 15804 1600 15820 1664
rect 15884 1600 15890 1664
rect 15574 1599 15890 1600
rect 23164 1664 23480 1665
rect 23164 1600 23170 1664
rect 23234 1600 23250 1664
rect 23314 1600 23330 1664
rect 23394 1600 23410 1664
rect 23474 1600 23480 1664
rect 23164 1599 23480 1600
rect 30754 1664 31070 1665
rect 30754 1600 30760 1664
rect 30824 1600 30840 1664
rect 30904 1600 30920 1664
rect 30984 1600 31000 1664
rect 31064 1600 31070 1664
rect 30754 1599 31070 1600
rect 1117 1458 1183 1461
rect 5165 1458 5231 1461
rect 1117 1456 5231 1458
rect 1117 1400 1122 1456
rect 1178 1400 5170 1456
rect 5226 1400 5231 1456
rect 1117 1398 5231 1400
rect 1117 1395 1183 1398
rect 5165 1395 5231 1398
rect 19425 1458 19491 1461
rect 25589 1458 25655 1461
rect 19425 1456 25655 1458
rect 19425 1400 19430 1456
rect 19486 1400 25594 1456
rect 25650 1400 25655 1456
rect 19425 1398 25655 1400
rect 19425 1395 19491 1398
rect 25589 1395 25655 1398
rect 4061 1322 4127 1325
rect 6729 1324 6795 1325
rect 4061 1320 6562 1322
rect 4061 1264 4066 1320
rect 4122 1264 6562 1320
rect 4061 1262 6562 1264
rect 4061 1259 4127 1262
rect 6502 1186 6562 1262
rect 6678 1260 6684 1324
rect 6748 1322 6795 1324
rect 18229 1322 18295 1325
rect 6748 1320 6840 1322
rect 6790 1264 6840 1320
rect 6748 1262 6840 1264
rect 8158 1320 18295 1322
rect 8158 1264 18234 1320
rect 18290 1264 18295 1320
rect 8158 1262 18295 1264
rect 6748 1260 6795 1262
rect 6729 1259 6795 1260
rect 8158 1186 8218 1262
rect 18229 1259 18295 1262
rect 18873 1322 18939 1325
rect 25681 1322 25747 1325
rect 29453 1322 29519 1325
rect 18873 1320 25747 1322
rect 18873 1264 18878 1320
rect 18934 1264 25686 1320
rect 25742 1264 25747 1320
rect 18873 1262 25747 1264
rect 18873 1259 18939 1262
rect 25681 1259 25747 1262
rect 25822 1320 29519 1322
rect 25822 1264 29458 1320
rect 29514 1264 29519 1320
rect 25822 1262 29519 1264
rect 6502 1126 8218 1186
rect 8293 1186 8359 1189
rect 9305 1186 9371 1189
rect 8293 1184 9371 1186
rect 8293 1128 8298 1184
rect 8354 1128 9310 1184
rect 9366 1128 9371 1184
rect 8293 1126 9371 1128
rect 8293 1123 8359 1126
rect 9305 1123 9371 1126
rect 23790 1124 23796 1188
rect 23860 1186 23866 1188
rect 25822 1186 25882 1262
rect 29453 1259 29519 1262
rect 23860 1126 25882 1186
rect 23860 1124 23866 1126
rect 4189 1120 4505 1121
rect 4189 1056 4195 1120
rect 4259 1056 4275 1120
rect 4339 1056 4355 1120
rect 4419 1056 4435 1120
rect 4499 1056 4505 1120
rect 4189 1055 4505 1056
rect 11779 1120 12095 1121
rect 11779 1056 11785 1120
rect 11849 1056 11865 1120
rect 11929 1056 11945 1120
rect 12009 1056 12025 1120
rect 12089 1056 12095 1120
rect 11779 1055 12095 1056
rect 19369 1120 19685 1121
rect 19369 1056 19375 1120
rect 19439 1056 19455 1120
rect 19519 1056 19535 1120
rect 19599 1056 19615 1120
rect 19679 1056 19685 1120
rect 19369 1055 19685 1056
rect 26959 1120 27275 1121
rect 26959 1056 26965 1120
rect 27029 1056 27045 1120
rect 27109 1056 27125 1120
rect 27189 1056 27205 1120
rect 27269 1056 27275 1120
rect 26959 1055 27275 1056
rect 6637 1050 6703 1053
rect 11421 1050 11487 1053
rect 6637 1048 11487 1050
rect 6637 992 6642 1048
rect 6698 992 11426 1048
rect 11482 992 11487 1048
rect 6637 990 11487 992
rect 6637 987 6703 990
rect 11421 987 11487 990
rect 20713 1050 20779 1053
rect 25681 1050 25747 1053
rect 20713 1048 25747 1050
rect 20713 992 20718 1048
rect 20774 992 25686 1048
rect 25742 992 25747 1048
rect 20713 990 25747 992
rect 20713 987 20779 990
rect 25681 987 25747 990
rect 11789 914 11855 917
rect 23473 914 23539 917
rect 11789 912 23539 914
rect 11789 856 11794 912
rect 11850 856 23478 912
rect 23534 856 23539 912
rect 11789 854 23539 856
rect 11789 851 11855 854
rect 23473 851 23539 854
rect 24710 852 24716 916
rect 24780 852 24786 916
rect 22001 778 22067 781
rect 23933 778 23999 781
rect 22001 776 23999 778
rect 22001 720 22006 776
rect 22062 720 23938 776
rect 23994 720 23999 776
rect 22001 718 23999 720
rect 24718 778 24778 852
rect 28993 778 29059 781
rect 24718 776 29059 778
rect 24718 720 28998 776
rect 29054 720 29059 776
rect 24718 718 29059 720
rect 22001 715 22067 718
rect 23933 715 23999 718
rect 28993 715 29059 718
rect 7984 576 8300 577
rect 7984 512 7990 576
rect 8054 512 8070 576
rect 8134 512 8150 576
rect 8214 512 8230 576
rect 8294 512 8300 576
rect 7984 511 8300 512
rect 15574 576 15890 577
rect 15574 512 15580 576
rect 15644 512 15660 576
rect 15724 512 15740 576
rect 15804 512 15820 576
rect 15884 512 15890 576
rect 15574 511 15890 512
rect 23164 576 23480 577
rect 23164 512 23170 576
rect 23234 512 23250 576
rect 23314 512 23330 576
rect 23394 512 23410 576
rect 23474 512 23480 576
rect 23164 511 23480 512
rect 30754 576 31070 577
rect 30754 512 30760 576
rect 30824 512 30840 576
rect 30904 512 30920 576
rect 30984 512 31000 576
rect 31064 512 31070 576
rect 30754 511 31070 512
rect 4245 370 4311 373
rect 29913 370 29979 373
rect 4245 368 29979 370
rect 4245 312 4250 368
rect 4306 312 29918 368
rect 29974 312 29979 368
rect 4245 310 29979 312
rect 4245 307 4311 310
rect 29913 307 29979 310
<< via3 >>
rect 10180 22068 10244 22132
rect 14412 22068 14476 22132
rect 8708 21932 8772 21996
rect 12572 21932 12636 21996
rect 13860 21992 13924 21996
rect 13860 21936 13874 21992
rect 13874 21936 13924 21992
rect 13860 21932 13924 21936
rect 9260 21796 9324 21860
rect 23612 21856 23676 21860
rect 23612 21800 23626 21856
rect 23626 21800 23676 21856
rect 23612 21796 23676 21800
rect 4195 21788 4259 21792
rect 4195 21732 4199 21788
rect 4199 21732 4255 21788
rect 4255 21732 4259 21788
rect 4195 21728 4259 21732
rect 4275 21788 4339 21792
rect 4275 21732 4279 21788
rect 4279 21732 4335 21788
rect 4335 21732 4339 21788
rect 4275 21728 4339 21732
rect 4355 21788 4419 21792
rect 4355 21732 4359 21788
rect 4359 21732 4415 21788
rect 4415 21732 4419 21788
rect 4355 21728 4419 21732
rect 4435 21788 4499 21792
rect 4435 21732 4439 21788
rect 4439 21732 4495 21788
rect 4495 21732 4499 21788
rect 4435 21728 4499 21732
rect 11785 21788 11849 21792
rect 11785 21732 11789 21788
rect 11789 21732 11845 21788
rect 11845 21732 11849 21788
rect 11785 21728 11849 21732
rect 11865 21788 11929 21792
rect 11865 21732 11869 21788
rect 11869 21732 11925 21788
rect 11925 21732 11929 21788
rect 11865 21728 11929 21732
rect 11945 21788 12009 21792
rect 11945 21732 11949 21788
rect 11949 21732 12005 21788
rect 12005 21732 12009 21788
rect 11945 21728 12009 21732
rect 12025 21788 12089 21792
rect 12025 21732 12029 21788
rect 12029 21732 12085 21788
rect 12085 21732 12089 21788
rect 12025 21728 12089 21732
rect 19375 21788 19439 21792
rect 19375 21732 19379 21788
rect 19379 21732 19435 21788
rect 19435 21732 19439 21788
rect 19375 21728 19439 21732
rect 19455 21788 19519 21792
rect 19455 21732 19459 21788
rect 19459 21732 19515 21788
rect 19515 21732 19519 21788
rect 19455 21728 19519 21732
rect 19535 21788 19599 21792
rect 19535 21732 19539 21788
rect 19539 21732 19595 21788
rect 19595 21732 19599 21788
rect 19535 21728 19599 21732
rect 19615 21788 19679 21792
rect 19615 21732 19619 21788
rect 19619 21732 19675 21788
rect 19675 21732 19679 21788
rect 19615 21728 19679 21732
rect 26965 21788 27029 21792
rect 26965 21732 26969 21788
rect 26969 21732 27025 21788
rect 27025 21732 27029 21788
rect 26965 21728 27029 21732
rect 27045 21788 27109 21792
rect 27045 21732 27049 21788
rect 27049 21732 27105 21788
rect 27105 21732 27109 21788
rect 27045 21728 27109 21732
rect 27125 21788 27189 21792
rect 27125 21732 27129 21788
rect 27129 21732 27185 21788
rect 27185 21732 27189 21788
rect 27125 21728 27189 21732
rect 27205 21788 27269 21792
rect 27205 21732 27209 21788
rect 27209 21732 27265 21788
rect 27265 21732 27269 21788
rect 27205 21728 27269 21732
rect 11468 21524 11532 21588
rect 12204 21584 12268 21588
rect 12204 21528 12254 21584
rect 12254 21528 12268 21584
rect 12204 21524 12268 21528
rect 16988 21524 17052 21588
rect 13124 21252 13188 21316
rect 7990 21244 8054 21248
rect 7990 21188 7994 21244
rect 7994 21188 8050 21244
rect 8050 21188 8054 21244
rect 7990 21184 8054 21188
rect 8070 21244 8134 21248
rect 8070 21188 8074 21244
rect 8074 21188 8130 21244
rect 8130 21188 8134 21244
rect 8070 21184 8134 21188
rect 8150 21244 8214 21248
rect 8150 21188 8154 21244
rect 8154 21188 8210 21244
rect 8210 21188 8214 21244
rect 8150 21184 8214 21188
rect 8230 21244 8294 21248
rect 8230 21188 8234 21244
rect 8234 21188 8290 21244
rect 8290 21188 8294 21244
rect 8230 21184 8294 21188
rect 15580 21244 15644 21248
rect 15580 21188 15584 21244
rect 15584 21188 15640 21244
rect 15640 21188 15644 21244
rect 15580 21184 15644 21188
rect 15660 21244 15724 21248
rect 15660 21188 15664 21244
rect 15664 21188 15720 21244
rect 15720 21188 15724 21244
rect 15660 21184 15724 21188
rect 15740 21244 15804 21248
rect 15740 21188 15744 21244
rect 15744 21188 15800 21244
rect 15800 21188 15804 21244
rect 15740 21184 15804 21188
rect 15820 21244 15884 21248
rect 15820 21188 15824 21244
rect 15824 21188 15880 21244
rect 15880 21188 15884 21244
rect 15820 21184 15884 21188
rect 23170 21244 23234 21248
rect 23170 21188 23174 21244
rect 23174 21188 23230 21244
rect 23230 21188 23234 21244
rect 23170 21184 23234 21188
rect 23250 21244 23314 21248
rect 23250 21188 23254 21244
rect 23254 21188 23310 21244
rect 23310 21188 23314 21244
rect 23250 21184 23314 21188
rect 23330 21244 23394 21248
rect 23330 21188 23334 21244
rect 23334 21188 23390 21244
rect 23390 21188 23394 21244
rect 23330 21184 23394 21188
rect 23410 21244 23474 21248
rect 23410 21188 23414 21244
rect 23414 21188 23470 21244
rect 23470 21188 23474 21244
rect 23410 21184 23474 21188
rect 30760 21244 30824 21248
rect 30760 21188 30764 21244
rect 30764 21188 30820 21244
rect 30820 21188 30824 21244
rect 30760 21184 30824 21188
rect 30840 21244 30904 21248
rect 30840 21188 30844 21244
rect 30844 21188 30900 21244
rect 30900 21188 30904 21244
rect 30840 21184 30904 21188
rect 30920 21244 30984 21248
rect 30920 21188 30924 21244
rect 30924 21188 30980 21244
rect 30980 21188 30984 21244
rect 30920 21184 30984 21188
rect 31000 21244 31064 21248
rect 31000 21188 31004 21244
rect 31004 21188 31060 21244
rect 31060 21188 31064 21244
rect 31000 21184 31064 21188
rect 11284 21116 11348 21180
rect 26372 21116 26436 21180
rect 11100 20844 11164 20908
rect 23612 20844 23676 20908
rect 8892 20708 8956 20772
rect 4195 20700 4259 20704
rect 4195 20644 4199 20700
rect 4199 20644 4255 20700
rect 4255 20644 4259 20700
rect 4195 20640 4259 20644
rect 4275 20700 4339 20704
rect 4275 20644 4279 20700
rect 4279 20644 4335 20700
rect 4335 20644 4339 20700
rect 4275 20640 4339 20644
rect 4355 20700 4419 20704
rect 4355 20644 4359 20700
rect 4359 20644 4415 20700
rect 4415 20644 4419 20700
rect 4355 20640 4419 20644
rect 4435 20700 4499 20704
rect 4435 20644 4439 20700
rect 4439 20644 4495 20700
rect 4495 20644 4499 20700
rect 4435 20640 4499 20644
rect 11785 20700 11849 20704
rect 11785 20644 11789 20700
rect 11789 20644 11845 20700
rect 11845 20644 11849 20700
rect 11785 20640 11849 20644
rect 11865 20700 11929 20704
rect 11865 20644 11869 20700
rect 11869 20644 11925 20700
rect 11925 20644 11929 20700
rect 11865 20640 11929 20644
rect 11945 20700 12009 20704
rect 11945 20644 11949 20700
rect 11949 20644 12005 20700
rect 12005 20644 12009 20700
rect 11945 20640 12009 20644
rect 12025 20700 12089 20704
rect 12025 20644 12029 20700
rect 12029 20644 12085 20700
rect 12085 20644 12089 20700
rect 12025 20640 12089 20644
rect 19375 20700 19439 20704
rect 19375 20644 19379 20700
rect 19379 20644 19435 20700
rect 19435 20644 19439 20700
rect 19375 20640 19439 20644
rect 19455 20700 19519 20704
rect 19455 20644 19459 20700
rect 19459 20644 19515 20700
rect 19515 20644 19519 20700
rect 19455 20640 19519 20644
rect 19535 20700 19599 20704
rect 19535 20644 19539 20700
rect 19539 20644 19595 20700
rect 19595 20644 19599 20700
rect 19535 20640 19599 20644
rect 19615 20700 19679 20704
rect 19615 20644 19619 20700
rect 19619 20644 19675 20700
rect 19675 20644 19679 20700
rect 19615 20640 19679 20644
rect 26965 20700 27029 20704
rect 26965 20644 26969 20700
rect 26969 20644 27025 20700
rect 27025 20644 27029 20700
rect 26965 20640 27029 20644
rect 27045 20700 27109 20704
rect 27045 20644 27049 20700
rect 27049 20644 27105 20700
rect 27105 20644 27109 20700
rect 27045 20640 27109 20644
rect 27125 20700 27189 20704
rect 27125 20644 27129 20700
rect 27129 20644 27185 20700
rect 27185 20644 27189 20700
rect 27125 20640 27189 20644
rect 27205 20700 27269 20704
rect 27205 20644 27209 20700
rect 27209 20644 27265 20700
rect 27265 20644 27269 20700
rect 27205 20640 27269 20644
rect 10916 20632 10980 20636
rect 10916 20576 10966 20632
rect 10966 20576 10980 20632
rect 10916 20572 10980 20576
rect 13676 20572 13740 20636
rect 9812 20436 9876 20500
rect 16068 20436 16132 20500
rect 7990 20156 8054 20160
rect 7990 20100 7994 20156
rect 7994 20100 8050 20156
rect 8050 20100 8054 20156
rect 7990 20096 8054 20100
rect 8070 20156 8134 20160
rect 8070 20100 8074 20156
rect 8074 20100 8130 20156
rect 8130 20100 8134 20156
rect 8070 20096 8134 20100
rect 8150 20156 8214 20160
rect 8150 20100 8154 20156
rect 8154 20100 8210 20156
rect 8210 20100 8214 20156
rect 8150 20096 8214 20100
rect 8230 20156 8294 20160
rect 8230 20100 8234 20156
rect 8234 20100 8290 20156
rect 8290 20100 8294 20156
rect 8230 20096 8294 20100
rect 15580 20156 15644 20160
rect 15580 20100 15584 20156
rect 15584 20100 15640 20156
rect 15640 20100 15644 20156
rect 15580 20096 15644 20100
rect 15660 20156 15724 20160
rect 15660 20100 15664 20156
rect 15664 20100 15720 20156
rect 15720 20100 15724 20156
rect 15660 20096 15724 20100
rect 15740 20156 15804 20160
rect 15740 20100 15744 20156
rect 15744 20100 15800 20156
rect 15800 20100 15804 20156
rect 15740 20096 15804 20100
rect 15820 20156 15884 20160
rect 15820 20100 15824 20156
rect 15824 20100 15880 20156
rect 15880 20100 15884 20156
rect 15820 20096 15884 20100
rect 23170 20156 23234 20160
rect 23170 20100 23174 20156
rect 23174 20100 23230 20156
rect 23230 20100 23234 20156
rect 23170 20096 23234 20100
rect 23250 20156 23314 20160
rect 23250 20100 23254 20156
rect 23254 20100 23310 20156
rect 23310 20100 23314 20156
rect 23250 20096 23314 20100
rect 23330 20156 23394 20160
rect 23330 20100 23334 20156
rect 23334 20100 23390 20156
rect 23390 20100 23394 20156
rect 23330 20096 23394 20100
rect 23410 20156 23474 20160
rect 23410 20100 23414 20156
rect 23414 20100 23470 20156
rect 23470 20100 23474 20156
rect 23410 20096 23474 20100
rect 30760 20156 30824 20160
rect 30760 20100 30764 20156
rect 30764 20100 30820 20156
rect 30820 20100 30824 20156
rect 30760 20096 30824 20100
rect 30840 20156 30904 20160
rect 30840 20100 30844 20156
rect 30844 20100 30900 20156
rect 30900 20100 30904 20156
rect 30840 20096 30904 20100
rect 30920 20156 30984 20160
rect 30920 20100 30924 20156
rect 30924 20100 30980 20156
rect 30980 20100 30984 20156
rect 30920 20096 30984 20100
rect 31000 20156 31064 20160
rect 31000 20100 31004 20156
rect 31004 20100 31060 20156
rect 31060 20100 31064 20156
rect 31000 20096 31064 20100
rect 4195 19612 4259 19616
rect 4195 19556 4199 19612
rect 4199 19556 4255 19612
rect 4255 19556 4259 19612
rect 4195 19552 4259 19556
rect 4275 19612 4339 19616
rect 4275 19556 4279 19612
rect 4279 19556 4335 19612
rect 4335 19556 4339 19612
rect 4275 19552 4339 19556
rect 4355 19612 4419 19616
rect 4355 19556 4359 19612
rect 4359 19556 4415 19612
rect 4415 19556 4419 19612
rect 4355 19552 4419 19556
rect 4435 19612 4499 19616
rect 4435 19556 4439 19612
rect 4439 19556 4495 19612
rect 4495 19556 4499 19612
rect 4435 19552 4499 19556
rect 11785 19612 11849 19616
rect 11785 19556 11789 19612
rect 11789 19556 11845 19612
rect 11845 19556 11849 19612
rect 11785 19552 11849 19556
rect 11865 19612 11929 19616
rect 11865 19556 11869 19612
rect 11869 19556 11925 19612
rect 11925 19556 11929 19612
rect 11865 19552 11929 19556
rect 11945 19612 12009 19616
rect 11945 19556 11949 19612
rect 11949 19556 12005 19612
rect 12005 19556 12009 19612
rect 11945 19552 12009 19556
rect 12025 19612 12089 19616
rect 12025 19556 12029 19612
rect 12029 19556 12085 19612
rect 12085 19556 12089 19612
rect 12025 19552 12089 19556
rect 19375 19612 19439 19616
rect 19375 19556 19379 19612
rect 19379 19556 19435 19612
rect 19435 19556 19439 19612
rect 19375 19552 19439 19556
rect 19455 19612 19519 19616
rect 19455 19556 19459 19612
rect 19459 19556 19515 19612
rect 19515 19556 19519 19612
rect 19455 19552 19519 19556
rect 19535 19612 19599 19616
rect 19535 19556 19539 19612
rect 19539 19556 19595 19612
rect 19595 19556 19599 19612
rect 19535 19552 19599 19556
rect 19615 19612 19679 19616
rect 19615 19556 19619 19612
rect 19619 19556 19675 19612
rect 19675 19556 19679 19612
rect 19615 19552 19679 19556
rect 26965 19612 27029 19616
rect 26965 19556 26969 19612
rect 26969 19556 27025 19612
rect 27025 19556 27029 19612
rect 26965 19552 27029 19556
rect 27045 19612 27109 19616
rect 27045 19556 27049 19612
rect 27049 19556 27105 19612
rect 27105 19556 27109 19612
rect 27045 19552 27109 19556
rect 27125 19612 27189 19616
rect 27125 19556 27129 19612
rect 27129 19556 27185 19612
rect 27185 19556 27189 19612
rect 27125 19552 27189 19556
rect 27205 19612 27269 19616
rect 27205 19556 27209 19612
rect 27209 19556 27265 19612
rect 27265 19556 27269 19612
rect 27205 19552 27269 19556
rect 6684 19348 6748 19412
rect 15332 19212 15396 19276
rect 16436 19272 16500 19276
rect 16436 19216 16486 19272
rect 16486 19216 16500 19272
rect 16436 19212 16500 19216
rect 7990 19068 8054 19072
rect 7990 19012 7994 19068
rect 7994 19012 8050 19068
rect 8050 19012 8054 19068
rect 7990 19008 8054 19012
rect 8070 19068 8134 19072
rect 8070 19012 8074 19068
rect 8074 19012 8130 19068
rect 8130 19012 8134 19068
rect 8070 19008 8134 19012
rect 8150 19068 8214 19072
rect 8150 19012 8154 19068
rect 8154 19012 8210 19068
rect 8210 19012 8214 19068
rect 8150 19008 8214 19012
rect 8230 19068 8294 19072
rect 8230 19012 8234 19068
rect 8234 19012 8290 19068
rect 8290 19012 8294 19068
rect 8230 19008 8294 19012
rect 15580 19068 15644 19072
rect 15580 19012 15584 19068
rect 15584 19012 15640 19068
rect 15640 19012 15644 19068
rect 15580 19008 15644 19012
rect 15660 19068 15724 19072
rect 15660 19012 15664 19068
rect 15664 19012 15720 19068
rect 15720 19012 15724 19068
rect 15660 19008 15724 19012
rect 15740 19068 15804 19072
rect 15740 19012 15744 19068
rect 15744 19012 15800 19068
rect 15800 19012 15804 19068
rect 15740 19008 15804 19012
rect 15820 19068 15884 19072
rect 15820 19012 15824 19068
rect 15824 19012 15880 19068
rect 15880 19012 15884 19068
rect 15820 19008 15884 19012
rect 23170 19068 23234 19072
rect 23170 19012 23174 19068
rect 23174 19012 23230 19068
rect 23230 19012 23234 19068
rect 23170 19008 23234 19012
rect 23250 19068 23314 19072
rect 23250 19012 23254 19068
rect 23254 19012 23310 19068
rect 23310 19012 23314 19068
rect 23250 19008 23314 19012
rect 23330 19068 23394 19072
rect 23330 19012 23334 19068
rect 23334 19012 23390 19068
rect 23390 19012 23394 19068
rect 23330 19008 23394 19012
rect 23410 19068 23474 19072
rect 23410 19012 23414 19068
rect 23414 19012 23470 19068
rect 23470 19012 23474 19068
rect 23410 19008 23474 19012
rect 30760 19068 30824 19072
rect 30760 19012 30764 19068
rect 30764 19012 30820 19068
rect 30820 19012 30824 19068
rect 30760 19008 30824 19012
rect 30840 19068 30904 19072
rect 30840 19012 30844 19068
rect 30844 19012 30900 19068
rect 30900 19012 30904 19068
rect 30840 19008 30904 19012
rect 30920 19068 30984 19072
rect 30920 19012 30924 19068
rect 30924 19012 30980 19068
rect 30980 19012 30984 19068
rect 30920 19008 30984 19012
rect 31000 19068 31064 19072
rect 31000 19012 31004 19068
rect 31004 19012 31060 19068
rect 31060 19012 31064 19068
rect 31000 19008 31064 19012
rect 3740 18940 3804 19004
rect 10364 18668 10428 18732
rect 24716 18804 24780 18868
rect 25268 18668 25332 18732
rect 4195 18524 4259 18528
rect 4195 18468 4199 18524
rect 4199 18468 4255 18524
rect 4255 18468 4259 18524
rect 4195 18464 4259 18468
rect 4275 18524 4339 18528
rect 4275 18468 4279 18524
rect 4279 18468 4335 18524
rect 4335 18468 4339 18524
rect 4275 18464 4339 18468
rect 4355 18524 4419 18528
rect 4355 18468 4359 18524
rect 4359 18468 4415 18524
rect 4415 18468 4419 18524
rect 4355 18464 4419 18468
rect 4435 18524 4499 18528
rect 4435 18468 4439 18524
rect 4439 18468 4495 18524
rect 4495 18468 4499 18524
rect 4435 18464 4499 18468
rect 7788 18592 7852 18596
rect 7788 18536 7802 18592
rect 7802 18536 7852 18592
rect 7788 18532 7852 18536
rect 26188 18532 26252 18596
rect 11785 18524 11849 18528
rect 11785 18468 11789 18524
rect 11789 18468 11845 18524
rect 11845 18468 11849 18524
rect 11785 18464 11849 18468
rect 11865 18524 11929 18528
rect 11865 18468 11869 18524
rect 11869 18468 11925 18524
rect 11925 18468 11929 18524
rect 11865 18464 11929 18468
rect 11945 18524 12009 18528
rect 11945 18468 11949 18524
rect 11949 18468 12005 18524
rect 12005 18468 12009 18524
rect 11945 18464 12009 18468
rect 12025 18524 12089 18528
rect 12025 18468 12029 18524
rect 12029 18468 12085 18524
rect 12085 18468 12089 18524
rect 12025 18464 12089 18468
rect 19375 18524 19439 18528
rect 19375 18468 19379 18524
rect 19379 18468 19435 18524
rect 19435 18468 19439 18524
rect 19375 18464 19439 18468
rect 19455 18524 19519 18528
rect 19455 18468 19459 18524
rect 19459 18468 19515 18524
rect 19515 18468 19519 18524
rect 19455 18464 19519 18468
rect 19535 18524 19599 18528
rect 19535 18468 19539 18524
rect 19539 18468 19595 18524
rect 19595 18468 19599 18524
rect 19535 18464 19599 18468
rect 19615 18524 19679 18528
rect 19615 18468 19619 18524
rect 19619 18468 19675 18524
rect 19675 18468 19679 18524
rect 19615 18464 19679 18468
rect 26965 18524 27029 18528
rect 26965 18468 26969 18524
rect 26969 18468 27025 18524
rect 27025 18468 27029 18524
rect 26965 18464 27029 18468
rect 27045 18524 27109 18528
rect 27045 18468 27049 18524
rect 27049 18468 27105 18524
rect 27105 18468 27109 18524
rect 27045 18464 27109 18468
rect 27125 18524 27189 18528
rect 27125 18468 27129 18524
rect 27129 18468 27185 18524
rect 27185 18468 27189 18524
rect 27125 18464 27189 18468
rect 27205 18524 27269 18528
rect 27205 18468 27209 18524
rect 27209 18468 27265 18524
rect 27265 18468 27269 18524
rect 27205 18464 27269 18468
rect 25820 18396 25884 18460
rect 7052 18260 7116 18324
rect 10732 18260 10796 18324
rect 30052 18260 30116 18324
rect 4660 18124 4724 18188
rect 13492 18124 13556 18188
rect 3924 17988 3988 18052
rect 4844 17988 4908 18052
rect 5396 17988 5460 18052
rect 5948 18048 6012 18052
rect 5948 17992 5998 18048
rect 5998 17992 6012 18048
rect 5948 17988 6012 17992
rect 7788 17988 7852 18052
rect 7990 17980 8054 17984
rect 7990 17924 7994 17980
rect 7994 17924 8050 17980
rect 8050 17924 8054 17980
rect 7990 17920 8054 17924
rect 8070 17980 8134 17984
rect 8070 17924 8074 17980
rect 8074 17924 8130 17980
rect 8130 17924 8134 17980
rect 8070 17920 8134 17924
rect 8150 17980 8214 17984
rect 8150 17924 8154 17980
rect 8154 17924 8210 17980
rect 8210 17924 8214 17980
rect 8150 17920 8214 17924
rect 8230 17980 8294 17984
rect 8230 17924 8234 17980
rect 8234 17924 8290 17980
rect 8290 17924 8294 17980
rect 8230 17920 8294 17924
rect 15580 17980 15644 17984
rect 15580 17924 15584 17980
rect 15584 17924 15640 17980
rect 15640 17924 15644 17980
rect 15580 17920 15644 17924
rect 15660 17980 15724 17984
rect 15660 17924 15664 17980
rect 15664 17924 15720 17980
rect 15720 17924 15724 17980
rect 15660 17920 15724 17924
rect 15740 17980 15804 17984
rect 15740 17924 15744 17980
rect 15744 17924 15800 17980
rect 15800 17924 15804 17980
rect 15740 17920 15804 17924
rect 15820 17980 15884 17984
rect 15820 17924 15824 17980
rect 15824 17924 15880 17980
rect 15880 17924 15884 17980
rect 15820 17920 15884 17924
rect 23170 17980 23234 17984
rect 23170 17924 23174 17980
rect 23174 17924 23230 17980
rect 23230 17924 23234 17980
rect 23170 17920 23234 17924
rect 23250 17980 23314 17984
rect 23250 17924 23254 17980
rect 23254 17924 23310 17980
rect 23310 17924 23314 17980
rect 23250 17920 23314 17924
rect 23330 17980 23394 17984
rect 23330 17924 23334 17980
rect 23334 17924 23390 17980
rect 23390 17924 23394 17980
rect 23330 17920 23394 17924
rect 23410 17980 23474 17984
rect 23410 17924 23414 17980
rect 23414 17924 23470 17980
rect 23470 17924 23474 17980
rect 23410 17920 23474 17924
rect 30760 17980 30824 17984
rect 30760 17924 30764 17980
rect 30764 17924 30820 17980
rect 30820 17924 30824 17980
rect 30760 17920 30824 17924
rect 30840 17980 30904 17984
rect 30840 17924 30844 17980
rect 30844 17924 30900 17980
rect 30900 17924 30904 17980
rect 30840 17920 30904 17924
rect 30920 17980 30984 17984
rect 30920 17924 30924 17980
rect 30924 17924 30980 17980
rect 30980 17924 30984 17980
rect 30920 17920 30984 17924
rect 31000 17980 31064 17984
rect 31000 17924 31004 17980
rect 31004 17924 31060 17980
rect 31060 17924 31064 17980
rect 31000 17920 31064 17924
rect 11652 17912 11716 17916
rect 11652 17856 11702 17912
rect 11702 17856 11716 17912
rect 11652 17852 11716 17856
rect 8524 17444 8588 17508
rect 23612 17716 23676 17780
rect 4195 17436 4259 17440
rect 4195 17380 4199 17436
rect 4199 17380 4255 17436
rect 4255 17380 4259 17436
rect 4195 17376 4259 17380
rect 4275 17436 4339 17440
rect 4275 17380 4279 17436
rect 4279 17380 4335 17436
rect 4335 17380 4339 17436
rect 4275 17376 4339 17380
rect 4355 17436 4419 17440
rect 4355 17380 4359 17436
rect 4359 17380 4415 17436
rect 4415 17380 4419 17436
rect 4355 17376 4419 17380
rect 4435 17436 4499 17440
rect 4435 17380 4439 17436
rect 4439 17380 4495 17436
rect 4495 17380 4499 17436
rect 4435 17376 4499 17380
rect 11785 17436 11849 17440
rect 11785 17380 11789 17436
rect 11789 17380 11845 17436
rect 11845 17380 11849 17436
rect 11785 17376 11849 17380
rect 11865 17436 11929 17440
rect 11865 17380 11869 17436
rect 11869 17380 11925 17436
rect 11925 17380 11929 17436
rect 11865 17376 11929 17380
rect 11945 17436 12009 17440
rect 11945 17380 11949 17436
rect 11949 17380 12005 17436
rect 12005 17380 12009 17436
rect 11945 17376 12009 17380
rect 12025 17436 12089 17440
rect 12025 17380 12029 17436
rect 12029 17380 12085 17436
rect 12085 17380 12089 17436
rect 12025 17376 12089 17380
rect 19375 17436 19439 17440
rect 19375 17380 19379 17436
rect 19379 17380 19435 17436
rect 19435 17380 19439 17436
rect 19375 17376 19439 17380
rect 19455 17436 19519 17440
rect 19455 17380 19459 17436
rect 19459 17380 19515 17436
rect 19515 17380 19519 17436
rect 19455 17376 19519 17380
rect 19535 17436 19599 17440
rect 19535 17380 19539 17436
rect 19539 17380 19595 17436
rect 19595 17380 19599 17436
rect 19535 17376 19599 17380
rect 19615 17436 19679 17440
rect 19615 17380 19619 17436
rect 19619 17380 19675 17436
rect 19675 17380 19679 17436
rect 19615 17376 19679 17380
rect 26965 17436 27029 17440
rect 26965 17380 26969 17436
rect 26969 17380 27025 17436
rect 27025 17380 27029 17436
rect 26965 17376 27029 17380
rect 27045 17436 27109 17440
rect 27045 17380 27049 17436
rect 27049 17380 27105 17436
rect 27105 17380 27109 17436
rect 27045 17376 27109 17380
rect 27125 17436 27189 17440
rect 27125 17380 27129 17436
rect 27129 17380 27185 17436
rect 27185 17380 27189 17436
rect 27125 17376 27189 17380
rect 27205 17436 27269 17440
rect 27205 17380 27209 17436
rect 27209 17380 27265 17436
rect 27265 17380 27269 17436
rect 27205 17376 27269 17380
rect 10548 17308 10612 17372
rect 11468 17172 11532 17236
rect 7990 16892 8054 16896
rect 7990 16836 7994 16892
rect 7994 16836 8050 16892
rect 8050 16836 8054 16892
rect 7990 16832 8054 16836
rect 8070 16892 8134 16896
rect 8070 16836 8074 16892
rect 8074 16836 8130 16892
rect 8130 16836 8134 16892
rect 8070 16832 8134 16836
rect 8150 16892 8214 16896
rect 8150 16836 8154 16892
rect 8154 16836 8210 16892
rect 8210 16836 8214 16892
rect 8150 16832 8214 16836
rect 8230 16892 8294 16896
rect 8230 16836 8234 16892
rect 8234 16836 8290 16892
rect 8290 16836 8294 16892
rect 8230 16832 8294 16836
rect 15580 16892 15644 16896
rect 15580 16836 15584 16892
rect 15584 16836 15640 16892
rect 15640 16836 15644 16892
rect 15580 16832 15644 16836
rect 15660 16892 15724 16896
rect 15660 16836 15664 16892
rect 15664 16836 15720 16892
rect 15720 16836 15724 16892
rect 15660 16832 15724 16836
rect 15740 16892 15804 16896
rect 15740 16836 15744 16892
rect 15744 16836 15800 16892
rect 15800 16836 15804 16892
rect 15740 16832 15804 16836
rect 15820 16892 15884 16896
rect 15820 16836 15824 16892
rect 15824 16836 15880 16892
rect 15880 16836 15884 16892
rect 15820 16832 15884 16836
rect 23170 16892 23234 16896
rect 23170 16836 23174 16892
rect 23174 16836 23230 16892
rect 23230 16836 23234 16892
rect 23170 16832 23234 16836
rect 23250 16892 23314 16896
rect 23250 16836 23254 16892
rect 23254 16836 23310 16892
rect 23310 16836 23314 16892
rect 23250 16832 23314 16836
rect 23330 16892 23394 16896
rect 23330 16836 23334 16892
rect 23334 16836 23390 16892
rect 23390 16836 23394 16892
rect 23330 16832 23394 16836
rect 23410 16892 23474 16896
rect 23410 16836 23414 16892
rect 23414 16836 23470 16892
rect 23470 16836 23474 16892
rect 23410 16832 23474 16836
rect 30760 16892 30824 16896
rect 30760 16836 30764 16892
rect 30764 16836 30820 16892
rect 30820 16836 30824 16892
rect 30760 16832 30824 16836
rect 30840 16892 30904 16896
rect 30840 16836 30844 16892
rect 30844 16836 30900 16892
rect 30900 16836 30904 16892
rect 30840 16832 30904 16836
rect 30920 16892 30984 16896
rect 30920 16836 30924 16892
rect 30924 16836 30980 16892
rect 30980 16836 30984 16892
rect 30920 16832 30984 16836
rect 31000 16892 31064 16896
rect 31000 16836 31004 16892
rect 31004 16836 31060 16892
rect 31060 16836 31064 16892
rect 31000 16832 31064 16836
rect 4195 16348 4259 16352
rect 4195 16292 4199 16348
rect 4199 16292 4255 16348
rect 4255 16292 4259 16348
rect 4195 16288 4259 16292
rect 4275 16348 4339 16352
rect 4275 16292 4279 16348
rect 4279 16292 4335 16348
rect 4335 16292 4339 16348
rect 4275 16288 4339 16292
rect 4355 16348 4419 16352
rect 4355 16292 4359 16348
rect 4359 16292 4415 16348
rect 4415 16292 4419 16348
rect 4355 16288 4419 16292
rect 4435 16348 4499 16352
rect 4435 16292 4439 16348
rect 4439 16292 4495 16348
rect 4495 16292 4499 16348
rect 4435 16288 4499 16292
rect 11785 16348 11849 16352
rect 11785 16292 11789 16348
rect 11789 16292 11845 16348
rect 11845 16292 11849 16348
rect 11785 16288 11849 16292
rect 11865 16348 11929 16352
rect 11865 16292 11869 16348
rect 11869 16292 11925 16348
rect 11925 16292 11929 16348
rect 11865 16288 11929 16292
rect 11945 16348 12009 16352
rect 11945 16292 11949 16348
rect 11949 16292 12005 16348
rect 12005 16292 12009 16348
rect 11945 16288 12009 16292
rect 12025 16348 12089 16352
rect 12025 16292 12029 16348
rect 12029 16292 12085 16348
rect 12085 16292 12089 16348
rect 12025 16288 12089 16292
rect 19375 16348 19439 16352
rect 19375 16292 19379 16348
rect 19379 16292 19435 16348
rect 19435 16292 19439 16348
rect 19375 16288 19439 16292
rect 19455 16348 19519 16352
rect 19455 16292 19459 16348
rect 19459 16292 19515 16348
rect 19515 16292 19519 16348
rect 19455 16288 19519 16292
rect 19535 16348 19599 16352
rect 19535 16292 19539 16348
rect 19539 16292 19595 16348
rect 19595 16292 19599 16348
rect 19535 16288 19599 16292
rect 19615 16348 19679 16352
rect 19615 16292 19619 16348
rect 19619 16292 19675 16348
rect 19675 16292 19679 16348
rect 19615 16288 19679 16292
rect 26965 16348 27029 16352
rect 26965 16292 26969 16348
rect 26969 16292 27025 16348
rect 27025 16292 27029 16348
rect 26965 16288 27029 16292
rect 27045 16348 27109 16352
rect 27045 16292 27049 16348
rect 27049 16292 27105 16348
rect 27105 16292 27109 16348
rect 27045 16288 27109 16292
rect 27125 16348 27189 16352
rect 27125 16292 27129 16348
rect 27129 16292 27185 16348
rect 27185 16292 27189 16348
rect 27125 16288 27189 16292
rect 27205 16348 27269 16352
rect 27205 16292 27209 16348
rect 27209 16292 27265 16348
rect 27265 16292 27269 16348
rect 27205 16288 27269 16292
rect 7990 15804 8054 15808
rect 7990 15748 7994 15804
rect 7994 15748 8050 15804
rect 8050 15748 8054 15804
rect 7990 15744 8054 15748
rect 8070 15804 8134 15808
rect 8070 15748 8074 15804
rect 8074 15748 8130 15804
rect 8130 15748 8134 15804
rect 8070 15744 8134 15748
rect 8150 15804 8214 15808
rect 8150 15748 8154 15804
rect 8154 15748 8210 15804
rect 8210 15748 8214 15804
rect 8150 15744 8214 15748
rect 8230 15804 8294 15808
rect 8230 15748 8234 15804
rect 8234 15748 8290 15804
rect 8290 15748 8294 15804
rect 8230 15744 8294 15748
rect 15580 15804 15644 15808
rect 15580 15748 15584 15804
rect 15584 15748 15640 15804
rect 15640 15748 15644 15804
rect 15580 15744 15644 15748
rect 15660 15804 15724 15808
rect 15660 15748 15664 15804
rect 15664 15748 15720 15804
rect 15720 15748 15724 15804
rect 15660 15744 15724 15748
rect 15740 15804 15804 15808
rect 15740 15748 15744 15804
rect 15744 15748 15800 15804
rect 15800 15748 15804 15804
rect 15740 15744 15804 15748
rect 15820 15804 15884 15808
rect 15820 15748 15824 15804
rect 15824 15748 15880 15804
rect 15880 15748 15884 15804
rect 15820 15744 15884 15748
rect 23170 15804 23234 15808
rect 23170 15748 23174 15804
rect 23174 15748 23230 15804
rect 23230 15748 23234 15804
rect 23170 15744 23234 15748
rect 23250 15804 23314 15808
rect 23250 15748 23254 15804
rect 23254 15748 23310 15804
rect 23310 15748 23314 15804
rect 23250 15744 23314 15748
rect 23330 15804 23394 15808
rect 23330 15748 23334 15804
rect 23334 15748 23390 15804
rect 23390 15748 23394 15804
rect 23330 15744 23394 15748
rect 23410 15804 23474 15808
rect 23410 15748 23414 15804
rect 23414 15748 23470 15804
rect 23470 15748 23474 15804
rect 23410 15744 23474 15748
rect 30760 15804 30824 15808
rect 30760 15748 30764 15804
rect 30764 15748 30820 15804
rect 30820 15748 30824 15804
rect 30760 15744 30824 15748
rect 30840 15804 30904 15808
rect 30840 15748 30844 15804
rect 30844 15748 30900 15804
rect 30900 15748 30904 15804
rect 30840 15744 30904 15748
rect 30920 15804 30984 15808
rect 30920 15748 30924 15804
rect 30924 15748 30980 15804
rect 30980 15748 30984 15804
rect 30920 15744 30984 15748
rect 31000 15804 31064 15808
rect 31000 15748 31004 15804
rect 31004 15748 31060 15804
rect 31060 15748 31064 15804
rect 31000 15744 31064 15748
rect 9628 15676 9692 15740
rect 24164 15404 24228 15468
rect 26372 15268 26436 15332
rect 4195 15260 4259 15264
rect 4195 15204 4199 15260
rect 4199 15204 4255 15260
rect 4255 15204 4259 15260
rect 4195 15200 4259 15204
rect 4275 15260 4339 15264
rect 4275 15204 4279 15260
rect 4279 15204 4335 15260
rect 4335 15204 4339 15260
rect 4275 15200 4339 15204
rect 4355 15260 4419 15264
rect 4355 15204 4359 15260
rect 4359 15204 4415 15260
rect 4415 15204 4419 15260
rect 4355 15200 4419 15204
rect 4435 15260 4499 15264
rect 4435 15204 4439 15260
rect 4439 15204 4495 15260
rect 4495 15204 4499 15260
rect 4435 15200 4499 15204
rect 11785 15260 11849 15264
rect 11785 15204 11789 15260
rect 11789 15204 11845 15260
rect 11845 15204 11849 15260
rect 11785 15200 11849 15204
rect 11865 15260 11929 15264
rect 11865 15204 11869 15260
rect 11869 15204 11925 15260
rect 11925 15204 11929 15260
rect 11865 15200 11929 15204
rect 11945 15260 12009 15264
rect 11945 15204 11949 15260
rect 11949 15204 12005 15260
rect 12005 15204 12009 15260
rect 11945 15200 12009 15204
rect 12025 15260 12089 15264
rect 12025 15204 12029 15260
rect 12029 15204 12085 15260
rect 12085 15204 12089 15260
rect 12025 15200 12089 15204
rect 19375 15260 19439 15264
rect 19375 15204 19379 15260
rect 19379 15204 19435 15260
rect 19435 15204 19439 15260
rect 19375 15200 19439 15204
rect 19455 15260 19519 15264
rect 19455 15204 19459 15260
rect 19459 15204 19515 15260
rect 19515 15204 19519 15260
rect 19455 15200 19519 15204
rect 19535 15260 19599 15264
rect 19535 15204 19539 15260
rect 19539 15204 19595 15260
rect 19595 15204 19599 15260
rect 19535 15200 19599 15204
rect 19615 15260 19679 15264
rect 19615 15204 19619 15260
rect 19619 15204 19675 15260
rect 19675 15204 19679 15260
rect 19615 15200 19679 15204
rect 26965 15260 27029 15264
rect 26965 15204 26969 15260
rect 26969 15204 27025 15260
rect 27025 15204 27029 15260
rect 26965 15200 27029 15204
rect 27045 15260 27109 15264
rect 27045 15204 27049 15260
rect 27049 15204 27105 15260
rect 27105 15204 27109 15260
rect 27045 15200 27109 15204
rect 27125 15260 27189 15264
rect 27125 15204 27129 15260
rect 27129 15204 27185 15260
rect 27185 15204 27189 15260
rect 27125 15200 27189 15204
rect 27205 15260 27269 15264
rect 27205 15204 27209 15260
rect 27209 15204 27265 15260
rect 27265 15204 27269 15260
rect 27205 15200 27269 15204
rect 10548 15192 10612 15196
rect 10548 15136 10598 15192
rect 10598 15136 10612 15192
rect 10548 15132 10612 15136
rect 12204 14860 12268 14924
rect 29500 14860 29564 14924
rect 7990 14716 8054 14720
rect 7990 14660 7994 14716
rect 7994 14660 8050 14716
rect 8050 14660 8054 14716
rect 7990 14656 8054 14660
rect 8070 14716 8134 14720
rect 8070 14660 8074 14716
rect 8074 14660 8130 14716
rect 8130 14660 8134 14716
rect 8070 14656 8134 14660
rect 8150 14716 8214 14720
rect 8150 14660 8154 14716
rect 8154 14660 8210 14716
rect 8210 14660 8214 14716
rect 8150 14656 8214 14660
rect 8230 14716 8294 14720
rect 8230 14660 8234 14716
rect 8234 14660 8290 14716
rect 8290 14660 8294 14716
rect 8230 14656 8294 14660
rect 15580 14716 15644 14720
rect 15580 14660 15584 14716
rect 15584 14660 15640 14716
rect 15640 14660 15644 14716
rect 15580 14656 15644 14660
rect 15660 14716 15724 14720
rect 15660 14660 15664 14716
rect 15664 14660 15720 14716
rect 15720 14660 15724 14716
rect 15660 14656 15724 14660
rect 15740 14716 15804 14720
rect 15740 14660 15744 14716
rect 15744 14660 15800 14716
rect 15800 14660 15804 14716
rect 15740 14656 15804 14660
rect 15820 14716 15884 14720
rect 15820 14660 15824 14716
rect 15824 14660 15880 14716
rect 15880 14660 15884 14716
rect 15820 14656 15884 14660
rect 23170 14716 23234 14720
rect 23170 14660 23174 14716
rect 23174 14660 23230 14716
rect 23230 14660 23234 14716
rect 23170 14656 23234 14660
rect 23250 14716 23314 14720
rect 23250 14660 23254 14716
rect 23254 14660 23310 14716
rect 23310 14660 23314 14716
rect 23250 14656 23314 14660
rect 23330 14716 23394 14720
rect 23330 14660 23334 14716
rect 23334 14660 23390 14716
rect 23390 14660 23394 14716
rect 23330 14656 23394 14660
rect 23410 14716 23474 14720
rect 23410 14660 23414 14716
rect 23414 14660 23470 14716
rect 23470 14660 23474 14716
rect 23410 14656 23474 14660
rect 30760 14716 30824 14720
rect 30760 14660 30764 14716
rect 30764 14660 30820 14716
rect 30820 14660 30824 14716
rect 30760 14656 30824 14660
rect 30840 14716 30904 14720
rect 30840 14660 30844 14716
rect 30844 14660 30900 14716
rect 30900 14660 30904 14716
rect 30840 14656 30904 14660
rect 30920 14716 30984 14720
rect 30920 14660 30924 14716
rect 30924 14660 30980 14716
rect 30980 14660 30984 14716
rect 30920 14656 30984 14660
rect 31000 14716 31064 14720
rect 31000 14660 31004 14716
rect 31004 14660 31060 14716
rect 31060 14660 31064 14716
rect 31000 14656 31064 14660
rect 10364 14240 10428 14244
rect 10364 14184 10378 14240
rect 10378 14184 10428 14240
rect 10364 14180 10428 14184
rect 12204 14180 12268 14244
rect 4195 14172 4259 14176
rect 4195 14116 4199 14172
rect 4199 14116 4255 14172
rect 4255 14116 4259 14172
rect 4195 14112 4259 14116
rect 4275 14172 4339 14176
rect 4275 14116 4279 14172
rect 4279 14116 4335 14172
rect 4335 14116 4339 14172
rect 4275 14112 4339 14116
rect 4355 14172 4419 14176
rect 4355 14116 4359 14172
rect 4359 14116 4415 14172
rect 4415 14116 4419 14172
rect 4355 14112 4419 14116
rect 4435 14172 4499 14176
rect 4435 14116 4439 14172
rect 4439 14116 4495 14172
rect 4495 14116 4499 14172
rect 4435 14112 4499 14116
rect 11785 14172 11849 14176
rect 11785 14116 11789 14172
rect 11789 14116 11845 14172
rect 11845 14116 11849 14172
rect 11785 14112 11849 14116
rect 11865 14172 11929 14176
rect 11865 14116 11869 14172
rect 11869 14116 11925 14172
rect 11925 14116 11929 14172
rect 11865 14112 11929 14116
rect 11945 14172 12009 14176
rect 11945 14116 11949 14172
rect 11949 14116 12005 14172
rect 12005 14116 12009 14172
rect 11945 14112 12009 14116
rect 12025 14172 12089 14176
rect 12025 14116 12029 14172
rect 12029 14116 12085 14172
rect 12085 14116 12089 14172
rect 12025 14112 12089 14116
rect 1716 13832 1780 13836
rect 1716 13776 1730 13832
rect 1730 13776 1780 13832
rect 1716 13772 1780 13776
rect 6500 13636 6564 13700
rect 11100 13772 11164 13836
rect 19375 14172 19439 14176
rect 19375 14116 19379 14172
rect 19379 14116 19435 14172
rect 19435 14116 19439 14172
rect 19375 14112 19439 14116
rect 19455 14172 19519 14176
rect 19455 14116 19459 14172
rect 19459 14116 19515 14172
rect 19515 14116 19519 14172
rect 19455 14112 19519 14116
rect 19535 14172 19599 14176
rect 19535 14116 19539 14172
rect 19539 14116 19595 14172
rect 19595 14116 19599 14172
rect 19535 14112 19599 14116
rect 19615 14172 19679 14176
rect 19615 14116 19619 14172
rect 19619 14116 19675 14172
rect 19675 14116 19679 14172
rect 19615 14112 19679 14116
rect 26965 14172 27029 14176
rect 26965 14116 26969 14172
rect 26969 14116 27025 14172
rect 27025 14116 27029 14172
rect 26965 14112 27029 14116
rect 27045 14172 27109 14176
rect 27045 14116 27049 14172
rect 27049 14116 27105 14172
rect 27105 14116 27109 14172
rect 27045 14112 27109 14116
rect 27125 14172 27189 14176
rect 27125 14116 27129 14172
rect 27129 14116 27185 14172
rect 27185 14116 27189 14172
rect 27125 14112 27189 14116
rect 27205 14172 27269 14176
rect 27205 14116 27209 14172
rect 27209 14116 27265 14172
rect 27265 14116 27269 14172
rect 27205 14112 27269 14116
rect 30052 13772 30116 13836
rect 7990 13628 8054 13632
rect 7990 13572 7994 13628
rect 7994 13572 8050 13628
rect 8050 13572 8054 13628
rect 7990 13568 8054 13572
rect 8070 13628 8134 13632
rect 8070 13572 8074 13628
rect 8074 13572 8130 13628
rect 8130 13572 8134 13628
rect 8070 13568 8134 13572
rect 8150 13628 8214 13632
rect 8150 13572 8154 13628
rect 8154 13572 8210 13628
rect 8210 13572 8214 13628
rect 8150 13568 8214 13572
rect 8230 13628 8294 13632
rect 8230 13572 8234 13628
rect 8234 13572 8290 13628
rect 8290 13572 8294 13628
rect 8230 13568 8294 13572
rect 15580 13628 15644 13632
rect 15580 13572 15584 13628
rect 15584 13572 15640 13628
rect 15640 13572 15644 13628
rect 15580 13568 15644 13572
rect 15660 13628 15724 13632
rect 15660 13572 15664 13628
rect 15664 13572 15720 13628
rect 15720 13572 15724 13628
rect 15660 13568 15724 13572
rect 15740 13628 15804 13632
rect 15740 13572 15744 13628
rect 15744 13572 15800 13628
rect 15800 13572 15804 13628
rect 15740 13568 15804 13572
rect 15820 13628 15884 13632
rect 15820 13572 15824 13628
rect 15824 13572 15880 13628
rect 15880 13572 15884 13628
rect 15820 13568 15884 13572
rect 23170 13628 23234 13632
rect 23170 13572 23174 13628
rect 23174 13572 23230 13628
rect 23230 13572 23234 13628
rect 23170 13568 23234 13572
rect 23250 13628 23314 13632
rect 23250 13572 23254 13628
rect 23254 13572 23310 13628
rect 23310 13572 23314 13628
rect 23250 13568 23314 13572
rect 23330 13628 23394 13632
rect 23330 13572 23334 13628
rect 23334 13572 23390 13628
rect 23390 13572 23394 13628
rect 23330 13568 23394 13572
rect 23410 13628 23474 13632
rect 23410 13572 23414 13628
rect 23414 13572 23470 13628
rect 23470 13572 23474 13628
rect 23410 13568 23474 13572
rect 30760 13628 30824 13632
rect 30760 13572 30764 13628
rect 30764 13572 30820 13628
rect 30820 13572 30824 13628
rect 30760 13568 30824 13572
rect 30840 13628 30904 13632
rect 30840 13572 30844 13628
rect 30844 13572 30900 13628
rect 30900 13572 30904 13628
rect 30840 13568 30904 13572
rect 30920 13628 30984 13632
rect 30920 13572 30924 13628
rect 30924 13572 30980 13628
rect 30980 13572 30984 13628
rect 30920 13568 30984 13572
rect 31000 13628 31064 13632
rect 31000 13572 31004 13628
rect 31004 13572 31060 13628
rect 31060 13572 31064 13628
rect 31000 13568 31064 13572
rect 8524 13500 8588 13564
rect 7604 13228 7668 13292
rect 12388 13364 12452 13428
rect 22508 13228 22572 13292
rect 26372 13092 26436 13156
rect 4195 13084 4259 13088
rect 4195 13028 4199 13084
rect 4199 13028 4255 13084
rect 4255 13028 4259 13084
rect 4195 13024 4259 13028
rect 4275 13084 4339 13088
rect 4275 13028 4279 13084
rect 4279 13028 4335 13084
rect 4335 13028 4339 13084
rect 4275 13024 4339 13028
rect 4355 13084 4419 13088
rect 4355 13028 4359 13084
rect 4359 13028 4415 13084
rect 4415 13028 4419 13084
rect 4355 13024 4419 13028
rect 4435 13084 4499 13088
rect 4435 13028 4439 13084
rect 4439 13028 4495 13084
rect 4495 13028 4499 13084
rect 4435 13024 4499 13028
rect 11785 13084 11849 13088
rect 11785 13028 11789 13084
rect 11789 13028 11845 13084
rect 11845 13028 11849 13084
rect 11785 13024 11849 13028
rect 11865 13084 11929 13088
rect 11865 13028 11869 13084
rect 11869 13028 11925 13084
rect 11925 13028 11929 13084
rect 11865 13024 11929 13028
rect 11945 13084 12009 13088
rect 11945 13028 11949 13084
rect 11949 13028 12005 13084
rect 12005 13028 12009 13084
rect 11945 13024 12009 13028
rect 12025 13084 12089 13088
rect 12025 13028 12029 13084
rect 12029 13028 12085 13084
rect 12085 13028 12089 13084
rect 12025 13024 12089 13028
rect 19375 13084 19439 13088
rect 19375 13028 19379 13084
rect 19379 13028 19435 13084
rect 19435 13028 19439 13084
rect 19375 13024 19439 13028
rect 19455 13084 19519 13088
rect 19455 13028 19459 13084
rect 19459 13028 19515 13084
rect 19515 13028 19519 13084
rect 19455 13024 19519 13028
rect 19535 13084 19599 13088
rect 19535 13028 19539 13084
rect 19539 13028 19595 13084
rect 19595 13028 19599 13084
rect 19535 13024 19599 13028
rect 19615 13084 19679 13088
rect 19615 13028 19619 13084
rect 19619 13028 19675 13084
rect 19675 13028 19679 13084
rect 19615 13024 19679 13028
rect 26965 13084 27029 13088
rect 26965 13028 26969 13084
rect 26969 13028 27025 13084
rect 27025 13028 27029 13084
rect 26965 13024 27029 13028
rect 27045 13084 27109 13088
rect 27045 13028 27049 13084
rect 27049 13028 27105 13084
rect 27105 13028 27109 13084
rect 27045 13024 27109 13028
rect 27125 13084 27189 13088
rect 27125 13028 27129 13084
rect 27129 13028 27185 13084
rect 27185 13028 27189 13084
rect 27125 13024 27189 13028
rect 27205 13084 27269 13088
rect 27205 13028 27209 13084
rect 27209 13028 27265 13084
rect 27265 13028 27269 13084
rect 27205 13024 27269 13028
rect 11284 13016 11348 13020
rect 11284 12960 11298 13016
rect 11298 12960 11348 13016
rect 11284 12956 11348 12960
rect 11468 12956 11532 13020
rect 12388 12956 12452 13020
rect 21956 12820 22020 12884
rect 7990 12540 8054 12544
rect 7990 12484 7994 12540
rect 7994 12484 8050 12540
rect 8050 12484 8054 12540
rect 7990 12480 8054 12484
rect 8070 12540 8134 12544
rect 8070 12484 8074 12540
rect 8074 12484 8130 12540
rect 8130 12484 8134 12540
rect 8070 12480 8134 12484
rect 8150 12540 8214 12544
rect 8150 12484 8154 12540
rect 8154 12484 8210 12540
rect 8210 12484 8214 12540
rect 8150 12480 8214 12484
rect 8230 12540 8294 12544
rect 8230 12484 8234 12540
rect 8234 12484 8290 12540
rect 8290 12484 8294 12540
rect 8230 12480 8294 12484
rect 15580 12540 15644 12544
rect 15580 12484 15584 12540
rect 15584 12484 15640 12540
rect 15640 12484 15644 12540
rect 15580 12480 15644 12484
rect 15660 12540 15724 12544
rect 15660 12484 15664 12540
rect 15664 12484 15720 12540
rect 15720 12484 15724 12540
rect 15660 12480 15724 12484
rect 15740 12540 15804 12544
rect 15740 12484 15744 12540
rect 15744 12484 15800 12540
rect 15800 12484 15804 12540
rect 15740 12480 15804 12484
rect 15820 12540 15884 12544
rect 15820 12484 15824 12540
rect 15824 12484 15880 12540
rect 15880 12484 15884 12540
rect 15820 12480 15884 12484
rect 23170 12540 23234 12544
rect 23170 12484 23174 12540
rect 23174 12484 23230 12540
rect 23230 12484 23234 12540
rect 23170 12480 23234 12484
rect 23250 12540 23314 12544
rect 23250 12484 23254 12540
rect 23254 12484 23310 12540
rect 23310 12484 23314 12540
rect 23250 12480 23314 12484
rect 23330 12540 23394 12544
rect 23330 12484 23334 12540
rect 23334 12484 23390 12540
rect 23390 12484 23394 12540
rect 23330 12480 23394 12484
rect 23410 12540 23474 12544
rect 23410 12484 23414 12540
rect 23414 12484 23470 12540
rect 23470 12484 23474 12540
rect 23410 12480 23474 12484
rect 3740 12412 3804 12476
rect 13492 12412 13556 12476
rect 26188 12684 26252 12748
rect 30760 12540 30824 12544
rect 30760 12484 30764 12540
rect 30764 12484 30820 12540
rect 30820 12484 30824 12540
rect 30760 12480 30824 12484
rect 30840 12540 30904 12544
rect 30840 12484 30844 12540
rect 30844 12484 30900 12540
rect 30900 12484 30904 12540
rect 30840 12480 30904 12484
rect 30920 12540 30984 12544
rect 30920 12484 30924 12540
rect 30924 12484 30980 12540
rect 30980 12484 30984 12540
rect 30920 12480 30984 12484
rect 31000 12540 31064 12544
rect 31000 12484 31004 12540
rect 31004 12484 31060 12540
rect 31060 12484 31064 12540
rect 31000 12480 31064 12484
rect 29500 12472 29564 12476
rect 29500 12416 29550 12472
rect 29550 12416 29564 12472
rect 29500 12412 29564 12416
rect 8892 12276 8956 12340
rect 22876 12276 22940 12340
rect 6684 12140 6748 12204
rect 4195 11996 4259 12000
rect 4195 11940 4199 11996
rect 4199 11940 4255 11996
rect 4255 11940 4259 11996
rect 4195 11936 4259 11940
rect 4275 11996 4339 12000
rect 4275 11940 4279 11996
rect 4279 11940 4335 11996
rect 4335 11940 4339 11996
rect 4275 11936 4339 11940
rect 4355 11996 4419 12000
rect 4355 11940 4359 11996
rect 4359 11940 4415 11996
rect 4415 11940 4419 11996
rect 4355 11936 4419 11940
rect 4435 11996 4499 12000
rect 4435 11940 4439 11996
rect 4439 11940 4495 11996
rect 4495 11940 4499 11996
rect 4435 11936 4499 11940
rect 11785 11996 11849 12000
rect 11785 11940 11789 11996
rect 11789 11940 11845 11996
rect 11845 11940 11849 11996
rect 11785 11936 11849 11940
rect 11865 11996 11929 12000
rect 11865 11940 11869 11996
rect 11869 11940 11925 11996
rect 11925 11940 11929 11996
rect 11865 11936 11929 11940
rect 11945 11996 12009 12000
rect 11945 11940 11949 11996
rect 11949 11940 12005 11996
rect 12005 11940 12009 11996
rect 11945 11936 12009 11940
rect 12025 11996 12089 12000
rect 12025 11940 12029 11996
rect 12029 11940 12085 11996
rect 12085 11940 12089 11996
rect 12025 11936 12089 11940
rect 19375 11996 19439 12000
rect 19375 11940 19379 11996
rect 19379 11940 19435 11996
rect 19435 11940 19439 11996
rect 19375 11936 19439 11940
rect 19455 11996 19519 12000
rect 19455 11940 19459 11996
rect 19459 11940 19515 11996
rect 19515 11940 19519 11996
rect 19455 11936 19519 11940
rect 19535 11996 19599 12000
rect 19535 11940 19539 11996
rect 19539 11940 19595 11996
rect 19595 11940 19599 11996
rect 19535 11936 19599 11940
rect 19615 11996 19679 12000
rect 19615 11940 19619 11996
rect 19619 11940 19675 11996
rect 19675 11940 19679 11996
rect 19615 11936 19679 11940
rect 26965 11996 27029 12000
rect 26965 11940 26969 11996
rect 26969 11940 27025 11996
rect 27025 11940 27029 11996
rect 26965 11936 27029 11940
rect 27045 11996 27109 12000
rect 27045 11940 27049 11996
rect 27049 11940 27105 11996
rect 27105 11940 27109 11996
rect 27045 11936 27109 11940
rect 27125 11996 27189 12000
rect 27125 11940 27129 11996
rect 27129 11940 27185 11996
rect 27185 11940 27189 11996
rect 27125 11936 27189 11940
rect 27205 11996 27269 12000
rect 27205 11940 27209 11996
rect 27209 11940 27265 11996
rect 27265 11940 27269 11996
rect 27205 11936 27269 11940
rect 10732 11792 10796 11796
rect 10732 11736 10782 11792
rect 10782 11736 10796 11792
rect 10732 11732 10796 11736
rect 11652 11732 11716 11796
rect 7788 11596 7852 11660
rect 7990 11452 8054 11456
rect 7990 11396 7994 11452
rect 7994 11396 8050 11452
rect 8050 11396 8054 11452
rect 7990 11392 8054 11396
rect 8070 11452 8134 11456
rect 8070 11396 8074 11452
rect 8074 11396 8130 11452
rect 8130 11396 8134 11452
rect 8070 11392 8134 11396
rect 8150 11452 8214 11456
rect 8150 11396 8154 11452
rect 8154 11396 8210 11452
rect 8210 11396 8214 11452
rect 8150 11392 8214 11396
rect 8230 11452 8294 11456
rect 8230 11396 8234 11452
rect 8234 11396 8290 11452
rect 8290 11396 8294 11452
rect 8230 11392 8294 11396
rect 15580 11452 15644 11456
rect 15580 11396 15584 11452
rect 15584 11396 15640 11452
rect 15640 11396 15644 11452
rect 15580 11392 15644 11396
rect 15660 11452 15724 11456
rect 15660 11396 15664 11452
rect 15664 11396 15720 11452
rect 15720 11396 15724 11452
rect 15660 11392 15724 11396
rect 15740 11452 15804 11456
rect 15740 11396 15744 11452
rect 15744 11396 15800 11452
rect 15800 11396 15804 11452
rect 15740 11392 15804 11396
rect 15820 11452 15884 11456
rect 15820 11396 15824 11452
rect 15824 11396 15880 11452
rect 15880 11396 15884 11452
rect 15820 11392 15884 11396
rect 23170 11452 23234 11456
rect 23170 11396 23174 11452
rect 23174 11396 23230 11452
rect 23230 11396 23234 11452
rect 23170 11392 23234 11396
rect 23250 11452 23314 11456
rect 23250 11396 23254 11452
rect 23254 11396 23310 11452
rect 23310 11396 23314 11452
rect 23250 11392 23314 11396
rect 23330 11452 23394 11456
rect 23330 11396 23334 11452
rect 23334 11396 23390 11452
rect 23390 11396 23394 11452
rect 23330 11392 23394 11396
rect 23410 11452 23474 11456
rect 23410 11396 23414 11452
rect 23414 11396 23470 11452
rect 23470 11396 23474 11452
rect 23410 11392 23474 11396
rect 30760 11452 30824 11456
rect 30760 11396 30764 11452
rect 30764 11396 30820 11452
rect 30820 11396 30824 11452
rect 30760 11392 30824 11396
rect 30840 11452 30904 11456
rect 30840 11396 30844 11452
rect 30844 11396 30900 11452
rect 30900 11396 30904 11452
rect 30840 11392 30904 11396
rect 30920 11452 30984 11456
rect 30920 11396 30924 11452
rect 30924 11396 30980 11452
rect 30980 11396 30984 11452
rect 30920 11392 30984 11396
rect 31000 11452 31064 11456
rect 31000 11396 31004 11452
rect 31004 11396 31060 11452
rect 31060 11396 31064 11452
rect 31000 11392 31064 11396
rect 15148 11052 15212 11116
rect 4195 10908 4259 10912
rect 4195 10852 4199 10908
rect 4199 10852 4255 10908
rect 4255 10852 4259 10908
rect 4195 10848 4259 10852
rect 4275 10908 4339 10912
rect 4275 10852 4279 10908
rect 4279 10852 4335 10908
rect 4335 10852 4339 10908
rect 4275 10848 4339 10852
rect 4355 10908 4419 10912
rect 4355 10852 4359 10908
rect 4359 10852 4415 10908
rect 4415 10852 4419 10908
rect 4355 10848 4419 10852
rect 4435 10908 4499 10912
rect 4435 10852 4439 10908
rect 4439 10852 4495 10908
rect 4495 10852 4499 10908
rect 4435 10848 4499 10852
rect 11785 10908 11849 10912
rect 11785 10852 11789 10908
rect 11789 10852 11845 10908
rect 11845 10852 11849 10908
rect 11785 10848 11849 10852
rect 11865 10908 11929 10912
rect 11865 10852 11869 10908
rect 11869 10852 11925 10908
rect 11925 10852 11929 10908
rect 11865 10848 11929 10852
rect 11945 10908 12009 10912
rect 11945 10852 11949 10908
rect 11949 10852 12005 10908
rect 12005 10852 12009 10908
rect 11945 10848 12009 10852
rect 12025 10908 12089 10912
rect 12025 10852 12029 10908
rect 12029 10852 12085 10908
rect 12085 10852 12089 10908
rect 12025 10848 12089 10852
rect 19375 10908 19439 10912
rect 19375 10852 19379 10908
rect 19379 10852 19435 10908
rect 19435 10852 19439 10908
rect 19375 10848 19439 10852
rect 19455 10908 19519 10912
rect 19455 10852 19459 10908
rect 19459 10852 19515 10908
rect 19515 10852 19519 10908
rect 19455 10848 19519 10852
rect 19535 10908 19599 10912
rect 19535 10852 19539 10908
rect 19539 10852 19595 10908
rect 19595 10852 19599 10908
rect 19535 10848 19599 10852
rect 19615 10908 19679 10912
rect 19615 10852 19619 10908
rect 19619 10852 19675 10908
rect 19675 10852 19679 10908
rect 19615 10848 19679 10852
rect 26965 10908 27029 10912
rect 26965 10852 26969 10908
rect 26969 10852 27025 10908
rect 27025 10852 27029 10908
rect 26965 10848 27029 10852
rect 27045 10908 27109 10912
rect 27045 10852 27049 10908
rect 27049 10852 27105 10908
rect 27105 10852 27109 10908
rect 27045 10848 27109 10852
rect 27125 10908 27189 10912
rect 27125 10852 27129 10908
rect 27129 10852 27185 10908
rect 27185 10852 27189 10908
rect 27125 10848 27189 10852
rect 27205 10908 27269 10912
rect 27205 10852 27209 10908
rect 27209 10852 27265 10908
rect 27265 10852 27269 10908
rect 27205 10848 27269 10852
rect 9628 10644 9692 10708
rect 5580 10508 5644 10572
rect 7990 10364 8054 10368
rect 7990 10308 7994 10364
rect 7994 10308 8050 10364
rect 8050 10308 8054 10364
rect 7990 10304 8054 10308
rect 8070 10364 8134 10368
rect 8070 10308 8074 10364
rect 8074 10308 8130 10364
rect 8130 10308 8134 10364
rect 8070 10304 8134 10308
rect 8150 10364 8214 10368
rect 8150 10308 8154 10364
rect 8154 10308 8210 10364
rect 8210 10308 8214 10364
rect 8150 10304 8214 10308
rect 8230 10364 8294 10368
rect 8230 10308 8234 10364
rect 8234 10308 8290 10364
rect 8290 10308 8294 10364
rect 8230 10304 8294 10308
rect 15580 10364 15644 10368
rect 15580 10308 15584 10364
rect 15584 10308 15640 10364
rect 15640 10308 15644 10364
rect 15580 10304 15644 10308
rect 15660 10364 15724 10368
rect 15660 10308 15664 10364
rect 15664 10308 15720 10364
rect 15720 10308 15724 10364
rect 15660 10304 15724 10308
rect 15740 10364 15804 10368
rect 15740 10308 15744 10364
rect 15744 10308 15800 10364
rect 15800 10308 15804 10364
rect 15740 10304 15804 10308
rect 15820 10364 15884 10368
rect 15820 10308 15824 10364
rect 15824 10308 15880 10364
rect 15880 10308 15884 10364
rect 15820 10304 15884 10308
rect 23170 10364 23234 10368
rect 23170 10308 23174 10364
rect 23174 10308 23230 10364
rect 23230 10308 23234 10364
rect 23170 10304 23234 10308
rect 23250 10364 23314 10368
rect 23250 10308 23254 10364
rect 23254 10308 23310 10364
rect 23310 10308 23314 10364
rect 23250 10304 23314 10308
rect 23330 10364 23394 10368
rect 23330 10308 23334 10364
rect 23334 10308 23390 10364
rect 23390 10308 23394 10364
rect 23330 10304 23394 10308
rect 23410 10364 23474 10368
rect 23410 10308 23414 10364
rect 23414 10308 23470 10364
rect 23470 10308 23474 10364
rect 23410 10304 23474 10308
rect 30760 10364 30824 10368
rect 30760 10308 30764 10364
rect 30764 10308 30820 10364
rect 30820 10308 30824 10364
rect 30760 10304 30824 10308
rect 30840 10364 30904 10368
rect 30840 10308 30844 10364
rect 30844 10308 30900 10364
rect 30900 10308 30904 10364
rect 30840 10304 30904 10308
rect 30920 10364 30984 10368
rect 30920 10308 30924 10364
rect 30924 10308 30980 10364
rect 30980 10308 30984 10364
rect 30920 10304 30984 10308
rect 31000 10364 31064 10368
rect 31000 10308 31004 10364
rect 31004 10308 31060 10364
rect 31060 10308 31064 10364
rect 31000 10304 31064 10308
rect 3924 10100 3988 10164
rect 4195 9820 4259 9824
rect 4195 9764 4199 9820
rect 4199 9764 4255 9820
rect 4255 9764 4259 9820
rect 4195 9760 4259 9764
rect 4275 9820 4339 9824
rect 4275 9764 4279 9820
rect 4279 9764 4335 9820
rect 4335 9764 4339 9820
rect 4275 9760 4339 9764
rect 4355 9820 4419 9824
rect 4355 9764 4359 9820
rect 4359 9764 4415 9820
rect 4415 9764 4419 9820
rect 4355 9760 4419 9764
rect 4435 9820 4499 9824
rect 4435 9764 4439 9820
rect 4439 9764 4495 9820
rect 4495 9764 4499 9820
rect 4435 9760 4499 9764
rect 11785 9820 11849 9824
rect 11785 9764 11789 9820
rect 11789 9764 11845 9820
rect 11845 9764 11849 9820
rect 11785 9760 11849 9764
rect 11865 9820 11929 9824
rect 11865 9764 11869 9820
rect 11869 9764 11925 9820
rect 11925 9764 11929 9820
rect 11865 9760 11929 9764
rect 11945 9820 12009 9824
rect 11945 9764 11949 9820
rect 11949 9764 12005 9820
rect 12005 9764 12009 9820
rect 11945 9760 12009 9764
rect 12025 9820 12089 9824
rect 12025 9764 12029 9820
rect 12029 9764 12085 9820
rect 12085 9764 12089 9820
rect 12025 9760 12089 9764
rect 19375 9820 19439 9824
rect 19375 9764 19379 9820
rect 19379 9764 19435 9820
rect 19435 9764 19439 9820
rect 19375 9760 19439 9764
rect 19455 9820 19519 9824
rect 19455 9764 19459 9820
rect 19459 9764 19515 9820
rect 19515 9764 19519 9820
rect 19455 9760 19519 9764
rect 19535 9820 19599 9824
rect 19535 9764 19539 9820
rect 19539 9764 19595 9820
rect 19595 9764 19599 9820
rect 19535 9760 19599 9764
rect 19615 9820 19679 9824
rect 19615 9764 19619 9820
rect 19619 9764 19675 9820
rect 19675 9764 19679 9820
rect 19615 9760 19679 9764
rect 26965 9820 27029 9824
rect 26965 9764 26969 9820
rect 26969 9764 27025 9820
rect 27025 9764 27029 9820
rect 26965 9760 27029 9764
rect 27045 9820 27109 9824
rect 27045 9764 27049 9820
rect 27049 9764 27105 9820
rect 27105 9764 27109 9820
rect 27045 9760 27109 9764
rect 27125 9820 27189 9824
rect 27125 9764 27129 9820
rect 27129 9764 27185 9820
rect 27185 9764 27189 9820
rect 27125 9760 27189 9764
rect 27205 9820 27269 9824
rect 27205 9764 27209 9820
rect 27209 9764 27265 9820
rect 27265 9764 27269 9820
rect 27205 9760 27269 9764
rect 7990 9276 8054 9280
rect 7990 9220 7994 9276
rect 7994 9220 8050 9276
rect 8050 9220 8054 9276
rect 7990 9216 8054 9220
rect 8070 9276 8134 9280
rect 8070 9220 8074 9276
rect 8074 9220 8130 9276
rect 8130 9220 8134 9276
rect 8070 9216 8134 9220
rect 8150 9276 8214 9280
rect 8150 9220 8154 9276
rect 8154 9220 8210 9276
rect 8210 9220 8214 9276
rect 8150 9216 8214 9220
rect 8230 9276 8294 9280
rect 8230 9220 8234 9276
rect 8234 9220 8290 9276
rect 8290 9220 8294 9276
rect 8230 9216 8294 9220
rect 15580 9276 15644 9280
rect 15580 9220 15584 9276
rect 15584 9220 15640 9276
rect 15640 9220 15644 9276
rect 15580 9216 15644 9220
rect 15660 9276 15724 9280
rect 15660 9220 15664 9276
rect 15664 9220 15720 9276
rect 15720 9220 15724 9276
rect 15660 9216 15724 9220
rect 15740 9276 15804 9280
rect 15740 9220 15744 9276
rect 15744 9220 15800 9276
rect 15800 9220 15804 9276
rect 15740 9216 15804 9220
rect 15820 9276 15884 9280
rect 15820 9220 15824 9276
rect 15824 9220 15880 9276
rect 15880 9220 15884 9276
rect 15820 9216 15884 9220
rect 23170 9276 23234 9280
rect 23170 9220 23174 9276
rect 23174 9220 23230 9276
rect 23230 9220 23234 9276
rect 23170 9216 23234 9220
rect 23250 9276 23314 9280
rect 23250 9220 23254 9276
rect 23254 9220 23310 9276
rect 23310 9220 23314 9276
rect 23250 9216 23314 9220
rect 23330 9276 23394 9280
rect 23330 9220 23334 9276
rect 23334 9220 23390 9276
rect 23390 9220 23394 9276
rect 23330 9216 23394 9220
rect 23410 9276 23474 9280
rect 23410 9220 23414 9276
rect 23414 9220 23470 9276
rect 23470 9220 23474 9276
rect 23410 9216 23474 9220
rect 30760 9276 30824 9280
rect 30760 9220 30764 9276
rect 30764 9220 30820 9276
rect 30820 9220 30824 9276
rect 30760 9216 30824 9220
rect 30840 9276 30904 9280
rect 30840 9220 30844 9276
rect 30844 9220 30900 9276
rect 30900 9220 30904 9276
rect 30840 9216 30904 9220
rect 30920 9276 30984 9280
rect 30920 9220 30924 9276
rect 30924 9220 30980 9276
rect 30980 9220 30984 9276
rect 30920 9216 30984 9220
rect 31000 9276 31064 9280
rect 31000 9220 31004 9276
rect 31004 9220 31060 9276
rect 31060 9220 31064 9276
rect 31000 9216 31064 9220
rect 4195 8732 4259 8736
rect 4195 8676 4199 8732
rect 4199 8676 4255 8732
rect 4255 8676 4259 8732
rect 4195 8672 4259 8676
rect 4275 8732 4339 8736
rect 4275 8676 4279 8732
rect 4279 8676 4335 8732
rect 4335 8676 4339 8732
rect 4275 8672 4339 8676
rect 4355 8732 4419 8736
rect 4355 8676 4359 8732
rect 4359 8676 4415 8732
rect 4415 8676 4419 8732
rect 4355 8672 4419 8676
rect 4435 8732 4499 8736
rect 4435 8676 4439 8732
rect 4439 8676 4495 8732
rect 4495 8676 4499 8732
rect 4435 8672 4499 8676
rect 11785 8732 11849 8736
rect 11785 8676 11789 8732
rect 11789 8676 11845 8732
rect 11845 8676 11849 8732
rect 11785 8672 11849 8676
rect 11865 8732 11929 8736
rect 11865 8676 11869 8732
rect 11869 8676 11925 8732
rect 11925 8676 11929 8732
rect 11865 8672 11929 8676
rect 11945 8732 12009 8736
rect 11945 8676 11949 8732
rect 11949 8676 12005 8732
rect 12005 8676 12009 8732
rect 11945 8672 12009 8676
rect 12025 8732 12089 8736
rect 12025 8676 12029 8732
rect 12029 8676 12085 8732
rect 12085 8676 12089 8732
rect 12025 8672 12089 8676
rect 19375 8732 19439 8736
rect 19375 8676 19379 8732
rect 19379 8676 19435 8732
rect 19435 8676 19439 8732
rect 19375 8672 19439 8676
rect 19455 8732 19519 8736
rect 19455 8676 19459 8732
rect 19459 8676 19515 8732
rect 19515 8676 19519 8732
rect 19455 8672 19519 8676
rect 19535 8732 19599 8736
rect 19535 8676 19539 8732
rect 19539 8676 19595 8732
rect 19595 8676 19599 8732
rect 19535 8672 19599 8676
rect 19615 8732 19679 8736
rect 19615 8676 19619 8732
rect 19619 8676 19675 8732
rect 19675 8676 19679 8732
rect 19615 8672 19679 8676
rect 26965 8732 27029 8736
rect 26965 8676 26969 8732
rect 26969 8676 27025 8732
rect 27025 8676 27029 8732
rect 26965 8672 27029 8676
rect 27045 8732 27109 8736
rect 27045 8676 27049 8732
rect 27049 8676 27105 8732
rect 27105 8676 27109 8732
rect 27045 8672 27109 8676
rect 27125 8732 27189 8736
rect 27125 8676 27129 8732
rect 27129 8676 27185 8732
rect 27185 8676 27189 8732
rect 27125 8672 27189 8676
rect 27205 8732 27269 8736
rect 27205 8676 27209 8732
rect 27209 8676 27265 8732
rect 27265 8676 27269 8732
rect 27205 8672 27269 8676
rect 7990 8188 8054 8192
rect 7990 8132 7994 8188
rect 7994 8132 8050 8188
rect 8050 8132 8054 8188
rect 7990 8128 8054 8132
rect 8070 8188 8134 8192
rect 8070 8132 8074 8188
rect 8074 8132 8130 8188
rect 8130 8132 8134 8188
rect 8070 8128 8134 8132
rect 8150 8188 8214 8192
rect 8150 8132 8154 8188
rect 8154 8132 8210 8188
rect 8210 8132 8214 8188
rect 8150 8128 8214 8132
rect 8230 8188 8294 8192
rect 8230 8132 8234 8188
rect 8234 8132 8290 8188
rect 8290 8132 8294 8188
rect 8230 8128 8294 8132
rect 15580 8188 15644 8192
rect 15580 8132 15584 8188
rect 15584 8132 15640 8188
rect 15640 8132 15644 8188
rect 15580 8128 15644 8132
rect 15660 8188 15724 8192
rect 15660 8132 15664 8188
rect 15664 8132 15720 8188
rect 15720 8132 15724 8188
rect 15660 8128 15724 8132
rect 15740 8188 15804 8192
rect 15740 8132 15744 8188
rect 15744 8132 15800 8188
rect 15800 8132 15804 8188
rect 15740 8128 15804 8132
rect 15820 8188 15884 8192
rect 15820 8132 15824 8188
rect 15824 8132 15880 8188
rect 15880 8132 15884 8188
rect 15820 8128 15884 8132
rect 23170 8188 23234 8192
rect 23170 8132 23174 8188
rect 23174 8132 23230 8188
rect 23230 8132 23234 8188
rect 23170 8128 23234 8132
rect 23250 8188 23314 8192
rect 23250 8132 23254 8188
rect 23254 8132 23310 8188
rect 23310 8132 23314 8188
rect 23250 8128 23314 8132
rect 23330 8188 23394 8192
rect 23330 8132 23334 8188
rect 23334 8132 23390 8188
rect 23390 8132 23394 8188
rect 23330 8128 23394 8132
rect 23410 8188 23474 8192
rect 23410 8132 23414 8188
rect 23414 8132 23470 8188
rect 23470 8132 23474 8188
rect 23410 8128 23474 8132
rect 30760 8188 30824 8192
rect 30760 8132 30764 8188
rect 30764 8132 30820 8188
rect 30820 8132 30824 8188
rect 30760 8128 30824 8132
rect 30840 8188 30904 8192
rect 30840 8132 30844 8188
rect 30844 8132 30900 8188
rect 30900 8132 30904 8188
rect 30840 8128 30904 8132
rect 30920 8188 30984 8192
rect 30920 8132 30924 8188
rect 30924 8132 30980 8188
rect 30980 8132 30984 8188
rect 30920 8128 30984 8132
rect 31000 8188 31064 8192
rect 31000 8132 31004 8188
rect 31004 8132 31060 8188
rect 31060 8132 31064 8188
rect 31000 8128 31064 8132
rect 4195 7644 4259 7648
rect 4195 7588 4199 7644
rect 4199 7588 4255 7644
rect 4255 7588 4259 7644
rect 4195 7584 4259 7588
rect 4275 7644 4339 7648
rect 4275 7588 4279 7644
rect 4279 7588 4335 7644
rect 4335 7588 4339 7644
rect 4275 7584 4339 7588
rect 4355 7644 4419 7648
rect 4355 7588 4359 7644
rect 4359 7588 4415 7644
rect 4415 7588 4419 7644
rect 4355 7584 4419 7588
rect 4435 7644 4499 7648
rect 4435 7588 4439 7644
rect 4439 7588 4495 7644
rect 4495 7588 4499 7644
rect 4435 7584 4499 7588
rect 11785 7644 11849 7648
rect 11785 7588 11789 7644
rect 11789 7588 11845 7644
rect 11845 7588 11849 7644
rect 11785 7584 11849 7588
rect 11865 7644 11929 7648
rect 11865 7588 11869 7644
rect 11869 7588 11925 7644
rect 11925 7588 11929 7644
rect 11865 7584 11929 7588
rect 11945 7644 12009 7648
rect 11945 7588 11949 7644
rect 11949 7588 12005 7644
rect 12005 7588 12009 7644
rect 11945 7584 12009 7588
rect 12025 7644 12089 7648
rect 12025 7588 12029 7644
rect 12029 7588 12085 7644
rect 12085 7588 12089 7644
rect 12025 7584 12089 7588
rect 19375 7644 19439 7648
rect 19375 7588 19379 7644
rect 19379 7588 19435 7644
rect 19435 7588 19439 7644
rect 19375 7584 19439 7588
rect 19455 7644 19519 7648
rect 19455 7588 19459 7644
rect 19459 7588 19515 7644
rect 19515 7588 19519 7644
rect 19455 7584 19519 7588
rect 19535 7644 19599 7648
rect 19535 7588 19539 7644
rect 19539 7588 19595 7644
rect 19595 7588 19599 7644
rect 19535 7584 19599 7588
rect 19615 7644 19679 7648
rect 19615 7588 19619 7644
rect 19619 7588 19675 7644
rect 19675 7588 19679 7644
rect 19615 7584 19679 7588
rect 26965 7644 27029 7648
rect 26965 7588 26969 7644
rect 26969 7588 27025 7644
rect 27025 7588 27029 7644
rect 26965 7584 27029 7588
rect 27045 7644 27109 7648
rect 27045 7588 27049 7644
rect 27049 7588 27105 7644
rect 27105 7588 27109 7644
rect 27045 7584 27109 7588
rect 27125 7644 27189 7648
rect 27125 7588 27129 7644
rect 27129 7588 27185 7644
rect 27185 7588 27189 7644
rect 27125 7584 27189 7588
rect 27205 7644 27269 7648
rect 27205 7588 27209 7644
rect 27209 7588 27265 7644
rect 27265 7588 27269 7644
rect 27205 7584 27269 7588
rect 17908 7576 17972 7580
rect 17908 7520 17958 7576
rect 17958 7520 17972 7576
rect 17908 7516 17972 7520
rect 7990 7100 8054 7104
rect 7990 7044 7994 7100
rect 7994 7044 8050 7100
rect 8050 7044 8054 7100
rect 7990 7040 8054 7044
rect 8070 7100 8134 7104
rect 8070 7044 8074 7100
rect 8074 7044 8130 7100
rect 8130 7044 8134 7100
rect 8070 7040 8134 7044
rect 8150 7100 8214 7104
rect 8150 7044 8154 7100
rect 8154 7044 8210 7100
rect 8210 7044 8214 7100
rect 8150 7040 8214 7044
rect 8230 7100 8294 7104
rect 8230 7044 8234 7100
rect 8234 7044 8290 7100
rect 8290 7044 8294 7100
rect 8230 7040 8294 7044
rect 15580 7100 15644 7104
rect 15580 7044 15584 7100
rect 15584 7044 15640 7100
rect 15640 7044 15644 7100
rect 15580 7040 15644 7044
rect 15660 7100 15724 7104
rect 15660 7044 15664 7100
rect 15664 7044 15720 7100
rect 15720 7044 15724 7100
rect 15660 7040 15724 7044
rect 15740 7100 15804 7104
rect 15740 7044 15744 7100
rect 15744 7044 15800 7100
rect 15800 7044 15804 7100
rect 15740 7040 15804 7044
rect 15820 7100 15884 7104
rect 15820 7044 15824 7100
rect 15824 7044 15880 7100
rect 15880 7044 15884 7100
rect 15820 7040 15884 7044
rect 23170 7100 23234 7104
rect 23170 7044 23174 7100
rect 23174 7044 23230 7100
rect 23230 7044 23234 7100
rect 23170 7040 23234 7044
rect 23250 7100 23314 7104
rect 23250 7044 23254 7100
rect 23254 7044 23310 7100
rect 23310 7044 23314 7100
rect 23250 7040 23314 7044
rect 23330 7100 23394 7104
rect 23330 7044 23334 7100
rect 23334 7044 23390 7100
rect 23390 7044 23394 7100
rect 23330 7040 23394 7044
rect 23410 7100 23474 7104
rect 23410 7044 23414 7100
rect 23414 7044 23470 7100
rect 23470 7044 23474 7100
rect 23410 7040 23474 7044
rect 30760 7100 30824 7104
rect 30760 7044 30764 7100
rect 30764 7044 30820 7100
rect 30820 7044 30824 7100
rect 30760 7040 30824 7044
rect 30840 7100 30904 7104
rect 30840 7044 30844 7100
rect 30844 7044 30900 7100
rect 30900 7044 30904 7100
rect 30840 7040 30904 7044
rect 30920 7100 30984 7104
rect 30920 7044 30924 7100
rect 30924 7044 30980 7100
rect 30980 7044 30984 7100
rect 30920 7040 30984 7044
rect 31000 7100 31064 7104
rect 31000 7044 31004 7100
rect 31004 7044 31060 7100
rect 31060 7044 31064 7100
rect 31000 7040 31064 7044
rect 4195 6556 4259 6560
rect 4195 6500 4199 6556
rect 4199 6500 4255 6556
rect 4255 6500 4259 6556
rect 4195 6496 4259 6500
rect 4275 6556 4339 6560
rect 4275 6500 4279 6556
rect 4279 6500 4335 6556
rect 4335 6500 4339 6556
rect 4275 6496 4339 6500
rect 4355 6556 4419 6560
rect 4355 6500 4359 6556
rect 4359 6500 4415 6556
rect 4415 6500 4419 6556
rect 4355 6496 4419 6500
rect 4435 6556 4499 6560
rect 4435 6500 4439 6556
rect 4439 6500 4495 6556
rect 4495 6500 4499 6556
rect 4435 6496 4499 6500
rect 11785 6556 11849 6560
rect 11785 6500 11789 6556
rect 11789 6500 11845 6556
rect 11845 6500 11849 6556
rect 11785 6496 11849 6500
rect 11865 6556 11929 6560
rect 11865 6500 11869 6556
rect 11869 6500 11925 6556
rect 11925 6500 11929 6556
rect 11865 6496 11929 6500
rect 11945 6556 12009 6560
rect 11945 6500 11949 6556
rect 11949 6500 12005 6556
rect 12005 6500 12009 6556
rect 11945 6496 12009 6500
rect 12025 6556 12089 6560
rect 12025 6500 12029 6556
rect 12029 6500 12085 6556
rect 12085 6500 12089 6556
rect 12025 6496 12089 6500
rect 19375 6556 19439 6560
rect 19375 6500 19379 6556
rect 19379 6500 19435 6556
rect 19435 6500 19439 6556
rect 19375 6496 19439 6500
rect 19455 6556 19519 6560
rect 19455 6500 19459 6556
rect 19459 6500 19515 6556
rect 19515 6500 19519 6556
rect 19455 6496 19519 6500
rect 19535 6556 19599 6560
rect 19535 6500 19539 6556
rect 19539 6500 19595 6556
rect 19595 6500 19599 6556
rect 19535 6496 19599 6500
rect 19615 6556 19679 6560
rect 19615 6500 19619 6556
rect 19619 6500 19675 6556
rect 19675 6500 19679 6556
rect 19615 6496 19679 6500
rect 26965 6556 27029 6560
rect 26965 6500 26969 6556
rect 26969 6500 27025 6556
rect 27025 6500 27029 6556
rect 26965 6496 27029 6500
rect 27045 6556 27109 6560
rect 27045 6500 27049 6556
rect 27049 6500 27105 6556
rect 27105 6500 27109 6556
rect 27045 6496 27109 6500
rect 27125 6556 27189 6560
rect 27125 6500 27129 6556
rect 27129 6500 27185 6556
rect 27185 6500 27189 6556
rect 27125 6496 27189 6500
rect 27205 6556 27269 6560
rect 27205 6500 27209 6556
rect 27209 6500 27265 6556
rect 27265 6500 27269 6556
rect 27205 6496 27269 6500
rect 1716 6292 1780 6356
rect 7990 6012 8054 6016
rect 7990 5956 7994 6012
rect 7994 5956 8050 6012
rect 8050 5956 8054 6012
rect 7990 5952 8054 5956
rect 8070 6012 8134 6016
rect 8070 5956 8074 6012
rect 8074 5956 8130 6012
rect 8130 5956 8134 6012
rect 8070 5952 8134 5956
rect 8150 6012 8214 6016
rect 8150 5956 8154 6012
rect 8154 5956 8210 6012
rect 8210 5956 8214 6012
rect 8150 5952 8214 5956
rect 8230 6012 8294 6016
rect 8230 5956 8234 6012
rect 8234 5956 8290 6012
rect 8290 5956 8294 6012
rect 8230 5952 8294 5956
rect 15580 6012 15644 6016
rect 15580 5956 15584 6012
rect 15584 5956 15640 6012
rect 15640 5956 15644 6012
rect 15580 5952 15644 5956
rect 15660 6012 15724 6016
rect 15660 5956 15664 6012
rect 15664 5956 15720 6012
rect 15720 5956 15724 6012
rect 15660 5952 15724 5956
rect 15740 6012 15804 6016
rect 15740 5956 15744 6012
rect 15744 5956 15800 6012
rect 15800 5956 15804 6012
rect 15740 5952 15804 5956
rect 15820 6012 15884 6016
rect 15820 5956 15824 6012
rect 15824 5956 15880 6012
rect 15880 5956 15884 6012
rect 15820 5952 15884 5956
rect 23170 6012 23234 6016
rect 23170 5956 23174 6012
rect 23174 5956 23230 6012
rect 23230 5956 23234 6012
rect 23170 5952 23234 5956
rect 23250 6012 23314 6016
rect 23250 5956 23254 6012
rect 23254 5956 23310 6012
rect 23310 5956 23314 6012
rect 23250 5952 23314 5956
rect 23330 6012 23394 6016
rect 23330 5956 23334 6012
rect 23334 5956 23390 6012
rect 23390 5956 23394 6012
rect 23330 5952 23394 5956
rect 23410 6012 23474 6016
rect 23410 5956 23414 6012
rect 23414 5956 23470 6012
rect 23470 5956 23474 6012
rect 23410 5952 23474 5956
rect 30760 6012 30824 6016
rect 30760 5956 30764 6012
rect 30764 5956 30820 6012
rect 30820 5956 30824 6012
rect 30760 5952 30824 5956
rect 30840 6012 30904 6016
rect 30840 5956 30844 6012
rect 30844 5956 30900 6012
rect 30900 5956 30904 6012
rect 30840 5952 30904 5956
rect 30920 6012 30984 6016
rect 30920 5956 30924 6012
rect 30924 5956 30980 6012
rect 30980 5956 30984 6012
rect 30920 5952 30984 5956
rect 31000 6012 31064 6016
rect 31000 5956 31004 6012
rect 31004 5956 31060 6012
rect 31060 5956 31064 6012
rect 31000 5952 31064 5956
rect 6684 5476 6748 5540
rect 4195 5468 4259 5472
rect 4195 5412 4199 5468
rect 4199 5412 4255 5468
rect 4255 5412 4259 5468
rect 4195 5408 4259 5412
rect 4275 5468 4339 5472
rect 4275 5412 4279 5468
rect 4279 5412 4335 5468
rect 4335 5412 4339 5468
rect 4275 5408 4339 5412
rect 4355 5468 4419 5472
rect 4355 5412 4359 5468
rect 4359 5412 4415 5468
rect 4415 5412 4419 5468
rect 4355 5408 4419 5412
rect 4435 5468 4499 5472
rect 4435 5412 4439 5468
rect 4439 5412 4495 5468
rect 4495 5412 4499 5468
rect 4435 5408 4499 5412
rect 11785 5468 11849 5472
rect 11785 5412 11789 5468
rect 11789 5412 11845 5468
rect 11845 5412 11849 5468
rect 11785 5408 11849 5412
rect 11865 5468 11929 5472
rect 11865 5412 11869 5468
rect 11869 5412 11925 5468
rect 11925 5412 11929 5468
rect 11865 5408 11929 5412
rect 11945 5468 12009 5472
rect 11945 5412 11949 5468
rect 11949 5412 12005 5468
rect 12005 5412 12009 5468
rect 11945 5408 12009 5412
rect 12025 5468 12089 5472
rect 12025 5412 12029 5468
rect 12029 5412 12085 5468
rect 12085 5412 12089 5468
rect 12025 5408 12089 5412
rect 19375 5468 19439 5472
rect 19375 5412 19379 5468
rect 19379 5412 19435 5468
rect 19435 5412 19439 5468
rect 19375 5408 19439 5412
rect 19455 5468 19519 5472
rect 19455 5412 19459 5468
rect 19459 5412 19515 5468
rect 19515 5412 19519 5468
rect 19455 5408 19519 5412
rect 19535 5468 19599 5472
rect 19535 5412 19539 5468
rect 19539 5412 19595 5468
rect 19595 5412 19599 5468
rect 19535 5408 19599 5412
rect 19615 5468 19679 5472
rect 19615 5412 19619 5468
rect 19619 5412 19675 5468
rect 19675 5412 19679 5468
rect 19615 5408 19679 5412
rect 26965 5468 27029 5472
rect 26965 5412 26969 5468
rect 26969 5412 27025 5468
rect 27025 5412 27029 5468
rect 26965 5408 27029 5412
rect 27045 5468 27109 5472
rect 27045 5412 27049 5468
rect 27049 5412 27105 5468
rect 27105 5412 27109 5468
rect 27045 5408 27109 5412
rect 27125 5468 27189 5472
rect 27125 5412 27129 5468
rect 27129 5412 27185 5468
rect 27185 5412 27189 5468
rect 27125 5408 27189 5412
rect 27205 5468 27269 5472
rect 27205 5412 27209 5468
rect 27209 5412 27265 5468
rect 27265 5412 27269 5468
rect 27205 5408 27269 5412
rect 7990 4924 8054 4928
rect 7990 4868 7994 4924
rect 7994 4868 8050 4924
rect 8050 4868 8054 4924
rect 7990 4864 8054 4868
rect 8070 4924 8134 4928
rect 8070 4868 8074 4924
rect 8074 4868 8130 4924
rect 8130 4868 8134 4924
rect 8070 4864 8134 4868
rect 8150 4924 8214 4928
rect 8150 4868 8154 4924
rect 8154 4868 8210 4924
rect 8210 4868 8214 4924
rect 8150 4864 8214 4868
rect 8230 4924 8294 4928
rect 8230 4868 8234 4924
rect 8234 4868 8290 4924
rect 8290 4868 8294 4924
rect 8230 4864 8294 4868
rect 15580 4924 15644 4928
rect 15580 4868 15584 4924
rect 15584 4868 15640 4924
rect 15640 4868 15644 4924
rect 15580 4864 15644 4868
rect 15660 4924 15724 4928
rect 15660 4868 15664 4924
rect 15664 4868 15720 4924
rect 15720 4868 15724 4924
rect 15660 4864 15724 4868
rect 15740 4924 15804 4928
rect 15740 4868 15744 4924
rect 15744 4868 15800 4924
rect 15800 4868 15804 4924
rect 15740 4864 15804 4868
rect 15820 4924 15884 4928
rect 15820 4868 15824 4924
rect 15824 4868 15880 4924
rect 15880 4868 15884 4924
rect 15820 4864 15884 4868
rect 23170 4924 23234 4928
rect 23170 4868 23174 4924
rect 23174 4868 23230 4924
rect 23230 4868 23234 4924
rect 23170 4864 23234 4868
rect 23250 4924 23314 4928
rect 23250 4868 23254 4924
rect 23254 4868 23310 4924
rect 23310 4868 23314 4924
rect 23250 4864 23314 4868
rect 23330 4924 23394 4928
rect 23330 4868 23334 4924
rect 23334 4868 23390 4924
rect 23390 4868 23394 4924
rect 23330 4864 23394 4868
rect 23410 4924 23474 4928
rect 23410 4868 23414 4924
rect 23414 4868 23470 4924
rect 23470 4868 23474 4924
rect 23410 4864 23474 4868
rect 30760 4924 30824 4928
rect 30760 4868 30764 4924
rect 30764 4868 30820 4924
rect 30820 4868 30824 4924
rect 30760 4864 30824 4868
rect 30840 4924 30904 4928
rect 30840 4868 30844 4924
rect 30844 4868 30900 4924
rect 30900 4868 30904 4924
rect 30840 4864 30904 4868
rect 30920 4924 30984 4928
rect 30920 4868 30924 4924
rect 30924 4868 30980 4924
rect 30980 4868 30984 4924
rect 30920 4864 30984 4868
rect 31000 4924 31064 4928
rect 31000 4868 31004 4924
rect 31004 4868 31060 4924
rect 31060 4868 31064 4924
rect 31000 4864 31064 4868
rect 23796 4660 23860 4724
rect 4195 4380 4259 4384
rect 4195 4324 4199 4380
rect 4199 4324 4255 4380
rect 4255 4324 4259 4380
rect 4195 4320 4259 4324
rect 4275 4380 4339 4384
rect 4275 4324 4279 4380
rect 4279 4324 4335 4380
rect 4335 4324 4339 4380
rect 4275 4320 4339 4324
rect 4355 4380 4419 4384
rect 4355 4324 4359 4380
rect 4359 4324 4415 4380
rect 4415 4324 4419 4380
rect 4355 4320 4419 4324
rect 4435 4380 4499 4384
rect 4435 4324 4439 4380
rect 4439 4324 4495 4380
rect 4495 4324 4499 4380
rect 4435 4320 4499 4324
rect 11785 4380 11849 4384
rect 11785 4324 11789 4380
rect 11789 4324 11845 4380
rect 11845 4324 11849 4380
rect 11785 4320 11849 4324
rect 11865 4380 11929 4384
rect 11865 4324 11869 4380
rect 11869 4324 11925 4380
rect 11925 4324 11929 4380
rect 11865 4320 11929 4324
rect 11945 4380 12009 4384
rect 11945 4324 11949 4380
rect 11949 4324 12005 4380
rect 12005 4324 12009 4380
rect 11945 4320 12009 4324
rect 12025 4380 12089 4384
rect 12025 4324 12029 4380
rect 12029 4324 12085 4380
rect 12085 4324 12089 4380
rect 12025 4320 12089 4324
rect 19375 4380 19439 4384
rect 19375 4324 19379 4380
rect 19379 4324 19435 4380
rect 19435 4324 19439 4380
rect 19375 4320 19439 4324
rect 19455 4380 19519 4384
rect 19455 4324 19459 4380
rect 19459 4324 19515 4380
rect 19515 4324 19519 4380
rect 19455 4320 19519 4324
rect 19535 4380 19599 4384
rect 19535 4324 19539 4380
rect 19539 4324 19595 4380
rect 19595 4324 19599 4380
rect 19535 4320 19599 4324
rect 19615 4380 19679 4384
rect 19615 4324 19619 4380
rect 19619 4324 19675 4380
rect 19675 4324 19679 4380
rect 19615 4320 19679 4324
rect 26965 4380 27029 4384
rect 26965 4324 26969 4380
rect 26969 4324 27025 4380
rect 27025 4324 27029 4380
rect 26965 4320 27029 4324
rect 27045 4380 27109 4384
rect 27045 4324 27049 4380
rect 27049 4324 27105 4380
rect 27105 4324 27109 4380
rect 27045 4320 27109 4324
rect 27125 4380 27189 4384
rect 27125 4324 27129 4380
rect 27129 4324 27185 4380
rect 27185 4324 27189 4380
rect 27125 4320 27189 4324
rect 27205 4380 27269 4384
rect 27205 4324 27209 4380
rect 27209 4324 27265 4380
rect 27265 4324 27269 4380
rect 27205 4320 27269 4324
rect 17908 4252 17972 4316
rect 7990 3836 8054 3840
rect 7990 3780 7994 3836
rect 7994 3780 8050 3836
rect 8050 3780 8054 3836
rect 7990 3776 8054 3780
rect 8070 3836 8134 3840
rect 8070 3780 8074 3836
rect 8074 3780 8130 3836
rect 8130 3780 8134 3836
rect 8070 3776 8134 3780
rect 8150 3836 8214 3840
rect 8150 3780 8154 3836
rect 8154 3780 8210 3836
rect 8210 3780 8214 3836
rect 8150 3776 8214 3780
rect 8230 3836 8294 3840
rect 8230 3780 8234 3836
rect 8234 3780 8290 3836
rect 8290 3780 8294 3836
rect 8230 3776 8294 3780
rect 15580 3836 15644 3840
rect 15580 3780 15584 3836
rect 15584 3780 15640 3836
rect 15640 3780 15644 3836
rect 15580 3776 15644 3780
rect 15660 3836 15724 3840
rect 15660 3780 15664 3836
rect 15664 3780 15720 3836
rect 15720 3780 15724 3836
rect 15660 3776 15724 3780
rect 15740 3836 15804 3840
rect 15740 3780 15744 3836
rect 15744 3780 15800 3836
rect 15800 3780 15804 3836
rect 15740 3776 15804 3780
rect 15820 3836 15884 3840
rect 15820 3780 15824 3836
rect 15824 3780 15880 3836
rect 15880 3780 15884 3836
rect 15820 3776 15884 3780
rect 23170 3836 23234 3840
rect 23170 3780 23174 3836
rect 23174 3780 23230 3836
rect 23230 3780 23234 3836
rect 23170 3776 23234 3780
rect 23250 3836 23314 3840
rect 23250 3780 23254 3836
rect 23254 3780 23310 3836
rect 23310 3780 23314 3836
rect 23250 3776 23314 3780
rect 23330 3836 23394 3840
rect 23330 3780 23334 3836
rect 23334 3780 23390 3836
rect 23390 3780 23394 3836
rect 23330 3776 23394 3780
rect 23410 3836 23474 3840
rect 23410 3780 23414 3836
rect 23414 3780 23470 3836
rect 23470 3780 23474 3836
rect 23410 3776 23474 3780
rect 30760 3836 30824 3840
rect 30760 3780 30764 3836
rect 30764 3780 30820 3836
rect 30820 3780 30824 3836
rect 30760 3776 30824 3780
rect 30840 3836 30904 3840
rect 30840 3780 30844 3836
rect 30844 3780 30900 3836
rect 30900 3780 30904 3836
rect 30840 3776 30904 3780
rect 30920 3836 30984 3840
rect 30920 3780 30924 3836
rect 30924 3780 30980 3836
rect 30980 3780 30984 3836
rect 30920 3776 30984 3780
rect 31000 3836 31064 3840
rect 31000 3780 31004 3836
rect 31004 3780 31060 3836
rect 31060 3780 31064 3836
rect 31000 3776 31064 3780
rect 4195 3292 4259 3296
rect 4195 3236 4199 3292
rect 4199 3236 4255 3292
rect 4255 3236 4259 3292
rect 4195 3232 4259 3236
rect 4275 3292 4339 3296
rect 4275 3236 4279 3292
rect 4279 3236 4335 3292
rect 4335 3236 4339 3292
rect 4275 3232 4339 3236
rect 4355 3292 4419 3296
rect 4355 3236 4359 3292
rect 4359 3236 4415 3292
rect 4415 3236 4419 3292
rect 4355 3232 4419 3236
rect 4435 3292 4499 3296
rect 4435 3236 4439 3292
rect 4439 3236 4495 3292
rect 4495 3236 4499 3292
rect 4435 3232 4499 3236
rect 11785 3292 11849 3296
rect 11785 3236 11789 3292
rect 11789 3236 11845 3292
rect 11845 3236 11849 3292
rect 11785 3232 11849 3236
rect 11865 3292 11929 3296
rect 11865 3236 11869 3292
rect 11869 3236 11925 3292
rect 11925 3236 11929 3292
rect 11865 3232 11929 3236
rect 11945 3292 12009 3296
rect 11945 3236 11949 3292
rect 11949 3236 12005 3292
rect 12005 3236 12009 3292
rect 11945 3232 12009 3236
rect 12025 3292 12089 3296
rect 12025 3236 12029 3292
rect 12029 3236 12085 3292
rect 12085 3236 12089 3292
rect 12025 3232 12089 3236
rect 19375 3292 19439 3296
rect 19375 3236 19379 3292
rect 19379 3236 19435 3292
rect 19435 3236 19439 3292
rect 19375 3232 19439 3236
rect 19455 3292 19519 3296
rect 19455 3236 19459 3292
rect 19459 3236 19515 3292
rect 19515 3236 19519 3292
rect 19455 3232 19519 3236
rect 19535 3292 19599 3296
rect 19535 3236 19539 3292
rect 19539 3236 19595 3292
rect 19595 3236 19599 3292
rect 19535 3232 19599 3236
rect 19615 3292 19679 3296
rect 19615 3236 19619 3292
rect 19619 3236 19675 3292
rect 19675 3236 19679 3292
rect 19615 3232 19679 3236
rect 26965 3292 27029 3296
rect 26965 3236 26969 3292
rect 26969 3236 27025 3292
rect 27025 3236 27029 3292
rect 26965 3232 27029 3236
rect 27045 3292 27109 3296
rect 27045 3236 27049 3292
rect 27049 3236 27105 3292
rect 27105 3236 27109 3292
rect 27045 3232 27109 3236
rect 27125 3292 27189 3296
rect 27125 3236 27129 3292
rect 27129 3236 27185 3292
rect 27185 3236 27189 3292
rect 27125 3232 27189 3236
rect 27205 3292 27269 3296
rect 27205 3236 27209 3292
rect 27209 3236 27265 3292
rect 27265 3236 27269 3292
rect 27205 3232 27269 3236
rect 15148 3028 15212 3092
rect 7990 2748 8054 2752
rect 7990 2692 7994 2748
rect 7994 2692 8050 2748
rect 8050 2692 8054 2748
rect 7990 2688 8054 2692
rect 8070 2748 8134 2752
rect 8070 2692 8074 2748
rect 8074 2692 8130 2748
rect 8130 2692 8134 2748
rect 8070 2688 8134 2692
rect 8150 2748 8214 2752
rect 8150 2692 8154 2748
rect 8154 2692 8210 2748
rect 8210 2692 8214 2748
rect 8150 2688 8214 2692
rect 8230 2748 8294 2752
rect 8230 2692 8234 2748
rect 8234 2692 8290 2748
rect 8290 2692 8294 2748
rect 8230 2688 8294 2692
rect 15580 2748 15644 2752
rect 15580 2692 15584 2748
rect 15584 2692 15640 2748
rect 15640 2692 15644 2748
rect 15580 2688 15644 2692
rect 15660 2748 15724 2752
rect 15660 2692 15664 2748
rect 15664 2692 15720 2748
rect 15720 2692 15724 2748
rect 15660 2688 15724 2692
rect 15740 2748 15804 2752
rect 15740 2692 15744 2748
rect 15744 2692 15800 2748
rect 15800 2692 15804 2748
rect 15740 2688 15804 2692
rect 15820 2748 15884 2752
rect 15820 2692 15824 2748
rect 15824 2692 15880 2748
rect 15880 2692 15884 2748
rect 15820 2688 15884 2692
rect 23170 2748 23234 2752
rect 23170 2692 23174 2748
rect 23174 2692 23230 2748
rect 23230 2692 23234 2748
rect 23170 2688 23234 2692
rect 23250 2748 23314 2752
rect 23250 2692 23254 2748
rect 23254 2692 23310 2748
rect 23310 2692 23314 2748
rect 23250 2688 23314 2692
rect 23330 2748 23394 2752
rect 23330 2692 23334 2748
rect 23334 2692 23390 2748
rect 23390 2692 23394 2748
rect 23330 2688 23394 2692
rect 23410 2748 23474 2752
rect 23410 2692 23414 2748
rect 23414 2692 23470 2748
rect 23470 2692 23474 2748
rect 23410 2688 23474 2692
rect 30760 2748 30824 2752
rect 30760 2692 30764 2748
rect 30764 2692 30820 2748
rect 30820 2692 30824 2748
rect 30760 2688 30824 2692
rect 30840 2748 30904 2752
rect 30840 2692 30844 2748
rect 30844 2692 30900 2748
rect 30900 2692 30904 2748
rect 30840 2688 30904 2692
rect 30920 2748 30984 2752
rect 30920 2692 30924 2748
rect 30924 2692 30980 2748
rect 30980 2692 30984 2748
rect 30920 2688 30984 2692
rect 31000 2748 31064 2752
rect 31000 2692 31004 2748
rect 31004 2692 31060 2748
rect 31060 2692 31064 2748
rect 31000 2688 31064 2692
rect 24716 2484 24780 2548
rect 15148 2348 15212 2412
rect 4195 2204 4259 2208
rect 4195 2148 4199 2204
rect 4199 2148 4255 2204
rect 4255 2148 4259 2204
rect 4195 2144 4259 2148
rect 4275 2204 4339 2208
rect 4275 2148 4279 2204
rect 4279 2148 4335 2204
rect 4335 2148 4339 2204
rect 4275 2144 4339 2148
rect 4355 2204 4419 2208
rect 4355 2148 4359 2204
rect 4359 2148 4415 2204
rect 4415 2148 4419 2204
rect 4355 2144 4419 2148
rect 4435 2204 4499 2208
rect 4435 2148 4439 2204
rect 4439 2148 4495 2204
rect 4495 2148 4499 2204
rect 4435 2144 4499 2148
rect 11785 2204 11849 2208
rect 11785 2148 11789 2204
rect 11789 2148 11845 2204
rect 11845 2148 11849 2204
rect 11785 2144 11849 2148
rect 11865 2204 11929 2208
rect 11865 2148 11869 2204
rect 11869 2148 11925 2204
rect 11925 2148 11929 2204
rect 11865 2144 11929 2148
rect 11945 2204 12009 2208
rect 11945 2148 11949 2204
rect 11949 2148 12005 2204
rect 12005 2148 12009 2204
rect 11945 2144 12009 2148
rect 12025 2204 12089 2208
rect 12025 2148 12029 2204
rect 12029 2148 12085 2204
rect 12085 2148 12089 2204
rect 12025 2144 12089 2148
rect 19375 2204 19439 2208
rect 19375 2148 19379 2204
rect 19379 2148 19435 2204
rect 19435 2148 19439 2204
rect 19375 2144 19439 2148
rect 19455 2204 19519 2208
rect 19455 2148 19459 2204
rect 19459 2148 19515 2204
rect 19515 2148 19519 2204
rect 19455 2144 19519 2148
rect 19535 2204 19599 2208
rect 19535 2148 19539 2204
rect 19539 2148 19595 2204
rect 19595 2148 19599 2204
rect 19535 2144 19599 2148
rect 19615 2204 19679 2208
rect 19615 2148 19619 2204
rect 19619 2148 19675 2204
rect 19675 2148 19679 2204
rect 19615 2144 19679 2148
rect 26965 2204 27029 2208
rect 26965 2148 26969 2204
rect 26969 2148 27025 2204
rect 27025 2148 27029 2204
rect 26965 2144 27029 2148
rect 27045 2204 27109 2208
rect 27045 2148 27049 2204
rect 27049 2148 27105 2204
rect 27105 2148 27109 2204
rect 27045 2144 27109 2148
rect 27125 2204 27189 2208
rect 27125 2148 27129 2204
rect 27129 2148 27185 2204
rect 27185 2148 27189 2204
rect 27125 2144 27189 2148
rect 27205 2204 27269 2208
rect 27205 2148 27209 2204
rect 27209 2148 27265 2204
rect 27265 2148 27269 2204
rect 27205 2144 27269 2148
rect 5580 2000 5644 2004
rect 5580 1944 5594 2000
rect 5594 1944 5644 2000
rect 5580 1940 5644 1944
rect 7990 1660 8054 1664
rect 7990 1604 7994 1660
rect 7994 1604 8050 1660
rect 8050 1604 8054 1660
rect 7990 1600 8054 1604
rect 8070 1660 8134 1664
rect 8070 1604 8074 1660
rect 8074 1604 8130 1660
rect 8130 1604 8134 1660
rect 8070 1600 8134 1604
rect 8150 1660 8214 1664
rect 8150 1604 8154 1660
rect 8154 1604 8210 1660
rect 8210 1604 8214 1660
rect 8150 1600 8214 1604
rect 8230 1660 8294 1664
rect 8230 1604 8234 1660
rect 8234 1604 8290 1660
rect 8290 1604 8294 1660
rect 8230 1600 8294 1604
rect 15580 1660 15644 1664
rect 15580 1604 15584 1660
rect 15584 1604 15640 1660
rect 15640 1604 15644 1660
rect 15580 1600 15644 1604
rect 15660 1660 15724 1664
rect 15660 1604 15664 1660
rect 15664 1604 15720 1660
rect 15720 1604 15724 1660
rect 15660 1600 15724 1604
rect 15740 1660 15804 1664
rect 15740 1604 15744 1660
rect 15744 1604 15800 1660
rect 15800 1604 15804 1660
rect 15740 1600 15804 1604
rect 15820 1660 15884 1664
rect 15820 1604 15824 1660
rect 15824 1604 15880 1660
rect 15880 1604 15884 1660
rect 15820 1600 15884 1604
rect 23170 1660 23234 1664
rect 23170 1604 23174 1660
rect 23174 1604 23230 1660
rect 23230 1604 23234 1660
rect 23170 1600 23234 1604
rect 23250 1660 23314 1664
rect 23250 1604 23254 1660
rect 23254 1604 23310 1660
rect 23310 1604 23314 1660
rect 23250 1600 23314 1604
rect 23330 1660 23394 1664
rect 23330 1604 23334 1660
rect 23334 1604 23390 1660
rect 23390 1604 23394 1660
rect 23330 1600 23394 1604
rect 23410 1660 23474 1664
rect 23410 1604 23414 1660
rect 23414 1604 23470 1660
rect 23470 1604 23474 1660
rect 23410 1600 23474 1604
rect 30760 1660 30824 1664
rect 30760 1604 30764 1660
rect 30764 1604 30820 1660
rect 30820 1604 30824 1660
rect 30760 1600 30824 1604
rect 30840 1660 30904 1664
rect 30840 1604 30844 1660
rect 30844 1604 30900 1660
rect 30900 1604 30904 1660
rect 30840 1600 30904 1604
rect 30920 1660 30984 1664
rect 30920 1604 30924 1660
rect 30924 1604 30980 1660
rect 30980 1604 30984 1660
rect 30920 1600 30984 1604
rect 31000 1660 31064 1664
rect 31000 1604 31004 1660
rect 31004 1604 31060 1660
rect 31060 1604 31064 1660
rect 31000 1600 31064 1604
rect 6684 1320 6748 1324
rect 6684 1264 6734 1320
rect 6734 1264 6748 1320
rect 6684 1260 6748 1264
rect 23796 1124 23860 1188
rect 4195 1116 4259 1120
rect 4195 1060 4199 1116
rect 4199 1060 4255 1116
rect 4255 1060 4259 1116
rect 4195 1056 4259 1060
rect 4275 1116 4339 1120
rect 4275 1060 4279 1116
rect 4279 1060 4335 1116
rect 4335 1060 4339 1116
rect 4275 1056 4339 1060
rect 4355 1116 4419 1120
rect 4355 1060 4359 1116
rect 4359 1060 4415 1116
rect 4415 1060 4419 1116
rect 4355 1056 4419 1060
rect 4435 1116 4499 1120
rect 4435 1060 4439 1116
rect 4439 1060 4495 1116
rect 4495 1060 4499 1116
rect 4435 1056 4499 1060
rect 11785 1116 11849 1120
rect 11785 1060 11789 1116
rect 11789 1060 11845 1116
rect 11845 1060 11849 1116
rect 11785 1056 11849 1060
rect 11865 1116 11929 1120
rect 11865 1060 11869 1116
rect 11869 1060 11925 1116
rect 11925 1060 11929 1116
rect 11865 1056 11929 1060
rect 11945 1116 12009 1120
rect 11945 1060 11949 1116
rect 11949 1060 12005 1116
rect 12005 1060 12009 1116
rect 11945 1056 12009 1060
rect 12025 1116 12089 1120
rect 12025 1060 12029 1116
rect 12029 1060 12085 1116
rect 12085 1060 12089 1116
rect 12025 1056 12089 1060
rect 19375 1116 19439 1120
rect 19375 1060 19379 1116
rect 19379 1060 19435 1116
rect 19435 1060 19439 1116
rect 19375 1056 19439 1060
rect 19455 1116 19519 1120
rect 19455 1060 19459 1116
rect 19459 1060 19515 1116
rect 19515 1060 19519 1116
rect 19455 1056 19519 1060
rect 19535 1116 19599 1120
rect 19535 1060 19539 1116
rect 19539 1060 19595 1116
rect 19595 1060 19599 1116
rect 19535 1056 19599 1060
rect 19615 1116 19679 1120
rect 19615 1060 19619 1116
rect 19619 1060 19675 1116
rect 19675 1060 19679 1116
rect 19615 1056 19679 1060
rect 26965 1116 27029 1120
rect 26965 1060 26969 1116
rect 26969 1060 27025 1116
rect 27025 1060 27029 1116
rect 26965 1056 27029 1060
rect 27045 1116 27109 1120
rect 27045 1060 27049 1116
rect 27049 1060 27105 1116
rect 27105 1060 27109 1116
rect 27045 1056 27109 1060
rect 27125 1116 27189 1120
rect 27125 1060 27129 1116
rect 27129 1060 27185 1116
rect 27185 1060 27189 1116
rect 27125 1056 27189 1060
rect 27205 1116 27269 1120
rect 27205 1060 27209 1116
rect 27209 1060 27265 1116
rect 27265 1060 27269 1116
rect 27205 1056 27269 1060
rect 24716 852 24780 916
rect 7990 572 8054 576
rect 7990 516 7994 572
rect 7994 516 8050 572
rect 8050 516 8054 572
rect 7990 512 8054 516
rect 8070 572 8134 576
rect 8070 516 8074 572
rect 8074 516 8130 572
rect 8130 516 8134 572
rect 8070 512 8134 516
rect 8150 572 8214 576
rect 8150 516 8154 572
rect 8154 516 8210 572
rect 8210 516 8214 572
rect 8150 512 8214 516
rect 8230 572 8294 576
rect 8230 516 8234 572
rect 8234 516 8290 572
rect 8290 516 8294 572
rect 8230 512 8294 516
rect 15580 572 15644 576
rect 15580 516 15584 572
rect 15584 516 15640 572
rect 15640 516 15644 572
rect 15580 512 15644 516
rect 15660 572 15724 576
rect 15660 516 15664 572
rect 15664 516 15720 572
rect 15720 516 15724 572
rect 15660 512 15724 516
rect 15740 572 15804 576
rect 15740 516 15744 572
rect 15744 516 15800 572
rect 15800 516 15804 572
rect 15740 512 15804 516
rect 15820 572 15884 576
rect 15820 516 15824 572
rect 15824 516 15880 572
rect 15880 516 15884 572
rect 15820 512 15884 516
rect 23170 572 23234 576
rect 23170 516 23174 572
rect 23174 516 23230 572
rect 23230 516 23234 572
rect 23170 512 23234 516
rect 23250 572 23314 576
rect 23250 516 23254 572
rect 23254 516 23310 572
rect 23310 516 23314 572
rect 23250 512 23314 516
rect 23330 572 23394 576
rect 23330 516 23334 572
rect 23334 516 23390 572
rect 23390 516 23394 572
rect 23330 512 23394 516
rect 23410 572 23474 576
rect 23410 516 23414 572
rect 23414 516 23470 572
rect 23470 516 23474 572
rect 23410 512 23474 516
rect 30760 572 30824 576
rect 30760 516 30764 572
rect 30764 516 30820 572
rect 30820 516 30824 572
rect 30760 512 30824 516
rect 30840 572 30904 576
rect 30840 516 30844 572
rect 30844 516 30900 572
rect 30900 516 30904 572
rect 30840 512 30904 516
rect 30920 572 30984 576
rect 30920 516 30924 572
rect 30924 516 30980 572
rect 30980 516 30984 572
rect 30920 512 30984 516
rect 31000 572 31064 576
rect 31000 516 31004 572
rect 31004 516 31060 572
rect 31060 516 31064 572
rect 31000 512 31064 516
<< metal4 >>
rect 4294 22130 4354 22304
rect 4478 22174 4722 22234
rect 4478 22130 4538 22174
rect 4294 22070 4538 22130
rect 4187 21792 4507 21808
rect 4187 21728 4195 21792
rect 4259 21728 4275 21792
rect 4339 21728 4355 21792
rect 4419 21728 4435 21792
rect 4499 21728 4507 21792
rect 4187 20704 4507 21728
rect 4187 20640 4195 20704
rect 4259 20640 4275 20704
rect 4339 20640 4355 20704
rect 4419 20640 4435 20704
rect 4499 20640 4507 20704
rect 4187 19616 4507 20640
rect 4187 19552 4195 19616
rect 4259 19552 4275 19616
rect 4339 19552 4355 19616
rect 4419 19552 4435 19616
rect 4499 19552 4507 19616
rect 3739 19004 3805 19005
rect 3739 18940 3740 19004
rect 3804 18940 3805 19004
rect 3739 18939 3805 18940
rect 1715 13836 1781 13837
rect 1715 13772 1716 13836
rect 1780 13772 1781 13836
rect 1715 13771 1781 13772
rect 1718 6357 1778 13771
rect 3742 12477 3802 18939
rect 4187 18528 4507 19552
rect 4187 18464 4195 18528
rect 4259 18464 4275 18528
rect 4339 18464 4355 18528
rect 4419 18464 4435 18528
rect 4499 18464 4507 18528
rect 3923 18052 3989 18053
rect 3923 17988 3924 18052
rect 3988 17988 3989 18052
rect 3923 17987 3989 17988
rect 3739 12476 3805 12477
rect 3739 12412 3740 12476
rect 3804 12412 3805 12476
rect 3739 12411 3805 12412
rect 3926 10165 3986 17987
rect 4187 17440 4507 18464
rect 4662 18189 4722 22174
rect 4659 18188 4725 18189
rect 4659 18124 4660 18188
rect 4724 18124 4725 18188
rect 4659 18123 4725 18124
rect 4846 18053 4906 22304
rect 5398 18053 5458 22304
rect 5950 18053 6010 22304
rect 4843 18052 4909 18053
rect 4843 17988 4844 18052
rect 4908 17988 4909 18052
rect 4843 17987 4909 17988
rect 5395 18052 5461 18053
rect 5395 17988 5396 18052
rect 5460 17988 5461 18052
rect 5395 17987 5461 17988
rect 5947 18052 6013 18053
rect 5947 17988 5948 18052
rect 6012 17988 6013 18052
rect 5947 17987 6013 17988
rect 4187 17376 4195 17440
rect 4259 17376 4275 17440
rect 4339 17376 4355 17440
rect 4419 17376 4435 17440
rect 4499 17376 4507 17440
rect 4187 16352 4507 17376
rect 4187 16288 4195 16352
rect 4259 16288 4275 16352
rect 4339 16288 4355 16352
rect 4419 16288 4435 16352
rect 4499 16288 4507 16352
rect 4187 15264 4507 16288
rect 4187 15200 4195 15264
rect 4259 15200 4275 15264
rect 4339 15200 4355 15264
rect 4419 15200 4435 15264
rect 4499 15200 4507 15264
rect 4187 14176 4507 15200
rect 4187 14112 4195 14176
rect 4259 14112 4275 14176
rect 4339 14112 4355 14176
rect 4419 14112 4435 14176
rect 4499 14112 4507 14176
rect 4187 13088 4507 14112
rect 6502 13701 6562 22304
rect 6683 19412 6749 19413
rect 6683 19348 6684 19412
rect 6748 19348 6749 19412
rect 6683 19347 6749 19348
rect 6499 13700 6565 13701
rect 6499 13636 6500 13700
rect 6564 13636 6565 13700
rect 6499 13635 6565 13636
rect 4187 13024 4195 13088
rect 4259 13024 4275 13088
rect 4339 13024 4355 13088
rect 4419 13024 4435 13088
rect 4499 13024 4507 13088
rect 4187 12000 4507 13024
rect 6686 12205 6746 19347
rect 7054 18325 7114 22304
rect 7051 18324 7117 18325
rect 7051 18260 7052 18324
rect 7116 18260 7117 18324
rect 7051 18259 7117 18260
rect 7606 13293 7666 22304
rect 7790 22174 8034 22234
rect 7790 18597 7850 22174
rect 7974 22130 8034 22174
rect 8158 22130 8218 22304
rect 7974 22070 8218 22130
rect 8710 21997 8770 22304
rect 8707 21996 8773 21997
rect 8707 21932 8708 21996
rect 8772 21932 8773 21996
rect 8707 21931 8773 21932
rect 9262 21861 9322 22304
rect 9259 21860 9325 21861
rect 7982 21248 8302 21808
rect 9259 21796 9260 21860
rect 9324 21796 9325 21860
rect 9259 21795 9325 21796
rect 7982 21184 7990 21248
rect 8054 21184 8070 21248
rect 8134 21184 8150 21248
rect 8214 21184 8230 21248
rect 8294 21184 8302 21248
rect 7982 20160 8302 21184
rect 8891 20772 8957 20773
rect 8891 20708 8892 20772
rect 8956 20708 8957 20772
rect 8891 20707 8957 20708
rect 7982 20096 7990 20160
rect 8054 20096 8070 20160
rect 8134 20096 8150 20160
rect 8214 20096 8230 20160
rect 8294 20096 8302 20160
rect 7982 19072 8302 20096
rect 7982 19008 7990 19072
rect 8054 19008 8070 19072
rect 8134 19008 8150 19072
rect 8214 19008 8230 19072
rect 8294 19008 8302 19072
rect 7787 18596 7853 18597
rect 7787 18532 7788 18596
rect 7852 18532 7853 18596
rect 7787 18531 7853 18532
rect 7787 18052 7853 18053
rect 7787 17988 7788 18052
rect 7852 17988 7853 18052
rect 7787 17987 7853 17988
rect 7603 13292 7669 13293
rect 7603 13228 7604 13292
rect 7668 13228 7669 13292
rect 7603 13227 7669 13228
rect 6683 12204 6749 12205
rect 6683 12140 6684 12204
rect 6748 12140 6749 12204
rect 6683 12139 6749 12140
rect 4187 11936 4195 12000
rect 4259 11936 4275 12000
rect 4339 11936 4355 12000
rect 4419 11936 4435 12000
rect 4499 11936 4507 12000
rect 4187 10912 4507 11936
rect 7790 11661 7850 17987
rect 7982 17984 8302 19008
rect 7982 17920 7990 17984
rect 8054 17920 8070 17984
rect 8134 17920 8150 17984
rect 8214 17920 8230 17984
rect 8294 17920 8302 17984
rect 7982 16896 8302 17920
rect 8523 17508 8589 17509
rect 8523 17444 8524 17508
rect 8588 17444 8589 17508
rect 8523 17443 8589 17444
rect 7982 16832 7990 16896
rect 8054 16832 8070 16896
rect 8134 16832 8150 16896
rect 8214 16832 8230 16896
rect 8294 16832 8302 16896
rect 7982 15808 8302 16832
rect 7982 15744 7990 15808
rect 8054 15744 8070 15808
rect 8134 15744 8150 15808
rect 8214 15744 8230 15808
rect 8294 15744 8302 15808
rect 7982 14720 8302 15744
rect 7982 14656 7990 14720
rect 8054 14656 8070 14720
rect 8134 14656 8150 14720
rect 8214 14656 8230 14720
rect 8294 14656 8302 14720
rect 7982 13632 8302 14656
rect 7982 13568 7990 13632
rect 8054 13568 8070 13632
rect 8134 13568 8150 13632
rect 8214 13568 8230 13632
rect 8294 13568 8302 13632
rect 7982 12544 8302 13568
rect 8526 13565 8586 17443
rect 8523 13564 8589 13565
rect 8523 13500 8524 13564
rect 8588 13500 8589 13564
rect 8523 13499 8589 13500
rect 7982 12480 7990 12544
rect 8054 12480 8070 12544
rect 8134 12480 8150 12544
rect 8214 12480 8230 12544
rect 8294 12480 8302 12544
rect 7787 11660 7853 11661
rect 7787 11596 7788 11660
rect 7852 11596 7853 11660
rect 7787 11595 7853 11596
rect 4187 10848 4195 10912
rect 4259 10848 4275 10912
rect 4339 10848 4355 10912
rect 4419 10848 4435 10912
rect 4499 10848 4507 10912
rect 3923 10164 3989 10165
rect 3923 10100 3924 10164
rect 3988 10100 3989 10164
rect 3923 10099 3989 10100
rect 4187 9824 4507 10848
rect 7982 11456 8302 12480
rect 8894 12341 8954 20707
rect 9814 20501 9874 22304
rect 10179 22132 10245 22133
rect 10179 22068 10180 22132
rect 10244 22130 10245 22132
rect 10366 22130 10426 22304
rect 10244 22070 10426 22130
rect 10244 22068 10245 22070
rect 10179 22067 10245 22068
rect 10918 20637 10978 22304
rect 11470 21589 11530 22304
rect 12022 22130 12082 22304
rect 12022 22070 12266 22130
rect 11777 21792 12097 21808
rect 11777 21728 11785 21792
rect 11849 21728 11865 21792
rect 11929 21728 11945 21792
rect 12009 21728 12025 21792
rect 12089 21728 12097 21792
rect 11467 21588 11533 21589
rect 11467 21524 11468 21588
rect 11532 21524 11533 21588
rect 11467 21523 11533 21524
rect 11283 21180 11349 21181
rect 11283 21116 11284 21180
rect 11348 21116 11349 21180
rect 11283 21115 11349 21116
rect 11099 20908 11165 20909
rect 11099 20844 11100 20908
rect 11164 20844 11165 20908
rect 11099 20843 11165 20844
rect 10915 20636 10981 20637
rect 10915 20572 10916 20636
rect 10980 20572 10981 20636
rect 10915 20571 10981 20572
rect 9811 20500 9877 20501
rect 9811 20436 9812 20500
rect 9876 20436 9877 20500
rect 9811 20435 9877 20436
rect 10363 18732 10429 18733
rect 10363 18668 10364 18732
rect 10428 18668 10429 18732
rect 10363 18667 10429 18668
rect 9627 15740 9693 15741
rect 9627 15676 9628 15740
rect 9692 15676 9693 15740
rect 9627 15675 9693 15676
rect 8891 12340 8957 12341
rect 8891 12276 8892 12340
rect 8956 12276 8957 12340
rect 8891 12275 8957 12276
rect 7982 11392 7990 11456
rect 8054 11392 8070 11456
rect 8134 11392 8150 11456
rect 8214 11392 8230 11456
rect 8294 11392 8302 11456
rect 5579 10572 5645 10573
rect 5579 10508 5580 10572
rect 5644 10508 5645 10572
rect 5579 10507 5645 10508
rect 4187 9760 4195 9824
rect 4259 9760 4275 9824
rect 4339 9760 4355 9824
rect 4419 9760 4435 9824
rect 4499 9760 4507 9824
rect 4187 8736 4507 9760
rect 4187 8672 4195 8736
rect 4259 8672 4275 8736
rect 4339 8672 4355 8736
rect 4419 8672 4435 8736
rect 4499 8672 4507 8736
rect 4187 7648 4507 8672
rect 4187 7584 4195 7648
rect 4259 7584 4275 7648
rect 4339 7584 4355 7648
rect 4419 7584 4435 7648
rect 4499 7584 4507 7648
rect 4187 6560 4507 7584
rect 4187 6496 4195 6560
rect 4259 6496 4275 6560
rect 4339 6496 4355 6560
rect 4419 6496 4435 6560
rect 4499 6496 4507 6560
rect 1715 6356 1781 6357
rect 1715 6292 1716 6356
rect 1780 6292 1781 6356
rect 1715 6291 1781 6292
rect 4187 5472 4507 6496
rect 4187 5408 4195 5472
rect 4259 5408 4275 5472
rect 4339 5408 4355 5472
rect 4419 5408 4435 5472
rect 4499 5408 4507 5472
rect 4187 4384 4507 5408
rect 4187 4320 4195 4384
rect 4259 4320 4275 4384
rect 4339 4320 4355 4384
rect 4419 4320 4435 4384
rect 4499 4320 4507 4384
rect 4187 3296 4507 4320
rect 4187 3232 4195 3296
rect 4259 3232 4275 3296
rect 4339 3232 4355 3296
rect 4419 3232 4435 3296
rect 4499 3232 4507 3296
rect 4187 2208 4507 3232
rect 4187 2144 4195 2208
rect 4259 2144 4275 2208
rect 4339 2144 4355 2208
rect 4419 2144 4435 2208
rect 4499 2144 4507 2208
rect 4187 1120 4507 2144
rect 5582 2005 5642 10507
rect 7982 10368 8302 11392
rect 9630 10709 9690 15675
rect 10366 14245 10426 18667
rect 10731 18324 10797 18325
rect 10731 18260 10732 18324
rect 10796 18260 10797 18324
rect 10731 18259 10797 18260
rect 10547 17372 10613 17373
rect 10547 17308 10548 17372
rect 10612 17308 10613 17372
rect 10547 17307 10613 17308
rect 10550 15197 10610 17307
rect 10547 15196 10613 15197
rect 10547 15132 10548 15196
rect 10612 15132 10613 15196
rect 10547 15131 10613 15132
rect 10363 14244 10429 14245
rect 10363 14180 10364 14244
rect 10428 14180 10429 14244
rect 10363 14179 10429 14180
rect 10734 11797 10794 18259
rect 11102 13837 11162 20843
rect 11099 13836 11165 13837
rect 11099 13772 11100 13836
rect 11164 13772 11165 13836
rect 11099 13771 11165 13772
rect 11286 13021 11346 21115
rect 11777 20704 12097 21728
rect 12206 21589 12266 22070
rect 12574 21997 12634 22304
rect 12571 21996 12637 21997
rect 12571 21932 12572 21996
rect 12636 21932 12637 21996
rect 12571 21931 12637 21932
rect 12203 21588 12269 21589
rect 12203 21524 12204 21588
rect 12268 21524 12269 21588
rect 12203 21523 12269 21524
rect 13126 21317 13186 22304
rect 13123 21316 13189 21317
rect 13123 21252 13124 21316
rect 13188 21252 13189 21316
rect 13123 21251 13189 21252
rect 11777 20640 11785 20704
rect 11849 20640 11865 20704
rect 11929 20640 11945 20704
rect 12009 20640 12025 20704
rect 12089 20640 12097 20704
rect 11777 19616 12097 20640
rect 13678 20637 13738 22304
rect 13862 22174 14106 22234
rect 13862 21997 13922 22174
rect 14046 22130 14106 22174
rect 14230 22130 14290 22304
rect 14046 22070 14290 22130
rect 14411 22132 14477 22133
rect 14411 22068 14412 22132
rect 14476 22130 14477 22132
rect 14782 22130 14842 22304
rect 14476 22070 14842 22130
rect 14476 22068 14477 22070
rect 14411 22067 14477 22068
rect 13859 21996 13925 21997
rect 13859 21932 13860 21996
rect 13924 21932 13925 21996
rect 13859 21931 13925 21932
rect 13675 20636 13741 20637
rect 13675 20572 13676 20636
rect 13740 20572 13741 20636
rect 13675 20571 13741 20572
rect 11777 19552 11785 19616
rect 11849 19552 11865 19616
rect 11929 19552 11945 19616
rect 12009 19552 12025 19616
rect 12089 19552 12097 19616
rect 11777 18528 12097 19552
rect 15334 19277 15394 22304
rect 15886 22130 15946 22304
rect 15886 22070 16130 22130
rect 15572 21248 15892 21808
rect 15572 21184 15580 21248
rect 15644 21184 15660 21248
rect 15724 21184 15740 21248
rect 15804 21184 15820 21248
rect 15884 21184 15892 21248
rect 15572 20160 15892 21184
rect 16070 20501 16130 22070
rect 16067 20500 16133 20501
rect 16067 20436 16068 20500
rect 16132 20436 16133 20500
rect 16067 20435 16133 20436
rect 15572 20096 15580 20160
rect 15644 20096 15660 20160
rect 15724 20096 15740 20160
rect 15804 20096 15820 20160
rect 15884 20096 15892 20160
rect 15331 19276 15397 19277
rect 15331 19212 15332 19276
rect 15396 19212 15397 19276
rect 15331 19211 15397 19212
rect 11777 18464 11785 18528
rect 11849 18464 11865 18528
rect 11929 18464 11945 18528
rect 12009 18464 12025 18528
rect 12089 18464 12097 18528
rect 11651 17916 11717 17917
rect 11651 17852 11652 17916
rect 11716 17852 11717 17916
rect 11651 17851 11717 17852
rect 11467 17236 11533 17237
rect 11467 17172 11468 17236
rect 11532 17172 11533 17236
rect 11467 17171 11533 17172
rect 11470 13021 11530 17171
rect 11283 13020 11349 13021
rect 11283 12956 11284 13020
rect 11348 12956 11349 13020
rect 11283 12955 11349 12956
rect 11467 13020 11533 13021
rect 11467 12956 11468 13020
rect 11532 12956 11533 13020
rect 11467 12955 11533 12956
rect 11654 11797 11714 17851
rect 11777 17440 12097 18464
rect 15572 19072 15892 20096
rect 16438 19277 16498 22304
rect 16990 21589 17050 22304
rect 17542 22104 17602 22304
rect 18094 22104 18154 22304
rect 18646 22104 18706 22304
rect 19198 22104 19258 22304
rect 19750 22104 19810 22304
rect 20302 22104 20362 22304
rect 20854 22104 20914 22304
rect 21406 22104 21466 22304
rect 19367 21792 19687 21808
rect 19367 21728 19375 21792
rect 19439 21728 19455 21792
rect 19519 21728 19535 21792
rect 19599 21728 19615 21792
rect 19679 21728 19687 21792
rect 16987 21588 17053 21589
rect 16987 21524 16988 21588
rect 17052 21524 17053 21588
rect 16987 21523 17053 21524
rect 19367 20704 19687 21728
rect 19367 20640 19375 20704
rect 19439 20640 19455 20704
rect 19519 20640 19535 20704
rect 19599 20640 19615 20704
rect 19679 20640 19687 20704
rect 19367 19616 19687 20640
rect 19367 19552 19375 19616
rect 19439 19552 19455 19616
rect 19519 19552 19535 19616
rect 19599 19552 19615 19616
rect 19679 19552 19687 19616
rect 16435 19276 16501 19277
rect 16435 19212 16436 19276
rect 16500 19212 16501 19276
rect 16435 19211 16501 19212
rect 15572 19008 15580 19072
rect 15644 19008 15660 19072
rect 15724 19008 15740 19072
rect 15804 19008 15820 19072
rect 15884 19008 15892 19072
rect 13491 18188 13557 18189
rect 13491 18124 13492 18188
rect 13556 18124 13557 18188
rect 13491 18123 13557 18124
rect 11777 17376 11785 17440
rect 11849 17376 11865 17440
rect 11929 17376 11945 17440
rect 12009 17376 12025 17440
rect 12089 17376 12097 17440
rect 11777 16352 12097 17376
rect 11777 16288 11785 16352
rect 11849 16288 11865 16352
rect 11929 16288 11945 16352
rect 12009 16288 12025 16352
rect 12089 16288 12097 16352
rect 11777 15264 12097 16288
rect 11777 15200 11785 15264
rect 11849 15200 11865 15264
rect 11929 15200 11945 15264
rect 12009 15200 12025 15264
rect 12089 15200 12097 15264
rect 11777 14176 12097 15200
rect 12203 14924 12269 14925
rect 12203 14860 12204 14924
rect 12268 14860 12269 14924
rect 12203 14859 12269 14860
rect 12206 14245 12266 14859
rect 12203 14244 12269 14245
rect 12203 14180 12204 14244
rect 12268 14180 12269 14244
rect 12203 14179 12269 14180
rect 11777 14112 11785 14176
rect 11849 14112 11865 14176
rect 11929 14112 11945 14176
rect 12009 14112 12025 14176
rect 12089 14112 12097 14176
rect 11777 13088 12097 14112
rect 12387 13428 12453 13429
rect 12387 13364 12388 13428
rect 12452 13364 12453 13428
rect 12387 13363 12453 13364
rect 11777 13024 11785 13088
rect 11849 13024 11865 13088
rect 11929 13024 11945 13088
rect 12009 13024 12025 13088
rect 12089 13024 12097 13088
rect 11777 12000 12097 13024
rect 12390 13021 12450 13363
rect 12387 13020 12453 13021
rect 12387 12956 12388 13020
rect 12452 12956 12453 13020
rect 12387 12955 12453 12956
rect 13494 12477 13554 18123
rect 15572 17984 15892 19008
rect 15572 17920 15580 17984
rect 15644 17920 15660 17984
rect 15724 17920 15740 17984
rect 15804 17920 15820 17984
rect 15884 17920 15892 17984
rect 15572 16896 15892 17920
rect 15572 16832 15580 16896
rect 15644 16832 15660 16896
rect 15724 16832 15740 16896
rect 15804 16832 15820 16896
rect 15884 16832 15892 16896
rect 15572 15808 15892 16832
rect 15572 15744 15580 15808
rect 15644 15744 15660 15808
rect 15724 15744 15740 15808
rect 15804 15744 15820 15808
rect 15884 15744 15892 15808
rect 15572 14720 15892 15744
rect 15572 14656 15580 14720
rect 15644 14656 15660 14720
rect 15724 14656 15740 14720
rect 15804 14656 15820 14720
rect 15884 14656 15892 14720
rect 15572 13632 15892 14656
rect 15572 13568 15580 13632
rect 15644 13568 15660 13632
rect 15724 13568 15740 13632
rect 15804 13568 15820 13632
rect 15884 13568 15892 13632
rect 15572 12544 15892 13568
rect 15572 12480 15580 12544
rect 15644 12480 15660 12544
rect 15724 12480 15740 12544
rect 15804 12480 15820 12544
rect 15884 12480 15892 12544
rect 13491 12476 13557 12477
rect 13491 12412 13492 12476
rect 13556 12412 13557 12476
rect 13491 12411 13557 12412
rect 11777 11936 11785 12000
rect 11849 11936 11865 12000
rect 11929 11936 11945 12000
rect 12009 11936 12025 12000
rect 12089 11936 12097 12000
rect 10731 11796 10797 11797
rect 10731 11732 10732 11796
rect 10796 11732 10797 11796
rect 10731 11731 10797 11732
rect 11651 11796 11717 11797
rect 11651 11732 11652 11796
rect 11716 11732 11717 11796
rect 11651 11731 11717 11732
rect 11777 10912 12097 11936
rect 15572 11456 15892 12480
rect 15572 11392 15580 11456
rect 15644 11392 15660 11456
rect 15724 11392 15740 11456
rect 15804 11392 15820 11456
rect 15884 11392 15892 11456
rect 15147 11116 15213 11117
rect 15147 11052 15148 11116
rect 15212 11052 15213 11116
rect 15147 11051 15213 11052
rect 11777 10848 11785 10912
rect 11849 10848 11865 10912
rect 11929 10848 11945 10912
rect 12009 10848 12025 10912
rect 12089 10848 12097 10912
rect 9627 10708 9693 10709
rect 9627 10644 9628 10708
rect 9692 10644 9693 10708
rect 9627 10643 9693 10644
rect 7982 10304 7990 10368
rect 8054 10304 8070 10368
rect 8134 10304 8150 10368
rect 8214 10304 8230 10368
rect 8294 10304 8302 10368
rect 7982 9280 8302 10304
rect 7982 9216 7990 9280
rect 8054 9216 8070 9280
rect 8134 9216 8150 9280
rect 8214 9216 8230 9280
rect 8294 9216 8302 9280
rect 7982 8192 8302 9216
rect 7982 8128 7990 8192
rect 8054 8128 8070 8192
rect 8134 8128 8150 8192
rect 8214 8128 8230 8192
rect 8294 8128 8302 8192
rect 7982 7104 8302 8128
rect 7982 7040 7990 7104
rect 8054 7040 8070 7104
rect 8134 7040 8150 7104
rect 8214 7040 8230 7104
rect 8294 7040 8302 7104
rect 7982 6016 8302 7040
rect 7982 5952 7990 6016
rect 8054 5952 8070 6016
rect 8134 5952 8150 6016
rect 8214 5952 8230 6016
rect 8294 5952 8302 6016
rect 6683 5540 6749 5541
rect 6683 5476 6684 5540
rect 6748 5476 6749 5540
rect 6683 5475 6749 5476
rect 5579 2004 5645 2005
rect 5579 1940 5580 2004
rect 5644 1940 5645 2004
rect 5579 1939 5645 1940
rect 6686 1325 6746 5475
rect 7982 4928 8302 5952
rect 7982 4864 7990 4928
rect 8054 4864 8070 4928
rect 8134 4864 8150 4928
rect 8214 4864 8230 4928
rect 8294 4864 8302 4928
rect 7982 3840 8302 4864
rect 7982 3776 7990 3840
rect 8054 3776 8070 3840
rect 8134 3776 8150 3840
rect 8214 3776 8230 3840
rect 8294 3776 8302 3840
rect 7982 2752 8302 3776
rect 7982 2688 7990 2752
rect 8054 2688 8070 2752
rect 8134 2688 8150 2752
rect 8214 2688 8230 2752
rect 8294 2688 8302 2752
rect 7982 1664 8302 2688
rect 7982 1600 7990 1664
rect 8054 1600 8070 1664
rect 8134 1600 8150 1664
rect 8214 1600 8230 1664
rect 8294 1600 8302 1664
rect 6683 1324 6749 1325
rect 6683 1260 6684 1324
rect 6748 1260 6749 1324
rect 6683 1259 6749 1260
rect 4187 1056 4195 1120
rect 4259 1056 4275 1120
rect 4339 1056 4355 1120
rect 4419 1056 4435 1120
rect 4499 1056 4507 1120
rect 4187 496 4507 1056
rect 7982 576 8302 1600
rect 7982 512 7990 576
rect 8054 512 8070 576
rect 8134 512 8150 576
rect 8214 512 8230 576
rect 8294 512 8302 576
rect 7982 496 8302 512
rect 11777 9824 12097 10848
rect 11777 9760 11785 9824
rect 11849 9760 11865 9824
rect 11929 9760 11945 9824
rect 12009 9760 12025 9824
rect 12089 9760 12097 9824
rect 11777 8736 12097 9760
rect 11777 8672 11785 8736
rect 11849 8672 11865 8736
rect 11929 8672 11945 8736
rect 12009 8672 12025 8736
rect 12089 8672 12097 8736
rect 11777 7648 12097 8672
rect 11777 7584 11785 7648
rect 11849 7584 11865 7648
rect 11929 7584 11945 7648
rect 12009 7584 12025 7648
rect 12089 7584 12097 7648
rect 11777 6560 12097 7584
rect 11777 6496 11785 6560
rect 11849 6496 11865 6560
rect 11929 6496 11945 6560
rect 12009 6496 12025 6560
rect 12089 6496 12097 6560
rect 11777 5472 12097 6496
rect 11777 5408 11785 5472
rect 11849 5408 11865 5472
rect 11929 5408 11945 5472
rect 12009 5408 12025 5472
rect 12089 5408 12097 5472
rect 11777 4384 12097 5408
rect 11777 4320 11785 4384
rect 11849 4320 11865 4384
rect 11929 4320 11945 4384
rect 12009 4320 12025 4384
rect 12089 4320 12097 4384
rect 11777 3296 12097 4320
rect 11777 3232 11785 3296
rect 11849 3232 11865 3296
rect 11929 3232 11945 3296
rect 12009 3232 12025 3296
rect 12089 3232 12097 3296
rect 11777 2208 12097 3232
rect 15150 3093 15210 11051
rect 15572 10368 15892 11392
rect 15572 10304 15580 10368
rect 15644 10304 15660 10368
rect 15724 10304 15740 10368
rect 15804 10304 15820 10368
rect 15884 10304 15892 10368
rect 15572 9280 15892 10304
rect 15572 9216 15580 9280
rect 15644 9216 15660 9280
rect 15724 9216 15740 9280
rect 15804 9216 15820 9280
rect 15884 9216 15892 9280
rect 15572 8192 15892 9216
rect 15572 8128 15580 8192
rect 15644 8128 15660 8192
rect 15724 8128 15740 8192
rect 15804 8128 15820 8192
rect 15884 8128 15892 8192
rect 15572 7104 15892 8128
rect 19367 18528 19687 19552
rect 19367 18464 19375 18528
rect 19439 18464 19455 18528
rect 19519 18464 19535 18528
rect 19599 18464 19615 18528
rect 19679 18464 19687 18528
rect 19367 17440 19687 18464
rect 19367 17376 19375 17440
rect 19439 17376 19455 17440
rect 19519 17376 19535 17440
rect 19599 17376 19615 17440
rect 19679 17376 19687 17440
rect 19367 16352 19687 17376
rect 19367 16288 19375 16352
rect 19439 16288 19455 16352
rect 19519 16288 19535 16352
rect 19599 16288 19615 16352
rect 19679 16288 19687 16352
rect 19367 15264 19687 16288
rect 19367 15200 19375 15264
rect 19439 15200 19455 15264
rect 19519 15200 19535 15264
rect 19599 15200 19615 15264
rect 19679 15200 19687 15264
rect 19367 14176 19687 15200
rect 19367 14112 19375 14176
rect 19439 14112 19455 14176
rect 19519 14112 19535 14176
rect 19599 14112 19615 14176
rect 19679 14112 19687 14176
rect 19367 13088 19687 14112
rect 19367 13024 19375 13088
rect 19439 13024 19455 13088
rect 19519 13024 19535 13088
rect 19599 13024 19615 13088
rect 19679 13024 19687 13088
rect 19367 12000 19687 13024
rect 21958 12885 22018 22304
rect 22510 13293 22570 22304
rect 23062 22130 23122 22304
rect 22878 22070 23122 22130
rect 22507 13292 22573 13293
rect 22507 13228 22508 13292
rect 22572 13228 22573 13292
rect 22507 13227 22573 13228
rect 21955 12884 22021 12885
rect 21955 12820 21956 12884
rect 22020 12820 22021 12884
rect 21955 12819 22021 12820
rect 22878 12341 22938 22070
rect 23614 21861 23674 22304
rect 23611 21860 23677 21861
rect 23162 21248 23482 21808
rect 23611 21796 23612 21860
rect 23676 21796 23677 21860
rect 23611 21795 23677 21796
rect 23162 21184 23170 21248
rect 23234 21184 23250 21248
rect 23314 21184 23330 21248
rect 23394 21184 23410 21248
rect 23474 21184 23482 21248
rect 23162 20160 23482 21184
rect 23611 20908 23677 20909
rect 23611 20844 23612 20908
rect 23676 20844 23677 20908
rect 23611 20843 23677 20844
rect 23162 20096 23170 20160
rect 23234 20096 23250 20160
rect 23314 20096 23330 20160
rect 23394 20096 23410 20160
rect 23474 20096 23482 20160
rect 23162 19072 23482 20096
rect 23162 19008 23170 19072
rect 23234 19008 23250 19072
rect 23314 19008 23330 19072
rect 23394 19008 23410 19072
rect 23474 19008 23482 19072
rect 23162 17984 23482 19008
rect 23162 17920 23170 17984
rect 23234 17920 23250 17984
rect 23314 17920 23330 17984
rect 23394 17920 23410 17984
rect 23474 17920 23482 17984
rect 23162 16896 23482 17920
rect 23614 17781 23674 20843
rect 23611 17780 23677 17781
rect 23611 17716 23612 17780
rect 23676 17716 23677 17780
rect 23611 17715 23677 17716
rect 23162 16832 23170 16896
rect 23234 16832 23250 16896
rect 23314 16832 23330 16896
rect 23394 16832 23410 16896
rect 23474 16832 23482 16896
rect 23162 15808 23482 16832
rect 23162 15744 23170 15808
rect 23234 15744 23250 15808
rect 23314 15744 23330 15808
rect 23394 15744 23410 15808
rect 23474 15744 23482 15808
rect 23162 14720 23482 15744
rect 24166 15469 24226 22304
rect 24718 18869 24778 22304
rect 24715 18868 24781 18869
rect 24715 18804 24716 18868
rect 24780 18804 24781 18868
rect 24715 18803 24781 18804
rect 25270 18733 25330 22304
rect 25267 18732 25333 18733
rect 25267 18668 25268 18732
rect 25332 18668 25333 18732
rect 25267 18667 25333 18668
rect 25822 18461 25882 22304
rect 26374 21181 26434 22304
rect 26926 22104 26986 22304
rect 27478 22104 27538 22304
rect 26957 21792 27277 21808
rect 26957 21728 26965 21792
rect 27029 21728 27045 21792
rect 27109 21728 27125 21792
rect 27189 21728 27205 21792
rect 27269 21728 27277 21792
rect 26371 21180 26437 21181
rect 26371 21116 26372 21180
rect 26436 21116 26437 21180
rect 26371 21115 26437 21116
rect 26957 20704 27277 21728
rect 26957 20640 26965 20704
rect 27029 20640 27045 20704
rect 27109 20640 27125 20704
rect 27189 20640 27205 20704
rect 27269 20640 27277 20704
rect 26957 19616 27277 20640
rect 26957 19552 26965 19616
rect 27029 19552 27045 19616
rect 27109 19552 27125 19616
rect 27189 19552 27205 19616
rect 27269 19552 27277 19616
rect 26187 18596 26253 18597
rect 26187 18532 26188 18596
rect 26252 18532 26253 18596
rect 26187 18531 26253 18532
rect 25819 18460 25885 18461
rect 25819 18396 25820 18460
rect 25884 18396 25885 18460
rect 25819 18395 25885 18396
rect 24163 15468 24229 15469
rect 24163 15404 24164 15468
rect 24228 15404 24229 15468
rect 24163 15403 24229 15404
rect 23162 14656 23170 14720
rect 23234 14656 23250 14720
rect 23314 14656 23330 14720
rect 23394 14656 23410 14720
rect 23474 14656 23482 14720
rect 23162 13632 23482 14656
rect 23162 13568 23170 13632
rect 23234 13568 23250 13632
rect 23314 13568 23330 13632
rect 23394 13568 23410 13632
rect 23474 13568 23482 13632
rect 23162 12544 23482 13568
rect 26190 12749 26250 18531
rect 26957 18528 27277 19552
rect 26957 18464 26965 18528
rect 27029 18464 27045 18528
rect 27109 18464 27125 18528
rect 27189 18464 27205 18528
rect 27269 18464 27277 18528
rect 26957 17440 27277 18464
rect 30752 21248 31072 21808
rect 30752 21184 30760 21248
rect 30824 21184 30840 21248
rect 30904 21184 30920 21248
rect 30984 21184 31000 21248
rect 31064 21184 31072 21248
rect 30752 20160 31072 21184
rect 30752 20096 30760 20160
rect 30824 20096 30840 20160
rect 30904 20096 30920 20160
rect 30984 20096 31000 20160
rect 31064 20096 31072 20160
rect 30752 19072 31072 20096
rect 30752 19008 30760 19072
rect 30824 19008 30840 19072
rect 30904 19008 30920 19072
rect 30984 19008 31000 19072
rect 31064 19008 31072 19072
rect 30051 18324 30117 18325
rect 30051 18260 30052 18324
rect 30116 18260 30117 18324
rect 30051 18259 30117 18260
rect 26957 17376 26965 17440
rect 27029 17376 27045 17440
rect 27109 17376 27125 17440
rect 27189 17376 27205 17440
rect 27269 17376 27277 17440
rect 26957 16352 27277 17376
rect 26957 16288 26965 16352
rect 27029 16288 27045 16352
rect 27109 16288 27125 16352
rect 27189 16288 27205 16352
rect 27269 16288 27277 16352
rect 26371 15332 26437 15333
rect 26371 15268 26372 15332
rect 26436 15268 26437 15332
rect 26371 15267 26437 15268
rect 26374 13157 26434 15267
rect 26957 15264 27277 16288
rect 26957 15200 26965 15264
rect 27029 15200 27045 15264
rect 27109 15200 27125 15264
rect 27189 15200 27205 15264
rect 27269 15200 27277 15264
rect 26957 14176 27277 15200
rect 29499 14924 29565 14925
rect 29499 14860 29500 14924
rect 29564 14860 29565 14924
rect 29499 14859 29565 14860
rect 26957 14112 26965 14176
rect 27029 14112 27045 14176
rect 27109 14112 27125 14176
rect 27189 14112 27205 14176
rect 27269 14112 27277 14176
rect 26371 13156 26437 13157
rect 26371 13092 26372 13156
rect 26436 13092 26437 13156
rect 26371 13091 26437 13092
rect 26957 13088 27277 14112
rect 26957 13024 26965 13088
rect 27029 13024 27045 13088
rect 27109 13024 27125 13088
rect 27189 13024 27205 13088
rect 27269 13024 27277 13088
rect 26187 12748 26253 12749
rect 26187 12684 26188 12748
rect 26252 12684 26253 12748
rect 26187 12683 26253 12684
rect 23162 12480 23170 12544
rect 23234 12480 23250 12544
rect 23314 12480 23330 12544
rect 23394 12480 23410 12544
rect 23474 12480 23482 12544
rect 22875 12340 22941 12341
rect 22875 12276 22876 12340
rect 22940 12276 22941 12340
rect 22875 12275 22941 12276
rect 19367 11936 19375 12000
rect 19439 11936 19455 12000
rect 19519 11936 19535 12000
rect 19599 11936 19615 12000
rect 19679 11936 19687 12000
rect 19367 10912 19687 11936
rect 19367 10848 19375 10912
rect 19439 10848 19455 10912
rect 19519 10848 19535 10912
rect 19599 10848 19615 10912
rect 19679 10848 19687 10912
rect 19367 9824 19687 10848
rect 19367 9760 19375 9824
rect 19439 9760 19455 9824
rect 19519 9760 19535 9824
rect 19599 9760 19615 9824
rect 19679 9760 19687 9824
rect 19367 8736 19687 9760
rect 19367 8672 19375 8736
rect 19439 8672 19455 8736
rect 19519 8672 19535 8736
rect 19599 8672 19615 8736
rect 19679 8672 19687 8736
rect 19367 7648 19687 8672
rect 19367 7584 19375 7648
rect 19439 7584 19455 7648
rect 19519 7584 19535 7648
rect 19599 7584 19615 7648
rect 19679 7584 19687 7648
rect 17907 7580 17973 7581
rect 17907 7516 17908 7580
rect 17972 7516 17973 7580
rect 17907 7515 17973 7516
rect 15572 7040 15580 7104
rect 15644 7040 15660 7104
rect 15724 7040 15740 7104
rect 15804 7040 15820 7104
rect 15884 7040 15892 7104
rect 15572 6016 15892 7040
rect 15572 5952 15580 6016
rect 15644 5952 15660 6016
rect 15724 5952 15740 6016
rect 15804 5952 15820 6016
rect 15884 5952 15892 6016
rect 15572 4928 15892 5952
rect 15572 4864 15580 4928
rect 15644 4864 15660 4928
rect 15724 4864 15740 4928
rect 15804 4864 15820 4928
rect 15884 4864 15892 4928
rect 15572 3840 15892 4864
rect 17910 4317 17970 7515
rect 19367 6560 19687 7584
rect 19367 6496 19375 6560
rect 19439 6496 19455 6560
rect 19519 6496 19535 6560
rect 19599 6496 19615 6560
rect 19679 6496 19687 6560
rect 19367 5472 19687 6496
rect 19367 5408 19375 5472
rect 19439 5408 19455 5472
rect 19519 5408 19535 5472
rect 19599 5408 19615 5472
rect 19679 5408 19687 5472
rect 19367 4384 19687 5408
rect 19367 4320 19375 4384
rect 19439 4320 19455 4384
rect 19519 4320 19535 4384
rect 19599 4320 19615 4384
rect 19679 4320 19687 4384
rect 17907 4316 17973 4317
rect 17907 4252 17908 4316
rect 17972 4252 17973 4316
rect 17907 4251 17973 4252
rect 15572 3776 15580 3840
rect 15644 3776 15660 3840
rect 15724 3776 15740 3840
rect 15804 3776 15820 3840
rect 15884 3776 15892 3840
rect 15147 3092 15213 3093
rect 15147 3028 15148 3092
rect 15212 3028 15213 3092
rect 15147 3027 15213 3028
rect 15150 2413 15210 3027
rect 15572 2752 15892 3776
rect 15572 2688 15580 2752
rect 15644 2688 15660 2752
rect 15724 2688 15740 2752
rect 15804 2688 15820 2752
rect 15884 2688 15892 2752
rect 15147 2412 15213 2413
rect 15147 2348 15148 2412
rect 15212 2348 15213 2412
rect 15147 2347 15213 2348
rect 11777 2144 11785 2208
rect 11849 2144 11865 2208
rect 11929 2144 11945 2208
rect 12009 2144 12025 2208
rect 12089 2144 12097 2208
rect 11777 1120 12097 2144
rect 11777 1056 11785 1120
rect 11849 1056 11865 1120
rect 11929 1056 11945 1120
rect 12009 1056 12025 1120
rect 12089 1056 12097 1120
rect 11777 496 12097 1056
rect 15572 1664 15892 2688
rect 15572 1600 15580 1664
rect 15644 1600 15660 1664
rect 15724 1600 15740 1664
rect 15804 1600 15820 1664
rect 15884 1600 15892 1664
rect 15572 576 15892 1600
rect 15572 512 15580 576
rect 15644 512 15660 576
rect 15724 512 15740 576
rect 15804 512 15820 576
rect 15884 512 15892 576
rect 15572 496 15892 512
rect 19367 3296 19687 4320
rect 19367 3232 19375 3296
rect 19439 3232 19455 3296
rect 19519 3232 19535 3296
rect 19599 3232 19615 3296
rect 19679 3232 19687 3296
rect 19367 2208 19687 3232
rect 19367 2144 19375 2208
rect 19439 2144 19455 2208
rect 19519 2144 19535 2208
rect 19599 2144 19615 2208
rect 19679 2144 19687 2208
rect 19367 1120 19687 2144
rect 19367 1056 19375 1120
rect 19439 1056 19455 1120
rect 19519 1056 19535 1120
rect 19599 1056 19615 1120
rect 19679 1056 19687 1120
rect 19367 496 19687 1056
rect 23162 11456 23482 12480
rect 23162 11392 23170 11456
rect 23234 11392 23250 11456
rect 23314 11392 23330 11456
rect 23394 11392 23410 11456
rect 23474 11392 23482 11456
rect 23162 10368 23482 11392
rect 23162 10304 23170 10368
rect 23234 10304 23250 10368
rect 23314 10304 23330 10368
rect 23394 10304 23410 10368
rect 23474 10304 23482 10368
rect 23162 9280 23482 10304
rect 23162 9216 23170 9280
rect 23234 9216 23250 9280
rect 23314 9216 23330 9280
rect 23394 9216 23410 9280
rect 23474 9216 23482 9280
rect 23162 8192 23482 9216
rect 23162 8128 23170 8192
rect 23234 8128 23250 8192
rect 23314 8128 23330 8192
rect 23394 8128 23410 8192
rect 23474 8128 23482 8192
rect 23162 7104 23482 8128
rect 23162 7040 23170 7104
rect 23234 7040 23250 7104
rect 23314 7040 23330 7104
rect 23394 7040 23410 7104
rect 23474 7040 23482 7104
rect 23162 6016 23482 7040
rect 23162 5952 23170 6016
rect 23234 5952 23250 6016
rect 23314 5952 23330 6016
rect 23394 5952 23410 6016
rect 23474 5952 23482 6016
rect 23162 4928 23482 5952
rect 23162 4864 23170 4928
rect 23234 4864 23250 4928
rect 23314 4864 23330 4928
rect 23394 4864 23410 4928
rect 23474 4864 23482 4928
rect 23162 3840 23482 4864
rect 26957 12000 27277 13024
rect 29502 12477 29562 14859
rect 30054 13837 30114 18259
rect 30752 17984 31072 19008
rect 30752 17920 30760 17984
rect 30824 17920 30840 17984
rect 30904 17920 30920 17984
rect 30984 17920 31000 17984
rect 31064 17920 31072 17984
rect 30752 16896 31072 17920
rect 30752 16832 30760 16896
rect 30824 16832 30840 16896
rect 30904 16832 30920 16896
rect 30984 16832 31000 16896
rect 31064 16832 31072 16896
rect 30752 15808 31072 16832
rect 30752 15744 30760 15808
rect 30824 15744 30840 15808
rect 30904 15744 30920 15808
rect 30984 15744 31000 15808
rect 31064 15744 31072 15808
rect 30752 14720 31072 15744
rect 30752 14656 30760 14720
rect 30824 14656 30840 14720
rect 30904 14656 30920 14720
rect 30984 14656 31000 14720
rect 31064 14656 31072 14720
rect 30051 13836 30117 13837
rect 30051 13772 30052 13836
rect 30116 13772 30117 13836
rect 30051 13771 30117 13772
rect 30752 13632 31072 14656
rect 30752 13568 30760 13632
rect 30824 13568 30840 13632
rect 30904 13568 30920 13632
rect 30984 13568 31000 13632
rect 31064 13568 31072 13632
rect 30752 12544 31072 13568
rect 30752 12480 30760 12544
rect 30824 12480 30840 12544
rect 30904 12480 30920 12544
rect 30984 12480 31000 12544
rect 31064 12480 31072 12544
rect 29499 12476 29565 12477
rect 29499 12412 29500 12476
rect 29564 12412 29565 12476
rect 29499 12411 29565 12412
rect 26957 11936 26965 12000
rect 27029 11936 27045 12000
rect 27109 11936 27125 12000
rect 27189 11936 27205 12000
rect 27269 11936 27277 12000
rect 26957 10912 27277 11936
rect 26957 10848 26965 10912
rect 27029 10848 27045 10912
rect 27109 10848 27125 10912
rect 27189 10848 27205 10912
rect 27269 10848 27277 10912
rect 26957 9824 27277 10848
rect 26957 9760 26965 9824
rect 27029 9760 27045 9824
rect 27109 9760 27125 9824
rect 27189 9760 27205 9824
rect 27269 9760 27277 9824
rect 26957 8736 27277 9760
rect 26957 8672 26965 8736
rect 27029 8672 27045 8736
rect 27109 8672 27125 8736
rect 27189 8672 27205 8736
rect 27269 8672 27277 8736
rect 26957 7648 27277 8672
rect 26957 7584 26965 7648
rect 27029 7584 27045 7648
rect 27109 7584 27125 7648
rect 27189 7584 27205 7648
rect 27269 7584 27277 7648
rect 26957 6560 27277 7584
rect 26957 6496 26965 6560
rect 27029 6496 27045 6560
rect 27109 6496 27125 6560
rect 27189 6496 27205 6560
rect 27269 6496 27277 6560
rect 26957 5472 27277 6496
rect 26957 5408 26965 5472
rect 27029 5408 27045 5472
rect 27109 5408 27125 5472
rect 27189 5408 27205 5472
rect 27269 5408 27277 5472
rect 23795 4724 23861 4725
rect 23795 4660 23796 4724
rect 23860 4660 23861 4724
rect 23795 4659 23861 4660
rect 23162 3776 23170 3840
rect 23234 3776 23250 3840
rect 23314 3776 23330 3840
rect 23394 3776 23410 3840
rect 23474 3776 23482 3840
rect 23162 2752 23482 3776
rect 23162 2688 23170 2752
rect 23234 2688 23250 2752
rect 23314 2688 23330 2752
rect 23394 2688 23410 2752
rect 23474 2688 23482 2752
rect 23162 1664 23482 2688
rect 23162 1600 23170 1664
rect 23234 1600 23250 1664
rect 23314 1600 23330 1664
rect 23394 1600 23410 1664
rect 23474 1600 23482 1664
rect 23162 576 23482 1600
rect 23798 1189 23858 4659
rect 26957 4384 27277 5408
rect 26957 4320 26965 4384
rect 27029 4320 27045 4384
rect 27109 4320 27125 4384
rect 27189 4320 27205 4384
rect 27269 4320 27277 4384
rect 26957 3296 27277 4320
rect 26957 3232 26965 3296
rect 27029 3232 27045 3296
rect 27109 3232 27125 3296
rect 27189 3232 27205 3296
rect 27269 3232 27277 3296
rect 24715 2548 24781 2549
rect 24715 2484 24716 2548
rect 24780 2484 24781 2548
rect 24715 2483 24781 2484
rect 23795 1188 23861 1189
rect 23795 1124 23796 1188
rect 23860 1124 23861 1188
rect 23795 1123 23861 1124
rect 24718 917 24778 2483
rect 26957 2208 27277 3232
rect 26957 2144 26965 2208
rect 27029 2144 27045 2208
rect 27109 2144 27125 2208
rect 27189 2144 27205 2208
rect 27269 2144 27277 2208
rect 26957 1120 27277 2144
rect 26957 1056 26965 1120
rect 27029 1056 27045 1120
rect 27109 1056 27125 1120
rect 27189 1056 27205 1120
rect 27269 1056 27277 1120
rect 24715 916 24781 917
rect 24715 852 24716 916
rect 24780 852 24781 916
rect 24715 851 24781 852
rect 23162 512 23170 576
rect 23234 512 23250 576
rect 23314 512 23330 576
rect 23394 512 23410 576
rect 23474 512 23482 576
rect 23162 496 23482 512
rect 26957 496 27277 1056
rect 30752 11456 31072 12480
rect 30752 11392 30760 11456
rect 30824 11392 30840 11456
rect 30904 11392 30920 11456
rect 30984 11392 31000 11456
rect 31064 11392 31072 11456
rect 30752 10368 31072 11392
rect 30752 10304 30760 10368
rect 30824 10304 30840 10368
rect 30904 10304 30920 10368
rect 30984 10304 31000 10368
rect 31064 10304 31072 10368
rect 30752 9280 31072 10304
rect 30752 9216 30760 9280
rect 30824 9216 30840 9280
rect 30904 9216 30920 9280
rect 30984 9216 31000 9280
rect 31064 9216 31072 9280
rect 30752 8192 31072 9216
rect 30752 8128 30760 8192
rect 30824 8128 30840 8192
rect 30904 8128 30920 8192
rect 30984 8128 31000 8192
rect 31064 8128 31072 8192
rect 30752 7104 31072 8128
rect 30752 7040 30760 7104
rect 30824 7040 30840 7104
rect 30904 7040 30920 7104
rect 30984 7040 31000 7104
rect 31064 7040 31072 7104
rect 30752 6016 31072 7040
rect 30752 5952 30760 6016
rect 30824 5952 30840 6016
rect 30904 5952 30920 6016
rect 30984 5952 31000 6016
rect 31064 5952 31072 6016
rect 30752 4928 31072 5952
rect 30752 4864 30760 4928
rect 30824 4864 30840 4928
rect 30904 4864 30920 4928
rect 30984 4864 31000 4928
rect 31064 4864 31072 4928
rect 30752 3840 31072 4864
rect 30752 3776 30760 3840
rect 30824 3776 30840 3840
rect 30904 3776 30920 3840
rect 30984 3776 31000 3840
rect 31064 3776 31072 3840
rect 30752 2752 31072 3776
rect 30752 2688 30760 2752
rect 30824 2688 30840 2752
rect 30904 2688 30920 2752
rect 30984 2688 31000 2752
rect 31064 2688 31072 2752
rect 30752 1664 31072 2688
rect 30752 1600 30760 1664
rect 30824 1600 30840 1664
rect 30904 1600 30920 1664
rect 30984 1600 31000 1664
rect 31064 1600 31072 1664
rect 30752 576 31072 1600
rect 30752 512 30760 576
rect 30824 512 30840 576
rect 30904 512 30920 576
rect 30984 512 31000 576
rect 31064 512 31072 576
rect 30752 496 31072 512
use sky130_fd_sc_hd__inv_2  _05_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 30360 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _06_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 21252 0 1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  _07_
timestamp 1693170804
transform 1 0 23828 0 1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _08_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 23000 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _09_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 23184 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _10_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 18676 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _11_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 19136 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 6532 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _21_
timestamp 1693170804
transform 1 0 13340 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _22_
timestamp 1693170804
transform 1 0 10304 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _23_
timestamp 1693170804
transform 1 0 12788 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _24_
timestamp 1693170804
transform 1 0 5980 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _25_
timestamp 1693170804
transform 1 0 3312 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _26_
timestamp 1693170804
transform 1 0 2576 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _27_
timestamp 1693170804
transform 1 0 2024 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1693170804
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1693170804
transform 1 0 29440 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1693170804
transform 1 0 20332 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1693170804
transform 1 0 17204 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1693170804
transform 1 0 15548 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1693170804
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1693170804
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1693170804
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1693170804
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1693170804
transform 1 0 19136 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1693170804
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1693170804
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1693170804
transform 1 0 19136 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1693170804
transform 1 0 19872 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1693170804
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1693170804
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1693170804
transform 1 0 3772 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1693170804
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1693170804
transform 1 0 13892 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1693170804
transform 1 0 4140 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1693170804
transform 1 0 3404 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1693170804
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1693170804
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1693170804
transform 1 0 3680 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2i_2  ct.cw.cc_test_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28980 0 1 19040
box -38 -48 1050 592
use sky130_ht_sc_tt05__mux2i_2  ct.cw.cc_test_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698890999
transform 1 0 28980 0 1 16864
box -38 -48 1050 592
use sky130_fd_sc_hd__maj3_2  ct.cw.cc_test_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 29808 0 1 20128
box -38 -48 866 592
use sky130_ht_sc_tt05__maj3_2  ct.cw.cc_test_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698890999
transform 1 0 28980 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dlrtp_1  ct.cw.cc_test_4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28980 0 1 17952
box -38 -48 1234 592
use sky130_ht_sc_tt05__dlrtp_1  ct.cw.cc_test_5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698890999
transform 1 0 28980 0 -1 19040
box -38 -48 1418 592
use sky130_fd_sc_hd__dfrtp_1  ct.cw.cc_test_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 27048 0 1 17952
box -38 -48 1878 592
use sky130_ht_sc_tt05__dfrtp_1  ct.cw.cc_test_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1698890999
transform 1 0 28612 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[0\].bits\[0\].cc_flop $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28612 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[0\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 16836 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[0\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 14260 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[0\].cc_clkbuf
timestamp 1693170804
transform 1 0 28152 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[1\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[1\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[1\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 21988 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[1\].cc_clkbuf
timestamp 1693170804
transform 1 0 28980 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[2\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[2\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 14260 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[2\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[2\].cc_clkbuf
timestamp 1693170804
transform 1 0 25760 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[3\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 26404 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[3\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 28612 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[3\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 16836 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[3\].cc_clkbuf
timestamp 1693170804
transform 1 0 26036 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[4\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 26404 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[4\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[4\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 21988 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[4\].cc_clkbuf
timestamp 1693170804
transform 1 0 23920 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[5\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 26404 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[5\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 26404 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[5\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 26956 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[5\].cc_clkbuf
timestamp 1693170804
transform 1 0 23828 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[6\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 24380 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[6\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 18768 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[6\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[6\].cc_clkbuf
timestamp 1693170804
transform 1 0 22724 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[7\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 20424 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[7\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 21252 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[7\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 19412 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[7\].cc_clkbuf
timestamp 1693170804
transform 1 0 20424 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[8\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 18676 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[8\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 18676 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[8\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 18676 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[8\].cc_clkbuf
timestamp 1693170804
transform 1 0 20424 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[9\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 16928 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[9\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 16928 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[9\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 18676 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[9\].cc_clkbuf
timestamp 1693170804
transform 1 0 18676 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[10\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 16560 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[10\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 16100 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[10\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 15916 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[10\].cc_clkbuf
timestamp 1693170804
transform 1 0 17848 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[11\].bits\[0\].cc_flop
timestamp 1693170804
transform 1 0 16100 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[11\].bits\[1\].cc_flop
timestamp 1693170804
transform 1 0 14260 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  ct.ic.frame\[11\].bits\[2\].cc_flop
timestamp 1693170804
transform 1 0 14260 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_4  ct.ic.frame\[11\].cc_clkbuf
timestamp 1693170804
transform 1 0 13708 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[0\].cc_scanflop $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 11224 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 12052 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 11132 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 8464 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 4416 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8004 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 12052 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[0\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 10948 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[0\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 12144 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[0\].cc_clkbuf
timestamp 1693170804
transform 1 0 13524 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[0\].rs_mbuf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 10672 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 10672 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 4968 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 4140 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 10580 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 5244 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[1\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 8924 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[1\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[1\].bits\[7\].rs_cbuf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 9200 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[1\].cc_clkbuf
timestamp 1693170804
transform 1 0 4692 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[1\].rs_mbuf
timestamp 1693170804
transform 1 0 10948 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 9292 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 8464 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 9936 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 8372 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 5520 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[2\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[2\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 6256 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 1104 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[2\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[2\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[2\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[2\].cc_clkbuf
timestamp 1693170804
transform 1 0 1472 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[2\].rs_mbuf
timestamp 1693170804
transform 1 0 3588 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 4692 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 3864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 5888 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[3\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 3312 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 1104 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 9200 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 9752 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 9476 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[3\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[3\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[3\].cc_clkbuf
timestamp 1693170804
transform 1 0 4140 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[3\].rs_mbuf
timestamp 1693170804
transform 1 0 920 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 5796 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 11500 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[4\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 5336 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[4\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[4\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 9016 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[4\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[4\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[4\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 8648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[4\].cc_clkbuf
timestamp 1693170804
transform 1 0 5796 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[4\].rs_mbuf
timestamp 1693170804
transform 1 0 3220 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 8648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3772 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 5060 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 10212 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3772 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 11868 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 1196 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11500 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[5\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[5\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[5\].cc_clkbuf
timestamp 1693170804
transform 1 0 3220 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[5\].rs_mbuf
timestamp 1693170804
transform 1 0 3220 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6348 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 6072 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 6348 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 9384 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 9016 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[6\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8556 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[6\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 8280 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[6\].cc_clkbuf
timestamp 1693170804
transform 1 0 5796 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[6\].rs_mbuf
timestamp 1693170804
transform 1 0 8832 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 12604 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 11040 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 11316 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 12328 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 11776 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11500 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 7452 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[7\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[7\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[7\].cc_clkbuf
timestamp 1693170804
transform 1 0 10948 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[7\].rs_mbuf
timestamp 1693170804
transform 1 0 11776 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 14168 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 15456 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 14628 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 15732 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 14168 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 16744 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 11500 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 14168 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10304 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 14352 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[8\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[8\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[8\].cc_clkbuf
timestamp 1693170804
transform 1 0 13524 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[8\].rs_mbuf
timestamp 1693170804
transform 1 0 14904 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 17848 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 18676 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 17112 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 17572 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 17020 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 19228 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 14352 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 16192 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 17112 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[9\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 17020 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[9\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 13984 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[9\].cc_clkbuf
timestamp 1693170804
transform 1 0 16100 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[9\].rs_mbuf
timestamp 1693170804
transform 1 0 18676 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 19780 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 20792 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 19964 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 19780 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 20240 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 20516 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 19688 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[10\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 20516 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[10\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 23276 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[10\].cc_clkbuf
timestamp 1693170804
transform 1 0 19228 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[10\].rs_mbuf
timestamp 1693170804
transform 1 0 20884 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 20608 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 19504 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 21344 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 24748 0 1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[11\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24748 0 1 17952
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[11\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[11\].cc_clkbuf
timestamp 1693170804
transform 1 0 22724 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[11\].rs_mbuf
timestamp 1693170804
transform 1 0 24196 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 30084 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 26036 0 1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 26036 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26772 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 29992 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 28244 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 24472 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 30360 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[12\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[12\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 29716 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[12\].cc_clkbuf
timestamp 1693170804
transform 1 0 25668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[12\].rs_mbuf
timestamp 1693170804
transform 1 0 28244 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 24012 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 23552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 26220 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 28336 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 29532 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 27784 0 -1 16864
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 30084 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[13\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 15776
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[13\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 29808 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[13\].cc_clkbuf
timestamp 1693170804
transform 1 0 28244 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[13\].rs_mbuf
timestamp 1693170804
transform 1 0 26036 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 21896 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 23368 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 23092 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 23920 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 28060 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 28612 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26588 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 29532 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 28152 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 29532 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[14\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[14\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 28336 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[14\].cc_clkbuf
timestamp 1693170804
transform 1 0 28980 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[14\].rs_mbuf
timestamp 1693170804
transform 1 0 25668 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 20332 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 20608 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 22356 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 22724 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 27600 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26128 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 23184 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 27600 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 29808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[15\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[15\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 29532 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[15\].cc_clkbuf
timestamp 1693170804
transform 1 0 26404 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[15\].rs_mbuf
timestamp 1693170804
transform 1 0 25760 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 18216 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 19688 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 19964 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26128 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 23552 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 23460 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[16\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[16\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[16\].cc_clkbuf
timestamp 1693170804
transform 1 0 25116 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[16\].rs_mbuf
timestamp 1693170804
transform 1 0 19136 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16744 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 16376 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16928 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 16928 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 16652 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 19964 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 20332 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26588 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 25944 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 22264 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 26036 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[17\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24380 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[17\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 25668 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[17\].cc_clkbuf
timestamp 1693170804
transform 1 0 19136 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[17\].rs_mbuf
timestamp 1693170804
transform 1 0 16192 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 17388 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 19136 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 18676 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 19872 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 19596 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 24104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[18\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[18\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 23276 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[18\].cc_clkbuf
timestamp 1693170804
transform 1 0 20608 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[18\].rs_mbuf
timestamp 1693170804
transform 1 0 16836 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 20792 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 18584 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[19\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 21436 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[19\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 21528 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[19\].cc_clkbuf
timestamp 1693170804
transform 1 0 19596 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[19\].rs_mbuf
timestamp 1693170804
transform 1 0 17572 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 27876 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 29808 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 27784 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 27508 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 27324 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26036 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 27048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21896 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 29532 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[20\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[20\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[20\].cc_clkbuf
timestamp 1693170804
transform 1 0 22632 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[20\].rs_mbuf
timestamp 1693170804
transform 1 0 25668 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 28612 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 14168 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 28428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[21\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 27508 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[21\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 27232 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26680 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[21\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 29164 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[21\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[21\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 29256 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[21\].cc_clkbuf
timestamp 1693170804
transform 1 0 27048 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[21\].rs_mbuf
timestamp 1693170804
transform 1 0 28980 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 28980 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18952 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 26404 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 26956 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 26220 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 26220 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[22\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 26680 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 29716 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[22\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[22\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 27048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[22\].cc_clkbuf
timestamp 1693170804
transform 1 0 27140 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[22\].rs_mbuf
timestamp 1693170804
transform 1 0 26588 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[23\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16376 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[23\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 26956 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 25024 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 24012 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 24748 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 24104 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 24196 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 24012 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 24472 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[23\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 27232 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[23\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 24288 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[23\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 25300 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[23\].cc_clkbuf
timestamp 1693170804
transform 1 0 25668 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[23\].rs_mbuf
timestamp 1693170804
transform 1 0 25668 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 26404 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 26036 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 23460 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 22908 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 23092 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 21896 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 22356 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 21988 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 22080 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21528 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 26680 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[24\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 23828 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[24\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 23184 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[24\].cc_clkbuf
timestamp 1693170804
transform 1 0 23460 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[24\].rs_mbuf
timestamp 1693170804
transform 1 0 22356 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 23092 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 23368 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 19964 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 21528 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 19872 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 20792 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 21252 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 23828 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[25\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 20884 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[25\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 21528 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[25\].cc_clkbuf
timestamp 1693170804
transform 1 0 23092 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[25\].rs_mbuf
timestamp 1693170804
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 20516 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 20792 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 19504 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 19228 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 18308 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 21252 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[26\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 18676 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[26\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 20792 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[26\].cc_clkbuf
timestamp 1693170804
transform 1 0 20516 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[26\].rs_mbuf
timestamp 1693170804
transform 1 0 19228 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 15824 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 18308 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 18124 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 18952 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 17296 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 15916 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 18676 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 18676 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[27\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 15916 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[27\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 18032 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[27\].cc_clkbuf
timestamp 1693170804
transform 1 0 18676 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[27\].rs_mbuf
timestamp 1693170804
transform 1 0 16744 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13616 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 11316 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 12604 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13708 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 12328 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11040 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[28\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 13708 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[28\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[28\].cc_clkbuf
timestamp 1693170804
transform 1 0 12880 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[28\].rs_mbuf
timestamp 1693170804
transform 1 0 13616 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 10304 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 11316 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 11040 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 11500 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 11316 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[29\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[29\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 9568 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[29\].cc_clkbuf
timestamp 1693170804
transform 1 0 11040 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[29\].rs_mbuf
timestamp 1693170804
transform 1 0 12052 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 8648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 9016 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 8924 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 9844 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10028 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[30\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[30\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 9292 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[30\].cc_clkbuf
timestamp 1693170804
transform 1 0 10948 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[30\].rs_mbuf
timestamp 1693170804
transform 1 0 10028 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 544
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16376 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 3588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 7820 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 6992 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 8648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 7820 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 8096 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[31\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[31\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 5152 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[31\].cc_clkbuf
timestamp 1693170804
transform 1 0 8372 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[31\].rs_mbuf
timestamp 1693170804
transform 1 0 7268 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[32\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[32\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 8648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 7176 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 5888 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 6900 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 6624 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 5888 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 6348 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[32\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[32\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 5888 0 1 1632
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[32\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 3404 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[32\].cc_clkbuf
timestamp 1693170804
transform 1 0 6256 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[32\].rs_mbuf
timestamp 1693170804
transform 1 0 5796 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 19040
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 9752 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 15732 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3680 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 5520 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 2208 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[33\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 12880 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[33\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[33\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[33\].cc_clkbuf
timestamp 1693170804
transform 1 0 8372 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[33\].rs_mbuf
timestamp 1693170804
transform 1 0 5796 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 15732 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 9844 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 1104 0 -1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 3808
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 6440 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 4896
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 7452 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[34\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 11776 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[34\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 2720
box -38 -48 2246 592
use sky130_fd_sc_hd__buf_1  ct.oc.frame\[34\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 11500 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[34\].cc_clkbuf
timestamp 1693170804
transform 1 0 8372 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[34\].rs_mbuf
timestamp 1693170804
transform 1 0 5796 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 1196 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 6072 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 5152 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 1104 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 6164 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[35\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[35\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 3220 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[35\].cc_clkbuf
timestamp 1693170804
transform 1 0 3220 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[35\].rs_mbuf
timestamp 1693170804
transform 1 0 1104 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 9384 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 7728 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 8372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 6716 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 9200 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 11224 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 9016 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[36\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[36\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 9108 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[36\].cc_clkbuf
timestamp 1693170804
transform 1 0 5796 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[36\].rs_mbuf
timestamp 1693170804
transform 1 0 8372 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 18124 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 16100 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 13708 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 15916 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 14536 0 1 5984
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 13616 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13892 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 14996 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11224 0 1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 12604 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11592 0 -1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 12880 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[37\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 12052 0 -1 7072
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[37\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[37\].cc_clkbuf
timestamp 1693170804
transform 1 0 10948 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[37\].rs_mbuf
timestamp 1693170804
transform 1 0 14260 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 13524 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13708 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13708 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 13800 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 16008 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 11132 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 12604 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 11132 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 10304 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[38\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 11132 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[38\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[38\].cc_clkbuf
timestamp 1693170804
transform 1 0 12052 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[38\].rs_mbuf
timestamp 1693170804
transform 1 0 12880 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 12604 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 13156 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 12512 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 12328 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 12604 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 13524 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 12788 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 12512 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 12880 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 8924 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 10396 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 9660 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 9292 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[39\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[39\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 10120 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[39\].cc_clkbuf
timestamp 1693170804
transform 1 0 11776 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[39\].rs_mbuf
timestamp 1693170804
transform 1 0 14812 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 9568 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 10396 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 9568 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 9568 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 10948 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 9660 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 10120 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 8648 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 9292 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 7636 0 -1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 7360 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[40\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[40\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 8004 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[40\].cc_clkbuf
timestamp 1693170804
transform 1 0 9108 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[40\].rs_mbuf
timestamp 1693170804
transform 1 0 8372 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 6440 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 6164 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 6624 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 6164 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 6624 0 -1 14688
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 7728 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 6716 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 8740 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 6072 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 6440 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 5428 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[41\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 5520 0 1 8160
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[41\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[41\].cc_clkbuf
timestamp 1693170804
transform 1 0 7728 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[41\].rs_mbuf
timestamp 1693170804
transform 1 0 5888 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 3680 0 1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 5796 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 4232 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 3864 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 3588 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 3496 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 3312 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 3312 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 3220 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 4876 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[42\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 3588 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[42\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 4600 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[42\].cc_clkbuf
timestamp 1693170804
transform 1 0 4508 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[42\].rs_mbuf
timestamp 1693170804
transform 1 0 3680 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[0\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 13600
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[0\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[1\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[1\].rs_cbuf
timestamp 1693170804
transform 1 0 920 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[2\].cc_scanflop
timestamp 1693170804
transform 1 0 1472 0 -1 11424
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[2\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[3\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[3\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[4\].cc_scanflop
timestamp 1693170804
transform 1 0 1288 0 -1 12512
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[4\].rs_cbuf
timestamp 1693170804
transform 1 0 1012 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[5\].cc_scanflop
timestamp 1693170804
transform 1 0 1104 0 -1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[5\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[6\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 10336
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[6\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_4  ct.oc.frame\[43\].bits\[7\].cc_scanflop
timestamp 1693170804
transform 1 0 920 0 1 9248
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_1  ct.oc.frame\[43\].bits\[7\].rs_cbuf
timestamp 1693170804
transform 1 0 828 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  ct.oc.frame\[43\].cc_clkbuf
timestamp 1693170804
transform 1 0 920 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  ct.oc.frame\[43\].rs_mbuf
timestamp 1693170804
transform 1 0 1656 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dlclkp_4  ct.ro.cc_clock_gate $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 22172 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_4  ct.ro.cc_clock_inv $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 23276 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  ct.ro.cc_ring_osc_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 21252 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  ct.ro.cc_ring_osc_1
timestamp 1693170804
transform 1 0 16376 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  ct.ro.cc_ring_osc_2
timestamp 1693170804
transform 1 0 23460 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[1\].cc_div_flop $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 18952 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[2\].cc_div_flop
timestamp 1693170804
transform 1 0 19228 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[3\].cc_div_flop
timestamp 1693170804
transform 1 0 21252 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[4\].cc_div_flop
timestamp 1693170804
transform 1 0 23460 0 -1 21216
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[5\].cc_div_flop
timestamp 1693170804
transform 1 0 22172 0 -1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[6\].cc_div_flop
timestamp 1693170804
transform 1 0 21528 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  ct.ro.count\[7\].cc_div_flop
timestamp 1693170804
transform 1 0 23828 0 1 20128
box -38 -48 2246 592
use sky130_fd_sc_hd__mux2i_2  cw.cc_test_0
timestamp 1693170804
transform 1 0 17848 0 -1 21216
box -38 -48 1050 592
use sky130_ht_sc_tt05__mux2i_2  cw.cc_test_1
timestamp 1698890999
transform 1 0 16100 0 -1 17952
box -38 -48 1050 592
use sky130_fd_sc_hd__maj3_2  cw.cc_test_2
timestamp 1693170804
transform 1 0 16100 0 -1 20128
box -38 -48 866 592
use sky130_ht_sc_tt05__maj3_2  cw.cc_test_3
timestamp 1698890999
transform 1 0 16100 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dlrtp_1  cw.cc_test_4
timestamp 1693170804
transform 1 0 7084 0 1 21216
box -38 -48 1234 592
use sky130_ht_sc_tt05__dlrtp_1  cw.cc_test_5
timestamp 1698890999
transform 1 0 8648 0 1 21216
box -38 -48 1418 592
use sky130_fd_sc_hd__dfrtp_1  cw.cc_test_6
timestamp 1693170804
transform 1 0 14260 0 1 20128
box -38 -48 1878 592
use sky130_ht_sc_tt05__dfrtp_1  cw.cc_test_7
timestamp 1698890999
transform 1 0 14076 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  fanout5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 8372 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout7
timestamp 1693170804
transform 1 0 11040 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout8
timestamp 1693170804
transform 1 0 28980 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout9
timestamp 1693170804
transform 1 0 30084 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout10
timestamp 1693170804
transform 1 0 8832 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout11
timestamp 1693170804
transform 1 0 11776 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout12
timestamp 1693170804
transform 1 0 13524 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 1693170804
transform 1 0 28336 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1693170804
transform 1 0 29532 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout15
timestamp 1693170804
transform 1 0 8924 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 1693170804
transform 1 0 12144 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout17
timestamp 1693170804
transform 1 0 13708 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 1693170804
transform 1 0 27508 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout19
timestamp 1693170804
transform 1 0 29992 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1693170804
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout21
timestamp 1693170804
transform 1 0 13064 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 1693170804
transform 1 0 13616 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1693170804
transform 1 0 25944 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1693170804
transform 1 0 29992 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1693170804
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout26
timestamp 1693170804
transform 1 0 16100 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 1693170804
transform 1 0 17664 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1693170804
transform 1 0 24656 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout29
timestamp 1693170804
transform 1 0 28980 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout30
timestamp 1693170804
transform 1 0 30084 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 1693170804
transform 1 0 8096 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout32
timestamp 1693170804
transform 1 0 12328 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout33
timestamp 1693170804
transform 1 0 5336 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout34
timestamp 1693170804
transform 1 0 28244 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout35
timestamp 1693170804
transform 1 0 27140 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1693170804
transform 1 0 29716 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout37
timestamp 1693170804
transform 1 0 10948 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 1693170804
transform 1 0 14720 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout39 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 10948 0 -1 20128
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout40
timestamp 1693170804
transform 1 0 28980 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout41
timestamp 1693170804
transform 1 0 26588 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 1693170804
transform 1 0 29348 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp 1693170804
transform 1 0 10856 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout44
timestamp 1693170804
transform 1 0 8096 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 1693170804
transform 1 0 12880 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout46
timestamp 1693170804
transform 1 0 29532 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout47
timestamp 1693170804
transform 1 0 25760 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout48
timestamp 1693170804
transform 1 0 28980 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1693170804
transform 1 0 13984 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp 1693170804
transform 1 0 13340 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 1693170804
transform 1 0 7728 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout52
timestamp 1693170804
transform 1 0 26956 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout53
timestamp 1693170804
transform 1 0 25668 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 1693170804
transform 1 0 24380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 828 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3220 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_33
timestamp 1693170804
transform 1 0 3588 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_37
timestamp 1693170804
transform 1 0 3956 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 4324 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_49
timestamp 1693170804
transform 1 0 5060 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_312
timestamp 1693170804
transform 1 0 29256 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_316
timestamp 1693170804
transform 1 0 29624 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_324 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 30360 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 1693170804
transform 1 0 828 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_63
timestamp 1693170804
transform 1 0 6348 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 1693170804
transform 1 0 10948 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1693170804
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1693170804
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_320 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 29992 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_326
timestamp 1693170804
transform 1 0 30544 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 1693170804
transform 1 0 828 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_56
timestamp 1693170804
transform 1 0 5704 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 1693170804
transform 1 0 8096 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_91
timestamp 1693170804
transform 1 0 8924 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_141
timestamp 1693170804
transform 1 0 13524 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1693170804
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_256
timestamp 1693170804
transform 1 0 24104 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_282
timestamp 1693170804
transform 1 0 26496 0 1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_312 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 29256 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_324
timestamp 1693170804
transform 1 0 30360 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_6
timestamp 1693170804
transform 1 0 1104 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_63
timestamp 1693170804
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_113
timestamp 1693170804
transform 1 0 10948 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1693170804
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_255
timestamp 1693170804
transform 1 0 24012 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_314
timestamp 1693170804
transform 1 0 29440 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_326
timestamp 1693170804
transform 1 0 30544 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_3
timestamp 1693170804
transform 1 0 828 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_29
timestamp 1693170804
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_91
timestamp 1693170804
transform 1 0 8924 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_141
timestamp 1693170804
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1693170804
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1693170804
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_277
timestamp 1693170804
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_306
timestamp 1693170804
transform 1 0 28704 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_315
timestamp 1693170804
transform 1 0 29532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_6
timestamp 1693170804
transform 1 0 1104 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_60
timestamp 1693170804
transform 1 0 6072 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_68
timestamp 1693170804
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_119
timestamp 1693170804
transform 1 0 11500 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1693170804
transform 1 0 21068 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1693170804
transform 1 0 26220 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_281
timestamp 1693170804
transform 1 0 26404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_295
timestamp 1693170804
transform 1 0 27692 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_321
timestamp 1693170804
transform 1 0 30084 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 1693170804
transform 1 0 828 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 1693170804
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1693170804
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_91
timestamp 1693170804
transform 1 0 8924 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_141
timestamp 1693170804
transform 1 0 13524 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_209
timestamp 1693170804
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_235
timestamp 1693170804
transform 1 0 22172 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_249
timestamp 1693170804
transform 1 0 23460 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1693170804
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_303 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 28428 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1693170804
transform 1 0 28796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1693170804
transform 1 0 28980 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_321
timestamp 1693170804
transform 1 0 30084 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_30
timestamp 1693170804
transform 1 0 3312 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_57
timestamp 1693170804
transform 1 0 5796 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_116
timestamp 1693170804
transform 1 0 11224 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1693170804
transform 1 0 21068 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_231
timestamp 1693170804
transform 1 0 21804 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_272
timestamp 1693170804
transform 1 0 25576 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_284
timestamp 1693170804
transform 1 0 26680 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_291
timestamp 1693170804
transform 1 0 27324 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_295
timestamp 1693170804
transform 1 0 27692 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_320
timestamp 1693170804
transform 1 0 29992 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_326
timestamp 1693170804
transform 1 0 30544 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1693170804
transform 1 0 828 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_35
timestamp 1693170804
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_91
timestamp 1693170804
transform 1 0 8924 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_141
timestamp 1693170804
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_191
timestamp 1693170804
transform 1 0 18124 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_248
timestamp 1693170804
transform 1 0 23368 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_277
timestamp 1693170804
transform 1 0 26036 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_283
timestamp 1693170804
transform 1 0 26588 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_315
timestamp 1693170804
transform 1 0 29532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_6
timestamp 1693170804
transform 1 0 1104 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_78
timestamp 1693170804
transform 1 0 7728 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 1693170804
transform 1 0 10948 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1693170804
transform 1 0 21068 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_231
timestamp 1693170804
transform 1 0 21804 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_317
timestamp 1693170804
transform 1 0 29716 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_325
timestamp 1693170804
transform 1 0 30452 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 1693170804
transform 1 0 828 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 1693170804
transform 1 0 3220 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_118
timestamp 1693170804
transform 1 0 11408 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_141
timestamp 1693170804
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_191
timestamp 1693170804
transform 1 0 18124 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_209
timestamp 1693170804
transform 1 0 19780 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_246
timestamp 1693170804
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1693170804
transform 1 0 23552 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_253
timestamp 1693170804
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_279
timestamp 1693170804
transform 1 0 26220 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_283
timestamp 1693170804
transform 1 0 26588 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_312
timestamp 1693170804
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_324
timestamp 1693170804
transform 1 0 30360 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1693170804
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_63
timestamp 1693170804
transform 1 0 6348 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_155
timestamp 1693170804
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_164
timestamp 1693170804
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_220
timestamp 1693170804
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_231
timestamp 1693170804
transform 1 0 21804 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_284
timestamp 1693170804
transform 1 0 26680 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_318
timestamp 1693170804
transform 1 0 29808 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_326
timestamp 1693170804
transform 1 0 30544 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 1693170804
transform 1 0 828 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_59
timestamp 1693170804
transform 1 0 5980 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_91
timestamp 1693170804
transform 1 0 8924 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_141
timestamp 1693170804
transform 1 0 13524 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_221
timestamp 1693170804
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_225
timestamp 1693170804
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1693170804
transform 1 0 23644 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1693170804
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_318
timestamp 1693170804
transform 1 0 29808 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_326
timestamp 1693170804
transform 1 0 30544 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_6
timestamp 1693170804
transform 1 0 1104 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_31
timestamp 1693170804
transform 1 0 3404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_63
timestamp 1693170804
transform 1 0 6348 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_119
timestamp 1693170804
transform 1 0 11500 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1693170804
transform 1 0 21068 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1693170804
transform 1 0 26220 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_284
timestamp 1693170804
transform 1 0 26680 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_321
timestamp 1693170804
transform 1 0 30084 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_3
timestamp 1693170804
transform 1 0 828 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_53
timestamp 1693170804
transform 1 0 5428 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_91
timestamp 1693170804
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_123
timestamp 1693170804
transform 1 0 11868 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 1693170804
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1693170804
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_221
timestamp 1693170804
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_280
timestamp 1693170804
transform 1 0 26312 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_321
timestamp 1693170804
transform 1 0 30084 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_42
timestamp 1693170804
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_60
timestamp 1693170804
transform 1 0 6072 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_73
timestamp 1693170804
transform 1 0 7268 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_104
timestamp 1693170804
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1693170804
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_143
timestamp 1693170804
transform 1 0 13708 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_175
timestamp 1693170804
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_213
timestamp 1693170804
transform 1 0 20148 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1693170804
transform 1 0 20516 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1693170804
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1693170804
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_324
timestamp 1693170804
transform 1 0 30360 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 1693170804
transform 1 0 828 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_29
timestamp 1693170804
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_89
timestamp 1693170804
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1693170804
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_141
timestamp 1693170804
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_167
timestamp 1693170804
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_245
timestamp 1693170804
transform 1 0 23092 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1693170804
transform 1 0 23552 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1693170804
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_315
timestamp 1693170804
transform 1 0 29532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1693170804
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1693170804
transform 1 0 5796 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 1693170804
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_139
timestamp 1693170804
transform 1 0 13340 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_143
timestamp 1693170804
transform 1 0 13708 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_169
timestamp 1693170804
transform 1 0 16100 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_200
timestamp 1693170804
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_205
timestamp 1693170804
transform 1 0 19412 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_213
timestamp 1693170804
transform 1 0 20148 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_249
timestamp 1693170804
transform 1 0 23460 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_274
timestamp 1693170804
transform 1 0 25760 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_324
timestamp 1693170804
transform 1 0 30360 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_3
timestamp 1693170804
transform 1 0 828 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_53
timestamp 1693170804
transform 1 0 5428 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_171
timestamp 1693170804
transform 1 0 16284 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_200
timestamp 1693170804
transform 1 0 18952 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_204
timestamp 1693170804
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_208
timestamp 1693170804
transform 1 0 19688 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_235
timestamp 1693170804
transform 1 0 22172 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_239
timestamp 1693170804
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_244
timestamp 1693170804
transform 1 0 23000 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_248
timestamp 1693170804
transform 1 0 23368 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_277
timestamp 1693170804
transform 1 0 26036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_321
timestamp 1693170804
transform 1 0 30084 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_3
timestamp 1693170804
transform 1 0 828 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1693170804
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_57
timestamp 1693170804
transform 1 0 5796 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_65
timestamp 1693170804
transform 1 0 6532 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_103
timestamp 1693170804
transform 1 0 10028 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 1693170804
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_163
timestamp 1693170804
transform 1 0 15548 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1693170804
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_169
timestamp 1693170804
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_208
timestamp 1693170804
transform 1 0 19688 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_212
timestamp 1693170804
transform 1 0 20056 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_228
timestamp 1693170804
transform 1 0 21528 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_236
timestamp 1693170804
transform 1 0 22264 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_261
timestamp 1693170804
transform 1 0 24564 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_266
timestamp 1693170804
transform 1 0 25024 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_273
timestamp 1693170804
transform 1 0 25668 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_324
timestamp 1693170804
transform 1 0 30360 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_3
timestamp 1693170804
transform 1 0 828 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_29
timestamp 1693170804
transform 1 0 3220 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_91
timestamp 1693170804
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_165
timestamp 1693170804
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_169
timestamp 1693170804
transform 1 0 16100 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_245
timestamp 1693170804
transform 1 0 23092 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_253
timestamp 1693170804
transform 1 0 23828 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_318
timestamp 1693170804
transform 1 0 29808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_326
timestamp 1693170804
transform 1 0 30544 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1693170804
transform 1 0 828 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_60
timestamp 1693170804
transform 1 0 6072 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_161
timestamp 1693170804
transform 1 0 15364 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 1693170804
transform 1 0 15732 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_169
timestamp 1693170804
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_173
timestamp 1693170804
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_214
timestamp 1693170804
transform 1 0 20240 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1693170804
transform 1 0 26220 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_297
timestamp 1693170804
transform 1 0 27876 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_323
timestamp 1693170804
transform 1 0 30268 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_3
timestamp 1693170804
transform 1 0 828 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_29
timestamp 1693170804
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_189
timestamp 1693170804
transform 1 0 17940 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1693170804
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1693170804
transform 1 0 23644 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1693170804
transform 1 0 28796 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp 1693170804
transform 1 0 828 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_60
timestamp 1693170804
transform 1 0 6072 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_103
timestamp 1693170804
transform 1 0 10028 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_110
timestamp 1693170804
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_128
timestamp 1693170804
transform 1 0 12328 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_154
timestamp 1693170804
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_169
timestamp 1693170804
transform 1 0 16100 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_175
timestamp 1693170804
transform 1 0 16652 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_179
timestamp 1693170804
transform 1 0 17020 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_183
timestamp 1693170804
transform 1 0 17388 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_191
timestamp 1693170804
transform 1 0 18124 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_217
timestamp 1693170804
transform 1 0 20516 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_225
timestamp 1693170804
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_3
timestamp 1693170804
transform 1 0 828 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_29
timestamp 1693170804
transform 1 0 3220 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_33
timestamp 1693170804
transform 1 0 3588 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_58
timestamp 1693170804
transform 1 0 5888 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_91
timestamp 1693170804
transform 1 0 8924 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_147
timestamp 1693170804
transform 1 0 14076 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_200
timestamp 1693170804
transform 1 0 18952 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_204
timestamp 1693170804
transform 1 0 19320 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_253
timestamp 1693170804
transform 1 0 23828 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_282
timestamp 1693170804
transform 1 0 26496 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_3
timestamp 1693170804
transform 1 0 828 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_31
timestamp 1693170804
transform 1 0 3404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1693170804
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_113
timestamp 1693170804
transform 1 0 10948 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_178
timestamp 1693170804
transform 1 0 16928 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_206
timestamp 1693170804
transform 1 0 19504 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1693170804
transform 1 0 21068 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_249
timestamp 1693170804
transform 1 0 23460 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_3
timestamp 1693170804
transform 1 0 828 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_59
timestamp 1693170804
transform 1 0 5980 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_85
timestamp 1693170804
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_111
timestamp 1693170804
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_147
timestamp 1693170804
transform 1 0 14076 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1693170804
transform 1 0 28796 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_3
timestamp 1693170804
transform 1 0 828 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_7
timestamp 1693170804
transform 1 0 1196 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1693170804
transform 1 0 10764 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_119
timestamp 1693170804
transform 1 0 11500 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_175
timestamp 1693170804
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_204
timestamp 1693170804
transform 1 0 19320 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_273
timestamp 1693170804
transform 1 0 25668 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_3
timestamp 1693170804
transform 1 0 828 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_59
timestamp 1693170804
transform 1 0 5980 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_85
timestamp 1693170804
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_111
timestamp 1693170804
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_141
timestamp 1693170804
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_149
timestamp 1693170804
transform 1 0 14260 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_227
timestamp 1693170804
transform 1 0 21436 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1693170804
transform 1 0 28796 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_325
timestamp 1693170804
transform 1 0 30452 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_3
timestamp 1693170804
transform 1 0 828 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1693170804
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_113
timestamp 1693170804
transform 1 0 10948 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_169
timestamp 1693170804
transform 1 0 16100 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_173
timestamp 1693170804
transform 1 0 16468 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_177
timestamp 1693170804
transform 1 0 16836 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_203
timestamp 1693170804
transform 1 0 19228 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1693170804
transform 1 0 26220 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_281
timestamp 1693170804
transform 1 0 26404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_295
timestamp 1693170804
transform 1 0 27692 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_326
timestamp 1693170804
transform 1 0 30544 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_3
timestamp 1693170804
transform 1 0 828 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_35
timestamp 1693170804
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_147
timestamp 1693170804
transform 1 0 14076 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_197
timestamp 1693170804
transform 1 0 18676 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 1693170804
transform 1 0 23552 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_256
timestamp 1693170804
transform 1 0 24104 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_306
timestamp 1693170804
transform 1 0 28704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_326
timestamp 1693170804
transform 1 0 30544 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_3
timestamp 1693170804
transform 1 0 828 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_63
timestamp 1693170804
transform 1 0 6348 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_143
timestamp 1693170804
transform 1 0 13708 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_147
timestamp 1693170804
transform 1 0 14076 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_204
timestamp 1693170804
transform 1 0 19320 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_254
timestamp 1693170804
transform 1 0 23920 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_326
timestamp 1693170804
transform 1 0 30544 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_3
timestamp 1693170804
transform 1 0 828 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_53
timestamp 1693170804
transform 1 0 5428 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_85
timestamp 1693170804
transform 1 0 8372 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_141
timestamp 1693170804
transform 1 0 13524 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_148
timestamp 1693170804
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_216
timestamp 1693170804
transform 1 0 20424 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_287
timestamp 1693170804
transform 1 0 26956 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_322
timestamp 1693170804
transform 1 0 30176 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_3
timestamp 1693170804
transform 1 0 828 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_32
timestamp 1693170804
transform 1 0 3496 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_51
timestamp 1693170804
transform 1 0 5244 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_57
timestamp 1693170804
transform 1 0 5796 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1693170804
transform 1 0 20976 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_284
timestamp 1693170804
transform 1 0 26680 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_3
timestamp 1693170804
transform 1 0 828 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_29
timestamp 1693170804
transform 1 0 3220 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_109
timestamp 1693170804
transform 1 0 10580 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_165
timestamp 1693170804
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_253
timestamp 1693170804
transform 1 0 23828 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_320
timestamp 1693170804
transform 1 0 29992 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_30
timestamp 1693170804
transform 1 0 3312 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_81
timestamp 1693170804
transform 1 0 8004 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_110
timestamp 1693170804
transform 1 0 10672 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_123
timestamp 1693170804
transform 1 0 11868 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_222
timestamp 1693170804
transform 1 0 20976 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_234
timestamp 1693170804
transform 1 0 22080 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_278
timestamp 1693170804
transform 1 0 26128 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_300
timestamp 1693170804
transform 1 0 28152 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_326
timestamp 1693170804
transform 1 0 30544 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_3
timestamp 1693170804
transform 1 0 828 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_29
timestamp 1693170804
transform 1 0 3220 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1693170804
transform 1 0 13340 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_141
timestamp 1693170804
transform 1 0 13524 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_194
timestamp 1693170804
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_227
timestamp 1693170804
transform 1 0 21436 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_283
timestamp 1693170804
transform 1 0 26588 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 1693170804
transform 1 0 5520 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_105
timestamp 1693170804
transform 1 0 10212 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_113
timestamp 1693170804
transform 1 0 10948 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_145
timestamp 1693170804
transform 1 0 13892 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_199
timestamp 1693170804
transform 1 0 18860 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1693170804
transform 1 0 26220 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_300
timestamp 1693170804
transform 1 0 28152 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_325
timestamp 1693170804
transform 1 0 30452 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_3
timestamp 1693170804
transform 1 0 828 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_57
timestamp 1693170804
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_103
timestamp 1693170804
transform 1 0 10028 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_147
timestamp 1693170804
transform 1 0 14076 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 1693170804
transform 1 0 28704 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_315
timestamp 1693170804
transform 1 0 29532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_323
timestamp 1693170804
transform 1 0 30268 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1693170804
transform 1 0 16836 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1693170804
transform 1 0 30360 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1693170804
transform 1 0 30084 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1693170804
transform 1 0 29808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_39
timestamp 1693170804
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1693170804
transform -1 0 30912 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_40
timestamp 1693170804
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1693170804
transform -1 0 30912 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_41
timestamp 1693170804
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1693170804
transform -1 0 30912 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_42
timestamp 1693170804
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1693170804
transform -1 0 30912 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_43
timestamp 1693170804
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1693170804
transform -1 0 30912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_44
timestamp 1693170804
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1693170804
transform -1 0 30912 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_45
timestamp 1693170804
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1693170804
transform -1 0 30912 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_46
timestamp 1693170804
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1693170804
transform -1 0 30912 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_47
timestamp 1693170804
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1693170804
transform -1 0 30912 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_48
timestamp 1693170804
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1693170804
transform -1 0 30912 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_49
timestamp 1693170804
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1693170804
transform -1 0 30912 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_50
timestamp 1693170804
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1693170804
transform -1 0 30912 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_51
timestamp 1693170804
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1693170804
transform -1 0 30912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_52
timestamp 1693170804
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1693170804
transform -1 0 30912 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_53
timestamp 1693170804
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1693170804
transform -1 0 30912 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_54
timestamp 1693170804
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1693170804
transform -1 0 30912 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_55
timestamp 1693170804
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1693170804
transform -1 0 30912 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_56
timestamp 1693170804
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1693170804
transform -1 0 30912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_57
timestamp 1693170804
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1693170804
transform -1 0 30912 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_58
timestamp 1693170804
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1693170804
transform -1 0 30912 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_59
timestamp 1693170804
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1693170804
transform -1 0 30912 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_60
timestamp 1693170804
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1693170804
transform -1 0 30912 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_61
timestamp 1693170804
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1693170804
transform -1 0 30912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_62
timestamp 1693170804
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1693170804
transform -1 0 30912 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_63
timestamp 1693170804
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1693170804
transform -1 0 30912 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_64
timestamp 1693170804
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1693170804
transform -1 0 30912 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_65
timestamp 1693170804
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1693170804
transform -1 0 30912 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_66
timestamp 1693170804
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1693170804
transform -1 0 30912 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_67
timestamp 1693170804
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1693170804
transform -1 0 30912 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_68
timestamp 1693170804
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1693170804
transform -1 0 30912 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_69
timestamp 1693170804
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1693170804
transform -1 0 30912 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_70
timestamp 1693170804
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1693170804
transform -1 0 30912 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_71
timestamp 1693170804
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1693170804
transform -1 0 30912 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_72
timestamp 1693170804
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1693170804
transform -1 0 30912 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_73
timestamp 1693170804
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1693170804
transform -1 0 30912 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_74
timestamp 1693170804
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1693170804
transform -1 0 30912 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_75
timestamp 1693170804
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1693170804
transform -1 0 30912 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_76
timestamp 1693170804
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1693170804
transform -1 0 30912 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_77
timestamp 1693170804
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1693170804
transform -1 0 30912 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_78 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_79
timestamp 1693170804
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_80
timestamp 1693170804
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_81
timestamp 1693170804
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_82
timestamp 1693170804
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_83
timestamp 1693170804
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_84
timestamp 1693170804
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_85
timestamp 1693170804
transform 1 0 21160 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_86
timestamp 1693170804
transform 1 0 23736 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_87
timestamp 1693170804
transform 1 0 26312 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1693170804
transform 1 0 28888 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_89
timestamp 1693170804
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_90
timestamp 1693170804
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_91
timestamp 1693170804
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_92
timestamp 1693170804
transform 1 0 21160 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_93
timestamp 1693170804
transform 1 0 26312 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_94
timestamp 1693170804
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_95
timestamp 1693170804
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_96
timestamp 1693170804
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_97
timestamp 1693170804
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_98
timestamp 1693170804
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_99
timestamp 1693170804
transform 1 0 28888 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_100
timestamp 1693170804
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_101
timestamp 1693170804
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_102
timestamp 1693170804
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_103
timestamp 1693170804
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_104
timestamp 1693170804
transform 1 0 26312 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 1693170804
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 1693170804
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 1693170804
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_108
timestamp 1693170804
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_109
timestamp 1693170804
transform 1 0 23736 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_110
timestamp 1693170804
transform 1 0 28888 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_111
timestamp 1693170804
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_112
timestamp 1693170804
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_113
timestamp 1693170804
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_114
timestamp 1693170804
transform 1 0 21160 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_115
timestamp 1693170804
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_116
timestamp 1693170804
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_117
timestamp 1693170804
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_118
timestamp 1693170804
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_119
timestamp 1693170804
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_120
timestamp 1693170804
transform 1 0 23736 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_121
timestamp 1693170804
transform 1 0 28888 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_122
timestamp 1693170804
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_123
timestamp 1693170804
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_124
timestamp 1693170804
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_125
timestamp 1693170804
transform 1 0 21160 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_126
timestamp 1693170804
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_127
timestamp 1693170804
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_128
timestamp 1693170804
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_129
timestamp 1693170804
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_130
timestamp 1693170804
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_131
timestamp 1693170804
transform 1 0 23736 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_132
timestamp 1693170804
transform 1 0 28888 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_133
timestamp 1693170804
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_134
timestamp 1693170804
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_135
timestamp 1693170804
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_136
timestamp 1693170804
transform 1 0 21160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_137
timestamp 1693170804
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_138
timestamp 1693170804
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_139
timestamp 1693170804
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_140
timestamp 1693170804
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 1693170804
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_142
timestamp 1693170804
transform 1 0 23736 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_143
timestamp 1693170804
transform 1 0 28888 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp 1693170804
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp 1693170804
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_146
timestamp 1693170804
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_147
timestamp 1693170804
transform 1 0 21160 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_148
timestamp 1693170804
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_149
timestamp 1693170804
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_150
timestamp 1693170804
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_151
timestamp 1693170804
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_152
timestamp 1693170804
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_153
timestamp 1693170804
transform 1 0 23736 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_154
timestamp 1693170804
transform 1 0 28888 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_155
timestamp 1693170804
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_156
timestamp 1693170804
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_157
timestamp 1693170804
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_158
timestamp 1693170804
transform 1 0 21160 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_159
timestamp 1693170804
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_160
timestamp 1693170804
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_161
timestamp 1693170804
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_162
timestamp 1693170804
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_163
timestamp 1693170804
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_164
timestamp 1693170804
transform 1 0 23736 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_165
timestamp 1693170804
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_166
timestamp 1693170804
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_167
timestamp 1693170804
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_168
timestamp 1693170804
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_169
timestamp 1693170804
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_170
timestamp 1693170804
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_171
timestamp 1693170804
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_172
timestamp 1693170804
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_173
timestamp 1693170804
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_174
timestamp 1693170804
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_175
timestamp 1693170804
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_176
timestamp 1693170804
transform 1 0 28888 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_177
timestamp 1693170804
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_178
timestamp 1693170804
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_179
timestamp 1693170804
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_180
timestamp 1693170804
transform 1 0 21160 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_181
timestamp 1693170804
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_182
timestamp 1693170804
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_183
timestamp 1693170804
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_184
timestamp 1693170804
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 1693170804
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_186
timestamp 1693170804
transform 1 0 23736 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_187
timestamp 1693170804
transform 1 0 28888 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_188
timestamp 1693170804
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_189
timestamp 1693170804
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_190
timestamp 1693170804
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_191
timestamp 1693170804
transform 1 0 21160 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_192
timestamp 1693170804
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_193
timestamp 1693170804
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_194
timestamp 1693170804
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_195
timestamp 1693170804
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_196
timestamp 1693170804
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_197
timestamp 1693170804
transform 1 0 23736 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_198
timestamp 1693170804
transform 1 0 28888 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_199
timestamp 1693170804
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_200
timestamp 1693170804
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_201
timestamp 1693170804
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_202
timestamp 1693170804
transform 1 0 21160 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_203
timestamp 1693170804
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_204
timestamp 1693170804
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_205
timestamp 1693170804
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_206
timestamp 1693170804
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_207
timestamp 1693170804
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_208
timestamp 1693170804
transform 1 0 23736 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_209
timestamp 1693170804
transform 1 0 28888 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_210
timestamp 1693170804
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_211
timestamp 1693170804
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_212
timestamp 1693170804
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_213
timestamp 1693170804
transform 1 0 21160 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_214
timestamp 1693170804
transform 1 0 26312 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_215
timestamp 1693170804
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_216
timestamp 1693170804
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_217
timestamp 1693170804
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_218
timestamp 1693170804
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_219
timestamp 1693170804
transform 1 0 23736 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_220
timestamp 1693170804
transform 1 0 28888 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_221
timestamp 1693170804
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_222
timestamp 1693170804
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_223
timestamp 1693170804
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_224
timestamp 1693170804
transform 1 0 21160 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_225
timestamp 1693170804
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_226
timestamp 1693170804
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_227
timestamp 1693170804
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_228
timestamp 1693170804
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_229
timestamp 1693170804
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_230
timestamp 1693170804
transform 1 0 23736 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_231
timestamp 1693170804
transform 1 0 28888 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_232
timestamp 1693170804
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_233
timestamp 1693170804
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_234
timestamp 1693170804
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_235
timestamp 1693170804
transform 1 0 21160 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_236
timestamp 1693170804
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_237
timestamp 1693170804
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_238
timestamp 1693170804
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_239
timestamp 1693170804
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_240
timestamp 1693170804
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_241
timestamp 1693170804
transform 1 0 23736 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_242
timestamp 1693170804
transform 1 0 28888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_243
timestamp 1693170804
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_244
timestamp 1693170804
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_245
timestamp 1693170804
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_246
timestamp 1693170804
transform 1 0 21160 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_247
timestamp 1693170804
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_248
timestamp 1693170804
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_249
timestamp 1693170804
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_250
timestamp 1693170804
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_251
timestamp 1693170804
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_252
timestamp 1693170804
transform 1 0 23736 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 1693170804
transform 1 0 28888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_254
timestamp 1693170804
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_255
timestamp 1693170804
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_256
timestamp 1693170804
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_257
timestamp 1693170804
transform 1 0 21160 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 1693170804
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_259
timestamp 1693170804
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_260
timestamp 1693170804
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_261
timestamp 1693170804
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_262
timestamp 1693170804
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 1693170804
transform 1 0 23736 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 1693170804
transform 1 0 28888 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_265
timestamp 1693170804
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_266
timestamp 1693170804
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_267
timestamp 1693170804
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 1693170804
transform 1 0 21160 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 1693170804
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_270
timestamp 1693170804
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_271
timestamp 1693170804
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_272
timestamp 1693170804
transform 1 0 13432 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 1693170804
transform 1 0 18584 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 1693170804
transform 1 0 23736 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1693170804
transform 1 0 28888 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_276
timestamp 1693170804
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_277
timestamp 1693170804
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 1693170804
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 1693170804
transform 1 0 21160 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1693170804
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_281
timestamp 1693170804
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_282
timestamp 1693170804
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 1693170804
transform 1 0 13432 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 1693170804
transform 1 0 18584 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1693170804
transform 1 0 23736 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 1693170804
transform 1 0 28888 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_287
timestamp 1693170804
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 1693170804
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 1693170804
transform 1 0 16008 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1693170804
transform 1 0 21160 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 1693170804
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_292
timestamp 1693170804
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 1693170804
transform 1 0 5704 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 1693170804
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1693170804
transform 1 0 10856 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 1693170804
transform 1 0 13432 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 1693170804
transform 1 0 16008 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_298
timestamp 1693170804
transform 1 0 18584 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_299
timestamp 1693170804
transform 1 0 21160 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_300
timestamp 1693170804
transform 1 0 23736 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_301
timestamp 1693170804
transform 1 0 26312 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_302
timestamp 1693170804
transform 1 0 28888 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1693170804
transform 1 0 12328 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_56
timestamp 1693170804
transform 1 0 13800 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_57
timestamp 1693170804
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_58
timestamp 1693170804
transform 1 0 9476 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_59
timestamp 1693170804
transform 1 0 5980 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_60
timestamp 1693170804
transform 1 0 11500 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_61
timestamp 1693170804
transform 1 0 12052 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_htfab_cell_tester_62
timestamp 1693170804
transform 1 0 12880 0 1 13600
box -38 -48 314 592
<< labels >>
flabel metal4 s 7982 496 8302 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15572 496 15892 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 23162 496 23482 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 30752 496 31072 21808 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4187 496 4507 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11777 496 12097 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19367 496 19687 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26957 496 27277 21808 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 26926 22104 26986 22304 0 FreeSans 480 90 0 0 clk
port 2 nsew signal input
flabel metal4 s 27478 22104 27538 22304 0 FreeSans 480 90 0 0 ena
port 3 nsew signal input
flabel metal4 s 26374 22104 26434 22304 0 FreeSans 480 90 0 0 rst_n
port 4 nsew signal input
flabel metal4 s 25822 22104 25882 22304 0 FreeSans 480 90 0 0 ui_in[0]
port 5 nsew signal input
flabel metal4 s 25270 22104 25330 22304 0 FreeSans 480 90 0 0 ui_in[1]
port 6 nsew signal input
flabel metal4 s 24718 22104 24778 22304 0 FreeSans 480 90 0 0 ui_in[2]
port 7 nsew signal input
flabel metal4 s 24166 22104 24226 22304 0 FreeSans 480 90 0 0 ui_in[3]
port 8 nsew signal input
flabel metal4 s 23614 22104 23674 22304 0 FreeSans 480 90 0 0 ui_in[4]
port 9 nsew signal input
flabel metal4 s 23062 22104 23122 22304 0 FreeSans 480 90 0 0 ui_in[5]
port 10 nsew signal input
flabel metal4 s 22510 22104 22570 22304 0 FreeSans 480 90 0 0 ui_in[6]
port 11 nsew signal input
flabel metal4 s 21958 22104 22018 22304 0 FreeSans 480 90 0 0 ui_in[7]
port 12 nsew signal input
flabel metal4 s 21406 22104 21466 22304 0 FreeSans 480 90 0 0 uio_in[0]
port 13 nsew signal input
flabel metal4 s 20854 22104 20914 22304 0 FreeSans 480 90 0 0 uio_in[1]
port 14 nsew signal input
flabel metal4 s 20302 22104 20362 22304 0 FreeSans 480 90 0 0 uio_in[2]
port 15 nsew signal input
flabel metal4 s 19750 22104 19810 22304 0 FreeSans 480 90 0 0 uio_in[3]
port 16 nsew signal input
flabel metal4 s 19198 22104 19258 22304 0 FreeSans 480 90 0 0 uio_in[4]
port 17 nsew signal input
flabel metal4 s 18646 22104 18706 22304 0 FreeSans 480 90 0 0 uio_in[5]
port 18 nsew signal input
flabel metal4 s 18094 22104 18154 22304 0 FreeSans 480 90 0 0 uio_in[6]
port 19 nsew signal input
flabel metal4 s 17542 22104 17602 22304 0 FreeSans 480 90 0 0 uio_in[7]
port 20 nsew signal input
flabel metal4 s 8158 22104 8218 22304 0 FreeSans 480 90 0 0 uio_oe[0]
port 21 nsew signal tristate
flabel metal4 s 7606 22104 7666 22304 0 FreeSans 480 90 0 0 uio_oe[1]
port 22 nsew signal tristate
flabel metal4 s 7054 22104 7114 22304 0 FreeSans 480 90 0 0 uio_oe[2]
port 23 nsew signal tristate
flabel metal4 s 6502 22104 6562 22304 0 FreeSans 480 90 0 0 uio_oe[3]
port 24 nsew signal tristate
flabel metal4 s 5950 22104 6010 22304 0 FreeSans 480 90 0 0 uio_oe[4]
port 25 nsew signal tristate
flabel metal4 s 5398 22104 5458 22304 0 FreeSans 480 90 0 0 uio_oe[5]
port 26 nsew signal tristate
flabel metal4 s 4846 22104 4906 22304 0 FreeSans 480 90 0 0 uio_oe[6]
port 27 nsew signal tristate
flabel metal4 s 4294 22104 4354 22304 0 FreeSans 480 90 0 0 uio_oe[7]
port 28 nsew signal tristate
flabel metal4 s 12574 22104 12634 22304 0 FreeSans 480 90 0 0 uio_out[0]
port 29 nsew signal tristate
flabel metal4 s 12022 22104 12082 22304 0 FreeSans 480 90 0 0 uio_out[1]
port 30 nsew signal tristate
flabel metal4 s 11470 22104 11530 22304 0 FreeSans 480 90 0 0 uio_out[2]
port 31 nsew signal tristate
flabel metal4 s 10918 22104 10978 22304 0 FreeSans 480 90 0 0 uio_out[3]
port 32 nsew signal tristate
flabel metal4 s 10366 22104 10426 22304 0 FreeSans 480 90 0 0 uio_out[4]
port 33 nsew signal tristate
flabel metal4 s 9814 22104 9874 22304 0 FreeSans 480 90 0 0 uio_out[5]
port 34 nsew signal tristate
flabel metal4 s 9262 22104 9322 22304 0 FreeSans 480 90 0 0 uio_out[6]
port 35 nsew signal tristate
flabel metal4 s 8710 22104 8770 22304 0 FreeSans 480 90 0 0 uio_out[7]
port 36 nsew signal tristate
flabel metal4 s 16990 22104 17050 22304 0 FreeSans 480 90 0 0 uo_out[0]
port 37 nsew signal tristate
flabel metal4 s 16438 22104 16498 22304 0 FreeSans 480 90 0 0 uo_out[1]
port 38 nsew signal tristate
flabel metal4 s 15886 22104 15946 22304 0 FreeSans 480 90 0 0 uo_out[2]
port 39 nsew signal tristate
flabel metal4 s 15334 22104 15394 22304 0 FreeSans 480 90 0 0 uo_out[3]
port 40 nsew signal tristate
flabel metal4 s 14782 22104 14842 22304 0 FreeSans 480 90 0 0 uo_out[4]
port 41 nsew signal tristate
flabel metal4 s 14230 22104 14290 22304 0 FreeSans 480 90 0 0 uo_out[5]
port 42 nsew signal tristate
flabel metal4 s 13678 22104 13738 22304 0 FreeSans 480 90 0 0 uo_out[6]
port 43 nsew signal tristate
flabel metal4 s 13126 22104 13186 22304 0 FreeSans 480 90 0 0 uo_out[7]
port 44 nsew signal tristate
rlabel via1 15812 21216 15812 21216 0 VGND
rlabel metal1 15732 21760 15732 21760 0 VPWR
rlabel metal1 30912 12954 30912 12954 0 _00_
rlabel metal1 23230 18938 23230 18938 0 _01_
rlabel metal1 23046 18802 23046 18802 0 _02_
rlabel metal1 22908 18666 22908 18666 0 _03_
rlabel metal1 19228 21454 19228 21454 0 _04_
rlabel metal1 30084 17102 30084 17102 0 ct.cw.source\[0\]
rlabel metal1 18492 16150 18492 16150 0 ct.cw.source\[1\]
rlabel metal1 16422 17646 16422 17646 0 ct.cw.source\[2\]
rlabel metal2 2254 14637 2254 14637 0 ct.cw.target\[0\]
rlabel metal2 2576 12036 2576 12036 0 ct.cw.target\[1\]
rlabel metal3 23644 14484 23644 14484 0 ct.cw.target\[2\]
rlabel metal1 1432 12809 1432 12809 0 ct.cw.target\[3\]
rlabel metal2 1978 12257 1978 12257 0 ct.cw.target\[4\]
rlabel metal1 14076 15946 14076 15946 0 ct.cw.target\[5\]
rlabel metal2 13662 17153 13662 17153 0 ct.cw.target\[6\]
rlabel metal1 11132 16626 11132 16626 0 ct.cw.target\[7\]
rlabel metal1 17158 13362 17158 13362 0 ct.ic.data_chain\[10\]
rlabel metal1 19412 15470 19412 15470 0 ct.ic.data_chain\[11\]
rlabel metal2 27416 21148 27416 21148 0 ct.ic.data_chain\[12\]
rlabel metal1 21068 21658 21068 21658 0 ct.ic.data_chain\[13\]
rlabel metal2 19274 21692 19274 21692 0 ct.ic.data_chain\[14\]
rlabel metal1 27278 21454 27278 21454 0 ct.ic.data_chain\[15\]
rlabel metal1 21390 21420 21390 21420 0 ct.ic.data_chain\[16\]
rlabel metal1 22632 14994 22632 14994 0 ct.ic.data_chain\[17\]
rlabel metal1 26404 19890 26404 19890 0 ct.ic.data_chain\[18\]
rlabel metal1 20470 17238 20470 17238 0 ct.ic.data_chain\[19\]
rlabel metal2 22770 16966 22770 16966 0 ct.ic.data_chain\[20\]
rlabel metal2 24702 19652 24702 19652 0 ct.ic.data_chain\[21\]
rlabel metal2 20746 17884 20746 17884 0 ct.ic.data_chain\[22\]
rlabel metal1 20286 16626 20286 16626 0 ct.ic.data_chain\[23\]
rlabel metal1 20516 18938 20516 18938 0 ct.ic.data_chain\[24\]
rlabel metal1 20332 18326 20332 18326 0 ct.ic.data_chain\[25\]
rlabel metal1 19780 17714 19780 17714 0 ct.ic.data_chain\[26\]
rlabel metal1 18814 18802 18814 18802 0 ct.ic.data_chain\[27\]
rlabel metal1 18814 18258 18814 18258 0 ct.ic.data_chain\[28\]
rlabel metal1 19550 19822 19550 19822 0 ct.ic.data_chain\[29\]
rlabel metal1 17480 18734 17480 18734 0 ct.ic.data_chain\[30\]
rlabel metal1 17388 19890 17388 19890 0 ct.ic.data_chain\[31\]
rlabel metal1 18906 19278 18906 19278 0 ct.ic.data_chain\[32\]
rlabel metal1 17066 18258 17066 18258 0 ct.ic.data_chain\[33\]
rlabel metal1 16146 18938 16146 18938 0 ct.ic.data_chain\[34\]
rlabel metal1 16054 19346 16054 19346 0 ct.ic.data_chain\[35\]
rlabel metal1 29486 9010 29486 9010 0 ct.ic.data_chain\[3\]
rlabel metal2 21390 11033 21390 11033 0 ct.ic.data_chain\[4\]
rlabel metal2 21758 14807 21758 14807 0 ct.ic.data_chain\[5\]
rlabel metal1 29486 13158 29486 13158 0 ct.ic.data_chain\[6\]
rlabel metal1 18906 20570 18906 20570 0 ct.ic.data_chain\[7\]
rlabel metal1 22264 13906 22264 13906 0 ct.ic.data_chain\[8\]
rlabel metal1 28474 13362 28474 13362 0 ct.ic.data_chain\[9\]
rlabel metal1 28290 21488 28290 21488 0 ct.ic.trig_chain\[0\]
rlabel metal1 18078 20298 18078 20298 0 ct.ic.trig_chain\[10\]
rlabel metal1 17204 20434 17204 20434 0 ct.ic.trig_chain\[11\]
rlabel metal1 14168 20570 14168 20570 0 ct.ic.trig_chain\[12\]
rlabel metal2 16882 16269 16882 16269 0 ct.ic.trig_chain\[1\]
rlabel metal1 26174 21386 26174 21386 0 ct.ic.trig_chain\[2\]
rlabel via2 19366 22083 19366 22083 0 ct.ic.trig_chain\[3\]
rlabel metal1 16882 21930 16882 21930 0 ct.ic.trig_chain\[4\]
rlabel metal1 19734 22168 19734 22168 0 ct.ic.trig_chain\[5\]
rlabel metal1 26634 19822 26634 19822 0 ct.ic.trig_chain\[6\]
rlabel metal1 20608 19890 20608 19890 0 ct.ic.trig_chain\[7\]
rlabel metal1 20516 18802 20516 18802 0 ct.ic.trig_chain\[8\]
rlabel metal1 18722 18666 18722 18666 0 ct.ic.trig_chain\[9\]
rlabel metal1 11684 19278 11684 19278 0 ct.oc.capture_buffer\[0\]
rlabel metal1 28060 20366 28060 20366 0 ct.oc.capture_buffer\[100\]
rlabel metal1 29854 14586 29854 14586 0 ct.oc.capture_buffer\[101\]
rlabel metal1 29762 13702 29762 13702 0 ct.oc.capture_buffer\[102\]
rlabel metal1 29762 18836 29762 18836 0 ct.oc.capture_buffer\[103\]
rlabel metal1 24748 13906 24748 13906 0 ct.oc.capture_buffer\[104\]
rlabel metal1 24564 14450 24564 14450 0 ct.oc.capture_buffer\[105\]
rlabel metal1 25208 13362 25208 13362 0 ct.oc.capture_buffer\[106\]
rlabel metal1 27554 13362 27554 13362 0 ct.oc.capture_buffer\[107\]
rlabel metal2 29578 16932 29578 16932 0 ct.oc.capture_buffer\[108\]
rlabel metal1 29164 14042 29164 14042 0 ct.oc.capture_buffer\[109\]
rlabel metal1 6716 20230 6716 20230 0 ct.oc.capture_buffer\[10\]
rlabel metal2 30130 15283 30130 15283 0 ct.oc.capture_buffer\[110\]
rlabel metal1 29762 14042 29762 14042 0 ct.oc.capture_buffer\[111\]
rlabel metal1 22356 13362 22356 13362 0 ct.oc.capture_buffer\[112\]
rlabel metal1 24291 12750 24291 12750 0 ct.oc.capture_buffer\[113\]
rlabel metal2 23506 12614 23506 12614 0 ct.oc.capture_buffer\[114\]
rlabel metal1 24543 11662 24543 11662 0 ct.oc.capture_buffer\[115\]
rlabel metal1 28750 11866 28750 11866 0 ct.oc.capture_buffer\[116\]
rlabel metal1 28474 12818 28474 12818 0 ct.oc.capture_buffer\[117\]
rlabel metal1 29118 14382 29118 14382 0 ct.oc.capture_buffer\[118\]
rlabel metal2 27508 13838 27508 13838 0 ct.oc.capture_buffer\[119\]
rlabel metal1 6302 18394 6302 18394 0 ct.oc.capture_buffer\[11\]
rlabel metal1 21712 12274 21712 12274 0 ct.oc.capture_buffer\[120\]
rlabel metal1 21620 11730 21620 11730 0 ct.oc.capture_buffer\[121\]
rlabel metal1 20838 12682 20838 12682 0 ct.oc.capture_buffer\[122\]
rlabel metal2 22816 10778 22816 10778 0 ct.oc.capture_buffer\[123\]
rlabel metal1 28842 7922 28842 7922 0 ct.oc.capture_buffer\[124\]
rlabel metal1 26588 11662 26588 11662 0 ct.oc.capture_buffer\[125\]
rlabel metal1 29026 6834 29026 6834 0 ct.oc.capture_buffer\[126\]
rlabel metal1 28106 8398 28106 8398 0 ct.oc.capture_buffer\[127\]
rlabel metal1 19044 12954 19044 12954 0 ct.oc.capture_buffer\[128\]
rlabel metal1 19596 12410 19596 12410 0 ct.oc.capture_buffer\[129\]
rlabel metal3 7751 20740 7751 20740 0 ct.oc.capture_buffer\[12\]
rlabel metal1 19550 13294 19550 13294 0 ct.oc.capture_buffer\[130\]
rlabel metal2 22034 10540 22034 10540 0 ct.oc.capture_buffer\[131\]
rlabel metal1 27968 10642 27968 10642 0 ct.oc.capture_buffer\[132\]
rlabel metal1 24426 10030 24426 10030 0 ct.oc.capture_buffer\[133\]
rlabel metal1 28336 9350 28336 9350 0 ct.oc.capture_buffer\[134\]
rlabel metal1 28796 9690 28796 9690 0 ct.oc.capture_buffer\[135\]
rlabel metal1 17204 10098 17204 10098 0 ct.oc.capture_buffer\[136\]
rlabel metal1 17388 12274 17388 12274 0 ct.oc.capture_buffer\[137\]
rlabel metal1 17388 11186 17388 11186 0 ct.oc.capture_buffer\[138\]
rlabel metal1 20562 10234 20562 10234 0 ct.oc.capture_buffer\[139\]
rlabel metal3 6647 19380 6647 19380 0 ct.oc.capture_buffer\[13\]
rlabel metal1 26358 9146 26358 9146 0 ct.oc.capture_buffer\[140\]
rlabel metal2 24610 10506 24610 10506 0 ct.oc.capture_buffer\[141\]
rlabel metal1 26312 8602 26312 8602 0 ct.oc.capture_buffer\[142\]
rlabel metal1 25576 9146 25576 9146 0 ct.oc.capture_buffer\[143\]
rlabel metal2 18170 9452 18170 9452 0 ct.oc.capture_buffer\[144\]
rlabel metal1 17756 9486 17756 9486 0 ct.oc.capture_buffer\[145\]
rlabel metal1 19090 7514 19090 7514 0 ct.oc.capture_buffer\[146\]
rlabel metal1 21344 9486 21344 9486 0 ct.oc.capture_buffer\[147\]
rlabel metal1 24288 8398 24288 8398 0 ct.oc.capture_buffer\[148\]
rlabel metal1 21988 8942 21988 8942 0 ct.oc.capture_buffer\[149\]
rlabel metal2 8970 13855 8970 13855 0 ct.oc.capture_buffer\[14\]
rlabel metal1 24380 7310 24380 7310 0 ct.oc.capture_buffer\[150\]
rlabel metal2 24242 9078 24242 9078 0 ct.oc.capture_buffer\[151\]
rlabel metal1 18722 6426 18722 6426 0 ct.oc.capture_buffer\[152\]
rlabel metal1 20010 7378 20010 7378 0 ct.oc.capture_buffer\[153\]
rlabel metal2 20838 8228 20838 8228 0 ct.oc.capture_buffer\[154\]
rlabel metal2 20562 6324 20562 6324 0 ct.oc.capture_buffer\[155\]
rlabel metal1 21666 8432 21666 8432 0 ct.oc.capture_buffer\[156\]
rlabel metal1 21436 6970 21436 6970 0 ct.oc.capture_buffer\[157\]
rlabel metal1 21482 6392 21482 6392 0 ct.oc.capture_buffer\[158\]
rlabel metal2 22218 6970 22218 6970 0 ct.oc.capture_buffer\[159\]
rlabel metal1 9292 13498 9292 13498 0 ct.oc.capture_buffer\[15\]
rlabel metal1 29256 3570 29256 3570 0 ct.oc.capture_buffer\[160\]
rlabel metal1 28750 4658 28750 4658 0 ct.oc.capture_buffer\[161\]
rlabel metal1 28060 5746 28060 5746 0 ct.oc.capture_buffer\[162\]
rlabel metal1 26634 6970 26634 6970 0 ct.oc.capture_buffer\[163\]
rlabel metal2 27462 6460 27462 6460 0 ct.oc.capture_buffer\[164\]
rlabel metal1 25254 6834 25254 6834 0 ct.oc.capture_buffer\[165\]
rlabel metal1 29302 6698 29302 6698 0 ct.oc.capture_buffer\[166\]
rlabel metal1 28014 6290 28014 6290 0 ct.oc.capture_buffer\[167\]
rlabel metal3 15479 11084 15479 11084 0 ct.oc.capture_buffer\[168\]
rlabel metal2 17802 7905 17802 7905 0 ct.oc.capture_buffer\[169\]
rlabel metal1 9384 14042 9384 14042 0 ct.oc.capture_buffer\[16\]
rlabel via2 14950 4029 14950 4029 0 ct.oc.capture_buffer\[170\]
rlabel metal2 29072 1836 29072 1836 0 ct.oc.capture_buffer\[171\]
rlabel metal1 28244 1326 28244 1326 0 ct.oc.capture_buffer\[172\]
rlabel metal1 28382 1938 28382 1938 0 ct.oc.capture_buffer\[173\]
rlabel metal2 17618 8381 17618 8381 0 ct.oc.capture_buffer\[174\]
rlabel metal1 20838 5304 20838 5304 0 ct.oc.capture_buffer\[175\]
rlabel metal3 12420 1904 12420 1904 0 ct.oc.capture_buffer\[176\]
rlabel metal2 5382 1921 5382 1921 0 ct.oc.capture_buffer\[177\]
rlabel metal1 20240 850 20240 850 0 ct.oc.capture_buffer\[178\]
rlabel metal1 27140 2482 27140 2482 0 ct.oc.capture_buffer\[179\]
rlabel metal2 9982 16388 9982 16388 0 ct.oc.capture_buffer\[17\]
rlabel metal1 26910 4114 26910 4114 0 ct.oc.capture_buffer\[180\]
rlabel metal1 26910 3026 26910 3026 0 ct.oc.capture_buffer\[181\]
rlabel metal1 2231 782 2231 782 0 ct.oc.capture_buffer\[182\]
rlabel metal2 21666 4352 21666 4352 0 ct.oc.capture_buffer\[183\]
rlabel metal1 21482 1904 21482 1904 0 ct.oc.capture_buffer\[184\]
rlabel metal1 20838 884 20838 884 0 ct.oc.capture_buffer\[185\]
rlabel metal2 24978 4454 24978 4454 0 ct.oc.capture_buffer\[186\]
rlabel metal2 24794 5508 24794 5508 0 ct.oc.capture_buffer\[187\]
rlabel metal1 24472 4794 24472 4794 0 ct.oc.capture_buffer\[188\]
rlabel metal1 24748 4114 24748 4114 0 ct.oc.capture_buffer\[189\]
rlabel metal1 8418 19346 8418 19346 0 ct.oc.capture_buffer\[18\]
rlabel metal2 22954 1122 22954 1122 0 ct.oc.capture_buffer\[190\]
rlabel metal2 25070 2349 25070 2349 0 ct.oc.capture_buffer\[191\]
rlabel metal1 24242 1360 24242 1360 0 ct.oc.capture_buffer\[192\]
rlabel metal1 25346 850 25346 850 0 ct.oc.capture_buffer\[193\]
rlabel metal1 24196 3570 24196 3570 0 ct.oc.capture_buffer\[194\]
rlabel metal1 24288 5134 24288 5134 0 ct.oc.capture_buffer\[195\]
rlabel metal1 22632 5746 22632 5746 0 ct.oc.capture_buffer\[196\]
rlabel metal1 22770 4624 22770 4624 0 ct.oc.capture_buffer\[197\]
rlabel metal1 23046 782 23046 782 0 ct.oc.capture_buffer\[198\]
rlabel metal1 24518 3026 24518 3026 0 ct.oc.capture_buffer\[199\]
rlabel metal1 9338 17714 9338 17714 0 ct.oc.capture_buffer\[19\]
rlabel metal1 17802 19414 17802 19414 0 ct.oc.capture_buffer\[1\]
rlabel metal1 23138 1972 23138 1972 0 ct.oc.capture_buffer\[200\]
rlabel metal2 22862 1530 22862 1530 0 ct.oc.capture_buffer\[201\]
rlabel metal1 21942 3570 21942 3570 0 ct.oc.capture_buffer\[202\]
rlabel metal1 20930 4114 20930 4114 0 ct.oc.capture_buffer\[203\]
rlabel metal1 20746 5882 20746 5882 0 ct.oc.capture_buffer\[204\]
rlabel metal2 21666 5406 21666 5406 0 ct.oc.capture_buffer\[205\]
rlabel metal2 22034 2244 22034 2244 0 ct.oc.capture_buffer\[206\]
rlabel metal1 21620 3026 21620 3026 0 ct.oc.capture_buffer\[207\]
rlabel metal1 20010 1530 20010 1530 0 ct.oc.capture_buffer\[208\]
rlabel metal1 19964 1326 19964 1326 0 ct.oc.capture_buffer\[209\]
rlabel metal2 12006 13481 12006 13481 0 ct.oc.capture_buffer\[20\]
rlabel metal2 19090 4012 19090 4012 0 ct.oc.capture_buffer\[210\]
rlabel metal1 19320 5746 19320 5746 0 ct.oc.capture_buffer\[211\]
rlabel metal1 19137 5134 19137 5134 0 ct.oc.capture_buffer\[212\]
rlabel metal2 19090 5372 19090 5372 0 ct.oc.capture_buffer\[213\]
rlabel metal2 21298 1632 21298 1632 0 ct.oc.capture_buffer\[214\]
rlabel metal1 19780 3026 19780 3026 0 ct.oc.capture_buffer\[215\]
rlabel metal1 17480 1938 17480 1938 0 ct.oc.capture_buffer\[216\]
rlabel metal1 16514 986 16514 986 0 ct.oc.capture_buffer\[217\]
rlabel metal1 17526 3162 17526 3162 0 ct.oc.capture_buffer\[218\]
rlabel metal1 17388 4590 17388 4590 0 ct.oc.capture_buffer\[219\]
rlabel metal1 4508 19822 4508 19822 0 ct.oc.capture_buffer\[21\]
rlabel metal1 17112 5746 17112 5746 0 ct.oc.capture_buffer\[220\]
rlabel metal1 17572 5134 17572 5134 0 ct.oc.capture_buffer\[221\]
rlabel metal1 18262 986 18262 986 0 ct.oc.capture_buffer\[222\]
rlabel metal1 18032 2074 18032 2074 0 ct.oc.capture_buffer\[223\]
rlabel metal1 13984 986 13984 986 0 ct.oc.capture_buffer\[224\]
rlabel metal1 14582 1360 14582 1360 0 ct.oc.capture_buffer\[225\]
rlabel metal1 14536 3570 14536 3570 0 ct.oc.capture_buffer\[226\]
rlabel metal1 14490 5746 14490 5746 0 ct.oc.capture_buffer\[227\]
rlabel metal1 14164 5134 14164 5134 0 ct.oc.capture_buffer\[228\]
rlabel metal1 14490 4590 14490 4590 0 ct.oc.capture_buffer\[229\]
rlabel metal2 1886 20961 1886 20961 0 ct.oc.capture_buffer\[22\]
rlabel metal1 13110 2380 13110 2380 0 ct.oc.capture_buffer\[230\]
rlabel metal1 14398 3026 14398 3026 0 ct.oc.capture_buffer\[231\]
rlabel metal1 9384 646 9384 646 0 ct.oc.capture_buffer\[232\]
rlabel metal1 12374 2448 12374 2448 0 ct.oc.capture_buffer\[233\]
rlabel metal1 11868 3570 11868 3570 0 ct.oc.capture_buffer\[234\]
rlabel metal1 12052 5746 12052 5746 0 ct.oc.capture_buffer\[235\]
rlabel metal1 11776 5134 11776 5134 0 ct.oc.capture_buffer\[236\]
rlabel metal1 12328 4658 12328 4658 0 ct.oc.capture_buffer\[237\]
rlabel metal2 10994 1530 10994 1530 0 ct.oc.capture_buffer\[238\]
rlabel metal1 11914 3026 11914 3026 0 ct.oc.capture_buffer\[239\]
rlabel metal2 13386 13889 13386 13889 0 ct.oc.capture_buffer\[23\]
rlabel metal1 6486 986 6486 986 0 ct.oc.capture_buffer\[240\]
rlabel metal2 9338 6086 9338 6086 0 ct.oc.capture_buffer\[241\]
rlabel metal1 9384 2482 9384 2482 0 ct.oc.capture_buffer\[242\]
rlabel metal1 10212 4590 10212 4590 0 ct.oc.capture_buffer\[243\]
rlabel metal1 9752 5202 9752 5202 0 ct.oc.capture_buffer\[244\]
rlabel metal1 10350 4046 10350 4046 0 ct.oc.capture_buffer\[245\]
rlabel metal1 6026 646 6026 646 0 ct.oc.capture_buffer\[246\]
rlabel metal1 9568 2958 9568 2958 0 ct.oc.capture_buffer\[247\]
rlabel metal1 6808 850 6808 850 0 ct.oc.capture_buffer\[248\]
rlabel metal3 4876 2516 4876 2516 0 ct.oc.capture_buffer\[249\]
rlabel metal1 6762 17170 6762 17170 0 ct.oc.capture_buffer\[24\]
rlabel metal1 6808 3434 6808 3434 0 ct.oc.capture_buffer\[250\]
rlabel metal1 8510 3502 8510 3502 0 ct.oc.capture_buffer\[251\]
rlabel metal1 7314 5202 7314 5202 0 ct.oc.capture_buffer\[252\]
rlabel metal1 8142 4556 8142 4556 0 ct.oc.capture_buffer\[253\]
rlabel metal1 7866 1258 7866 1258 0 ct.oc.capture_buffer\[254\]
rlabel metal1 5244 986 5244 986 0 ct.oc.capture_buffer\[255\]
rlabel metal1 17204 7854 17204 7854 0 ct.oc.capture_buffer\[256\]
rlabel metal1 2162 1938 2162 1938 0 ct.oc.capture_buffer\[257\]
rlabel metal1 4830 3570 4830 3570 0 ct.oc.capture_buffer\[258\]
rlabel metal1 6716 4114 6716 4114 0 ct.oc.capture_buffer\[259\]
rlabel metal1 6624 17714 6624 17714 0 ct.oc.capture_buffer\[25\]
rlabel metal1 5060 5134 5060 5134 0 ct.oc.capture_buffer\[260\]
rlabel metal1 6624 4658 6624 4658 0 ct.oc.capture_buffer\[261\]
rlabel metal2 2070 884 2070 884 0 ct.oc.capture_buffer\[262\]
rlabel metal1 6440 1870 6440 1870 0 ct.oc.capture_buffer\[263\]
rlabel metal2 19826 10965 19826 10965 0 ct.oc.capture_buffer\[264\]
rlabel via3 1725 13804 1725 13804 0 ct.oc.capture_buffer\[265\]
rlabel metal2 2438 3842 2438 3842 0 ct.oc.capture_buffer\[266\]
rlabel metal2 5842 4148 5842 4148 0 ct.oc.capture_buffer\[267\]
rlabel metal1 5060 4046 5060 4046 0 ct.oc.capture_buffer\[268\]
rlabel metal1 3358 2006 3358 2006 0 ct.oc.capture_buffer\[269\]
rlabel metal1 6578 18802 6578 18802 0 ct.oc.capture_buffer\[26\]
rlabel metal1 13064 6426 13064 6426 0 ct.oc.capture_buffer\[270\]
rlabel metal2 16146 6477 16146 6477 0 ct.oc.capture_buffer\[271\]
rlabel metal1 15824 12954 15824 12954 0 ct.oc.capture_buffer\[272\]
rlabel metal2 6854 4726 6854 4726 0 ct.oc.capture_buffer\[273\]
rlabel metal1 1840 4046 1840 4046 0 ct.oc.capture_buffer\[274\]
rlabel metal1 1058 3706 1058 3706 0 ct.oc.capture_buffer\[275\]
rlabel metal1 1150 2618 1150 2618 0 ct.oc.capture_buffer\[276\]
rlabel via1 4094 5219 4094 5219 0 ct.oc.capture_buffer\[277\]
rlabel metal1 11454 6698 11454 6698 0 ct.oc.capture_buffer\[278\]
rlabel metal2 11730 6273 11730 6273 0 ct.oc.capture_buffer\[279\]
rlabel metal1 6532 18190 6532 18190 0 ct.oc.capture_buffer\[27\]
rlabel metal1 1426 5882 1426 5882 0 ct.oc.capture_buffer\[280\]
rlabel metal1 6118 6936 6118 6936 0 ct.oc.capture_buffer\[281\]
rlabel metal1 1380 4794 1380 4794 0 ct.oc.capture_buffer\[282\]
rlabel metal1 4968 6290 4968 6290 0 ct.oc.capture_buffer\[283\]
rlabel metal1 4646 6834 4646 6834 0 ct.oc.capture_buffer\[284\]
rlabel metal2 5842 7412 5842 7412 0 ct.oc.capture_buffer\[285\]
rlabel metal1 2323 6766 2323 6766 0 ct.oc.capture_buffer\[286\]
rlabel metal1 4089 7310 4089 7310 0 ct.oc.capture_buffer\[287\]
rlabel metal2 9384 7854 9384 7854 0 ct.oc.capture_buffer\[288\]
rlabel metal1 7314 7378 7314 7378 0 ct.oc.capture_buffer\[289\]
rlabel metal2 2024 19822 2024 19822 0 ct.oc.capture_buffer\[28\]
rlabel metal2 7222 7684 7222 7684 0 ct.oc.capture_buffer\[290\]
rlabel metal1 7176 7922 7176 7922 0 ct.oc.capture_buffer\[291\]
rlabel metal2 6854 7548 6854 7548 0 ct.oc.capture_buffer\[292\]
rlabel metal1 10396 6290 10396 6290 0 ct.oc.capture_buffer\[293\]
rlabel metal1 10810 6698 10810 6698 0 ct.oc.capture_buffer\[294\]
rlabel metal1 9476 6834 9476 6834 0 ct.oc.capture_buffer\[295\]
rlabel metal1 16376 7922 16376 7922 0 ct.oc.capture_buffer\[296\]
rlabel metal2 13754 6970 13754 6970 0 ct.oc.capture_buffer\[297\]
rlabel metal1 13432 6426 13432 6426 0 ct.oc.capture_buffer\[298\]
rlabel metal1 14999 6222 14999 6222 0 ct.oc.capture_buffer\[299\]
rlabel metal1 9890 13498 9890 13498 0 ct.oc.capture_buffer\[29\]
rlabel metal1 13386 21046 13386 21046 0 ct.oc.capture_buffer\[2\]
rlabel metal1 14858 6970 14858 6970 0 ct.oc.capture_buffer\[300\]
rlabel metal1 12696 6426 12696 6426 0 ct.oc.capture_buffer\[301\]
rlabel metal2 12742 8092 12742 8092 0 ct.oc.capture_buffer\[302\]
rlabel metal1 13018 6834 13018 6834 0 ct.oc.capture_buffer\[303\]
rlabel metal2 14582 10438 14582 10438 0 ct.oc.capture_buffer\[304\]
rlabel metal2 16146 10132 16146 10132 0 ct.oc.capture_buffer\[305\]
rlabel metal1 14674 8466 14674 8466 0 ct.oc.capture_buffer\[306\]
rlabel metal1 15318 9146 15318 9146 0 ct.oc.capture_buffer\[307\]
rlabel metal1 15318 9010 15318 9010 0 ct.oc.capture_buffer\[308\]
rlabel metal1 12604 8262 12604 8262 0 ct.oc.capture_buffer\[309\]
rlabel metal3 7314 17748 7314 17748 0 ct.oc.capture_buffer\[30\]
rlabel metal1 11500 9010 11500 9010 0 ct.oc.capture_buffer\[310\]
rlabel metal1 11270 9146 11270 9146 0 ct.oc.capture_buffer\[311\]
rlabel metal2 13202 12517 13202 12517 0 ct.oc.capture_buffer\[312\]
rlabel metal2 13294 11509 13294 11509 0 ct.oc.capture_buffer\[313\]
rlabel metal1 13984 12750 13984 12750 0 ct.oc.capture_buffer\[314\]
rlabel metal1 13984 11662 13984 11662 0 ct.oc.capture_buffer\[315\]
rlabel metal1 13110 12954 13110 12954 0 ct.oc.capture_buffer\[316\]
rlabel metal1 10074 9554 10074 9554 0 ct.oc.capture_buffer\[317\]
rlabel metal1 10212 8398 10212 8398 0 ct.oc.capture_buffer\[318\]
rlabel metal1 9798 10098 9798 10098 0 ct.oc.capture_buffer\[319\]
rlabel metal3 2484 3740 2484 3740 0 ct.oc.capture_buffer\[31\]
rlabel metal1 10396 12818 10396 12818 0 ct.oc.capture_buffer\[320\]
rlabel metal1 10534 10642 10534 10642 0 ct.oc.capture_buffer\[321\]
rlabel metal1 10672 13498 10672 13498 0 ct.oc.capture_buffer\[322\]
rlabel metal2 10258 12954 10258 12954 0 ct.oc.capture_buffer\[323\]
rlabel metal1 9384 12274 9384 12274 0 ct.oc.capture_buffer\[324\]
rlabel metal1 7958 11526 7958 11526 0 ct.oc.capture_buffer\[325\]
rlabel metal1 7268 9146 7268 9146 0 ct.oc.capture_buffer\[326\]
rlabel metal1 7820 8602 7820 8602 0 ct.oc.capture_buffer\[327\]
rlabel metal2 7222 12138 7222 12138 0 ct.oc.capture_buffer\[328\]
rlabel metal1 7360 11186 7360 11186 0 ct.oc.capture_buffer\[329\]
rlabel metal1 12972 21590 12972 21590 0 ct.oc.capture_buffer\[32\]
rlabel metal1 7636 11866 7636 11866 0 ct.oc.capture_buffer\[330\]
rlabel metal1 8142 12954 8142 12954 0 ct.oc.capture_buffer\[331\]
rlabel metal1 6808 12818 6808 12818 0 ct.oc.capture_buffer\[332\]
rlabel metal1 6072 9690 6072 9690 0 ct.oc.capture_buffer\[333\]
rlabel metal1 6256 11662 6256 11662 0 ct.oc.capture_buffer\[334\]
rlabel metal1 6256 8398 6256 8398 0 ct.oc.capture_buffer\[335\]
rlabel metal1 5060 13294 5060 13294 0 ct.oc.capture_buffer\[336\]
rlabel metal1 5520 13498 5520 13498 0 ct.oc.capture_buffer\[337\]
rlabel metal1 4186 11322 4186 11322 0 ct.oc.capture_buffer\[338\]
rlabel metal1 4416 12750 4416 12750 0 ct.oc.capture_buffer\[339\]
rlabel metal1 11454 11050 11454 11050 0 ct.oc.capture_buffer\[33\]
rlabel metal1 3726 14042 3726 14042 0 ct.oc.capture_buffer\[340\]
rlabel metal2 5750 8772 5750 8772 0 ct.oc.capture_buffer\[341\]
rlabel metal2 4922 9860 4922 9860 0 ct.oc.capture_buffer\[342\]
rlabel metal1 4508 9146 4508 9146 0 ct.oc.capture_buffer\[343\]
rlabel metal1 1751 13362 1751 13362 0 ct.oc.capture_buffer\[344\]
rlabel metal1 1104 15334 1104 15334 0 ct.oc.capture_buffer\[345\]
rlabel metal1 1656 11186 1656 11186 0 ct.oc.capture_buffer\[346\]
rlabel metal1 1656 12750 1656 12750 0 ct.oc.capture_buffer\[347\]
rlabel metal2 2070 12138 2070 12138 0 ct.oc.capture_buffer\[348\]
rlabel metal2 874 9418 874 9418 0 ct.oc.capture_buffer\[349\]
rlabel metal1 4784 17646 4784 17646 0 ct.oc.capture_buffer\[34\]
rlabel metal1 1196 6630 1196 6630 0 ct.oc.capture_buffer\[350\]
rlabel metal1 1288 8058 1288 8058 0 ct.oc.capture_buffer\[351\]
rlabel metal1 4830 16626 4830 16626 0 ct.oc.capture_buffer\[35\]
rlabel metal1 8142 11798 8142 11798 0 ct.oc.capture_buffer\[36\]
rlabel metal2 2438 17153 2438 17153 0 ct.oc.capture_buffer\[37\]
rlabel metal2 2070 16813 2070 16813 0 ct.oc.capture_buffer\[38\]
rlabel metal1 8418 11866 8418 11866 0 ct.oc.capture_buffer\[39\]
rlabel metal2 874 21335 874 21335 0 ct.oc.capture_buffer\[3\]
rlabel metal1 8602 14042 8602 14042 0 ct.oc.capture_buffer\[40\]
rlabel metal1 4830 11322 4830 11322 0 ct.oc.capture_buffer\[41\]
rlabel metal1 9269 14314 9269 14314 0 ct.oc.capture_buffer\[42\]
rlabel metal1 506 17408 506 17408 0 ct.oc.capture_buffer\[43\]
rlabel metal1 6762 13192 6762 13192 0 ct.oc.capture_buffer\[44\]
rlabel metal1 8694 11560 8694 11560 0 ct.oc.capture_buffer\[45\]
rlabel metal2 7590 12801 7590 12801 0 ct.oc.capture_buffer\[46\]
rlabel metal1 3726 16116 3726 16116 0 ct.oc.capture_buffer\[47\]
rlabel metal1 6854 13872 6854 13872 0 ct.oc.capture_buffer\[48\]
rlabel metal1 6026 14586 6026 14586 0 ct.oc.capture_buffer\[49\]
rlabel metal1 4508 18666 4508 18666 0 ct.oc.capture_buffer\[4\]
rlabel metal1 6440 14314 6440 14314 0 ct.oc.capture_buffer\[50\]
rlabel metal1 8050 14042 8050 14042 0 ct.oc.capture_buffer\[51\]
rlabel metal1 9384 14586 9384 14586 0 ct.oc.capture_buffer\[52\]
rlabel metal1 9154 14042 9154 14042 0 ct.oc.capture_buffer\[53\]
rlabel metal2 9706 14756 9706 14756 0 ct.oc.capture_buffer\[54\]
rlabel metal1 9016 16626 9016 16626 0 ct.oc.capture_buffer\[55\]
rlabel metal1 12604 14042 12604 14042 0 ct.oc.capture_buffer\[56\]
rlabel metal1 11178 14586 11178 14586 0 ct.oc.capture_buffer\[57\]
rlabel metal1 11684 14586 11684 14586 0 ct.oc.capture_buffer\[58\]
rlabel metal2 12374 14178 12374 14178 0 ct.oc.capture_buffer\[59\]
rlabel metal3 9706 21012 9706 21012 0 ct.oc.capture_buffer\[5\]
rlabel metal2 12926 16932 12926 16932 0 ct.oc.capture_buffer\[60\]
rlabel metal1 11684 17102 11684 17102 0 ct.oc.capture_buffer\[61\]
rlabel metal1 11730 17714 11730 17714 0 ct.oc.capture_buffer\[62\]
rlabel metal1 12328 16558 12328 16558 0 ct.oc.capture_buffer\[63\]
rlabel metal1 15364 13498 15364 13498 0 ct.oc.capture_buffer\[64\]
rlabel metal1 15778 13464 15778 13464 0 ct.oc.capture_buffer\[65\]
rlabel metal1 16790 13464 16790 13464 0 ct.oc.capture_buffer\[66\]
rlabel metal1 15640 14382 15640 14382 0 ct.oc.capture_buffer\[67\]
rlabel metal1 14628 16558 14628 16558 0 ct.oc.capture_buffer\[68\]
rlabel metal2 14950 17034 14950 17034 0 ct.oc.capture_buffer\[69\]
rlabel metal3 7337 18020 7337 18020 0 ct.oc.capture_buffer\[6\]
rlabel metal1 12650 16184 12650 16184 0 ct.oc.capture_buffer\[70\]
rlabel metal2 14582 17663 14582 17663 0 ct.oc.capture_buffer\[71\]
rlabel metal1 17710 13498 17710 13498 0 ct.oc.capture_buffer\[72\]
rlabel metal1 18354 14042 18354 14042 0 ct.oc.capture_buffer\[73\]
rlabel metal1 17756 13226 17756 13226 0 ct.oc.capture_buffer\[74\]
rlabel metal1 18538 14382 18538 14382 0 ct.oc.capture_buffer\[75\]
rlabel metal1 15548 15878 15548 15878 0 ct.oc.capture_buffer\[76\]
rlabel metal1 19182 16012 19182 16012 0 ct.oc.capture_buffer\[77\]
rlabel metal1 18124 17714 18124 17714 0 ct.oc.capture_buffer\[78\]
rlabel metal1 17756 16558 17756 16558 0 ct.oc.capture_buffer\[79\]
rlabel metal1 12098 11866 12098 11866 0 ct.oc.capture_buffer\[7\]
rlabel metal1 20654 13906 20654 13906 0 ct.oc.capture_buffer\[80\]
rlabel metal1 20102 14586 20102 14586 0 ct.oc.capture_buffer\[81\]
rlabel metal1 20286 14552 20286 14552 0 ct.oc.capture_buffer\[82\]
rlabel metal1 21666 14450 21666 14450 0 ct.oc.capture_buffer\[83\]
rlabel metal2 22954 18122 22954 18122 0 ct.oc.capture_buffer\[84\]
rlabel metal1 19826 14586 19826 14586 0 ct.oc.capture_buffer\[85\]
rlabel metal1 22954 16694 22954 16694 0 ct.oc.capture_buffer\[86\]
rlabel metal1 21689 17170 21689 17170 0 ct.oc.capture_buffer\[87\]
rlabel metal2 20654 13651 20654 13651 0 ct.oc.capture_buffer\[88\]
rlabel via2 19550 13957 19550 13957 0 ct.oc.capture_buffer\[89\]
rlabel metal1 8694 16762 8694 16762 0 ct.oc.capture_buffer\[8\]
rlabel metal1 21022 13498 21022 13498 0 ct.oc.capture_buffer\[90\]
rlabel metal1 21666 13158 21666 13158 0 ct.oc.capture_buffer\[91\]
rlabel metal1 30406 18088 30406 18088 0 ct.oc.capture_buffer\[92\]
rlabel metal1 27879 17646 27879 17646 0 ct.oc.capture_buffer\[93\]
rlabel metal1 25990 17170 25990 17170 0 ct.oc.capture_buffer\[94\]
rlabel metal1 26266 18190 26266 18190 0 ct.oc.capture_buffer\[95\]
rlabel metal1 29348 15130 29348 15130 0 ct.oc.capture_buffer\[96\]
rlabel metal1 29900 13498 29900 13498 0 ct.oc.capture_buffer\[97\]
rlabel metal1 28934 16081 28934 16081 0 ct.oc.capture_buffer\[98\]
rlabel metal1 29854 15674 29854 15674 0 ct.oc.capture_buffer\[99\]
rlabel metal1 11132 18190 11132 18190 0 ct.oc.capture_buffer\[9\]
rlabel metal2 12466 20009 12466 20009 0 ct.oc.data_chain\[0\]
rlabel metal1 24725 17646 24725 17646 0 ct.oc.data_chain\[100\]
rlabel via1 26911 17646 26911 17646 0 ct.oc.data_chain\[101\]
rlabel viali 25255 17168 25255 17168 0 ct.oc.data_chain\[102\]
rlabel metal1 25645 18258 25645 18258 0 ct.oc.data_chain\[103\]
rlabel metal1 26358 13770 26358 13770 0 ct.oc.data_chain\[104\]
rlabel viali 26545 14985 26545 14985 0 ct.oc.data_chain\[105\]
rlabel metal1 26451 16082 26451 16082 0 ct.oc.data_chain\[106\]
rlabel metal1 27393 18734 27393 18734 0 ct.oc.data_chain\[107\]
rlabel metal1 27991 20434 27991 20434 0 ct.oc.data_chain\[108\]
rlabel metal1 28865 20910 28865 20910 0 ct.oc.data_chain\[109\]
rlabel metal1 10488 20570 10488 20570 0 ct.oc.data_chain\[10\]
rlabel metal1 25875 19346 25875 19346 0 ct.oc.data_chain\[110\]
rlabel metal1 24104 16218 24104 16218 0 ct.oc.data_chain\[111\]
rlabel metal1 24381 13906 24381 13906 0 ct.oc.data_chain\[112\]
rlabel metal1 25185 14382 25185 14382 0 ct.oc.data_chain\[113\]
rlabel metal1 25001 13294 25001 13294 0 ct.oc.data_chain\[114\]
rlabel metal1 26036 11866 26036 11866 0 ct.oc.data_chain\[115\]
rlabel metal2 29118 16796 29118 16796 0 ct.oc.data_chain\[116\]
rlabel metal1 28405 16558 28405 16558 0 ct.oc.data_chain\[117\]
rlabel metal1 28589 19346 28589 19346 0 ct.oc.data_chain\[118\]
rlabel metal2 22034 15827 22034 15827 0 ct.oc.data_chain\[119\]
rlabel metal1 13663 19346 13663 19346 0 ct.oc.data_chain\[11\]
rlabel metal1 22517 13294 22517 13294 0 ct.oc.data_chain\[120\]
rlabel metal1 24289 12818 24289 12818 0 ct.oc.data_chain\[121\]
rlabel via1 23967 12206 23967 12206 0 ct.oc.data_chain\[122\]
rlabel viali 24472 11729 24472 11729 0 ct.oc.data_chain\[123\]
rlabel metal1 28681 12206 28681 12206 0 ct.oc.data_chain\[124\]
rlabel metal1 27209 12818 27209 12818 0 ct.oc.data_chain\[125\]
rlabel metal1 30590 14382 30590 14382 0 ct.oc.data_chain\[126\]
rlabel metal2 27416 13124 27416 13124 0 ct.oc.data_chain\[127\]
rlabel metal1 20930 11594 20930 11594 0 ct.oc.data_chain\[128\]
rlabel metal1 21069 11730 21069 11730 0 ct.oc.data_chain\[129\]
rlabel via1 8971 19822 8971 19822 0 ct.oc.data_chain\[12\]
rlabel metal1 20885 12818 20885 12818 0 ct.oc.data_chain\[130\]
rlabel viali 22865 11119 22865 11119 0 ct.oc.data_chain\[131\]
rlabel metal1 28155 7854 28155 7854 0 ct.oc.data_chain\[132\]
rlabel viali 26680 11729 26680 11729 0 ct.oc.data_chain\[133\]
rlabel metal1 28198 11050 28198 11050 0 ct.oc.data_chain\[134\]
rlabel metal1 27761 8466 27761 8466 0 ct.oc.data_chain\[135\]
rlabel metal1 19185 11695 19185 11695 0 ct.oc.data_chain\[136\]
rlabel metal1 19137 12818 19137 12818 0 ct.oc.data_chain\[137\]
rlabel via1 18815 13294 18815 13294 0 ct.oc.data_chain\[138\]
rlabel via1 21759 10030 21759 10030 0 ct.oc.data_chain\[139\]
rlabel metal2 7866 20536 7866 20536 0 ct.oc.data_chain\[13\]
rlabel metal1 26749 10642 26749 10642 0 ct.oc.data_chain\[140\]
rlabel metal1 24173 10030 24173 10030 0 ct.oc.data_chain\[141\]
rlabel viali 26953 11136 26953 11136 0 ct.oc.data_chain\[142\]
rlabel metal1 26680 9690 26680 9690 0 ct.oc.data_chain\[143\]
rlabel metal2 18814 9418 18814 9418 0 ct.oc.data_chain\[144\]
rlabel metal1 17779 12206 17779 12206 0 ct.oc.data_chain\[145\]
rlabel metal1 19021 11118 19021 11118 0 ct.oc.data_chain\[146\]
rlabel metal2 22770 10166 22770 10166 0 ct.oc.data_chain\[147\]
rlabel metal1 26497 9554 26497 9554 0 ct.oc.data_chain\[148\]
rlabel metal1 23046 9146 23046 9146 0 ct.oc.data_chain\[149\]
rlabel metal1 6877 20434 6877 20434 0 ct.oc.data_chain\[14\]
rlabel metal1 26404 7514 26404 7514 0 ct.oc.data_chain\[150\]
rlabel via1 24887 9554 24887 9554 0 ct.oc.data_chain\[151\]
rlabel metal1 19067 8942 19067 8942 0 ct.oc.data_chain\[152\]
rlabel metal1 20240 7174 20240 7174 0 ct.oc.data_chain\[153\]
rlabel metal1 19918 8602 19918 8602 0 ct.oc.data_chain\[154\]
rlabel metal1 21253 9554 21253 9554 0 ct.oc.data_chain\[155\]
rlabel metal1 24013 8466 24013 8466 0 ct.oc.data_chain\[156\]
rlabel viali 21806 8944 21806 8944 0 ct.oc.data_chain\[157\]
rlabel metal1 24863 7378 24863 7378 0 ct.oc.data_chain\[158\]
rlabel metal1 23782 7514 23782 7514 0 ct.oc.data_chain\[159\]
rlabel via1 11455 21522 11455 21522 0 ct.oc.data_chain\[15\]
rlabel metal1 20562 8806 20562 8806 0 ct.oc.data_chain\[160\]
rlabel metal1 20240 7310 20240 7310 0 ct.oc.data_chain\[161\]
rlabel metal2 19274 8415 19274 8415 0 ct.oc.data_chain\[162\]
rlabel via2 20746 6851 20746 6851 0 ct.oc.data_chain\[163\]
rlabel metal1 22747 8466 22747 8466 0 ct.oc.data_chain\[164\]
rlabel metal1 21794 7889 21794 7889 0 ct.oc.data_chain\[165\]
rlabel metal2 23966 7412 23966 7412 0 ct.oc.data_chain\[166\]
rlabel metal1 23782 7276 23782 7276 0 ct.oc.data_chain\[167\]
rlabel via2 6026 2907 6026 2907 0 ct.oc.data_chain\[168\]
rlabel metal2 18538 9707 18538 9707 0 ct.oc.data_chain\[169\]
rlabel metal1 10534 18768 10534 18768 0 ct.oc.data_chain\[16\]
rlabel metal2 22402 5117 22402 5117 0 ct.oc.data_chain\[170\]
rlabel metal2 28566 1873 28566 1873 0 ct.oc.data_chain\[171\]
rlabel metal1 28290 2074 28290 2074 0 ct.oc.data_chain\[172\]
rlabel metal2 28658 4284 28658 4284 0 ct.oc.data_chain\[173\]
rlabel metal2 18446 11288 18446 11288 0 ct.oc.data_chain\[174\]
rlabel metal1 20838 6664 20838 6664 0 ct.oc.data_chain\[175\]
rlabel metal1 5014 2074 5014 2074 0 ct.oc.data_chain\[176\]
rlabel via2 16606 10659 16606 10659 0 ct.oc.data_chain\[177\]
rlabel metal2 20378 748 20378 748 0 ct.oc.data_chain\[178\]
rlabel metal1 27761 850 27761 850 0 ct.oc.data_chain\[179\]
rlabel metal1 10903 18258 10903 18258 0 ct.oc.data_chain\[17\]
rlabel metal1 28060 1326 28060 1326 0 ct.oc.data_chain\[180\]
rlabel metal1 27301 1938 27301 1938 0 ct.oc.data_chain\[181\]
rlabel via1 16883 11730 16883 11730 0 ct.oc.data_chain\[182\]
rlabel metal1 16997 6766 16997 6766 0 ct.oc.data_chain\[183\]
rlabel metal2 14490 544 14490 544 0 ct.oc.data_chain\[184\]
rlabel metal2 18262 1105 18262 1105 0 ct.oc.data_chain\[185\]
rlabel metal2 19550 646 19550 646 0 ct.oc.data_chain\[186\]
rlabel metal1 26819 2414 26819 2414 0 ct.oc.data_chain\[187\]
rlabel metal1 26451 4114 26451 4114 0 ct.oc.data_chain\[188\]
rlabel metal1 26405 3026 26405 3026 0 ct.oc.data_chain\[189\]
rlabel metal1 9591 20434 9591 20434 0 ct.oc.data_chain\[18\]
rlabel metal1 1518 306 1518 306 0 ct.oc.data_chain\[190\]
rlabel metal2 19734 3519 19734 3519 0 ct.oc.data_chain\[191\]
rlabel metal2 19458 1309 19458 1309 0 ct.oc.data_chain\[192\]
rlabel via2 20746 1003 20746 1003 0 ct.oc.data_chain\[193\]
rlabel metal1 24656 2414 24656 2414 0 ct.oc.data_chain\[194\]
rlabel metal1 24863 6290 24863 6290 0 ct.oc.data_chain\[195\]
rlabel viali 24611 5678 24611 5678 0 ct.oc.data_chain\[196\]
rlabel metal1 24427 4114 24427 4114 0 ct.oc.data_chain\[197\]
rlabel metal2 23506 935 23506 935 0 ct.oc.data_chain\[198\]
rlabel via1 24795 1938 24795 1938 0 ct.oc.data_chain\[199\]
rlabel metal1 10902 17850 10902 17850 0 ct.oc.data_chain\[19\]
rlabel metal1 13708 20978 13708 20978 0 ct.oc.data_chain\[1\]
rlabel via1 23967 1326 23967 1326 0 ct.oc.data_chain\[200\]
rlabel metal1 23967 850 23967 850 0 ct.oc.data_chain\[201\]
rlabel metal1 23969 3537 23969 3537 0 ct.oc.data_chain\[202\]
rlabel metal1 23967 5202 23967 5202 0 ct.oc.data_chain\[203\]
rlabel metal1 22405 5715 22405 5715 0 ct.oc.data_chain\[204\]
rlabel metal1 22609 4590 22609 4590 0 ct.oc.data_chain\[205\]
rlabel metal1 22563 850 22563 850 0 ct.oc.data_chain\[206\]
rlabel metal1 23691 3026 23691 3026 0 ct.oc.data_chain\[207\]
rlabel metal1 21115 1938 21115 1938 0 ct.oc.data_chain\[208\]
rlabel metal1 21575 1326 21575 1326 0 ct.oc.data_chain\[209\]
rlabel viali 6303 20910 6303 20910 0 ct.oc.data_chain\[20\]
rlabel viali 21761 3511 21761 3511 0 ct.oc.data_chain\[210\]
rlabel metal1 20425 4114 20425 4114 0 ct.oc.data_chain\[211\]
rlabel metal1 20585 6290 20585 6290 0 ct.oc.data_chain\[212\]
rlabel viali 21399 5184 21399 5184 0 ct.oc.data_chain\[213\]
rlabel metal1 21713 2414 21713 2414 0 ct.oc.data_chain\[214\]
rlabel metal1 21115 3026 21115 3026 0 ct.oc.data_chain\[215\]
rlabel via1 19183 1938 19183 1938 0 ct.oc.data_chain\[216\]
rlabel viali 18815 1326 18815 1326 0 ct.oc.data_chain\[217\]
rlabel metal1 18817 3537 18817 3537 0 ct.oc.data_chain\[218\]
rlabel metal1 18492 4794 18492 4794 0 ct.oc.data_chain\[219\]
rlabel viali 6303 19822 6303 19822 0 ct.oc.data_chain\[21\]
rlabel metal1 18677 5202 18677 5202 0 ct.oc.data_chain\[220\]
rlabel viali 18823 4608 18823 4608 0 ct.oc.data_chain\[221\]
rlabel viali 18815 2414 18815 2414 0 ct.oc.data_chain\[222\]
rlabel metal1 18631 3026 18631 3026 0 ct.oc.data_chain\[223\]
rlabel metal1 16055 1938 16055 1938 0 ct.oc.data_chain\[224\]
rlabel viali 16607 1326 16607 1326 0 ct.oc.data_chain\[225\]
rlabel metal1 16609 3537 16609 3537 0 ct.oc.data_chain\[226\]
rlabel metal1 16721 4590 16721 4590 0 ct.oc.data_chain\[227\]
rlabel metal1 16192 5338 16192 5338 0 ct.oc.data_chain\[228\]
rlabel metal1 16285 5202 16285 5202 0 ct.oc.data_chain\[229\]
rlabel metal1 5659 19346 5659 19346 0 ct.oc.data_chain\[22\]
rlabel viali 16607 2414 16607 2414 0 ct.oc.data_chain\[230\]
rlabel metal1 16147 3026 16147 3026 0 ct.oc.data_chain\[231\]
rlabel metal1 14177 1938 14177 1938 0 ct.oc.data_chain\[232\]
rlabel metal1 14169 1326 14169 1326 0 ct.oc.data_chain\[233\]
rlabel metal1 14309 3537 14309 3537 0 ct.oc.data_chain\[234\]
rlabel metal1 14309 5713 14309 5713 0 ct.oc.data_chain\[235\]
rlabel metal1 14077 5202 14077 5202 0 ct.oc.data_chain\[236\]
rlabel metal1 14309 4625 14309 4625 0 ct.oc.data_chain\[237\]
rlabel metal1 13708 2074 13708 2074 0 ct.oc.data_chain\[238\]
rlabel metal1 13801 3026 13801 3026 0 ct.oc.data_chain\[239\]
rlabel metal1 4761 20434 4761 20434 0 ct.oc.data_chain\[23\]
rlabel metal1 11455 1326 11455 1326 0 ct.oc.data_chain\[240\]
rlabel metal1 11178 646 11178 646 0 ct.oc.data_chain\[241\]
rlabel metal1 11362 2278 11362 2278 0 ct.oc.data_chain\[242\]
rlabel metal1 10994 4794 10994 4794 0 ct.oc.data_chain\[243\]
rlabel metal1 11455 5202 11455 5202 0 ct.oc.data_chain\[244\]
rlabel metal1 12052 4250 12052 4250 0 ct.oc.data_chain\[245\]
rlabel metal1 11455 1938 11455 1938 0 ct.oc.data_chain\[246\]
rlabel metal1 11455 3026 11455 3026 0 ct.oc.data_chain\[247\]
rlabel metal1 8694 986 8694 986 0 ct.oc.data_chain\[248\]
rlabel metal2 7314 1564 7314 1564 0 ct.oc.data_chain\[249\]
rlabel metal1 9157 17136 9157 17136 0 ct.oc.data_chain\[24\]
rlabel viali 9155 2414 9155 2414 0 ct.oc.data_chain\[250\]
rlabel metal1 9269 4590 9269 4590 0 ct.oc.data_chain\[251\]
rlabel metal1 9479 5202 9479 5202 0 ct.oc.data_chain\[252\]
rlabel metal1 10259 4114 10259 4114 0 ct.oc.data_chain\[253\]
rlabel via1 9523 1938 9523 1938 0 ct.oc.data_chain\[254\]
rlabel metal1 8879 3026 8879 3026 0 ct.oc.data_chain\[255\]
rlabel metal4 17940 5916 17940 5916 0 ct.oc.data_chain\[256\]
rlabel metal1 3496 2074 3496 2074 0 ct.oc.data_chain\[257\]
rlabel metal1 6949 2449 6949 2449 0 ct.oc.data_chain\[258\]
rlabel metal1 8189 3502 8189 3502 0 ct.oc.data_chain\[259\]
rlabel metal1 8741 18258 8741 18258 0 ct.oc.data_chain\[25\]
rlabel metal1 6303 5202 6303 5202 0 ct.oc.data_chain\[260\]
rlabel metal1 8188 4794 8188 4794 0 ct.oc.data_chain\[261\]
rlabel viali 6947 1344 6947 1344 0 ct.oc.data_chain\[262\]
rlabel metal1 7222 2074 7222 2074 0 ct.oc.data_chain\[263\]
rlabel via1 16607 7854 16607 7854 0 ct.oc.data_chain\[264\]
rlabel metal1 1817 1870 1817 1870 0 ct.oc.data_chain\[265\]
rlabel metal1 3934 3504 3934 3504 0 ct.oc.data_chain\[266\]
rlabel metal1 5981 4114 5981 4114 0 ct.oc.data_chain\[267\]
rlabel metal1 5083 5202 5083 5202 0 ct.oc.data_chain\[268\]
rlabel metal1 6693 4590 6693 4590 0 ct.oc.data_chain\[269\]
rlabel metal1 8741 19346 8741 19346 0 ct.oc.data_chain\[26\]
rlabel metal1 1840 1361 1840 1361 0 ct.oc.data_chain\[270\]
rlabel metal1 6026 2346 6026 2346 0 ct.oc.data_chain\[271\]
rlabel metal2 1978 18122 1978 18122 0 ct.oc.data_chain\[272\]
rlabel metal1 2323 13906 2323 13906 0 ct.oc.data_chain\[273\]
rlabel metal1 1978 3536 1978 3536 0 ct.oc.data_chain\[274\]
rlabel via1 4003 4590 4003 4590 0 ct.oc.data_chain\[275\]
rlabel metal1 4531 4114 4531 4114 0 ct.oc.data_chain\[276\]
rlabel metal1 3542 5338 3542 5338 0 ct.oc.data_chain\[277\]
rlabel metal1 2829 8942 2829 8942 0 ct.oc.data_chain\[278\]
rlabel metal1 2323 3026 2323 3026 0 ct.oc.data_chain\[279\]
rlabel metal1 9157 17681 9157 17681 0 ct.oc.data_chain\[27\]
rlabel via2 3358 7939 3358 7939 0 ct.oc.data_chain\[280\]
rlabel metal1 2254 4591 2254 4591 0 ct.oc.data_chain\[281\]
rlabel viali 1462 4105 1462 4105 0 ct.oc.data_chain\[282\]
rlabel metal1 1978 5712 1978 5712 0 ct.oc.data_chain\[283\]
rlabel metal1 2116 6290 2116 6290 0 ct.oc.data_chain\[284\]
rlabel metal1 1610 5168 1610 5168 0 ct.oc.data_chain\[285\]
rlabel metal1 3589 8466 3589 8466 0 ct.oc.data_chain\[286\]
rlabel metal1 1840 2449 1840 2449 0 ct.oc.data_chain\[287\]
rlabel metal1 1886 7888 1886 7888 0 ct.oc.data_chain\[288\]
rlabel metal1 2231 7378 2231 7378 0 ct.oc.data_chain\[289\]
rlabel metal1 3496 20026 3496 20026 0 ct.oc.data_chain\[28\]
rlabel metal1 3358 8432 3358 8432 0 ct.oc.data_chain\[290\]
rlabel metal1 3933 6290 3933 6290 0 ct.oc.data_chain\[291\]
rlabel metal1 5037 6766 5037 6766 0 ct.oc.data_chain\[292\]
rlabel metal1 4117 7854 4117 7854 0 ct.oc.data_chain\[293\]
rlabel via2 1794 6749 1794 6749 0 ct.oc.data_chain\[294\]
rlabel metal1 5083 7378 5083 7378 0 ct.oc.data_chain\[295\]
rlabel metal1 13386 7752 13386 7752 0 ct.oc.data_chain\[296\]
rlabel via2 17986 7429 17986 7429 0 ct.oc.data_chain\[297\]
rlabel via2 18078 8347 18078 8347 0 ct.oc.data_chain\[298\]
rlabel metal2 14490 7123 14490 7123 0 ct.oc.data_chain\[299\]
rlabel metal1 4120 19822 4120 19822 0 ct.oc.data_chain\[29\]
rlabel metal1 10442 21080 10442 21080 0 ct.oc.data_chain\[2\]
rlabel metal2 13570 6324 13570 6324 0 ct.oc.data_chain\[300\]
rlabel metal1 9821 6290 9821 6290 0 ct.oc.data_chain\[301\]
rlabel metal2 13478 7616 13478 7616 0 ct.oc.data_chain\[302\]
rlabel metal1 11914 6698 11914 6698 0 ct.oc.data_chain\[303\]
rlabel metal1 14697 7854 14697 7854 0 ct.oc.data_chain\[304\]
rlabel viali 16609 7377 16609 7377 0 ct.oc.data_chain\[305\]
rlabel metal1 16147 8466 16147 8466 0 ct.oc.data_chain\[306\]
rlabel metal1 15249 6290 15249 6290 0 ct.oc.data_chain\[307\]
rlabel via1 14399 7378 14399 7378 0 ct.oc.data_chain\[308\]
rlabel metal2 12374 8636 12374 8636 0 ct.oc.data_chain\[309\]
rlabel metal2 1794 20740 1794 20740 0 ct.oc.data_chain\[30\]
rlabel metal2 13018 8330 13018 8330 0 ct.oc.data_chain\[310\]
rlabel viali 12561 6767 12561 6767 0 ct.oc.data_chain\[311\]
rlabel metal1 14421 10030 14421 10030 0 ct.oc.data_chain\[312\]
rlabel viali 14309 10641 14309 10641 0 ct.oc.data_chain\[313\]
rlabel metal1 14812 12614 14812 12614 0 ct.oc.data_chain\[314\]
rlabel metal1 14605 9554 14605 9554 0 ct.oc.data_chain\[315\]
rlabel metal2 14398 12789 14398 12789 0 ct.oc.data_chain\[316\]
rlabel metal2 10994 9894 10994 9894 0 ct.oc.data_chain\[317\]
rlabel viali 11639 8944 11639 8944 0 ct.oc.data_chain\[318\]
rlabel metal1 11363 9554 11363 9554 0 ct.oc.data_chain\[319\]
rlabel metal1 3405 21522 3405 21522 0 ct.oc.data_chain\[31\]
rlabel viali 13121 12208 13121 12208 0 ct.oc.data_chain\[320\]
rlabel metal2 13018 10948 13018 10948 0 ct.oc.data_chain\[321\]
rlabel metal1 13939 12818 13939 12818 0 ct.oc.data_chain\[322\]
rlabel metal1 13202 11764 13202 11764 0 ct.oc.data_chain\[323\]
rlabel metal1 10764 12138 10764 12138 0 ct.oc.data_chain\[324\]
rlabel viali 9431 9552 9431 9552 0 ct.oc.data_chain\[325\]
rlabel metal1 9914 8466 9914 8466 0 ct.oc.data_chain\[326\]
rlabel metal1 9157 10065 9157 10065 0 ct.oc.data_chain\[327\]
rlabel metal2 10212 12580 10212 12580 0 ct.oc.data_chain\[328\]
rlabel metal1 9983 10642 9983 10642 0 ct.oc.data_chain\[329\]
rlabel metal1 6303 17170 6303 17170 0 ct.oc.data_chain\[32\]
rlabel metal1 9983 13906 9983 13906 0 ct.oc.data_chain\[330\]
rlabel metal1 9384 13430 9384 13430 0 ct.oc.data_chain\[331\]
rlabel metal1 8971 12206 8971 12206 0 ct.oc.data_chain\[332\]
rlabel via1 8143 8942 8143 8942 0 ct.oc.data_chain\[333\]
rlabel metal1 6785 9554 6785 9554 0 ct.oc.data_chain\[334\]
rlabel viali 6949 10031 6949 10031 0 ct.oc.data_chain\[335\]
rlabel viali 6947 12206 6947 12206 0 ct.oc.data_chain\[336\]
rlabel metal1 6625 11118 6625 11118 0 ct.oc.data_chain\[337\]
rlabel metal2 7084 12580 7084 12580 0 ct.oc.data_chain\[338\]
rlabel metal1 6578 12954 6578 12954 0 ct.oc.data_chain\[339\]
rlabel viali 6949 17647 6949 17647 0 ct.oc.data_chain\[33\]
rlabel metal1 6119 12818 6119 12818 0 ct.oc.data_chain\[340\]
rlabel metal1 5751 10642 5751 10642 0 ct.oc.data_chain\[341\]
rlabel metal1 5935 11730 5935 11730 0 ct.oc.data_chain\[342\]
rlabel metal1 5843 8466 5843 8466 0 ct.oc.data_chain\[343\]
rlabel metal1 4005 13329 4005 13329 0 ct.oc.data_chain\[344\]
rlabel metal1 4071 13906 4071 13906 0 ct.oc.data_chain\[345\]
rlabel metal1 3727 11730 3727 11730 0 ct.oc.data_chain\[346\]
rlabel metal1 4325 12818 4325 12818 0 ct.oc.data_chain\[347\]
rlabel viali 4005 12207 4005 12207 0 ct.oc.data_chain\[348\]
rlabel viali 3819 10030 3819 10030 0 ct.oc.data_chain\[349\]
rlabel metal1 5980 17850 5980 17850 0 ct.oc.data_chain\[34\]
rlabel metal1 3405 10642 3405 10642 0 ct.oc.data_chain\[350\]
rlabel metal1 3589 9554 3589 9554 0 ct.oc.data_chain\[351\]
rlabel metal1 6119 18258 6119 18258 0 ct.oc.data_chain\[35\]
rlabel metal1 1800 19856 1800 19856 0 ct.oc.data_chain\[36\]
rlabel metal1 3635 18258 3635 18258 0 ct.oc.data_chain\[37\]
rlabel metal2 3266 18598 3266 18598 0 ct.oc.data_chain\[38\]
rlabel metal2 2806 18870 2806 18870 0 ct.oc.data_chain\[39\]
rlabel metal1 13340 20366 13340 20366 0 ct.oc.data_chain\[3\]
rlabel viali 4416 17169 4416 17169 0 ct.oc.data_chain\[40\]
rlabel metal1 6118 15130 6118 15130 0 ct.oc.data_chain\[41\]
rlabel metal1 4120 17646 4120 17646 0 ct.oc.data_chain\[42\]
rlabel viali 4005 16559 4005 16559 0 ct.oc.data_chain\[43\]
rlabel metal2 2806 16150 2806 16150 0 ct.oc.data_chain\[44\]
rlabel metal1 1978 17680 1978 17680 0 ct.oc.data_chain\[45\]
rlabel metal1 1978 16592 1978 16592 0 ct.oc.data_chain\[46\]
rlabel metal2 2990 17238 2990 17238 0 ct.oc.data_chain\[47\]
rlabel metal1 4117 15470 4117 15470 0 ct.oc.data_chain\[48\]
rlabel metal1 5313 14994 5313 14994 0 ct.oc.data_chain\[49\]
rlabel metal1 6118 21522 6118 21522 0 ct.oc.data_chain\[4\]
rlabel metal1 4117 14382 4117 14382 0 ct.oc.data_chain\[50\]
rlabel metal1 5221 16082 5221 16082 0 ct.oc.data_chain\[51\]
rlabel metal2 2990 15215 2990 15215 0 ct.oc.data_chain\[52\]
rlabel metal1 1978 15504 1978 15504 0 ct.oc.data_chain\[53\]
rlabel metal1 1886 14416 1886 14416 0 ct.oc.data_chain\[54\]
rlabel metal1 10442 17068 10442 17068 0 ct.oc.data_chain\[55\]
rlabel via2 11086 15317 11086 15317 0 ct.oc.data_chain\[56\]
rlabel metal2 13110 15776 13110 15776 0 ct.oc.data_chain\[57\]
rlabel via2 13110 15045 13110 15045 0 ct.oc.data_chain\[58\]
rlabel metal2 13478 15079 13478 15079 0 ct.oc.data_chain\[59\]
rlabel metal1 3634 20366 3634 20366 0 ct.oc.data_chain\[5\]
rlabel metal2 13846 17221 13846 17221 0 ct.oc.data_chain\[60\]
rlabel metal2 11546 16694 11546 16694 0 ct.oc.data_chain\[61\]
rlabel metal1 11270 17544 11270 17544 0 ct.oc.data_chain\[62\]
rlabel via2 12834 16779 12834 16779 0 ct.oc.data_chain\[63\]
rlabel metal1 12213 15470 12213 15470 0 ct.oc.data_chain\[64\]
rlabel metal1 14490 16150 14490 16150 0 ct.oc.data_chain\[65\]
rlabel metal1 14306 14892 14306 14892 0 ct.oc.data_chain\[66\]
rlabel metal1 12213 14382 12213 14382 0 ct.oc.data_chain\[67\]
rlabel metal1 12397 18734 12397 18734 0 ct.oc.data_chain\[68\]
rlabel metal1 11270 17238 11270 17238 0 ct.oc.data_chain\[69\]
rlabel metal1 2714 21488 2714 21488 0 ct.oc.data_chain\[6\]
rlabel metal1 13938 17748 13938 17748 0 ct.oc.data_chain\[70\]
rlabel metal1 12134 16593 12134 16593 0 ct.oc.data_chain\[71\]
rlabel metal1 15157 14994 15157 14994 0 ct.oc.data_chain\[72\]
rlabel metal1 15137 16047 15137 16047 0 ct.oc.data_chain\[73\]
rlabel metal1 14789 13906 14789 13906 0 ct.oc.data_chain\[74\]
rlabel metal1 14421 14382 14421 14382 0 ct.oc.data_chain\[75\]
rlabel viali 14307 16560 14307 16560 0 ct.oc.data_chain\[76\]
rlabel metal1 15571 17170 15571 17170 0 ct.oc.data_chain\[77\]
rlabel metal1 15847 18258 15847 18258 0 ct.oc.data_chain\[78\]
rlabel metal1 15663 15470 15663 15470 0 ct.oc.data_chain\[79\]
rlabel metal2 2162 21658 2162 21658 0 ct.oc.data_chain\[7\]
rlabel metal1 18101 13906 18101 13906 0 ct.oc.data_chain\[80\]
rlabel metal2 21850 15759 21850 15759 0 ct.oc.data_chain\[81\]
rlabel metal2 20746 15232 20746 15232 0 ct.oc.data_chain\[82\]
rlabel metal2 17526 14433 17526 14433 0 ct.oc.data_chain\[83\]
rlabel metal1 19734 17238 19734 17238 0 ct.oc.data_chain\[84\]
rlabel metal1 20654 16150 20654 16150 0 ct.oc.data_chain\[85\]
rlabel metal1 20930 17544 20930 17544 0 ct.oc.data_chain\[86\]
rlabel metal2 19550 16779 19550 16779 0 ct.oc.data_chain\[87\]
rlabel metal2 20470 14399 20470 14399 0 ct.oc.data_chain\[88\]
rlabel metal1 23046 15504 23046 15504 0 ct.oc.data_chain\[89\]
rlabel metal1 11271 19346 11271 19346 0 ct.oc.data_chain\[8\]
rlabel metal1 21758 14892 21758 14892 0 ct.oc.data_chain\[90\]
rlabel metal1 22701 14382 22701 14382 0 ct.oc.data_chain\[91\]
rlabel viali 21794 17672 21794 17672 0 ct.oc.data_chain\[92\]
rlabel metal1 21137 18258 21137 18258 0 ct.oc.data_chain\[93\]
rlabel metal1 22839 16558 22839 16558 0 ct.oc.data_chain\[94\]
rlabel metal2 21206 17731 21206 17731 0 ct.oc.data_chain\[95\]
rlabel viali 24380 16081 24380 16081 0 ct.oc.data_chain\[96\]
rlabel metal1 24021 16558 24021 16558 0 ct.oc.data_chain\[97\]
rlabel metal1 25231 14994 25231 14994 0 ct.oc.data_chain\[98\]
rlabel viali 23969 15471 23969 15471 0 ct.oc.data_chain\[99\]
rlabel via1 12559 19822 12559 19822 0 ct.oc.data_chain\[9\]
rlabel metal1 13779 19278 13779 19278 0 ct.oc.mode_buffer\[0\]
rlabel via1 20289 14790 20289 14790 0 ct.oc.mode_buffer\[10\]
rlabel metal1 25717 18054 25717 18054 0 ct.oc.mode_buffer\[11\]
rlabel via1 27073 20366 27073 20366 0 ct.oc.mode_buffer\[12\]
rlabel metal1 28637 19822 28637 19822 0 ct.oc.mode_buffer\[13\]
rlabel metal1 27465 13702 27465 13702 0 ct.oc.mode_buffer\[14\]
rlabel metal1 26843 8466 26843 8466 0 ct.oc.mode_buffer\[15\]
rlabel metal1 21485 10234 21485 10234 0 ct.oc.mode_buffer\[16\]
rlabel metal1 24659 9350 24659 9350 0 ct.oc.mode_buffer\[17\]
rlabel metal1 17158 9112 17158 9112 0 ct.oc.mode_buffer\[18\]
rlabel metal1 18885 6766 18885 6766 0 ct.oc.mode_buffer\[19\]
rlabel metal1 8789 20230 8789 20230 0 ct.oc.mode_buffer\[1\]
rlabel metal1 24428 6834 24428 6834 0 ct.oc.mode_buffer\[20\]
rlabel metal1 14769 3910 14769 3910 0 ct.oc.mode_buffer\[21\]
rlabel metal1 15272 2278 15272 2278 0 ct.oc.mode_buffer\[22\]
rlabel metal1 16907 782 16907 782 0 ct.oc.mode_buffer\[23\]
rlabel metal1 24153 646 24153 646 0 ct.oc.mode_buffer\[24\]
rlabel metal1 20771 5202 20771 5202 0 ct.oc.mode_buffer\[25\]
rlabel metal1 18955 4998 18955 4998 0 ct.oc.mode_buffer\[26\]
rlabel via1 16609 2618 16609 2618 0 ct.oc.mode_buffer\[27\]
rlabel metal1 14263 2618 14263 2618 0 ct.oc.mode_buffer\[28\]
rlabel metal1 11917 2618 11917 2618 0 ct.oc.mode_buffer\[29\]
rlabel via1 3889 19822 3889 19822 0 ct.oc.mode_buffer\[2\]
rlabel metal1 10031 3910 10031 3910 0 ct.oc.mode_buffer\[30\]
rlabel metal1 8421 3706 8421 3706 0 ct.oc.mode_buffer\[31\]
rlabel metal1 13938 4216 13938 4216 0 ct.oc.mode_buffer\[32\]
rlabel metal1 4211 4046 4211 4046 0 ct.oc.mode_buffer\[33\]
rlabel metal2 1656 2380 1656 2380 0 ct.oc.mode_buffer\[34\]
rlabel via1 1429 8262 1429 8262 0 ct.oc.mode_buffer\[35\]
rlabel via1 9409 7310 9409 7310 0 ct.oc.mode_buffer\[36\]
rlabel metal1 16517 7174 16517 7174 0 ct.oc.mode_buffer\[37\]
rlabel metal1 13018 10506 13018 10506 0 ct.oc.mode_buffer\[38\]
rlabel via1 9341 10234 9341 10234 0 ct.oc.mode_buffer\[39\]
rlabel metal1 1705 20026 1705 20026 0 ct.oc.mode_buffer\[3\]
rlabel metal1 7041 9350 7041 9350 0 ct.oc.mode_buffer\[40\]
rlabel via1 5913 8398 5913 8398 0 ct.oc.mode_buffer\[41\]
rlabel via1 3981 9486 3981 9486 0 ct.oc.mode_buffer\[42\]
rlabel via1 1681 13294 1681 13294 0 ct.oc.mode_buffer\[43\]
rlabel metal1 5158 16762 5158 16762 0 ct.oc.mode_buffer\[4\]
rlabel metal1 1543 15538 1543 15538 0 ct.oc.mode_buffer\[5\]
rlabel metal1 6535 14790 6535 14790 0 ct.oc.mode_buffer\[6\]
rlabel metal1 12101 17850 12101 17850 0 ct.oc.mode_buffer\[7\]
rlabel metal1 14699 17102 14699 17102 0 ct.oc.mode_buffer\[8\]
rlabel metal1 16839 14790 16839 14790 0 ct.oc.mode_buffer\[9\]
rlabel metal1 19366 14960 19366 14960 0 ct.oc.trig_chain\[10\]
rlabel metal2 19826 14382 19826 14382 0 ct.oc.trig_chain\[11\]
rlabel metal2 25806 17136 25806 17136 0 ct.oc.trig_chain\[12\]
rlabel metal1 26680 20434 26680 20434 0 ct.oc.trig_chain\[13\]
rlabel metal1 28014 19822 28014 19822 0 ct.oc.trig_chain\[14\]
rlabel metal1 23782 12750 23782 12750 0 ct.oc.trig_chain\[15\]
rlabel metal1 27738 7854 27738 7854 0 ct.oc.trig_chain\[16\]
rlabel metal1 21206 10098 21206 10098 0 ct.oc.trig_chain\[17\]
rlabel metal1 20010 10506 20010 10506 0 ct.oc.trig_chain\[18\]
rlabel metal1 17250 9010 17250 9010 0 ct.oc.trig_chain\[19\]
rlabel metal1 5520 20366 5520 20366 0 ct.oc.trig_chain\[1\]
rlabel metal1 21482 7242 21482 7242 0 ct.oc.trig_chain\[20\]
rlabel metal1 22494 6290 22494 6290 0 ct.oc.trig_chain\[21\]
rlabel metal1 14122 4046 14122 4046 0 ct.oc.trig_chain\[22\]
rlabel metal1 25760 1394 25760 1394 0 ct.oc.trig_chain\[23\]
rlabel metal1 16422 748 16422 748 0 ct.oc.trig_chain\[24\]
rlabel metal1 21988 4658 21988 4658 0 ct.oc.trig_chain\[25\]
rlabel metal1 21068 2482 21068 2482 0 ct.oc.trig_chain\[26\]
rlabel metal1 18446 2414 18446 2414 0 ct.oc.trig_chain\[27\]
rlabel metal1 16100 2414 16100 2414 0 ct.oc.trig_chain\[28\]
rlabel metal1 13110 2618 13110 2618 0 ct.oc.trig_chain\[29\]
rlabel metal1 10626 20332 10626 20332 0 ct.oc.trig_chain\[2\]
rlabel metal1 11454 2414 11454 2414 0 ct.oc.trig_chain\[30\]
rlabel metal1 8694 2346 8694 2346 0 ct.oc.trig_chain\[31\]
rlabel metal2 7866 4590 7866 4590 0 ct.oc.trig_chain\[32\]
rlabel metal2 15226 6205 15226 6205 0 ct.oc.trig_chain\[33\]
rlabel metal1 966 13974 966 13974 0 ct.oc.trig_chain\[34\]
rlabel metal1 1150 2550 1150 2550 0 ct.oc.trig_chain\[35\]
rlabel metal1 4738 7922 4738 7922 0 ct.oc.trig_chain\[36\]
rlabel metal1 9108 7922 9108 7922 0 ct.oc.trig_chain\[37\]
rlabel metal1 15640 7310 15640 7310 0 ct.oc.trig_chain\[38\]
rlabel metal1 13800 9486 13800 9486 0 ct.oc.trig_chain\[39\]
rlabel metal1 1334 20910 1334 20910 0 ct.oc.trig_chain\[3\]
rlabel metal1 13064 12070 13064 12070 0 ct.oc.trig_chain\[40\]
rlabel metal2 7728 9010 7728 9010 0 ct.oc.trig_chain\[41\]
rlabel metal2 5566 9029 5566 9029 0 ct.oc.trig_chain\[42\]
rlabel metal2 1610 11390 1610 11390 0 ct.oc.trig_chain\[43\]
rlabel metal1 1150 12750 1150 12750 0 ct.oc.trig_chain\[44\]
rlabel metal1 5888 17714 5888 17714 0 ct.oc.trig_chain\[4\]
rlabel metal1 1334 16694 1334 16694 0 ct.oc.trig_chain\[5\]
rlabel metal1 1334 15402 1334 15402 0 ct.oc.trig_chain\[6\]
rlabel metal1 9982 16184 9982 16184 0 ct.oc.trig_chain\[7\]
rlabel metal1 13018 14824 13018 14824 0 ct.oc.trig_chain\[8\]
rlabel metal1 14306 17170 14306 17170 0 ct.oc.trig_chain\[9\]
rlabel metal2 21482 21726 21482 21726 0 ct.ro.counter\[0\]
rlabel metal1 21298 21386 21298 21386 0 ct.ro.counter\[1\]
rlabel metal1 21574 20230 21574 20230 0 ct.ro.counter\[2\]
rlabel metal2 22218 21284 22218 21284 0 ct.ro.counter\[3\]
rlabel metal1 24058 21386 24058 21386 0 ct.ro.counter\[4\]
rlabel metal1 23921 21522 23921 21522 0 ct.ro.counter\[5\]
rlabel metal1 23920 20230 23920 20230 0 ct.ro.counter\[6\]
rlabel metal1 25254 20230 25254 20230 0 ct.ro.counter\[7\]
rlabel metal1 18998 20842 18998 20842 0 ct.ro.counter_n\[0\]
rlabel metal1 20148 20910 20148 20910 0 ct.ro.counter_n\[1\]
rlabel metal1 20422 20434 20422 20434 0 ct.ro.counter_n\[2\]
rlabel metal1 23322 20944 23322 20944 0 ct.ro.counter_n\[3\]
rlabel metal1 23690 20910 23690 20910 0 ct.ro.counter_n\[4\]
rlabel metal1 22816 19822 22816 19822 0 ct.ro.counter_n\[5\]
rlabel metal1 23598 20400 23598 20400 0 ct.ro.counter_n\[6\]
rlabel metal1 25898 20400 25898 20400 0 ct.ro.counter_n\[7\]
rlabel metal1 19918 21658 19918 21658 0 ct.ro.gate
rlabel metal1 23421 19278 23421 19278 0 ct.ro.ring\[0\]
rlabel metal1 19458 21420 19458 21420 0 ct.ro.ring\[1\]
rlabel metal2 16790 21131 16790 21131 0 ct.ro.ring\[2\]
rlabel metal2 16882 15640 16882 15640 0 net1
rlabel metal2 12926 6596 12926 6596 0 net10
rlabel metal2 6026 612 6026 612 0 net11
rlabel metal2 7682 18666 7682 18666 0 net12
rlabel metal1 29486 2482 29486 2482 0 net13
rlabel metal1 18538 18292 18538 18292 0 net14
rlabel metal1 7866 10438 7866 10438 0 net15
rlabel metal2 12604 10132 12604 10132 0 net16
rlabel metal1 12006 21318 12006 21318 0 net17
rlabel metal1 18906 6188 18906 6188 0 net18
rlabel metal2 16606 14059 16606 14059 0 net19
rlabel metal1 29486 12070 29486 12070 0 net2
rlabel metal1 5658 6222 5658 6222 0 net20
rlabel via2 9154 6205 9154 6205 0 net21
rlabel metal3 7222 18904 7222 18904 0 net22
rlabel metal2 18538 5406 18538 5406 0 net23
rlabel metal1 30498 18190 30498 18190 0 net24
rlabel metal1 1058 3468 1058 3468 0 net25
rlabel metal1 1196 17714 1196 17714 0 net26
rlabel metal2 17986 18955 17986 18955 0 net27
rlabel metal1 21804 5746 21804 5746 0 net28
rlabel metal1 29164 13838 29164 13838 0 net29
rlabel metal2 28796 17204 28796 17204 0 net3
rlabel metal1 16100 14450 16100 14450 0 net30
rlabel metal1 874 19890 874 19890 0 net31
rlabel metal2 12834 4250 12834 4250 0 net32
rlabel metal2 9614 18649 9614 18649 0 net33
rlabel metal1 17020 11118 17020 11118 0 net34
rlabel metal1 18446 13396 18446 13396 0 net35
rlabel metal1 21022 13158 21022 13158 0 net36
rlabel metal1 10166 14416 10166 14416 0 net37
rlabel metal1 15318 11118 15318 11118 0 net38
rlabel metal1 11362 19822 11362 19822 0 net39
rlabel metal1 23782 18734 23782 18734 0 net4
rlabel metal2 21068 2380 21068 2380 0 net40
rlabel metal2 20194 14331 20194 14331 0 net41
rlabel metal3 20102 12444 20102 12444 0 net42
rlabel metal1 8234 16558 8234 16558 0 net43
rlabel metal2 8510 19822 8510 19822 0 net44
rlabel metal2 1104 2244 1104 2244 0 net45
rlabel metal2 20746 1615 20746 1615 0 net46
rlabel metal1 15686 13328 15686 13328 0 net47
rlabel metal2 12650 17442 12650 17442 0 net48
rlabel metal2 13662 5100 13662 5100 0 net49
rlabel via2 16330 6851 16330 6851 0 net5
rlabel metal1 13800 6834 13800 6834 0 net50
rlabel metal1 966 21522 966 21522 0 net51
rlabel metal1 19872 2482 19872 2482 0 net52
rlabel metal1 18906 21896 18906 21896 0 net53
rlabel metal1 18998 14926 18998 14926 0 net54
rlabel metal4 7912 22204 7912 22204 0 net55
rlabel metal2 13846 13481 13846 13481 0 net56
rlabel metal1 9890 14518 9890 14518 0 net57
rlabel metal1 9430 13294 9430 13294 0 net58
rlabel metal4 5980 20097 5980 20097 0 net59
rlabel metal1 9246 8500 9246 8500 0 net6
rlabel metal1 11730 13294 11730 13294 0 net60
rlabel metal2 12098 13651 12098 13651 0 net61
rlabel metal2 12926 13617 12926 13617 0 net62
rlabel metal1 8464 9486 8464 9486 0 net7
rlabel metal2 18262 2244 18262 2244 0 net8
rlabel metal2 16422 18207 16422 18207 0 net9
rlabel metal1 25031 20978 25031 20978 0 rst_n
rlabel metal2 16698 17884 16698 17884 0 ui_in[0]
rlabel metal1 16606 18802 16606 18802 0 ui_in[1]
rlabel metal1 16836 18734 16836 18734 0 ui_in[2]
rlabel metal1 19366 15606 19366 15606 0 ui_in[3]
rlabel metal2 20562 21590 20562 21590 0 ui_in[4]
rlabel metal4 23092 22137 23092 22137 0 ui_in[5]
rlabel metal4 22540 17717 22540 17717 0 ui_in[6]
rlabel metal2 29854 12801 29854 12801 0 ui_in[7]
rlabel metal2 6946 21760 6946 21760 0 uio_out[0]
rlabel metal1 12926 20808 12926 20808 0 uio_out[1]
rlabel metal1 10902 21046 10902 21046 0 uio_out[2]
rlabel metal4 10948 21389 10948 21389 0 uio_out[3]
rlabel metal1 6440 21658 6440 21658 0 uio_out[4]
rlabel metal1 4002 20230 4002 20230 0 uio_out[5]
rlabel metal1 3220 21386 3220 21386 0 uio_out[6]
rlabel metal1 2484 21658 2484 21658 0 uio_out[7]
rlabel metal1 18400 21114 18400 21114 0 uo_out[0]
rlabel metal1 16790 17850 16790 17850 0 uo_out[1]
rlabel metal1 16698 20026 16698 20026 0 uo_out[2]
rlabel metal1 16790 18904 16790 18904 0 uo_out[3]
rlabel metal4 14812 22137 14812 22137 0 uo_out[4]
rlabel metal4 14260 22137 14260 22137 0 uo_out[5]
rlabel metal1 15640 20570 15640 20570 0 uo_out[6]
rlabel metal1 14904 20774 14904 20774 0 uo_out[7]
<< properties >>
string FIXED_BBOX 0 0 31464 22304
<< end >>
