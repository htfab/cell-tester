magic
tech sky130A
magscale 1 2
timestamp 1699069426
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 827 203
rect 29 -17 63 21
<< scnmos >>
rect 605 47 635 177
rect 709 47 739 177
rect 509 47 539 131
rect 425 47 455 131
rect 341 47 371 131
rect 257 47 287 131
rect 173 47 203 131
rect 81 47 111 131
<< scpmoshvt >>
rect 81 369 111 497
rect 173 369 203 497
rect 257 369 287 497
rect 341 369 371 497
rect 425 369 455 497
rect 509 369 539 497
rect 605 297 635 497
rect 709 297 739 497
<< ndiff >>
rect 739 47 791 59
rect 739 59 749 93
rect 783 59 791 93
rect 739 93 791 127
rect 739 127 749 161
rect 783 127 791 161
rect 739 161 791 177
rect 539 47 605 59
rect 539 59 561 93
rect 595 59 605 93
rect 539 93 605 131
rect 554 131 605 177
rect 635 47 709 59
rect 635 59 665 93
rect 699 59 709 93
rect 635 93 709 127
rect 635 127 665 161
rect 699 127 709 161
rect 635 161 709 177
rect 111 47 173 131
rect 29 47 81 59
rect 29 59 37 93
rect 71 59 81 93
rect 29 93 81 131
rect 203 47 257 59
rect 203 59 213 93
rect 247 59 257 93
rect 203 93 257 131
rect 287 47 341 131
rect 371 47 425 59
rect 371 59 381 93
rect 415 59 425 93
rect 371 93 425 131
rect 455 47 509 131
<< pdiff >>
rect 635 297 709 315
rect 635 315 665 349
rect 699 315 709 349
rect 635 349 709 383
rect 635 383 665 417
rect 699 383 709 417
rect 635 417 709 451
rect 635 451 665 485
rect 699 451 709 485
rect 635 485 709 497
rect 554 297 605 369
rect 539 369 605 383
rect 539 383 561 417
rect 595 383 605 417
rect 539 417 605 451
rect 539 451 561 485
rect 595 451 605 485
rect 539 485 605 497
rect 455 369 509 497
rect 371 369 425 383
rect 371 383 381 417
rect 415 383 425 417
rect 371 417 425 451
rect 371 451 381 485
rect 415 451 425 485
rect 371 485 425 497
rect 287 369 341 497
rect 203 369 257 451
rect 203 451 213 485
rect 247 451 257 485
rect 203 485 257 497
rect 111 369 173 497
rect 29 369 81 383
rect 29 383 37 417
rect 71 383 81 417
rect 29 417 81 451
rect 29 451 37 485
rect 71 451 81 485
rect 29 485 81 497
rect 739 297 791 315
rect 739 315 749 349
rect 783 315 791 349
rect 739 349 791 383
rect 739 383 749 417
rect 783 383 791 417
rect 739 417 791 451
rect 739 451 749 485
rect 783 451 791 485
rect 739 485 791 497
<< ndiffc >>
rect 749 127 783 161
rect 665 127 699 161
rect 37 59 71 93
rect 665 59 699 93
rect 381 59 415 93
rect 749 59 783 93
rect 213 59 247 93
rect 561 59 595 93
<< pdiffc >>
rect 749 451 783 485
rect 381 451 415 485
rect 665 451 699 485
rect 213 451 247 485
rect 561 451 595 485
rect 37 451 71 485
rect 749 383 783 417
rect 381 383 415 417
rect 561 383 595 417
rect 37 383 71 417
rect 665 383 699 417
rect 749 315 783 349
rect 665 315 699 349
<< poly >>
rect 509 497 539 523
rect 425 497 455 523
rect 341 497 371 523
rect 81 497 111 523
rect 257 497 287 523
rect 173 497 203 523
rect 709 497 739 523
rect 605 497 635 523
rect 173 131 203 199
rect 257 131 287 199
rect 173 199 287 215
rect 173 215 211 249
rect 245 215 287 249
rect 173 249 287 265
rect 173 265 203 369
rect 257 265 287 369
rect 509 131 539 199
rect 497 199 551 215
rect 497 215 507 249
rect 541 215 551 249
rect 497 249 551 265
rect 509 265 539 369
rect 341 131 371 199
rect 425 131 455 199
rect 341 199 455 215
rect 341 215 379 249
rect 413 215 455 249
rect 341 249 455 265
rect 341 265 371 369
rect 425 265 455 369
rect 81 131 111 199
rect 77 199 131 215
rect 77 215 87 249
rect 121 215 131 249
rect 77 249 131 265
rect 81 265 111 369
rect 605 177 635 199
rect 709 177 739 199
rect 593 199 739 215
rect 593 215 603 249
rect 637 215 739 249
rect 593 249 739 265
rect 605 265 635 297
rect 709 265 739 297
rect 173 21 203 47
rect 81 21 111 47
rect 257 21 287 47
rect 341 21 371 47
rect 425 21 455 47
rect 509 21 539 47
rect 605 21 635 47
rect 709 21 739 47
<< polycont >>
rect 507 215 541 249
rect 87 215 121 249
rect 211 215 245 249
rect 379 215 413 249
rect 603 215 637 249
<< locali >>
rect 197 451 213 485
rect 247 451 263 485
rect 197 485 263 527
rect 155 527 213 561
rect 247 527 305 561
rect 799 527 828 561
rect 17 59 37 93
rect 71 59 87 93
rect 365 59 381 93
rect 415 59 431 93
rect 17 93 87 127
rect 365 93 431 127
rect 17 127 615 161
rect 17 161 51 199
rect 581 161 615 199
rect 17 199 51 215
rect 581 199 637 215
rect 17 215 51 249
rect 581 215 603 249
rect 17 249 51 265
rect 603 249 637 265
rect 17 265 51 383
rect 17 383 37 417
rect 71 383 381 417
rect 415 383 431 417
rect 17 417 87 451
rect 365 417 431 451
rect 17 451 37 485
rect 71 451 87 485
rect 365 451 381 485
rect 415 451 431 485
rect 649 59 665 93
rect 699 59 715 93
rect 649 93 715 127
rect 649 127 665 161
rect 699 127 715 161
rect 681 161 715 315
rect 649 315 665 349
rect 699 315 715 349
rect 649 349 715 383
rect 649 383 665 417
rect 699 383 715 417
rect 649 417 715 451
rect 649 451 665 485
rect 699 451 715 485
rect 749 417 783 451
rect 749 349 783 383
rect 87 199 149 215
rect 121 215 149 221
rect 121 221 155 249
rect 489 221 507 249
rect 87 249 155 265
rect 489 249 541 265
rect 121 265 155 315
rect 489 265 523 315
rect 121 315 523 349
rect 749 299 783 315
rect 413 221 431 249
rect 379 249 431 255
rect 379 255 413 265
rect 245 221 339 249
rect 211 249 339 255
rect 211 255 245 265
rect 379 199 413 215
rect 507 199 541 215
rect 211 199 245 215
rect 749 161 783 177
rect 749 93 783 127
rect 799 -17 828 17
rect 63 527 121 561
rect 0 527 29 561
rect 749 485 783 527
rect 707 527 765 561
rect 615 527 673 561
rect 545 383 561 417
rect 595 383 611 417
rect 545 417 611 451
rect 545 451 561 485
rect 595 451 611 485
rect 545 485 611 527
rect 523 527 581 561
rect 431 527 489 561
rect 339 527 397 561
rect 707 -17 765 17
rect 749 17 783 59
rect 523 -17 581 17
rect 615 -17 673 17
rect 545 17 611 59
rect 545 59 561 93
rect 595 59 611 93
rect 431 -17 489 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 197 17 263 59
rect 197 59 213 93
rect 247 59 263 93
rect 0 -17 29 17
rect 63 -17 121 17
<< viali >>
rect 305 527 339 561
rect 765 527 799 561
rect 213 527 247 561
rect 673 527 707 561
rect 121 527 155 561
rect 581 527 615 561
rect 29 527 63 561
rect 489 527 523 561
rect 397 527 431 561
rect 121 -17 155 17
rect 765 -17 799 17
rect 397 -17 431 17
rect 29 -17 63 17
rect 673 -17 707 17
rect 305 -17 339 17
rect 581 -17 615 17
rect 213 -17 247 17
rect 489 -17 523 17
<< metal1 >>
rect 0 496 828 527
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 561 828 592
rect 0 -48 828 -17
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 17 828 48
<< labels >>
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 489 289 523 323 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 673 85 707 119 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 0 -48 828 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 maj3_2
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ht_sc_tt05.gds
string GDS_START 7312
string GDS_END 13216
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
