magic
tech sky130A
magscale 1 2
timestamp 1698676622
<< nwell >>
rect -38 261 2154 582
<< pwell >>
rect 1 21 2115 203
rect 29 -17 63 21
<< locali >>
rect 1587 59 1745 85
rect 1587 85 1813 127
rect 1495 127 1837 161
rect 1495 161 1561 383
rect 1771 161 1837 383
rect 1495 383 1837 417
rect 1587 417 1745 485
rect 299 59 365 85
rect 299 85 433 127
rect 299 127 365 451
rect 115 451 549 485
rect 667 59 825 85
rect 667 85 893 127
rect 575 127 917 161
rect 575 161 641 383
rect 851 161 917 383
rect 575 383 917 417
rect 667 417 825 485
rect 1035 59 1285 85
rect 1035 85 1353 93
rect 1035 93 1101 127
rect 1219 93 1353 127
rect 1035 127 1101 161
rect 1219 127 1377 161
rect 1035 161 1101 383
rect 1311 161 1377 383
rect 1035 383 1101 417
rect 1219 383 1377 417
rect 1035 417 1101 451
rect 1219 417 1285 451
rect 1035 451 1285 485
<< obsli1 >>
rect 2087 527 2116 561
rect 2087 -17 2116 17
rect 1995 527 2053 561
rect 1903 527 1961 561
rect 1811 527 1869 561
rect 1719 527 1777 561
rect 1627 527 1685 561
rect 1535 527 1593 561
rect 1443 527 1501 561
rect 1351 527 1409 561
rect 1259 527 1317 561
rect 1167 527 1225 561
rect 1075 527 1133 561
rect 983 527 1041 561
rect 891 527 949 561
rect 799 527 857 561
rect 707 527 765 561
rect 615 527 673 561
rect 523 527 581 561
rect 431 527 489 561
rect 339 527 397 561
rect 247 527 305 561
rect 155 527 213 561
rect 63 527 121 561
rect 0 527 29 561
rect 1995 -17 2053 17
rect 1903 -17 1961 17
rect 1811 -17 1869 17
rect 1719 -17 1777 17
rect 1627 -17 1685 17
rect 1535 -17 1593 17
rect 1443 -17 1501 17
rect 1351 -17 1409 17
rect 1259 -17 1317 17
rect 1167 -17 1225 17
rect 1075 -17 1133 17
rect 983 -17 1041 17
rect 891 -17 949 17
rect 799 -17 857 17
rect 707 -17 765 17
rect 615 -17 673 17
rect 523 -17 581 17
rect 431 -17 489 17
rect 339 -17 397 17
rect 247 -17 305 17
rect 155 -17 213 17
rect 63 -17 121 17
rect 0 -17 29 17
<< obsli1c >>
rect 673 527 707 561
rect 2053 527 2087 561
rect 1501 527 1535 561
rect 1041 527 1075 561
rect 1777 527 1811 561
rect 29 527 63 561
rect 581 527 615 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1961 527 1995 561
rect 397 527 431 561
rect 949 527 983 561
rect 489 527 523 561
rect 857 527 891 561
rect 305 527 339 561
rect 1869 527 1903 561
rect 121 527 155 561
rect 1593 527 1627 561
rect 1225 527 1259 561
rect 1133 527 1167 561
rect 1685 527 1719 561
rect 213 527 247 561
rect 765 527 799 561
rect 1501 -17 1535 17
rect 2053 -17 2087 17
rect 1961 -17 1995 17
rect 1409 -17 1443 17
rect 1869 -17 1903 17
rect 1317 -17 1351 17
rect 1777 -17 1811 17
rect 1225 -17 1259 17
rect 1685 -17 1719 17
rect 1133 -17 1167 17
rect 1593 -17 1627 17
rect 305 -17 339 17
rect 1041 -17 1075 17
rect 213 -17 247 17
rect 949 -17 983 17
rect 121 -17 155 17
rect 857 -17 891 17
rect 29 -17 63 17
rect 765 -17 799 17
rect 673 -17 707 17
rect 581 -17 615 17
rect 489 -17 523 17
rect 397 -17 431 17
<< metal1 >>
rect 0 496 2116 527
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2116 561
rect 0 561 2116 592
rect 0 -48 2116 -17
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2116 17
rect 0 17 2116 48
<< obsm1 >>
rect 308 88 336 428
rect 124 428 520 456
rect 1044 88 1256 116
rect 1044 116 1072 156
rect 1228 116 1256 156
rect 1044 156 1072 184
rect 1228 156 1348 184
rect 1044 184 1072 360
rect 1320 184 1348 360
rect 1044 360 1072 388
rect 1228 360 1348 388
rect 1044 388 1072 428
rect 1228 388 1256 428
rect 1044 428 1256 456
rect 1596 88 1716 116
rect 1596 116 1624 156
rect 1688 116 1716 156
rect 1504 156 1624 184
rect 1688 156 1808 184
rect 1504 184 1532 360
rect 1780 184 1808 360
rect 1504 360 1624 388
rect 1688 360 1808 388
rect 1596 388 1624 428
rect 1688 388 1716 428
rect 1596 428 1716 456
rect 676 88 796 116
rect 676 116 704 156
rect 768 116 796 156
rect 584 156 704 184
rect 768 156 888 184
rect 584 184 612 360
rect 860 184 888 360
rect 584 360 704 388
rect 768 360 888 388
rect 676 388 704 428
rect 768 388 796 428
rect 676 428 796 456
<< labels >>
rlabel locali s 299 59 365 85 6 CLK
port 5 nsew signal input
rlabel locali s 299 85 433 127 6 CLK
port 5 nsew signal input
rlabel locali s 299 127 365 451 6 CLK
port 5 nsew signal input
rlabel locali s 115 451 549 485 6 CLK
port 5 nsew signal input
rlabel locali s 667 59 825 85 6 D
port 6 nsew signal input
rlabel locali s 667 85 893 127 6 D
port 6 nsew signal input
rlabel locali s 575 127 917 161 6 D
port 6 nsew signal input
rlabel locali s 575 161 641 383 6 D
port 6 nsew signal input
rlabel locali s 851 161 917 383 6 D
port 6 nsew signal input
rlabel locali s 575 383 917 417 6 D
port 6 nsew signal input
rlabel locali s 667 417 825 485 6 D
port 6 nsew signal input
rlabel locali s 1035 59 1285 85 6 RESET_B
port 7 nsew signal input
rlabel locali s 1035 85 1353 93 6 RESET_B
port 7 nsew signal input
rlabel locali s 1035 93 1101 127 6 RESET_B
port 7 nsew signal input
rlabel locali s 1219 93 1353 127 6 RESET_B
port 7 nsew signal input
rlabel locali s 1035 127 1101 161 6 RESET_B
port 7 nsew signal input
rlabel locali s 1219 127 1377 161 6 RESET_B
port 7 nsew signal input
rlabel locali s 1035 161 1101 383 6 RESET_B
port 7 nsew signal input
rlabel locali s 1311 161 1377 383 6 RESET_B
port 7 nsew signal input
rlabel locali s 1035 383 1101 417 6 RESET_B
port 7 nsew signal input
rlabel locali s 1219 383 1377 417 6 RESET_B
port 7 nsew signal input
rlabel locali s 1035 417 1101 451 6 RESET_B
port 7 nsew signal input
rlabel locali s 1219 417 1285 451 6 RESET_B
port 7 nsew signal input
rlabel locali s 1035 451 1285 485 6 RESET_B
port 7 nsew signal input
rlabel locali s 1587 59 1745 85 6 Q
port 8 nsew signal output
rlabel locali s 1587 85 1813 127 6 Q
port 8 nsew signal output
rlabel locali s 1495 127 1837 161 6 Q
port 8 nsew signal output
rlabel locali s 1495 161 1561 383 6 Q
port 8 nsew signal output
rlabel locali s 1771 161 1837 383 6 Q
port 8 nsew signal output
rlabel locali s 1495 383 1837 417 6 Q
port 8 nsew signal output
rlabel locali s 1587 417 1745 485 6 Q
port 8 nsew signal output
rlabel pwell s 30 -17 64 21 6 VNB
port 1 nsew ground bidirectional
rlabel pwell s 1 21 2115 203 6 VNB
port 1 nsew ground bidirectional
rlabel nwell s -38 261 2154 582 6 VPB
port 2 nsew power bidirectional
rlabel metal1 s 0 -48 2116 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2116 592 6 VPWR
port 4 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2116 544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_ht_sc_tt05.gds
string GDS_START 24132
string GDS_END 35092
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
<< end >>
